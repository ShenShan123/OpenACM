module sram_multiplier_system (clk,
    init_done,
    init_enable,
    pe_ce,
    rst_n,
    valid_out,
    data_in,
    data_out);
 input clk;
 output init_done;
 input init_enable;
 input pe_ce;
 input rst_n;
 output valid_out;
 input [15:0] data_in;
 output [31:0] data_out;

 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire \u_multiplier/pp_0 ;
 wire \u_multiplier/pp_30 ;
 wire \u_multiplier/s_0 ;
 wire \u_multiplier/s_30 ;
 wire \u_multiplier/STAGE1/_178_ ;
 wire \u_multiplier/STAGE1/_179_ ;
 wire \u_multiplier/STAGE1/_180_ ;
 wire \u_multiplier/STAGE1/_181_ ;
 wire \u_multiplier/STAGE1/_182_ ;
 wire \u_multiplier/STAGE1/_183_ ;
 wire \u_multiplier/STAGE1/_184_ ;
 wire \u_multiplier/STAGE1/_185_ ;
 wire \u_multiplier/STAGE1/_186_ ;
 wire \u_multiplier/STAGE1/_187_ ;
 wire \u_multiplier/STAGE1/_188_ ;
 wire \u_multiplier/STAGE1/_189_ ;
 wire \u_multiplier/STAGE1/_190_ ;
 wire \u_multiplier/STAGE1/_191_ ;
 wire \u_multiplier/STAGE1/_192_ ;
 wire \u_multiplier/STAGE1/_193_ ;
 wire \u_multiplier/STAGE1/_194_ ;
 wire \u_multiplier/STAGE1/_195_ ;
 wire \u_multiplier/STAGE1/_196_ ;
 wire \u_multiplier/STAGE1/_197_ ;
 wire \u_multiplier/STAGE1/_198_ ;
 wire \u_multiplier/STAGE1/_199_ ;
 wire \u_multiplier/STAGE1/_200_ ;
 wire \u_multiplier/STAGE1/_201_ ;
 wire \u_multiplier/STAGE1/_202_ ;
 wire \u_multiplier/STAGE1/_203_ ;
 wire \u_multiplier/STAGE1/_204_ ;
 wire \u_multiplier/STAGE1/_205_ ;
 wire \u_multiplier/STAGE1/_206_ ;
 wire \u_multiplier/STAGE1/_207_ ;
 wire \u_multiplier/STAGE1/_208_ ;
 wire \u_multiplier/STAGE1/_209_ ;
 wire \u_multiplier/STAGE1/_210_ ;
 wire \u_multiplier/STAGE1/_211_ ;
 wire \u_multiplier/STAGE1/_212_ ;
 wire \u_multiplier/STAGE1/_213_ ;
 wire \u_multiplier/STAGE1/_214_ ;
 wire \u_multiplier/STAGE1/_215_ ;
 wire \u_multiplier/STAGE1/_216_ ;
 wire \u_multiplier/STAGE1/_217_ ;
 wire \u_multiplier/STAGE1/_218_ ;
 wire \u_multiplier/STAGE1/_219_ ;
 wire \u_multiplier/STAGE1/_220_ ;
 wire \u_multiplier/STAGE1/_221_ ;
 wire \u_multiplier/STAGE1/_222_ ;
 wire \u_multiplier/STAGE1/_223_ ;
 wire \u_multiplier/STAGE1/_224_ ;
 wire \u_multiplier/STAGE1/_225_ ;
 wire \u_multiplier/STAGE1/_226_ ;
 wire \u_multiplier/STAGE1/_227_ ;
 wire \u_multiplier/STAGE1/_228_ ;
 wire \u_multiplier/STAGE1/_229_ ;
 wire \u_multiplier/STAGE1/_230_ ;
 wire \u_multiplier/STAGE1/_231_ ;
 wire \u_multiplier/STAGE1/_232_ ;
 wire \u_multiplier/STAGE1/_233_ ;
 wire \u_multiplier/STAGE1/_234_ ;
 wire \u_multiplier/STAGE1/_235_ ;
 wire \u_multiplier/STAGE1/_236_ ;
 wire \u_multiplier/STAGE1/_237_ ;
 wire \u_multiplier/STAGE1/_238_ ;
 wire \u_multiplier/STAGE1/_239_ ;
 wire \u_multiplier/STAGE1/_240_ ;
 wire \u_multiplier/STAGE1/_241_ ;
 wire \u_multiplier/STAGE1/_242_ ;
 wire \u_multiplier/STAGE1/_243_ ;
 wire \u_multiplier/STAGE1/_244_ ;
 wire \u_multiplier/STAGE1/_245_ ;
 wire \u_multiplier/STAGE1/_246_ ;
 wire \u_multiplier/STAGE1/_247_ ;
 wire \u_multiplier/STAGE1/_248_ ;
 wire \u_multiplier/STAGE1/_249_ ;
 wire \u_multiplier/STAGE1/_250_ ;
 wire \u_multiplier/STAGE1/_251_ ;
 wire \u_multiplier/STAGE1/_252_ ;
 wire \u_multiplier/STAGE1/_253_ ;
 wire \u_multiplier/STAGE1/_254_ ;
 wire \u_multiplier/STAGE1/_255_ ;
 wire \u_multiplier/STAGE1/_256_ ;
 wire \u_multiplier/STAGE1/_257_ ;
 wire \u_multiplier/STAGE1/_258_ ;
 wire \u_multiplier/STAGE1/_259_ ;
 wire \u_multiplier/STAGE1/_260_ ;
 wire \u_multiplier/STAGE1/_261_ ;
 wire \u_multiplier/STAGE1/_262_ ;
 wire \u_multiplier/STAGE1/_263_ ;
 wire \u_multiplier/STAGE1/_264_ ;
 wire \u_multiplier/STAGE1/_265_ ;
 wire \u_multiplier/STAGE1/_266_ ;
 wire \u_multiplier/STAGE1/_267_ ;
 wire \u_multiplier/STAGE1/_268_ ;
 wire \u_multiplier/STAGE1/_269_ ;
 wire \u_multiplier/STAGE1/_270_ ;
 wire \u_multiplier/STAGE1/_271_ ;
 wire \u_multiplier/STAGE1/_272_ ;
 wire \u_multiplier/STAGE1/_273_ ;
 wire \u_multiplier/STAGE1/_274_ ;
 wire \u_multiplier/STAGE1/_275_ ;
 wire \u_multiplier/STAGE1/_276_ ;
 wire \u_multiplier/STAGE1/_277_ ;
 wire \u_multiplier/STAGE1/_278_ ;
 wire \u_multiplier/STAGE1/_279_ ;
 wire \u_multiplier/STAGE1/_280_ ;
 wire \u_multiplier/STAGE1/_281_ ;
 wire \u_multiplier/STAGE1/_282_ ;
 wire \u_multiplier/STAGE1/_283_ ;
 wire \u_multiplier/STAGE1/_284_ ;
 wire \u_multiplier/STAGE1/_285_ ;
 wire \u_multiplier/STAGE1/_286_ ;
 wire \u_multiplier/STAGE1/_287_ ;
 wire \u_multiplier/STAGE1/_288_ ;
 wire \u_multiplier/STAGE1/_289_ ;
 wire \u_multiplier/STAGE1/_290_ ;
 wire \u_multiplier/STAGE1/_291_ ;
 wire \u_multiplier/STAGE1/_292_ ;
 wire \u_multiplier/STAGE1/_293_ ;
 wire \u_multiplier/STAGE1/_294_ ;
 wire \u_multiplier/STAGE1/_295_ ;
 wire \u_multiplier/STAGE1/_296_ ;
 wire \u_multiplier/STAGE1/_297_ ;
 wire \u_multiplier/STAGE1/_298_ ;
 wire \u_multiplier/STAGE1/_299_ ;
 wire \u_multiplier/STAGE1/_300_ ;
 wire \u_multiplier/STAGE1/_301_ ;
 wire \u_multiplier/STAGE1/_302_ ;
 wire \u_multiplier/STAGE1/_303_ ;
 wire \u_multiplier/STAGE1/_304_ ;
 wire \u_multiplier/STAGE1/_305_ ;
 wire \u_multiplier/STAGE1/_306_ ;
 wire \u_multiplier/STAGE1/_307_ ;
 wire \u_multiplier/STAGE1/_308_ ;
 wire \u_multiplier/STAGE1/_309_ ;
 wire \u_multiplier/STAGE1/_310_ ;
 wire \u_multiplier/STAGE1/_311_ ;
 wire \u_multiplier/STAGE1/_312_ ;
 wire \u_multiplier/STAGE1/_313_ ;
 wire \u_multiplier/STAGE1/_314_ ;
 wire \u_multiplier/STAGE1/_315_ ;
 wire \u_multiplier/STAGE1/_316_ ;
 wire \u_multiplier/STAGE1/_317_ ;
 wire \u_multiplier/STAGE1/_318_ ;
 wire \u_multiplier/STAGE1/_319_ ;
 wire \u_multiplier/STAGE1/_320_ ;
 wire \u_multiplier/STAGE1/_321_ ;
 wire \u_multiplier/STAGE1/_322_ ;
 wire \u_multiplier/STAGE1/_323_ ;
 wire \u_multiplier/STAGE1/pp_16_c2 ;
 wire \u_multiplier/STAGE1/pp_16_c4 ;
 wire \u_multiplier/STAGE1/pp_16_c6 ;
 wire \u_multiplier/STAGE1/pp_17_c2 ;
 wire \u_multiplier/STAGE1/pp_17_c4 ;
 wire \u_multiplier/STAGE1/pp_17_c6 ;
 wire \u_multiplier/STAGE1/pp_18_c2 ;
 wire \u_multiplier/STAGE1/pp_18_c4 ;
 wire \u_multiplier/STAGE1/pp_19_c2 ;
 wire \u_multiplier/STAGE1/pp_19_c4 ;
 wire \u_multiplier/STAGE1/pp_20_c2 ;
 wire \u_multiplier/STAGE1/pp_21_c2 ;
 wire net60;
 wire \u_multiplier/STAGE1/ACCI1_pp_10/_15_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_10/_16_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_10/_17_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_10/_18_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_10/_19_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_10/_20_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_11_1/_15_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_11_1/_16_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_11_1/_17_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_11_1/_18_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_11_1/_19_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_11_1/_20_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_11_2/_15_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_11_2/_16_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_11_2/_17_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_11_2/_18_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_11_2/_19_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_11_2/_20_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_12_1/_15_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_12_1/_16_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_12_1/_17_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_12_1/_18_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_12_1/_19_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_12_1/_20_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_12_2/_15_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_12_2/_16_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_12_2/_17_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_12_2/_18_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_12_2/_19_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_12_2/_20_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_13_1/_15_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_13_1/_16_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_13_1/_17_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_13_1/_18_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_13_1/_19_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_13_1/_20_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_13_2/_15_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_13_2/_16_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_13_2/_17_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_13_2/_18_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_13_2/_19_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_13_2/_20_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_13_3/_15_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_13_3/_16_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_13_3/_17_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_13_3/_18_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_13_3/_19_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_13_3/_20_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_14_1/_15_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_14_1/_16_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_14_1/_17_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_14_1/_18_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_14_1/_19_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_14_1/_20_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_14_2/_15_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_14_2/_16_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_14_2/_17_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_14_2/_18_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_14_2/_19_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_14_2/_20_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_14_3/_15_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_14_3/_16_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_14_3/_17_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_14_3/_18_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_14_3/_19_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_14_3/_20_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_15_1/_15_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_15_1/_16_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_15_1/_17_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_15_1/_18_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_15_1/_19_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_15_1/_20_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_15_2/_15_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_15_2/_16_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_15_2/_17_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_15_2/_18_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_15_2/_19_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_15_2/_20_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_15_3/_15_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_15_3/_16_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_15_3/_17_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_15_3/_18_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_15_3/_19_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_15_3/_20_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_15_4/_15_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_15_4/_16_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_15_4/_17_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_15_4/_18_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_15_4/_19_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_15_4/_20_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_9/_15_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_9/_16_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_9/_17_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_9/_18_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_9/_19_ ;
 wire \u_multiplier/STAGE1/ACCI1_pp_9/_20_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22/_17_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_16_4/_08_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_16_4/_09_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_16_4/_10_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_16_4/_11_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_19/_08_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_19/_09_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_19/_10_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_19/_11_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_21/_08_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_21/_09_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_21/_10_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_21/_11_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_23/_08_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_23/_09_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_23/_10_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_23/_11_ ;
 wire \u_multiplier/STAGE2/pp_16_c2 ;
 wire \u_multiplier/STAGE2/pp_16_c4 ;
 wire \u_multiplier/STAGE2/pp_17_c2 ;
 wire \u_multiplier/STAGE2/pp_17_c4 ;
 wire \u_multiplier/STAGE2/pp_18_c2 ;
 wire \u_multiplier/STAGE2/pp_18_c4 ;
 wire \u_multiplier/STAGE2/pp_19_c2 ;
 wire \u_multiplier/STAGE2/pp_19_c4 ;
 wire \u_multiplier/STAGE2/pp_20_c2 ;
 wire \u_multiplier/STAGE2/pp_20_c4 ;
 wire \u_multiplier/STAGE2/pp_21_c2 ;
 wire \u_multiplier/STAGE2/pp_21_c4 ;
 wire \u_multiplier/STAGE2/pp_22_c2 ;
 wire \u_multiplier/STAGE2/pp_22_c4 ;
 wire \u_multiplier/STAGE2/pp_23_c2 ;
 wire \u_multiplier/STAGE2/pp_23_c4 ;
 wire \u_multiplier/STAGE2/pp_24_c2 ;
 wire \u_multiplier/STAGE2/pp_24_c4 ;
 wire \u_multiplier/STAGE2/pp_25_c2 ;
 wire net64;
 wire \u_multiplier/STAGE2/ACCI1_pp_10_1/_15_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_10_1/_16_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_10_1/_17_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_10_1/_18_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_10_1/_19_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_10_1/_20_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_10_2/_15_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_10_2/_16_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_10_2/_17_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_10_2/_18_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_10_2/_19_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_10_2/_20_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_11_1/_15_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_11_1/_16_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_11_1/_17_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_11_1/_18_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_11_1/_19_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_11_1/_20_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_11_2/_15_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_11_2/_16_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_11_2/_17_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_11_2/_18_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_11_2/_19_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_11_2/_20_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_12_1/_15_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_12_1/_16_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_12_1/_17_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_12_1/_18_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_12_1/_19_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_12_1/_20_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_12_2/_15_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_12_2/_16_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_12_2/_17_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_12_2/_18_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_12_2/_19_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_12_2/_20_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_13_1/_15_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_13_1/_16_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_13_1/_17_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_13_1/_18_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_13_1/_19_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_13_1/_20_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_13_2/_15_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_13_2/_16_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_13_2/_17_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_13_2/_18_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_13_2/_19_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_13_2/_20_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_14_1/_15_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_14_1/_16_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_14_1/_17_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_14_1/_18_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_14_1/_19_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_14_1/_20_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_14_2/_15_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_14_2/_16_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_14_2/_17_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_14_2/_18_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_14_2/_19_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_14_2/_20_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_15_1/_15_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_15_1/_16_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_15_1/_17_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_15_1/_18_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_15_1/_19_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_15_1/_20_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_15_2/_15_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_15_2/_16_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_15_2/_17_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_15_2/_18_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_15_2/_19_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_15_2/_20_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_5/_15_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_5/_16_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_5/_17_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_5/_18_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_5/_19_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_5/_20_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_6/_15_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_6/_16_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_6/_17_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_6/_18_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_6/_19_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_6/_20_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_7_1/_15_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_7_1/_16_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_7_1/_17_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_7_1/_18_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_7_1/_19_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_7_1/_20_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_7_2/_15_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_7_2/_16_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_7_2/_17_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_7_2/_18_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_7_2/_19_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_7_2/_20_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_8_1/_15_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_8_1/_16_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_8_1/_17_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_8_1/_18_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_8_1/_19_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_8_1/_20_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_8_2/_15_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_8_2/_16_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_8_2/_17_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_8_2/_18_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_8_2/_19_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_8_2/_20_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_9_1/_15_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_9_1/_16_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_9_1/_17_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_9_1/_18_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_9_1/_19_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_9_1/_20_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_9_2/_15_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_9_2/_16_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_9_2/_17_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_9_2/_18_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_9_2/_19_ ;
 wire \u_multiplier/STAGE2/ACCI1_pp_9_2/_20_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_25_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_25_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_25_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_25_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_25_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_25_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_25_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_26_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_26_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_26_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_26_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_26_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_26_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_26_1/_17_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp_25/_08_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp_25/_09_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp_25/_10_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp_25/_11_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp_27/_08_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp_27/_09_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp_27/_10_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp_27/_11_ ;
 wire \u_multiplier/STAGE3/pp_10_c ;
 wire \u_multiplier/STAGE3/pp_10_s ;
 wire \u_multiplier/STAGE3/pp_11_c ;
 wire \u_multiplier/STAGE3/pp_11_s ;
 wire \u_multiplier/STAGE3/pp_12_c ;
 wire \u_multiplier/STAGE3/pp_12_s ;
 wire \u_multiplier/STAGE3/pp_13_c ;
 wire \u_multiplier/STAGE3/pp_13_s ;
 wire \u_multiplier/STAGE3/pp_14_c ;
 wire \u_multiplier/STAGE3/pp_14_s ;
 wire \u_multiplier/STAGE3/pp_15_c ;
 wire \u_multiplier/STAGE3/pp_15_s ;
 wire \u_multiplier/STAGE3/pp_16_c1 ;
 wire \u_multiplier/STAGE3/pp_16_c2 ;
 wire \u_multiplier/STAGE3/pp_16_s ;
 wire \u_multiplier/STAGE3/pp_17_c1 ;
 wire \u_multiplier/STAGE3/pp_17_c2 ;
 wire \u_multiplier/STAGE3/pp_17_s ;
 wire \u_multiplier/STAGE3/pp_18_c1 ;
 wire \u_multiplier/STAGE3/pp_18_c2 ;
 wire \u_multiplier/STAGE3/pp_18_s ;
 wire \u_multiplier/STAGE3/pp_19_c1 ;
 wire \u_multiplier/STAGE3/pp_19_c2 ;
 wire \u_multiplier/STAGE3/pp_19_s ;
 wire \u_multiplier/STAGE3/pp_20_c1 ;
 wire \u_multiplier/STAGE3/pp_20_c2 ;
 wire \u_multiplier/STAGE3/pp_20_s ;
 wire \u_multiplier/STAGE3/pp_21_c1 ;
 wire \u_multiplier/STAGE3/pp_21_c2 ;
 wire \u_multiplier/STAGE3/pp_21_s ;
 wire \u_multiplier/STAGE3/pp_22_c1 ;
 wire \u_multiplier/STAGE3/pp_22_c2 ;
 wire \u_multiplier/STAGE3/pp_22_s ;
 wire \u_multiplier/STAGE3/pp_23_c1 ;
 wire \u_multiplier/STAGE3/pp_23_c2 ;
 wire \u_multiplier/STAGE3/pp_23_s ;
 wire \u_multiplier/STAGE3/pp_24_c1 ;
 wire \u_multiplier/STAGE3/pp_24_c2 ;
 wire \u_multiplier/STAGE3/pp_24_s ;
 wire \u_multiplier/STAGE3/pp_25_c1 ;
 wire \u_multiplier/STAGE3/pp_25_c2 ;
 wire \u_multiplier/STAGE3/pp_25_s ;
 wire \u_multiplier/STAGE3/pp_26_c1 ;
 wire \u_multiplier/STAGE3/pp_26_c2 ;
 wire \u_multiplier/STAGE3/pp_26_s ;
 wire \u_multiplier/STAGE3/pp_27_c1 ;
 wire \u_multiplier/STAGE3/pp_27_c2 ;
 wire \u_multiplier/STAGE3/pp_27_s ;
 wire \u_multiplier/STAGE3/pp_28_c1 ;
 wire \u_multiplier/STAGE3/pp_28_c2 ;
 wire \u_multiplier/STAGE3/pp_28_s ;
 wire \u_multiplier/STAGE3/pp_29_c ;
 wire \u_multiplier/STAGE3/pp_29_s ;
 wire \u_multiplier/STAGE3/pp_2_c ;
 wire \u_multiplier/STAGE3/pp_2_s ;
 wire \u_multiplier/STAGE3/pp_3_c ;
 wire \u_multiplier/STAGE3/pp_3_s ;
 wire \u_multiplier/STAGE3/pp_4_c ;
 wire \u_multiplier/STAGE3/pp_4_s ;
 wire \u_multiplier/STAGE3/pp_5_c ;
 wire \u_multiplier/STAGE3/pp_5_s ;
 wire \u_multiplier/STAGE3/pp_6_c ;
 wire \u_multiplier/STAGE3/pp_6_s ;
 wire \u_multiplier/STAGE3/pp_7_c ;
 wire \u_multiplier/STAGE3/pp_7_s ;
 wire \u_multiplier/STAGE3/pp_8_c ;
 wire \u_multiplier/STAGE3/pp_8_s ;
 wire \u_multiplier/STAGE3/pp_9_c ;
 wire \u_multiplier/STAGE3/pp_9_s ;
 wire net77;
 wire \u_multiplier/STAGE3/ACCI1_pp_10_1/_15_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_10_1/_16_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_10_1/_17_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_10_1/_18_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_10_1/_19_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_10_1/_20_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_11_1/_15_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_11_1/_16_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_11_1/_17_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_11_1/_18_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_11_1/_19_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_11_1/_20_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_12_1/_15_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_12_1/_16_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_12_1/_17_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_12_1/_18_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_12_1/_19_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_12_1/_20_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_13_1/_15_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_13_1/_16_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_13_1/_17_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_13_1/_18_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_13_1/_19_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_13_1/_20_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_14_1/_15_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_14_1/_16_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_14_1/_17_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_14_1/_18_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_14_1/_19_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_14_1/_20_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_15_1/_15_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_15_1/_16_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_15_1/_17_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_15_1/_18_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_15_1/_19_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_15_1/_20_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_3/_15_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_3/_16_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_3/_17_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_3/_18_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_3/_19_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_3/_20_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_4/_15_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_4/_16_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_4/_17_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_4/_18_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_4/_19_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_4/_20_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_5/_15_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_5/_16_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_5/_17_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_5/_18_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_5/_19_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_5/_20_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_6/_15_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_6/_16_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_6/_17_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_6/_18_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_6/_19_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_6/_20_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_7/_15_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_7/_16_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_7/_17_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_7/_18_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_7/_19_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_7/_20_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_8/_15_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_8/_16_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_8/_17_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_8/_18_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_8/_19_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_8/_20_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_9/_15_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_9/_16_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_9/_17_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_9/_18_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_9/_19_ ;
 wire \u_multiplier/STAGE3/ACCI1_pp_9/_20_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_16_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_16_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_16_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_16_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_16_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_16_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_16_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_17_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_17_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_17_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_17_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_17_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_17_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_17_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_18_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_18_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_18_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_18_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_18_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_18_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_18_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_19_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_19_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_19_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_19_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_19_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_19_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_19_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_20_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_20_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_20_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_20_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_20_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_20_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_20_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_21_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_21_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_21_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_21_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_21_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_21_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_21_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_22_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_22_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_22_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_22_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_22_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_22_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_22_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_23_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_23_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_23_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_23_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_23_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_23_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_23_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_24_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_24_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_24_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_24_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_24_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_24_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_24_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_25_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_25_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_25_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_25_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_25_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_25_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_25_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_26_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_26_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_26_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_26_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_26_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_26_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_26_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_27_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_27_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_27_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_27_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_27_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_27_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_27_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_28_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_28_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_28_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_28_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_28_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_28_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_28_1/_17_ ;
 wire \u_multiplier/STAGE3/Final_add/Cout ;
 wire \u_multiplier/STAGE3/Final_add/c1 ;
 wire \u_multiplier/STAGE3/Final_add/cla1/c1 ;
 wire \u_multiplier/STAGE3/Final_add/cla1/c2 ;
 wire \u_multiplier/STAGE3/Final_add/cla1/c3 ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_25_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_26_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_27_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_28_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_29_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_30_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_31_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_32_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_33_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_34_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_35_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_36_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_37_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_38_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_39_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_25_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_26_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_27_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_28_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_29_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_30_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_31_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_32_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_33_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_34_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_35_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_36_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_37_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_38_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_39_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_25_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_26_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_27_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_28_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_29_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_30_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_31_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_32_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_33_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_34_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_35_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_36_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_37_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_38_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_39_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_25_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_26_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_27_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_28_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_29_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_30_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_31_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_32_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_33_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_34_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_35_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_36_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_37_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_38_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_39_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/c1 ;
 wire \u_multiplier/STAGE3/Final_add/cla2/c2 ;
 wire \u_multiplier/STAGE3/Final_add/cla2/c3 ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_25_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_26_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_27_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_28_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_29_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_30_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_31_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_32_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_33_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_34_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_35_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_36_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_37_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_38_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_39_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_25_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_26_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_27_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_28_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_29_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_30_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_31_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_32_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_33_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_34_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_35_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_36_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_37_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_38_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_39_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_25_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_26_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_27_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_28_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_29_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_30_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_31_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_32_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_33_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_34_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_35_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_36_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_37_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_38_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_39_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_25_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_26_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_27_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_28_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_29_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_30_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_31_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_32_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_33_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_34_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_35_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_36_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_37_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_38_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_39_ ;
 wire \u_multiplier/STAGE3/Full_adder_pp_29/_08_ ;
 wire \u_multiplier/STAGE3/Full_adder_pp_29/_09_ ;
 wire \u_multiplier/STAGE3/Full_adder_pp_29/_10_ ;
 wire \u_multiplier/STAGE3/Full_adder_pp_29/_11_ ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire valid_reg_out;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net61;
 wire net62;
 wire net63;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire clknet_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire [4:0] addr_ptr;
 wire [2:0] curr_state;
 wire [15:0] data_in_reg;
 wire [4:0] init_count;
 wire [31:0] product;
 wire [15:0] sram_rdata;
 wire [15:0] sram_rdata_reg;
 wire [1:0] \u_multiplier/pp_1 ;
 wire [7:0] \u_multiplier/pp_10 ;
 wire [7:0] \u_multiplier/pp_11 ;
 wire [7:0] \u_multiplier/pp_12 ;
 wire [7:0] \u_multiplier/pp_13 ;
 wire [7:0] \u_multiplier/pp_14 ;
 wire [7:0] \u_multiplier/pp_15 ;
 wire [7:0] \u_multiplier/pp_16 ;
 wire [7:0] \u_multiplier/pp_17 ;
 wire [7:0] \u_multiplier/pp_18 ;
 wire [7:0] \u_multiplier/pp_19 ;
 wire [2:0] \u_multiplier/pp_2 ;
 wire [7:0] \u_multiplier/pp_20 ;
 wire [7:0] \u_multiplier/pp_21 ;
 wire [7:0] \u_multiplier/pp_22 ;
 wire [7:0] \u_multiplier/pp_23 ;
 wire [7:0] \u_multiplier/pp_24 ;
 wire [5:0] \u_multiplier/pp_25 ;
 wire [4:0] \u_multiplier/pp_26 ;
 wire [3:0] \u_multiplier/pp_27 ;
 wire [2:0] \u_multiplier/pp_28 ;
 wire [1:0] \u_multiplier/pp_29 ;
 wire [3:0] \u_multiplier/pp_3 ;
 wire [4:0] \u_multiplier/pp_4 ;
 wire [5:0] \u_multiplier/pp_5 ;
 wire [6:0] \u_multiplier/pp_6 ;
 wire [7:0] \u_multiplier/pp_7 ;
 wire [7:0] \u_multiplier/pp_8 ;
 wire [7:0] \u_multiplier/pp_9 ;
 wire [1:0] \u_multiplier/s_1 ;
 wire [3:0] \u_multiplier/s_10 ;
 wire [3:0] \u_multiplier/s_11 ;
 wire [3:0] \u_multiplier/s_12 ;
 wire [3:0] \u_multiplier/s_13 ;
 wire [3:0] \u_multiplier/s_14 ;
 wire [3:0] \u_multiplier/s_15 ;
 wire [3:0] \u_multiplier/s_16 ;
 wire [3:0] \u_multiplier/s_17 ;
 wire [3:0] \u_multiplier/s_18 ;
 wire [3:0] \u_multiplier/s_19 ;
 wire [2:0] \u_multiplier/s_2 ;
 wire [3:0] \u_multiplier/s_20 ;
 wire [3:0] \u_multiplier/s_21 ;
 wire [3:0] \u_multiplier/s_22 ;
 wire [3:0] \u_multiplier/s_23 ;
 wire [3:0] \u_multiplier/s_24 ;
 wire [3:0] \u_multiplier/s_25 ;
 wire [3:0] \u_multiplier/s_26 ;
 wire [3:0] \u_multiplier/s_27 ;
 wire [3:0] \u_multiplier/s_28 ;
 wire [1:0] \u_multiplier/s_29 ;
 wire [3:0] \u_multiplier/s_3 ;
 wire [3:0] \u_multiplier/s_4 ;
 wire [3:0] \u_multiplier/s_5 ;
 wire [3:0] \u_multiplier/s_6 ;
 wire [3:0] \u_multiplier/s_7 ;
 wire [3:0] \u_multiplier/s_8 ;
 wire [3:0] \u_multiplier/s_9 ;

 INV_X1 _420_ (.A(net19),
    .ZN(_238_));
 INV_X1 _421_ (.A(net18),
    .ZN(_195_));
 INV_X1 _422_ (.A(curr_state[2]),
    .ZN(_239_));
 INV_X1 _423_ (.A(_408_),
    .ZN(_240_));
 INV_X1 _424_ (.A(addr_ptr[0]),
    .ZN(_241_));
 INV_X1 _425_ (.A(_401_),
    .ZN(_242_));
 AND2_X4 _426_ (.A1(net19),
    .A2(net20),
    .ZN(_191_));
 INV_X1 _427_ (.A(_191_),
    .ZN(_243_));
 NAND2_X1 _428_ (.A1(net19),
    .A2(net141),
    .ZN(_196_));
 NAND2_X1 _429_ (.A1(init_count[1]),
    .A2(init_count[0]),
    .ZN(_244_));
 AND3_X1 _430_ (.A1(init_count[1]),
    .A2(init_count[0]),
    .A3(init_count[2]),
    .ZN(_245_));
 AND4_X2 _431_ (.A1(init_count[1]),
    .A2(init_count[0]),
    .A3(init_count[3]),
    .A4(init_count[2]),
    .ZN(_246_));
 AND3_X1 _432_ (.A1(net18),
    .A2(init_count[4]),
    .A3(_246_),
    .ZN(_247_));
 NOR2_X1 _433_ (.A1(_191_),
    .A2(_247_),
    .ZN(_248_));
 AOI21_X1 _434_ (.A(_248_),
    .B1(_196_),
    .B2(_243_),
    .ZN(_193_));
 NOR2_X2 _435_ (.A1(_238_),
    .A2(_195_),
    .ZN(_249_));
 NAND2_X2 _436_ (.A1(net19),
    .A2(net18),
    .ZN(_250_));
 NAND3_X1 _437_ (.A1(net17),
    .A2(net105),
    .A3(_249_),
    .ZN(_251_));
 OAI21_X1 _438_ (.A(net106),
    .B1(_247_),
    .B2(_196_),
    .ZN(_194_));
 AOI22_X1 _439_ (.A1(net19),
    .A2(net79),
    .B1(_249_),
    .B2(net17),
    .ZN(_192_));
 AND2_X1 _440_ (.A1(net19),
    .A2(sram_rdata[0]),
    .ZN(_175_));
 AND2_X1 _441_ (.A1(net19),
    .A2(sram_rdata[1]),
    .ZN(_182_));
 AND2_X1 _442_ (.A1(net19),
    .A2(sram_rdata[2]),
    .ZN(_183_));
 AND2_X1 _443_ (.A1(net19),
    .A2(sram_rdata[3]),
    .ZN(_184_));
 AND2_X1 _444_ (.A1(net19),
    .A2(sram_rdata[4]),
    .ZN(_185_));
 AND2_X1 _445_ (.A1(net19),
    .A2(sram_rdata[5]),
    .ZN(_186_));
 AND2_X1 _446_ (.A1(net19),
    .A2(sram_rdata[6]),
    .ZN(_187_));
 AND2_X1 _447_ (.A1(net19),
    .A2(sram_rdata[7]),
    .ZN(_188_));
 AND2_X1 _448_ (.A1(net19),
    .A2(sram_rdata[8]),
    .ZN(_189_));
 AND2_X1 _449_ (.A1(net19),
    .A2(sram_rdata[9]),
    .ZN(_190_));
 AND2_X1 _450_ (.A1(net19),
    .A2(sram_rdata[10]),
    .ZN(_176_));
 AND2_X1 _451_ (.A1(net19),
    .A2(sram_rdata[11]),
    .ZN(_177_));
 AND2_X1 _452_ (.A1(net19),
    .A2(sram_rdata[12]),
    .ZN(_178_));
 AND2_X1 _453_ (.A1(net19),
    .A2(sram_rdata[13]),
    .ZN(_179_));
 AND2_X1 _454_ (.A1(net19),
    .A2(sram_rdata[14]),
    .ZN(_180_));
 AND2_X1 _455_ (.A1(net19),
    .A2(sram_rdata[15]),
    .ZN(_181_));
 AND2_X1 _456_ (.A1(product[0]),
    .A2(_191_),
    .ZN(_138_));
 AND2_X1 _457_ (.A1(product[1]),
    .A2(_191_),
    .ZN(_149_));
 AND2_X1 _458_ (.A1(product[2]),
    .A2(_191_),
    .ZN(_160_));
 AND2_X1 _459_ (.A1(product[3]),
    .A2(_191_),
    .ZN(_163_));
 AND2_X1 _460_ (.A1(product[4]),
    .A2(_191_),
    .ZN(_164_));
 AND2_X1 _461_ (.A1(product[5]),
    .A2(_191_),
    .ZN(_165_));
 AND2_X1 _462_ (.A1(product[6]),
    .A2(_191_),
    .ZN(_166_));
 AND2_X1 _463_ (.A1(product[7]),
    .A2(_191_),
    .ZN(_167_));
 AND2_X1 _464_ (.A1(product[8]),
    .A2(_191_),
    .ZN(_168_));
 AND2_X1 _465_ (.A1(product[9]),
    .A2(_191_),
    .ZN(_169_));
 AND2_X1 _466_ (.A1(product[10]),
    .A2(_191_),
    .ZN(_139_));
 AND2_X1 _467_ (.A1(product[11]),
    .A2(_191_),
    .ZN(_140_));
 AND2_X1 _468_ (.A1(product[12]),
    .A2(_191_),
    .ZN(_141_));
 AND2_X1 _469_ (.A1(product[13]),
    .A2(_191_),
    .ZN(_142_));
 AND2_X1 _470_ (.A1(product[14]),
    .A2(_191_),
    .ZN(_143_));
 AND2_X1 _471_ (.A1(product[15]),
    .A2(_191_),
    .ZN(_144_));
 AND2_X1 _472_ (.A1(product[16]),
    .A2(_191_),
    .ZN(_145_));
 AND2_X1 _473_ (.A1(product[17]),
    .A2(_191_),
    .ZN(_146_));
 AND2_X1 _474_ (.A1(product[18]),
    .A2(_191_),
    .ZN(_147_));
 AND2_X1 _475_ (.A1(product[19]),
    .A2(_191_),
    .ZN(_148_));
 AND2_X1 _476_ (.A1(product[20]),
    .A2(_191_),
    .ZN(_150_));
 AND2_X1 _477_ (.A1(product[21]),
    .A2(_191_),
    .ZN(_151_));
 AND2_X1 _478_ (.A1(product[22]),
    .A2(_191_),
    .ZN(_152_));
 AND2_X1 _479_ (.A1(product[23]),
    .A2(_191_),
    .ZN(_153_));
 AND2_X1 _480_ (.A1(product[24]),
    .A2(_191_),
    .ZN(_154_));
 AND2_X1 _481_ (.A1(product[25]),
    .A2(_191_),
    .ZN(_155_));
 AND2_X1 _482_ (.A1(product[26]),
    .A2(_191_),
    .ZN(_156_));
 AND2_X1 _483_ (.A1(product[27]),
    .A2(_191_),
    .ZN(_157_));
 AND2_X1 _484_ (.A1(product[28]),
    .A2(_191_),
    .ZN(_158_));
 AND2_X1 _485_ (.A1(product[29]),
    .A2(_191_),
    .ZN(_159_));
 AND2_X1 _486_ (.A1(product[30]),
    .A2(_191_),
    .ZN(_161_));
 AND2_X1 _487_ (.A1(product[31]),
    .A2(_191_),
    .ZN(_162_));
 AND2_X1 _488_ (.A1(net19),
    .A2(net1),
    .ZN(_122_));
 AND2_X1 _489_ (.A1(net19),
    .A2(net8),
    .ZN(_129_));
 AND2_X1 _490_ (.A1(net19),
    .A2(net9),
    .ZN(_130_));
 AND2_X1 _491_ (.A1(net19),
    .A2(net10),
    .ZN(_131_));
 AND2_X1 _492_ (.A1(net19),
    .A2(net11),
    .ZN(_132_));
 AND2_X1 _493_ (.A1(net19),
    .A2(net12),
    .ZN(_133_));
 AND2_X1 _494_ (.A1(net19),
    .A2(net13),
    .ZN(_134_));
 AND2_X1 _495_ (.A1(net19),
    .A2(net14),
    .ZN(_135_));
 AND2_X1 _496_ (.A1(net19),
    .A2(net15),
    .ZN(_136_));
 AND2_X1 _497_ (.A1(net19),
    .A2(net16),
    .ZN(_137_));
 AND2_X1 _498_ (.A1(net19),
    .A2(net2),
    .ZN(_123_));
 AND2_X1 _499_ (.A1(net19),
    .A2(net3),
    .ZN(_124_));
 AND2_X1 _500_ (.A1(net19),
    .A2(net4),
    .ZN(_125_));
 AND2_X1 _501_ (.A1(net19),
    .A2(net5),
    .ZN(_126_));
 AND2_X1 _502_ (.A1(net19),
    .A2(net6),
    .ZN(_127_));
 AND2_X1 _503_ (.A1(net19),
    .A2(net7),
    .ZN(_128_));
 NAND2_X2 _504_ (.A1(net19),
    .A2(_195_),
    .ZN(_252_));
 NAND2_X2 _505_ (.A1(_240_),
    .A2(_246_),
    .ZN(_253_));
 XNOR2_X1 _506_ (.A(net115),
    .B(_253_),
    .ZN(_254_));
 AOI22_X1 _507_ (.A1(init_count[0]),
    .A2(net20),
    .B1(_254_),
    .B2(curr_state[2]),
    .ZN(_255_));
 OAI22_X1 _508_ (.A1(net116),
    .A2(_252_),
    .B1(_255_),
    .B2(_250_),
    .ZN(_170_));
 XNOR2_X1 _509_ (.A(init_count[1]),
    .B(init_count[0]),
    .ZN(_256_));
 AOI21_X1 _510_ (.A(_239_),
    .B1(_253_),
    .B2(_256_),
    .ZN(_257_));
 AOI21_X1 _511_ (.A(_257_),
    .B1(net20),
    .B2(init_count[1]),
    .ZN(_258_));
 OAI22_X1 _512_ (.A1(net99),
    .A2(_252_),
    .B1(_258_),
    .B2(_250_),
    .ZN(_171_));
 XNOR2_X1 _513_ (.A(_406_),
    .B(_244_),
    .ZN(_259_));
 AOI21_X1 _514_ (.A(_239_),
    .B1(_253_),
    .B2(_259_),
    .ZN(_260_));
 AOI21_X1 _515_ (.A(_260_),
    .B1(net20),
    .B2(init_count[2]),
    .ZN(_261_));
 OAI22_X1 _516_ (.A1(net102),
    .A2(_252_),
    .B1(_261_),
    .B2(_250_),
    .ZN(_172_));
 OAI21_X1 _517_ (.A(curr_state[2]),
    .B1(_245_),
    .B2(init_count[3]),
    .ZN(_262_));
 AOI21_X1 _518_ (.A(_262_),
    .B1(_246_),
    .B2(_408_),
    .ZN(_263_));
 AOI21_X1 _519_ (.A(_263_),
    .B1(net20),
    .B2(init_count[3]),
    .ZN(_264_));
 OAI22_X1 _520_ (.A1(net77),
    .A2(_252_),
    .B1(_264_),
    .B2(_250_),
    .ZN(_173_));
 AND2_X1 _521_ (.A1(init_count[4]),
    .A2(net20),
    .ZN(_265_));
 OAI221_X1 _522_ (.A(_249_),
    .B1(_265_),
    .B2(curr_state[2]),
    .C1(_246_),
    .C2(init_count[4]),
    .ZN(_266_));
 OAI21_X1 _523_ (.A(_266_),
    .B1(_252_),
    .B2(net124),
    .ZN(_174_));
 AND2_X1 _524_ (.A1(curr_state[2]),
    .A2(net108),
    .ZN(_267_));
 AOI22_X1 _525_ (.A1(net20),
    .A2(_241_),
    .B1(_253_),
    .B2(_267_),
    .ZN(_268_));
 OAI22_X1 _526_ (.A1(net109),
    .A2(_252_),
    .B1(_268_),
    .B2(_250_),
    .ZN(_117_));
 AOI21_X2 _527_ (.A(_239_),
    .B1(_246_),
    .B2(init_count[4]),
    .ZN(_269_));
 AND2_X1 _528_ (.A1(addr_ptr[0]),
    .A2(addr_ptr[1]),
    .ZN(_270_));
 NOR2_X1 _529_ (.A1(_250_),
    .A2(_270_),
    .ZN(_271_));
 OAI221_X1 _530_ (.A(_271_),
    .B1(addr_ptr[1]),
    .B2(addr_ptr[0]),
    .C1(net20),
    .C2(_269_),
    .ZN(_272_));
 OAI21_X1 _531_ (.A(_272_),
    .B1(_252_),
    .B2(net94),
    .ZN(_118_));
 NAND4_X1 _532_ (.A1(addr_ptr[3]),
    .A2(addr_ptr[2]),
    .A3(addr_ptr[4]),
    .A4(_270_),
    .ZN(_273_));
 AOI21_X2 _533_ (.A(_269_),
    .B1(_273_),
    .B2(net20),
    .ZN(_274_));
 XNOR2_X1 _534_ (.A(net112),
    .B(_270_),
    .ZN(_275_));
 NAND2_X1 _535_ (.A1(_249_),
    .A2(_275_),
    .ZN(_276_));
 OAI22_X1 _536_ (.A1(net113),
    .A2(_252_),
    .B1(_274_),
    .B2(_276_),
    .ZN(_119_));
 NAND3_X1 _537_ (.A1(net18),
    .A2(_242_),
    .A3(_270_),
    .ZN(_277_));
 XNOR2_X1 _538_ (.A(net132),
    .B(_277_),
    .ZN(_278_));
 AOI211_X1 _539_ (.A(_238_),
    .B(net133),
    .C1(_274_),
    .C2(net18),
    .ZN(_120_));
 NAND4_X1 _540_ (.A1(net18),
    .A2(addr_ptr[3]),
    .A3(addr_ptr[2]),
    .A4(_270_),
    .ZN(_279_));
 XNOR2_X1 _541_ (.A(net96),
    .B(_279_),
    .ZN(_280_));
 AOI211_X1 _542_ (.A(_238_),
    .B(net97),
    .C1(_274_),
    .C2(net18),
    .ZN(_121_));
 DFF_X1 _543_ (.D(net80),
    .CK(clknet_3_2_0_clk),
    .Q(curr_state[0]),
    .QN(_331_));
 DFF_X2 _544_ (.D(_193_),
    .CK(clknet_3_2_0_clk),
    .Q(net20),
    .QN(_332_));
 DFF_X2 _545_ (.D(net107),
    .CK(clknet_3_2_0_clk),
    .Q(curr_state[2]),
    .QN(_333_));
 DFF_X1 _546_ (.D(_138_),
    .CK(clknet_3_7_0_clk),
    .Q(net21),
    .QN(_334_));
 DFF_X1 _547_ (.D(_149_),
    .CK(clknet_3_7_0_clk),
    .Q(net32),
    .QN(_335_));
 DFF_X1 _548_ (.D(_160_),
    .CK(clknet_3_7_0_clk),
    .Q(net43),
    .QN(_336_));
 DFF_X2 _549_ (.D(_163_),
    .CK(clknet_3_6_0_clk),
    .Q(net46),
    .QN(_337_));
 DFF_X2 _550_ (.D(_164_),
    .CK(clknet_3_3_0_clk),
    .Q(net47),
    .QN(_338_));
 DFF_X2 _551_ (.D(_165_),
    .CK(clknet_3_6_0_clk),
    .Q(net48),
    .QN(_339_));
 DFF_X1 _552_ (.D(_166_),
    .CK(clknet_3_3_0_clk),
    .Q(net49),
    .QN(_340_));
 DFF_X1 _553_ (.D(_167_),
    .CK(clknet_3_7_0_clk),
    .Q(net50),
    .QN(_341_));
 DFF_X2 _554_ (.D(_168_),
    .CK(clknet_3_7_0_clk),
    .Q(net51),
    .QN(_342_));
 DFF_X2 _555_ (.D(_169_),
    .CK(clknet_3_7_0_clk),
    .Q(net52),
    .QN(_343_));
 DFF_X2 _556_ (.D(_139_),
    .CK(clknet_3_7_0_clk),
    .Q(net22),
    .QN(_344_));
 DFF_X2 _557_ (.D(_140_),
    .CK(clknet_3_7_0_clk),
    .Q(net23),
    .QN(_345_));
 DFF_X2 _558_ (.D(_141_),
    .CK(clknet_3_3_0_clk),
    .Q(net24),
    .QN(_346_));
 DFF_X2 _559_ (.D(_142_),
    .CK(clknet_3_6_0_clk),
    .Q(net25),
    .QN(_347_));
 DFF_X2 _560_ (.D(_143_),
    .CK(clknet_3_6_0_clk),
    .Q(net26),
    .QN(_348_));
 DFF_X2 _561_ (.D(_144_),
    .CK(clknet_3_6_0_clk),
    .Q(net27),
    .QN(_349_));
 DFF_X2 _562_ (.D(_145_),
    .CK(clknet_3_3_0_clk),
    .Q(net28),
    .QN(_350_));
 DFF_X2 _563_ (.D(_146_),
    .CK(clknet_3_5_0_clk),
    .Q(net29),
    .QN(_351_));
 DFF_X1 _564_ (.D(_147_),
    .CK(clknet_3_2_0_clk),
    .Q(net30),
    .QN(_352_));
 DFF_X2 _565_ (.D(_148_),
    .CK(clknet_3_4_0_clk),
    .Q(net31),
    .QN(_353_));
 DFF_X2 _566_ (.D(_150_),
    .CK(clknet_3_0_0_clk),
    .Q(net33),
    .QN(_354_));
 DFF_X2 _567_ (.D(_151_),
    .CK(clknet_3_4_0_clk),
    .Q(net34),
    .QN(_355_));
 DFF_X2 _568_ (.D(_152_),
    .CK(clknet_3_5_0_clk),
    .Q(net35),
    .QN(_356_));
 DFF_X2 _569_ (.D(_153_),
    .CK(clknet_3_4_0_clk),
    .Q(net36),
    .QN(_357_));
 DFF_X2 _570_ (.D(_154_),
    .CK(clknet_3_6_0_clk),
    .Q(net37),
    .QN(_358_));
 DFF_X2 _571_ (.D(_155_),
    .CK(clknet_3_5_0_clk),
    .Q(net38),
    .QN(_359_));
 DFF_X2 _572_ (.D(_156_),
    .CK(clknet_3_5_0_clk),
    .Q(net39),
    .QN(_360_));
 DFF_X1 _573_ (.D(_157_),
    .CK(clknet_3_5_0_clk),
    .Q(net40),
    .QN(_361_));
 DFF_X1 _574_ (.D(_158_),
    .CK(clknet_3_5_0_clk),
    .Q(net41),
    .QN(_362_));
 DFF_X2 _575_ (.D(_159_),
    .CK(clknet_3_5_0_clk),
    .Q(net42),
    .QN(_363_));
 DFF_X2 _576_ (.D(_161_),
    .CK(clknet_3_4_0_clk),
    .Q(net44),
    .QN(_364_));
 DFF_X2 _577_ (.D(_162_),
    .CK(clknet_3_5_0_clk),
    .Q(net45),
    .QN(_365_));
 DFF_X2 _578_ (.D(_122_),
    .CK(clknet_3_7_0_clk),
    .Q(data_in_reg[0]),
    .QN(_366_));
 DFF_X2 _579_ (.D(_129_),
    .CK(clknet_3_3_0_clk),
    .Q(data_in_reg[1]),
    .QN(_367_));
 DFF_X2 _580_ (.D(_130_),
    .CK(clknet_3_5_0_clk),
    .Q(data_in_reg[2]),
    .QN(_368_));
 DFF_X2 _581_ (.D(_131_),
    .CK(clknet_3_6_0_clk),
    .Q(data_in_reg[3]),
    .QN(_369_));
 DFF_X2 _582_ (.D(_132_),
    .CK(clknet_3_3_0_clk),
    .Q(data_in_reg[4]),
    .QN(_370_));
 DFF_X2 _583_ (.D(_133_),
    .CK(clknet_3_4_0_clk),
    .Q(data_in_reg[5]),
    .QN(_371_));
 DFF_X2 _584_ (.D(_134_),
    .CK(clknet_3_5_0_clk),
    .Q(data_in_reg[6]),
    .QN(_372_));
 DFF_X2 _585_ (.D(_135_),
    .CK(clknet_3_7_0_clk),
    .Q(data_in_reg[7]),
    .QN(_373_));
 DFF_X2 _586_ (.D(_136_),
    .CK(clknet_3_2_0_clk),
    .Q(data_in_reg[8]),
    .QN(_374_));
 DFF_X2 _587_ (.D(_137_),
    .CK(clknet_3_3_0_clk),
    .Q(data_in_reg[9]),
    .QN(_375_));
 DFF_X2 _588_ (.D(_123_),
    .CK(clknet_3_4_0_clk),
    .Q(data_in_reg[10]),
    .QN(_376_));
 DFF_X2 _589_ (.D(_124_),
    .CK(clknet_3_6_0_clk),
    .Q(data_in_reg[11]),
    .QN(_377_));
 DFF_X2 _590_ (.D(_125_),
    .CK(clknet_3_6_0_clk),
    .Q(data_in_reg[12]),
    .QN(_378_));
 DFF_X2 _591_ (.D(_126_),
    .CK(clknet_3_4_0_clk),
    .Q(data_in_reg[13]),
    .QN(_379_));
 DFF_X2 _592_ (.D(_127_),
    .CK(clknet_3_1_0_clk),
    .Q(data_in_reg[14]),
    .QN(_380_));
 DFF_X2 _593_ (.D(_128_),
    .CK(clknet_3_0_0_clk),
    .Q(data_in_reg[15]),
    .QN(_381_));
 DFF_X2 _594_ (.D(_175_),
    .CK(clknet_3_0_0_clk),
    .Q(sram_rdata_reg[0]),
    .QN(_382_));
 DFF_X2 _595_ (.D(_182_),
    .CK(clknet_3_0_0_clk),
    .Q(sram_rdata_reg[1]),
    .QN(_383_));
 DFF_X2 _596_ (.D(_183_),
    .CK(clknet_3_0_0_clk),
    .Q(sram_rdata_reg[2]),
    .QN(_384_));
 DFF_X2 _597_ (.D(_184_),
    .CK(clknet_3_0_0_clk),
    .Q(sram_rdata_reg[3]),
    .QN(_385_));
 DFF_X2 _598_ (.D(_185_),
    .CK(clknet_3_0_0_clk),
    .Q(sram_rdata_reg[4]),
    .QN(_386_));
 DFF_X2 _599_ (.D(_186_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[5]),
    .QN(_387_));
 DFF_X2 _600_ (.D(_187_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[6]),
    .QN(_388_));
 DFF_X2 _601_ (.D(_188_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[7]),
    .QN(_389_));
 DFF_X2 _602_ (.D(_189_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[8]),
    .QN(_390_));
 DFF_X2 _603_ (.D(_190_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[9]),
    .QN(_391_));
 DFF_X2 _604_ (.D(_176_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[10]),
    .QN(_392_));
 DFF_X2 _605_ (.D(_177_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[11]),
    .QN(_393_));
 DFF_X2 _606_ (.D(_178_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[12]),
    .QN(_394_));
 DFF_X2 _607_ (.D(_179_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[13]),
    .QN(_395_));
 DFF_X2 _608_ (.D(_180_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[14]),
    .QN(_396_));
 DFF_X2 _609_ (.D(_181_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[15]),
    .QN(_397_));
 DFF_X1 _610_ (.D(_191_),
    .CK(clknet_3_7_0_clk),
    .Q(net53),
    .QN(_398_));
 DFF_X2 _611_ (.D(net110),
    .CK(clknet_3_2_0_clk),
    .Q(addr_ptr[0]),
    .QN(_399_));
 DFF_X1 _612_ (.D(net95),
    .CK(clknet_3_2_0_clk),
    .Q(addr_ptr[1]),
    .QN(_400_));
 DFF_X1 _613_ (.D(_119_),
    .CK(clknet_3_2_0_clk),
    .Q(addr_ptr[2]),
    .QN(_401_));
 DFF_X2 _614_ (.D(_120_),
    .CK(clknet_3_3_0_clk),
    .Q(addr_ptr[3]),
    .QN(_402_));
 DFF_X1 _615_ (.D(_121_),
    .CK(clknet_3_3_0_clk),
    .Q(addr_ptr[4]),
    .QN(_403_));
 DFF_X2 _616_ (.D(net117),
    .CK(clknet_3_2_0_clk),
    .Q(init_count[0]),
    .QN(_404_));
 DFF_X2 _617_ (.D(net100),
    .CK(clknet_3_2_0_clk),
    .Q(init_count[1]),
    .QN(_405_));
 DFF_X1 _618_ (.D(net103),
    .CK(clknet_3_2_0_clk),
    .Q(init_count[2]),
    .QN(_406_));
 DFF_X1 _619_ (.D(net78),
    .CK(clknet_3_2_0_clk),
    .Q(init_count[3]),
    .QN(_407_));
 DFF_X1 _620_ (.D(net125),
    .CK(clknet_3_2_0_clk),
    .Q(init_count[4]),
    .QN(_408_));
 SRAM_6T_CORE_32x16_MC_TB sram_inst (.ce_in(_195_),
    .we_in(_196_),
    .clk(clknet_3_0_0_clk),
    .addr_in({net127,
    net91,
    net89,
    net129,
    net92}),
    .rd_out({sram_rdata[15],
    sram_rdata[14],
    sram_rdata[13],
    sram_rdata[12],
    sram_rdata[11],
    sram_rdata[10],
    sram_rdata[9],
    sram_rdata[8],
    sram_rdata[7],
    sram_rdata[6],
    sram_rdata[5],
    sram_rdata[4],
    sram_rdata[3],
    sram_rdata[2],
    sram_rdata[1],
    sram_rdata[0]}),
    .wd_in({net122,
    net104,
    net111,
    net118,
    net121,
    net120,
    net143,
    net136,
    net145,
    net138,
    net119,
    net131,
    net134,
    net135,
    net114,
    net144}));
 NAND3_X1 \u_multiplier/STAGE1/ACCI1_pp_10/_21_  (.A1(\u_multiplier/STAGE1/_185_ ),
    .A2(\u_multiplier/STAGE1/_184_ ),
    .A3(\u_multiplier/STAGE1/_186_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_10/_18_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_10/_22_  (.A(\u_multiplier/STAGE1/_185_ ),
    .B(\u_multiplier/STAGE1/_184_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_10/_19_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_10/_23_  (.A(\u_multiplier/STAGE1/_186_ ),
    .B(\u_multiplier/STAGE1/_187_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_10/_20_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_10/_24_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_10/_19_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_10/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_10/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE1/ACCI1_pp_10/_25_  (.A(\u_multiplier/STAGE1/ACCI1_pp_10/_19_ ),
    .B(\u_multiplier/STAGE1/ACCI1_pp_10/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_10/_16_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_10/_26_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_10/_18_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_10/_16_ ),
    .ZN(\u_multiplier/pp_10 [1]));
 AOI22_X1 \u_multiplier/STAGE1/ACCI1_pp_10/_27_  (.A1(\u_multiplier/STAGE1/_185_ ),
    .A2(\u_multiplier/STAGE1/_184_ ),
    .B1(\u_multiplier/STAGE1/_186_ ),
    .B2(\u_multiplier/STAGE1/_187_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_10/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_10/_28_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_10/_15_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_10/_17_ ),
    .ZN(\u_multiplier/pp_11 [2]));
 NAND3_X1 \u_multiplier/STAGE1/ACCI1_pp_11_1/_21_  (.A1(\u_multiplier/STAGE1/_191_ ),
    .A2(\u_multiplier/STAGE1/_190_ ),
    .A3(\u_multiplier/STAGE1/_192_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_11_1/_18_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_11_1/_22_  (.A(\u_multiplier/STAGE1/_191_ ),
    .B(\u_multiplier/STAGE1/_190_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_11_1/_19_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_11_1/_23_  (.A(\u_multiplier/STAGE1/_192_ ),
    .B(\u_multiplier/STAGE1/_193_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_11_1/_20_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_11_1/_24_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_11_1/_19_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_11_1/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_11_1/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE1/ACCI1_pp_11_1/_25_  (.A(\u_multiplier/STAGE1/ACCI1_pp_11_1/_19_ ),
    .B(\u_multiplier/STAGE1/ACCI1_pp_11_1/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_11_1/_16_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_11_1/_26_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_11_1/_18_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_11_1/_16_ ),
    .ZN(\u_multiplier/pp_11 [1]));
 AOI22_X2 \u_multiplier/STAGE1/ACCI1_pp_11_1/_27_  (.A1(\u_multiplier/STAGE1/_191_ ),
    .A2(\u_multiplier/STAGE1/_190_ ),
    .B1(\u_multiplier/STAGE1/_192_ ),
    .B2(\u_multiplier/STAGE1/_193_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_11_1/_17_ ));
 NAND2_X2 \u_multiplier/STAGE1/ACCI1_pp_11_1/_28_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_11_1/_15_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_11_1/_17_ ),
    .ZN(\u_multiplier/pp_12 [2]));
 NAND3_X1 \u_multiplier/STAGE1/ACCI1_pp_11_2/_21_  (.A1(\u_multiplier/STAGE1/_195_ ),
    .A2(\u_multiplier/STAGE1/_194_ ),
    .A3(\u_multiplier/STAGE1/_196_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_11_2/_18_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_11_2/_22_  (.A(\u_multiplier/STAGE1/_195_ ),
    .B(\u_multiplier/STAGE1/_194_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_11_2/_19_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_11_2/_23_  (.A(\u_multiplier/STAGE1/_196_ ),
    .B(\u_multiplier/STAGE1/_197_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_11_2/_20_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_11_2/_24_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_11_2/_19_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_11_2/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_11_2/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE1/ACCI1_pp_11_2/_25_  (.A(\u_multiplier/STAGE1/ACCI1_pp_11_2/_19_ ),
    .B(\u_multiplier/STAGE1/ACCI1_pp_11_2/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_11_2/_16_ ));
 NAND2_X2 \u_multiplier/STAGE1/ACCI1_pp_11_2/_26_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_11_2/_18_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_11_2/_16_ ),
    .ZN(\u_multiplier/pp_11 [0]));
 AOI22_X1 \u_multiplier/STAGE1/ACCI1_pp_11_2/_27_  (.A1(\u_multiplier/STAGE1/_195_ ),
    .A2(\u_multiplier/STAGE1/_194_ ),
    .B1(\u_multiplier/STAGE1/_196_ ),
    .B2(\u_multiplier/STAGE1/_197_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_11_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_11_2/_28_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_11_2/_15_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_11_2/_17_ ),
    .ZN(\u_multiplier/pp_12 [3]));
 NAND3_X1 \u_multiplier/STAGE1/ACCI1_pp_12_1/_21_  (.A1(\u_multiplier/STAGE1/_199_ ),
    .A2(\u_multiplier/STAGE1/_198_ ),
    .A3(\u_multiplier/STAGE1/_200_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_12_1/_18_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_12_1/_22_  (.A(\u_multiplier/STAGE1/_199_ ),
    .B(\u_multiplier/STAGE1/_198_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_12_1/_19_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_12_1/_23_  (.A(\u_multiplier/STAGE1/_200_ ),
    .B(\u_multiplier/STAGE1/_201_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_12_1/_20_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_12_1/_24_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_12_1/_19_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_12_1/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_12_1/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE1/ACCI1_pp_12_1/_25_  (.A(\u_multiplier/STAGE1/ACCI1_pp_12_1/_19_ ),
    .B(\u_multiplier/STAGE1/ACCI1_pp_12_1/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_12_1/_16_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_12_1/_26_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_12_1/_18_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_12_1/_16_ ),
    .ZN(\u_multiplier/pp_12 [4]));
 AOI22_X2 \u_multiplier/STAGE1/ACCI1_pp_12_1/_27_  (.A1(\u_multiplier/STAGE1/_199_ ),
    .A2(\u_multiplier/STAGE1/_198_ ),
    .B1(\u_multiplier/STAGE1/_200_ ),
    .B2(\u_multiplier/STAGE1/_201_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_12_1/_17_ ));
 NAND2_X2 \u_multiplier/STAGE1/ACCI1_pp_12_1/_28_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_12_1/_15_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_12_1/_17_ ),
    .ZN(\u_multiplier/pp_13 [2]));
 NAND3_X1 \u_multiplier/STAGE1/ACCI1_pp_12_2/_21_  (.A1(\u_multiplier/STAGE1/_203_ ),
    .A2(\u_multiplier/STAGE1/_202_ ),
    .A3(\u_multiplier/STAGE1/_204_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_12_2/_18_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_12_2/_22_  (.A(\u_multiplier/STAGE1/_203_ ),
    .B(\u_multiplier/STAGE1/_202_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_12_2/_19_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_12_2/_23_  (.A(\u_multiplier/STAGE1/_204_ ),
    .B(\u_multiplier/STAGE1/_205_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_12_2/_20_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_12_2/_24_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_12_2/_19_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_12_2/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_12_2/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE1/ACCI1_pp_12_2/_25_  (.A(\u_multiplier/STAGE1/ACCI1_pp_12_2/_19_ ),
    .B(\u_multiplier/STAGE1/ACCI1_pp_12_2/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_12_2/_16_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_12_2/_26_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_12_2/_18_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_12_2/_16_ ),
    .ZN(\u_multiplier/pp_12 [1]));
 AOI22_X2 \u_multiplier/STAGE1/ACCI1_pp_12_2/_27_  (.A1(\u_multiplier/STAGE1/_203_ ),
    .A2(\u_multiplier/STAGE1/_202_ ),
    .B1(\u_multiplier/STAGE1/_204_ ),
    .B2(\u_multiplier/STAGE1/_205_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_12_2/_17_ ));
 NAND2_X2 \u_multiplier/STAGE1/ACCI1_pp_12_2/_28_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_12_2/_15_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_12_2/_17_ ),
    .ZN(\u_multiplier/pp_13 [3]));
 NAND3_X1 \u_multiplier/STAGE1/ACCI1_pp_13_1/_21_  (.A1(\u_multiplier/STAGE1/_209_ ),
    .A2(\u_multiplier/STAGE1/_208_ ),
    .A3(\u_multiplier/STAGE1/_210_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_13_1/_18_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_13_1/_22_  (.A(\u_multiplier/STAGE1/_209_ ),
    .B(\u_multiplier/STAGE1/_208_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_13_1/_19_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_13_1/_23_  (.A(\u_multiplier/STAGE1/_210_ ),
    .B(\u_multiplier/STAGE1/_211_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_13_1/_20_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_13_1/_24_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_13_1/_19_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_13_1/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_13_1/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE1/ACCI1_pp_13_1/_25_  (.A(\u_multiplier/STAGE1/ACCI1_pp_13_1/_19_ ),
    .B(\u_multiplier/STAGE1/ACCI1_pp_13_1/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_13_1/_16_ ));
 NAND2_X2 \u_multiplier/STAGE1/ACCI1_pp_13_1/_26_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_13_1/_18_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_13_1/_16_ ),
    .ZN(\u_multiplier/pp_13 [1]));
 AOI22_X2 \u_multiplier/STAGE1/ACCI1_pp_13_1/_27_  (.A1(\u_multiplier/STAGE1/_209_ ),
    .A2(\u_multiplier/STAGE1/_208_ ),
    .B1(\u_multiplier/STAGE1/_210_ ),
    .B2(\u_multiplier/STAGE1/_211_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_13_1/_17_ ));
 NAND2_X2 \u_multiplier/STAGE1/ACCI1_pp_13_1/_28_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_13_1/_15_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_13_1/_17_ ),
    .ZN(\u_multiplier/pp_14 [2]));
 NAND3_X1 \u_multiplier/STAGE1/ACCI1_pp_13_2/_21_  (.A1(\u_multiplier/STAGE1/_213_ ),
    .A2(\u_multiplier/STAGE1/_212_ ),
    .A3(\u_multiplier/STAGE1/_214_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_13_2/_18_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_13_2/_22_  (.A(\u_multiplier/STAGE1/_213_ ),
    .B(\u_multiplier/STAGE1/_212_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_13_2/_19_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_13_2/_23_  (.A(\u_multiplier/STAGE1/_214_ ),
    .B(\u_multiplier/STAGE1/_215_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_13_2/_20_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_13_2/_24_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_13_2/_19_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_13_2/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_13_2/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE1/ACCI1_pp_13_2/_25_  (.A(\u_multiplier/STAGE1/ACCI1_pp_13_2/_19_ ),
    .B(\u_multiplier/STAGE1/ACCI1_pp_13_2/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_13_2/_16_ ));
 NAND2_X2 \u_multiplier/STAGE1/ACCI1_pp_13_2/_26_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_13_2/_18_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_13_2/_16_ ),
    .ZN(\u_multiplier/pp_13 [0]));
 AOI22_X1 \u_multiplier/STAGE1/ACCI1_pp_13_2/_27_  (.A1(\u_multiplier/STAGE1/_213_ ),
    .A2(\u_multiplier/STAGE1/_212_ ),
    .B1(\u_multiplier/STAGE1/_214_ ),
    .B2(\u_multiplier/STAGE1/_215_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_13_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_13_2/_28_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_13_2/_15_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_13_2/_17_ ),
    .ZN(\u_multiplier/pp_14 [3]));
 NAND3_X1 \u_multiplier/STAGE1/ACCI1_pp_13_3/_21_  (.A1(\u_multiplier/STAGE1/_217_ ),
    .A2(\u_multiplier/STAGE1/_216_ ),
    .A3(\u_multiplier/STAGE1/_218_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_13_3/_18_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_13_3/_22_  (.A(\u_multiplier/STAGE1/_217_ ),
    .B(\u_multiplier/STAGE1/_216_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_13_3/_19_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_13_3/_23_  (.A(\u_multiplier/STAGE1/_218_ ),
    .B(\u_multiplier/STAGE1/_219_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_13_3/_20_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_13_3/_24_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_13_3/_19_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_13_3/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_13_3/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE1/ACCI1_pp_13_3/_25_  (.A(\u_multiplier/STAGE1/ACCI1_pp_13_3/_19_ ),
    .B(\u_multiplier/STAGE1/ACCI1_pp_13_3/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_13_3/_16_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_13_3/_26_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_13_3/_18_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_13_3/_16_ ),
    .ZN(\u_multiplier/pp_13 [4]));
 AOI22_X1 \u_multiplier/STAGE1/ACCI1_pp_13_3/_27_  (.A1(\u_multiplier/STAGE1/_217_ ),
    .A2(\u_multiplier/STAGE1/_216_ ),
    .B1(\u_multiplier/STAGE1/_218_ ),
    .B2(\u_multiplier/STAGE1/_219_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_13_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_13_3/_28_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_13_3/_15_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_13_3/_17_ ),
    .ZN(\u_multiplier/pp_14 [7]));
 NAND3_X1 \u_multiplier/STAGE1/ACCI1_pp_14_1/_21_  (.A1(\u_multiplier/STAGE1/_221_ ),
    .A2(\u_multiplier/STAGE1/_220_ ),
    .A3(\u_multiplier/STAGE1/_222_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_14_1/_18_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_14_1/_22_  (.A(\u_multiplier/STAGE1/_221_ ),
    .B(\u_multiplier/STAGE1/_220_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_14_1/_19_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_14_1/_23_  (.A(\u_multiplier/STAGE1/_222_ ),
    .B(\u_multiplier/STAGE1/_223_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_14_1/_20_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_14_1/_24_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_14_1/_19_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_14_1/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_14_1/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE1/ACCI1_pp_14_1/_25_  (.A(\u_multiplier/STAGE1/ACCI1_pp_14_1/_19_ ),
    .B(\u_multiplier/STAGE1/ACCI1_pp_14_1/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_14_1/_16_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_14_1/_26_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_14_1/_18_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_14_1/_16_ ),
    .ZN(\u_multiplier/pp_14 [1]));
 AOI22_X2 \u_multiplier/STAGE1/ACCI1_pp_14_1/_27_  (.A1(\u_multiplier/STAGE1/_221_ ),
    .A2(\u_multiplier/STAGE1/_220_ ),
    .B1(\u_multiplier/STAGE1/_222_ ),
    .B2(\u_multiplier/STAGE1/_223_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_14_1/_17_ ));
 NAND2_X2 \u_multiplier/STAGE1/ACCI1_pp_14_1/_28_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_14_1/_15_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_14_1/_17_ ),
    .ZN(\u_multiplier/pp_15 [2]));
 NAND3_X1 \u_multiplier/STAGE1/ACCI1_pp_14_2/_21_  (.A1(\u_multiplier/STAGE1/_225_ ),
    .A2(\u_multiplier/STAGE1/_224_ ),
    .A3(\u_multiplier/STAGE1/_226_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_14_2/_18_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_14_2/_22_  (.A(\u_multiplier/STAGE1/_225_ ),
    .B(\u_multiplier/STAGE1/_224_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_14_2/_19_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_14_2/_23_  (.A(\u_multiplier/STAGE1/_226_ ),
    .B(\u_multiplier/STAGE1/_227_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_14_2/_20_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_14_2/_24_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_14_2/_19_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_14_2/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_14_2/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE1/ACCI1_pp_14_2/_25_  (.A(\u_multiplier/STAGE1/ACCI1_pp_14_2/_19_ ),
    .B(\u_multiplier/STAGE1/ACCI1_pp_14_2/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_14_2/_16_ ));
 NAND2_X2 \u_multiplier/STAGE1/ACCI1_pp_14_2/_26_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_14_2/_18_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_14_2/_16_ ),
    .ZN(\u_multiplier/pp_14 [0]));
 AOI22_X1 \u_multiplier/STAGE1/ACCI1_pp_14_2/_27_  (.A1(\u_multiplier/STAGE1/_225_ ),
    .A2(\u_multiplier/STAGE1/_224_ ),
    .B1(\u_multiplier/STAGE1/_226_ ),
    .B2(\u_multiplier/STAGE1/_227_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_14_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_14_2/_28_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_14_2/_15_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_14_2/_17_ ),
    .ZN(\u_multiplier/pp_15 [3]));
 NAND3_X1 \u_multiplier/STAGE1/ACCI1_pp_14_3/_21_  (.A1(\u_multiplier/STAGE1/_229_ ),
    .A2(\u_multiplier/STAGE1/_228_ ),
    .A3(\u_multiplier/STAGE1/_230_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_14_3/_18_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_14_3/_22_  (.A(\u_multiplier/STAGE1/_229_ ),
    .B(\u_multiplier/STAGE1/_228_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_14_3/_19_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_14_3/_23_  (.A(\u_multiplier/STAGE1/_230_ ),
    .B(\u_multiplier/STAGE1/_231_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_14_3/_20_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_14_3/_24_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_14_3/_19_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_14_3/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_14_3/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE1/ACCI1_pp_14_3/_25_  (.A(\u_multiplier/STAGE1/ACCI1_pp_14_3/_19_ ),
    .B(\u_multiplier/STAGE1/ACCI1_pp_14_3/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_14_3/_16_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_14_3/_26_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_14_3/_18_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_14_3/_16_ ),
    .ZN(\u_multiplier/pp_14 [4]));
 AOI22_X2 \u_multiplier/STAGE1/ACCI1_pp_14_3/_27_  (.A1(\u_multiplier/STAGE1/_229_ ),
    .A2(\u_multiplier/STAGE1/_228_ ),
    .B1(\u_multiplier/STAGE1/_230_ ),
    .B2(\u_multiplier/STAGE1/_231_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_14_3/_17_ ));
 NAND2_X2 \u_multiplier/STAGE1/ACCI1_pp_14_3/_28_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_14_3/_15_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_14_3/_17_ ),
    .ZN(\u_multiplier/pp_15 [6]));
 NAND3_X1 \u_multiplier/STAGE1/ACCI1_pp_15_1/_21_  (.A1(\u_multiplier/STAGE1/_235_ ),
    .A2(\u_multiplier/STAGE1/_234_ ),
    .A3(\u_multiplier/STAGE1/_236_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_15_1/_18_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_15_1/_22_  (.A(\u_multiplier/STAGE1/_235_ ),
    .B(\u_multiplier/STAGE1/_234_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_15_1/_19_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_15_1/_23_  (.A(\u_multiplier/STAGE1/_236_ ),
    .B(\u_multiplier/STAGE1/_237_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_15_1/_20_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_15_1/_24_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_15_1/_19_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_15_1/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_15_1/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE1/ACCI1_pp_15_1/_25_  (.A(\u_multiplier/STAGE1/ACCI1_pp_15_1/_19_ ),
    .B(\u_multiplier/STAGE1/ACCI1_pp_15_1/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_15_1/_16_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_15_1/_26_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_15_1/_18_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_15_1/_16_ ),
    .ZN(\u_multiplier/pp_15 [1]));
 AOI22_X1 \u_multiplier/STAGE1/ACCI1_pp_15_1/_27_  (.A1(\u_multiplier/STAGE1/_235_ ),
    .A2(\u_multiplier/STAGE1/_234_ ),
    .B1(\u_multiplier/STAGE1/_236_ ),
    .B2(\u_multiplier/STAGE1/_237_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_15_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_15_1/_28_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_15_1/_15_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_15_1/_17_ ),
    .ZN(\u_multiplier/pp_16 [0]));
 NAND3_X1 \u_multiplier/STAGE1/ACCI1_pp_15_2/_21_  (.A1(\u_multiplier/STAGE1/_239_ ),
    .A2(\u_multiplier/STAGE1/_238_ ),
    .A3(\u_multiplier/STAGE1/_240_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_15_2/_18_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_15_2/_22_  (.A(\u_multiplier/STAGE1/_239_ ),
    .B(\u_multiplier/STAGE1/_238_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_15_2/_19_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_15_2/_23_  (.A(\u_multiplier/STAGE1/_240_ ),
    .B(\u_multiplier/STAGE1/_241_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_15_2/_20_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_15_2/_24_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_15_2/_19_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_15_2/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_15_2/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE1/ACCI1_pp_15_2/_25_  (.A(\u_multiplier/STAGE1/ACCI1_pp_15_2/_19_ ),
    .B(\u_multiplier/STAGE1/ACCI1_pp_15_2/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_15_2/_16_ ));
 NAND2_X2 \u_multiplier/STAGE1/ACCI1_pp_15_2/_26_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_15_2/_18_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_15_2/_16_ ),
    .ZN(\u_multiplier/pp_15 [0]));
 AOI22_X1 \u_multiplier/STAGE1/ACCI1_pp_15_2/_27_  (.A1(\u_multiplier/STAGE1/_239_ ),
    .A2(\u_multiplier/STAGE1/_238_ ),
    .B1(\u_multiplier/STAGE1/_240_ ),
    .B2(\u_multiplier/STAGE1/_241_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_15_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_15_2/_28_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_15_2/_15_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_15_2/_17_ ),
    .ZN(\u_multiplier/pp_16 [2]));
 NAND3_X1 \u_multiplier/STAGE1/ACCI1_pp_15_3/_21_  (.A1(\u_multiplier/STAGE1/_243_ ),
    .A2(\u_multiplier/STAGE1/_242_ ),
    .A3(\u_multiplier/STAGE1/_244_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_15_3/_18_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_15_3/_22_  (.A(\u_multiplier/STAGE1/_243_ ),
    .B(\u_multiplier/STAGE1/_242_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_15_3/_19_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_15_3/_23_  (.A(\u_multiplier/STAGE1/_244_ ),
    .B(\u_multiplier/STAGE1/_245_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_15_3/_20_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_15_3/_24_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_15_3/_19_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_15_3/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_15_3/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE1/ACCI1_pp_15_3/_25_  (.A(\u_multiplier/STAGE1/ACCI1_pp_15_3/_19_ ),
    .B(\u_multiplier/STAGE1/ACCI1_pp_15_3/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_15_3/_16_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_15_3/_26_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_15_3/_18_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_15_3/_16_ ),
    .ZN(\u_multiplier/pp_15 [4]));
 AOI22_X1 \u_multiplier/STAGE1/ACCI1_pp_15_3/_27_  (.A1(\u_multiplier/STAGE1/_243_ ),
    .A2(\u_multiplier/STAGE1/_242_ ),
    .B1(\u_multiplier/STAGE1/_244_ ),
    .B2(\u_multiplier/STAGE1/_245_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_15_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_15_3/_28_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_15_3/_15_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_15_3/_17_ ),
    .ZN(\u_multiplier/pp_16 [4]));
 NAND3_X1 \u_multiplier/STAGE1/ACCI1_pp_15_4/_21_  (.A1(\u_multiplier/STAGE1/_247_ ),
    .A2(\u_multiplier/STAGE1/_246_ ),
    .A3(\u_multiplier/STAGE1/_248_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_15_4/_18_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_15_4/_22_  (.A(\u_multiplier/STAGE1/_247_ ),
    .B(\u_multiplier/STAGE1/_246_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_15_4/_19_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_15_4/_23_  (.A(\u_multiplier/STAGE1/_248_ ),
    .B(\u_multiplier/STAGE1/_249_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_15_4/_20_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_15_4/_24_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_15_4/_19_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_15_4/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_15_4/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE1/ACCI1_pp_15_4/_25_  (.A(\u_multiplier/STAGE1/ACCI1_pp_15_4/_19_ ),
    .B(\u_multiplier/STAGE1/ACCI1_pp_15_4/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_15_4/_16_ ));
 NAND2_X2 \u_multiplier/STAGE1/ACCI1_pp_15_4/_26_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_15_4/_18_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_15_4/_16_ ),
    .ZN(\u_multiplier/pp_15 [5]));
 AOI22_X1 \u_multiplier/STAGE1/ACCI1_pp_15_4/_27_  (.A1(\u_multiplier/STAGE1/_247_ ),
    .A2(\u_multiplier/STAGE1/_246_ ),
    .B1(\u_multiplier/STAGE1/_248_ ),
    .B2(\u_multiplier/STAGE1/_249_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_15_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_15_4/_28_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_15_4/_15_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_15_4/_17_ ),
    .ZN(\u_multiplier/pp_16 [6]));
 NAND3_X1 \u_multiplier/STAGE1/ACCI1_pp_9/_21_  (.A1(\u_multiplier/STAGE1/_181_ ),
    .A2(\u_multiplier/STAGE1/_180_ ),
    .A3(\u_multiplier/STAGE1/_182_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_9/_18_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_9/_22_  (.A(\u_multiplier/STAGE1/_181_ ),
    .B(\u_multiplier/STAGE1/_180_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_9/_19_ ));
 XOR2_X2 \u_multiplier/STAGE1/ACCI1_pp_9/_23_  (.A(\u_multiplier/STAGE1/_182_ ),
    .B(\u_multiplier/STAGE1/_183_ ),
    .Z(\u_multiplier/STAGE1/ACCI1_pp_9/_20_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_9/_24_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_9/_19_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_9/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_9/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE1/ACCI1_pp_9/_25_  (.A(\u_multiplier/STAGE1/ACCI1_pp_9/_19_ ),
    .B(\u_multiplier/STAGE1/ACCI1_pp_9/_20_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_9/_16_ ));
 NAND2_X2 \u_multiplier/STAGE1/ACCI1_pp_9/_26_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_9/_18_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_9/_16_ ),
    .ZN(\u_multiplier/pp_9 [0]));
 AOI22_X1 \u_multiplier/STAGE1/ACCI1_pp_9/_27_  (.A1(\u_multiplier/STAGE1/_181_ ),
    .A2(\u_multiplier/STAGE1/_180_ ),
    .B1(\u_multiplier/STAGE1/_182_ ),
    .B2(\u_multiplier/STAGE1/_183_ ),
    .ZN(\u_multiplier/STAGE1/ACCI1_pp_9/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/ACCI1_pp_9/_28_  (.A1(\u_multiplier/STAGE1/ACCI1_pp_9/_15_ ),
    .A2(\u_multiplier/STAGE1/ACCI1_pp_9/_17_ ),
    .ZN(\u_multiplier/pp_10 [3]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_16_1/_18_  (.A(net54),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_1/_19_  (.A1(\u_multiplier/STAGE1/_251_ ),
    .A2(\u_multiplier/STAGE1/_250_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_1/_20_  (.A(\u_multiplier/STAGE1/_251_ ),
    .B(\u_multiplier/STAGE1/_250_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_16_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_1/_21_  (.A1(\u_multiplier/STAGE1/_252_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_16_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_1/_22_  (.A(\u_multiplier/STAGE1/_252_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_16_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_16_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_1/_23_  (.A1(\u_multiplier/STAGE1/_253_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_16_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_1/_24_  (.A(\u_multiplier/STAGE1/_253_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_16_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_1/_25_  (.A(net55),
    .B(\u_multiplier/STAGE1/E_4_2_pp_16_1/_16_ ),
    .ZN(\u_multiplier/pp_16 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_16_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_16_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_16_c2 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_16_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_16_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_16_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_16_1/_17_ ),
    .ZN(\u_multiplier/pp_17 [0]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_16_2/_18_  (.A(net56),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_2/_19_  (.A1(\u_multiplier/STAGE1/_255_ ),
    .A2(\u_multiplier/STAGE1/_254_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_2/_20_  (.A(\u_multiplier/STAGE1/_255_ ),
    .B(\u_multiplier/STAGE1/_254_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_16_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_2/_21_  (.A1(\u_multiplier/STAGE1/_256_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_16_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_2/_22_  (.A(\u_multiplier/STAGE1/_256_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_16_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_16_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_2/_23_  (.A1(\u_multiplier/STAGE1/_257_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_16_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_2/_24_  (.A(\u_multiplier/STAGE1/_257_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_16_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_2/_25_  (.A(net57),
    .B(\u_multiplier/STAGE1/E_4_2_pp_16_2/_16_ ),
    .ZN(\u_multiplier/pp_16 [3]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_16_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_16_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_16_c4 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_16_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_16_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_16_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_16_2/_17_ ),
    .ZN(\u_multiplier/pp_17 [2]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_16_3/_18_  (.A(net58),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_3/_19_  (.A1(\u_multiplier/STAGE1/_259_ ),
    .A2(\u_multiplier/STAGE1/_258_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_3/_20_  (.A(\u_multiplier/STAGE1/_259_ ),
    .B(\u_multiplier/STAGE1/_258_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_16_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_3/_21_  (.A1(\u_multiplier/STAGE1/_260_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_16_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_3/_22_  (.A(\u_multiplier/STAGE1/_260_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_16_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_16_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_3/_23_  (.A1(\u_multiplier/STAGE1/_261_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_16_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_3/_24_  (.A(\u_multiplier/STAGE1/_261_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_16_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_3/_25_  (.A(net59),
    .B(\u_multiplier/STAGE1/E_4_2_pp_16_3/_16_ ),
    .ZN(\u_multiplier/pp_16 [5]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_16_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_16_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_16_c6 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_16_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_16_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_16_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_16_3/_17_ ),
    .ZN(\u_multiplier/pp_17 [4]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_17_1/_18_  (.A(\u_multiplier/STAGE1/pp_16_c2 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_1/_19_  (.A1(\u_multiplier/STAGE1/_266_ ),
    .A2(\u_multiplier/STAGE1/_265_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_1/_20_  (.A(\u_multiplier/STAGE1/_266_ ),
    .B(\u_multiplier/STAGE1/_265_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_17_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_1/_21_  (.A1(\u_multiplier/STAGE1/_267_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_17_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_1/_22_  (.A(\u_multiplier/STAGE1/_267_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_17_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_17_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_1/_23_  (.A1(\u_multiplier/STAGE1/_268_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_17_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_1/_24_  (.A(\u_multiplier/STAGE1/_268_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_17_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_1/_25_  (.A(\u_multiplier/STAGE1/pp_16_c2 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_17_1/_16_ ),
    .ZN(\u_multiplier/pp_17 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_17_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_17_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_17_c2 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_17_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_17_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_17_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_17_1/_17_ ),
    .ZN(\u_multiplier/pp_18 [1]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_17_2/_18_  (.A(\u_multiplier/STAGE1/pp_16_c4 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_2/_19_  (.A1(\u_multiplier/STAGE1/_270_ ),
    .A2(\u_multiplier/STAGE1/_269_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_2/_20_  (.A(\u_multiplier/STAGE1/_270_ ),
    .B(\u_multiplier/STAGE1/_269_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_17_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_2/_21_  (.A1(\u_multiplier/STAGE1/_271_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_17_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_2/_22_  (.A(\u_multiplier/STAGE1/_271_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_17_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_17_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_2/_23_  (.A1(\u_multiplier/STAGE1/_272_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_17_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_2/_24_  (.A(\u_multiplier/STAGE1/_272_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_17_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_2/_25_  (.A(\u_multiplier/STAGE1/pp_16_c4 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_17_2/_16_ ),
    .ZN(\u_multiplier/pp_17 [3]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_17_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_17_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_17_c4 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_17_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_17_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_17_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_17_2/_17_ ),
    .ZN(\u_multiplier/pp_18 [3]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_17_3/_18_  (.A(\u_multiplier/STAGE1/pp_16_c6 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_3/_19_  (.A1(\u_multiplier/STAGE1/_274_ ),
    .A2(\u_multiplier/STAGE1/_273_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_3/_20_  (.A(\u_multiplier/STAGE1/_274_ ),
    .B(\u_multiplier/STAGE1/_273_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_17_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_3/_21_  (.A1(\u_multiplier/STAGE1/_275_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_17_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_3/_22_  (.A(\u_multiplier/STAGE1/_275_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_17_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_17_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_3/_23_  (.A1(\u_multiplier/STAGE1/_276_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_17_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_3/_24_  (.A(\u_multiplier/STAGE1/_276_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_17_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_3/_25_  (.A(\u_multiplier/STAGE1/pp_16_c6 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_17_3/_16_ ),
    .ZN(\u_multiplier/pp_17 [5]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_17_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_17_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_17_c6 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_17_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_17_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_17_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_17_3/_17_ ),
    .ZN(\u_multiplier/pp_18 [5]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_18_1/_18_  (.A(\u_multiplier/STAGE1/pp_17_c2 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_18_1/_19_  (.A1(\u_multiplier/STAGE1/_280_ ),
    .A2(\u_multiplier/STAGE1/_279_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_1/_20_  (.A(\u_multiplier/STAGE1/_280_ ),
    .B(\u_multiplier/STAGE1/_279_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_18_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_18_1/_21_  (.A1(\u_multiplier/STAGE1/_281_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_18_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_1/_22_  (.A(\u_multiplier/STAGE1/_281_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_18_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_18_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_18_1/_23_  (.A1(\u_multiplier/STAGE1/_282_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_18_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_1/_24_  (.A(\u_multiplier/STAGE1/_282_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_18_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_1/_25_  (.A(\u_multiplier/STAGE1/pp_17_c2 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_18_1/_16_ ),
    .ZN(\u_multiplier/pp_18 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_18_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_18_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_18_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_18_c2 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_18_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_18_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_18_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_18_1/_17_ ),
    .ZN(\u_multiplier/pp_19 [1]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_18_2/_18_  (.A(\u_multiplier/STAGE1/pp_17_c4 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_18_2/_19_  (.A1(\u_multiplier/STAGE1/_284_ ),
    .A2(\u_multiplier/STAGE1/_283_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_2/_20_  (.A(\u_multiplier/STAGE1/_284_ ),
    .B(\u_multiplier/STAGE1/_283_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_18_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_18_2/_21_  (.A1(\u_multiplier/STAGE1/_285_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_18_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_2/_22_  (.A(\u_multiplier/STAGE1/_285_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_18_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_18_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_18_2/_23_  (.A1(\u_multiplier/STAGE1/_286_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_18_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_2/_24_  (.A(\u_multiplier/STAGE1/_286_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_18_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_2/_25_  (.A(\u_multiplier/STAGE1/pp_17_c4 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_18_2/_16_ ),
    .ZN(\u_multiplier/pp_18 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_18_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_18_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_18_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_18_c4 ));
 OAI21_X1 \u_multiplier/STAGE1/E_4_2_pp_18_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_18_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_18_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_18_2/_17_ ),
    .ZN(\u_multiplier/pp_19 [3]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_18_3/_18_  (.A(\u_multiplier/STAGE1/pp_17_c6 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_18_3/_19_  (.A1(\u_multiplier/STAGE1/_288_ ),
    .A2(\u_multiplier/STAGE1/_287_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_3/_20_  (.A(\u_multiplier/STAGE1/_288_ ),
    .B(\u_multiplier/STAGE1/_287_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_18_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_18_3/_21_  (.A1(\u_multiplier/STAGE1/_289_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_18_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_3/_22_  (.A(\u_multiplier/STAGE1/_289_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_18_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_18_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_18_3/_23_  (.A1(\u_multiplier/STAGE1/_290_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_18_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_3/_24_  (.A(\u_multiplier/STAGE1/_290_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_18_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_3/_25_  (.A(\u_multiplier/STAGE1/pp_17_c6 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_18_3/_16_ ),
    .ZN(\u_multiplier/pp_18 [6]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_18_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_18_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_18_3/_13_ ),
    .ZN(\u_multiplier/pp_19 [6]));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_18_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_18_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_18_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_18_3/_17_ ),
    .ZN(\u_multiplier/pp_19 [4]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_19_1/_18_  (.A(\u_multiplier/STAGE1/pp_18_c2 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_19_1/_19_  (.A1(\u_multiplier/STAGE1/_292_ ),
    .A2(\u_multiplier/STAGE1/_291_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_19_1/_20_  (.A(\u_multiplier/STAGE1/_292_ ),
    .B(\u_multiplier/STAGE1/_291_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_19_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_19_1/_21_  (.A1(\u_multiplier/STAGE1/_293_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_19_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_19_1/_22_  (.A(\u_multiplier/STAGE1/_293_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_19_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_19_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_19_1/_23_  (.A1(\u_multiplier/STAGE1/_294_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_19_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_19_1/_24_  (.A(\u_multiplier/STAGE1/_294_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_19_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_19_1/_25_  (.A(\u_multiplier/STAGE1/pp_18_c2 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_19_1/_16_ ),
    .ZN(\u_multiplier/pp_19 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_19_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_19_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_19_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_19_c2 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_19_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_19_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_19_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_19_1/_17_ ),
    .ZN(\u_multiplier/pp_20 [1]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_19_2/_18_  (.A(\u_multiplier/STAGE1/pp_18_c4 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_19_2/_19_  (.A1(\u_multiplier/STAGE1/_296_ ),
    .A2(\u_multiplier/STAGE1/_295_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_19_2/_20_  (.A(\u_multiplier/STAGE1/_296_ ),
    .B(\u_multiplier/STAGE1/_295_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_19_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_19_2/_21_  (.A1(\u_multiplier/STAGE1/_297_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_19_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_19_2/_22_  (.A(\u_multiplier/STAGE1/_297_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_19_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_19_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_19_2/_23_  (.A1(\u_multiplier/STAGE1/_298_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_19_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_19_2/_24_  (.A(\u_multiplier/STAGE1/_298_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_19_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_19_2/_25_  (.A(\u_multiplier/STAGE1/pp_18_c4 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_19_2/_16_ ),
    .ZN(\u_multiplier/pp_19 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_19_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_19_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_19_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_19_c4 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_19_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_19_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_19_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_19_2/_17_ ),
    .ZN(\u_multiplier/pp_20 [3]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_20_1/_18_  (.A(\u_multiplier/STAGE1/pp_19_c2 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_20_1/_19_  (.A1(\u_multiplier/STAGE1/_303_ ),
    .A2(\u_multiplier/STAGE1/_302_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_20_1/_20_  (.A(\u_multiplier/STAGE1/_303_ ),
    .B(\u_multiplier/STAGE1/_302_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_20_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_20_1/_21_  (.A1(\u_multiplier/STAGE1/_304_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_20_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_20_1/_22_  (.A(\u_multiplier/STAGE1/_304_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_20_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_20_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_20_1/_23_  (.A1(\u_multiplier/STAGE1/_305_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_20_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_20_1/_24_  (.A(\u_multiplier/STAGE1/_305_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_20_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_20_1/_25_  (.A(\u_multiplier/STAGE1/pp_19_c2 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_20_1/_16_ ),
    .ZN(\u_multiplier/pp_20 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_20_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_20_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_20_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_20_c2 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_20_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_20_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_20_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_20_1/_17_ ),
    .ZN(\u_multiplier/pp_21 [1]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_20_2/_18_  (.A(\u_multiplier/STAGE1/pp_19_c4 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_20_2/_19_  (.A1(\u_multiplier/STAGE1/_307_ ),
    .A2(\u_multiplier/STAGE1/_306_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_20_2/_20_  (.A(\u_multiplier/STAGE1/_307_ ),
    .B(\u_multiplier/STAGE1/_306_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_20_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_20_2/_21_  (.A1(\u_multiplier/STAGE1/_308_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_20_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_20_2/_22_  (.A(\u_multiplier/STAGE1/_308_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_20_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_20_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_20_2/_23_  (.A1(\u_multiplier/STAGE1/_309_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_20_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_20_2/_24_  (.A(\u_multiplier/STAGE1/_309_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_20_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_20_2/_25_  (.A(\u_multiplier/STAGE1/pp_19_c4 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_20_2/_16_ ),
    .ZN(\u_multiplier/pp_20 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_20_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_20_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_20_2/_13_ ),
    .ZN(\u_multiplier/pp_21 [4]));
 OAI21_X1 \u_multiplier/STAGE1/E_4_2_pp_20_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_20_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_20_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_20_2/_17_ ),
    .ZN(\u_multiplier/pp_21 [3]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_21_1/_18_  (.A(\u_multiplier/STAGE1/pp_20_c2 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_21_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_21_1/_19_  (.A1(\u_multiplier/STAGE1/_311_ ),
    .A2(\u_multiplier/STAGE1/_310_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_21_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_21_1/_20_  (.A(\u_multiplier/STAGE1/_311_ ),
    .B(\u_multiplier/STAGE1/_310_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_21_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_21_1/_21_  (.A1(\u_multiplier/STAGE1/_312_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_21_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_21_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_21_1/_22_  (.A(\u_multiplier/STAGE1/_312_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_21_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_21_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_21_1/_23_  (.A1(\u_multiplier/STAGE1/_313_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_21_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_21_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_21_1/_24_  (.A(\u_multiplier/STAGE1/_313_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_21_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_21_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_21_1/_25_  (.A(\u_multiplier/STAGE1/pp_20_c2 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_21_1/_16_ ),
    .ZN(\u_multiplier/pp_21 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_21_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_21_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_21_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_21_c2 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_21_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_21_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_21_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_21_1/_17_ ),
    .ZN(\u_multiplier/pp_22 [1]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_22/_18_  (.A(\u_multiplier/STAGE1/pp_21_c2 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_22/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_22/_19_  (.A1(\u_multiplier/STAGE1/_318_ ),
    .A2(\u_multiplier/STAGE1/_317_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_22/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_22/_20_  (.A(\u_multiplier/STAGE1/_318_ ),
    .B(\u_multiplier/STAGE1/_317_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_22/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_22/_21_  (.A1(\u_multiplier/STAGE1/_319_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_22/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_22/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_22/_22_  (.A(\u_multiplier/STAGE1/_319_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_22/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_22/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_22/_23_  (.A1(\u_multiplier/STAGE1/_320_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_22/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_22/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_22/_24_  (.A(\u_multiplier/STAGE1/_320_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_22/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_22/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_22/_25_  (.A(\u_multiplier/STAGE1/pp_21_c2 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_22/_16_ ),
    .ZN(\u_multiplier/pp_22 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_22/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_22/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_22/_13_ ),
    .ZN(\u_multiplier/pp_23 [4]));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_22/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_22/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_22/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_22/_17_ ),
    .ZN(\u_multiplier/pp_23 [1]));
 INV_X1 \u_multiplier/STAGE1/Full_adder_pp_16_4/_12_  (.A(\u_multiplier/STAGE1/_264_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_16_4/_08_ ));
 NAND3_X1 \u_multiplier/STAGE1/Full_adder_pp_16_4/_13_  (.A1(\u_multiplier/STAGE1/_263_ ),
    .A2(\u_multiplier/STAGE1/_262_ ),
    .A3(\u_multiplier/STAGE1/_264_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_16_4/_09_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_16_4/_14_  (.A1(\u_multiplier/STAGE1/_263_ ),
    .A2(\u_multiplier/STAGE1/_262_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_16_4/_10_ ));
 AOI21_X1 \u_multiplier/STAGE1/Full_adder_pp_16_4/_15_  (.A(\u_multiplier/STAGE1/_264_ ),
    .B1(\u_multiplier/STAGE1/_262_ ),
    .B2(\u_multiplier/STAGE1/_263_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_16_4/_11_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_16_4/_16_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_16_4/_10_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_16_4/_11_ ),
    .ZN(\u_multiplier/pp_17 [6]));
 AOI22_X2 \u_multiplier/STAGE1/Full_adder_pp_16_4/_17_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_16_4/_08_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_16_4/_10_ ),
    .B1(\u_multiplier/pp_17 [6]),
    .B2(\u_multiplier/STAGE1/Full_adder_pp_16_4/_09_ ),
    .ZN(\u_multiplier/pp_16 [7]));
 INV_X1 \u_multiplier/STAGE1/Full_adder_pp_19/_12_  (.A(\u_multiplier/STAGE1/_301_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_19/_08_ ));
 NAND3_X2 \u_multiplier/STAGE1/Full_adder_pp_19/_13_  (.A1(\u_multiplier/STAGE1/_300_ ),
    .A2(\u_multiplier/STAGE1/_299_ ),
    .A3(\u_multiplier/STAGE1/_301_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_19/_09_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_19/_14_  (.A1(\u_multiplier/STAGE1/_300_ ),
    .A2(\u_multiplier/STAGE1/_299_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_19/_10_ ));
 AOI21_X1 \u_multiplier/STAGE1/Full_adder_pp_19/_15_  (.A(\u_multiplier/STAGE1/_301_ ),
    .B1(\u_multiplier/STAGE1/_299_ ),
    .B2(\u_multiplier/STAGE1/_300_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_19/_11_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_19/_16_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_19/_10_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_19/_11_ ),
    .ZN(\u_multiplier/pp_20 [4]));
 AOI22_X4 \u_multiplier/STAGE1/Full_adder_pp_19/_17_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_19/_08_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_19/_10_ ),
    .B1(\u_multiplier/pp_20 [4]),
    .B2(\u_multiplier/STAGE1/Full_adder_pp_19/_09_ ),
    .ZN(\u_multiplier/pp_19 [5]));
 INV_X1 \u_multiplier/STAGE1/Full_adder_pp_21/_12_  (.A(\u_multiplier/STAGE1/_316_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_21/_08_ ));
 NAND3_X2 \u_multiplier/STAGE1/Full_adder_pp_21/_13_  (.A1(\u_multiplier/STAGE1/_315_ ),
    .A2(\u_multiplier/STAGE1/_314_ ),
    .A3(\u_multiplier/STAGE1/_316_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_21/_09_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_21/_14_  (.A1(\u_multiplier/STAGE1/_315_ ),
    .A2(\u_multiplier/STAGE1/_314_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_21/_10_ ));
 AOI21_X1 \u_multiplier/STAGE1/Full_adder_pp_21/_15_  (.A(\u_multiplier/STAGE1/_316_ ),
    .B1(\u_multiplier/STAGE1/_314_ ),
    .B2(\u_multiplier/STAGE1/_315_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_21/_11_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_21/_16_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_21/_10_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_21/_11_ ),
    .ZN(\u_multiplier/pp_22 [4]));
 AOI22_X4 \u_multiplier/STAGE1/Full_adder_pp_21/_17_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_21/_08_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_21/_10_ ),
    .B1(\u_multiplier/pp_22 [4]),
    .B2(\u_multiplier/STAGE1/Full_adder_pp_21/_09_ ),
    .ZN(\u_multiplier/pp_21 [2]));
 INV_X1 \u_multiplier/STAGE1/Full_adder_pp_23/_12_  (.A(\u_multiplier/STAGE1/_323_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_23/_08_ ));
 NAND3_X2 \u_multiplier/STAGE1/Full_adder_pp_23/_13_  (.A1(\u_multiplier/STAGE1/_322_ ),
    .A2(\u_multiplier/STAGE1/_321_ ),
    .A3(\u_multiplier/STAGE1/_323_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_23/_09_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_23/_14_  (.A1(\u_multiplier/STAGE1/_322_ ),
    .A2(\u_multiplier/STAGE1/_321_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_23/_10_ ));
 AOI21_X1 \u_multiplier/STAGE1/Full_adder_pp_23/_15_  (.A(\u_multiplier/STAGE1/_323_ ),
    .B1(\u_multiplier/STAGE1/_321_ ),
    .B2(\u_multiplier/STAGE1/_322_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_23/_11_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_23/_16_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_23/_10_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_23/_11_ ),
    .ZN(\u_multiplier/pp_24 [0]));
 AOI22_X4 \u_multiplier/STAGE1/Full_adder_pp_23/_17_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_23/_08_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_23/_10_ ),
    .B1(\u_multiplier/pp_24 [0]),
    .B2(\u_multiplier/STAGE1/Full_adder_pp_23/_09_ ),
    .ZN(\u_multiplier/pp_23 [0]));
 AND2_X1 \u_multiplier/STAGE1/Half_adder_pp_10/_4_  (.A1(\u_multiplier/STAGE1/_189_ ),
    .A2(\u_multiplier/STAGE1/_188_ ),
    .ZN(\u_multiplier/pp_11 [3]));
 XOR2_X2 \u_multiplier/STAGE1/Half_adder_pp_10/_5_  (.A(\u_multiplier/STAGE1/_189_ ),
    .B(\u_multiplier/STAGE1/_188_ ),
    .Z(\u_multiplier/pp_10 [0]));
 AND2_X1 \u_multiplier/STAGE1/Half_adder_pp_12/_4_  (.A1(\u_multiplier/STAGE1/_207_ ),
    .A2(\u_multiplier/STAGE1/_206_ ),
    .ZN(\u_multiplier/pp_13 [7]));
 XOR2_X2 \u_multiplier/STAGE1/Half_adder_pp_12/_5_  (.A(\u_multiplier/STAGE1/_207_ ),
    .B(\u_multiplier/STAGE1/_206_ ),
    .Z(\u_multiplier/pp_12 [0]));
 AND2_X1 \u_multiplier/STAGE1/Half_adder_pp_14/_4_  (.A1(\u_multiplier/STAGE1/_233_ ),
    .A2(\u_multiplier/STAGE1/_232_ ),
    .ZN(\u_multiplier/pp_15 [7]));
 XOR2_X2 \u_multiplier/STAGE1/Half_adder_pp_14/_5_  (.A(\u_multiplier/STAGE1/_233_ ),
    .B(\u_multiplier/STAGE1/_232_ ),
    .Z(\u_multiplier/pp_14 [5]));
 AND2_X1 \u_multiplier/STAGE1/Half_adder_pp_17/_4_  (.A1(\u_multiplier/STAGE1/_278_ ),
    .A2(\u_multiplier/STAGE1/_277_ ),
    .ZN(\u_multiplier/pp_18 [4]));
 XOR2_X2 \u_multiplier/STAGE1/Half_adder_pp_17/_5_  (.A(\u_multiplier/STAGE1/_278_ ),
    .B(\u_multiplier/STAGE1/_277_ ),
    .Z(\u_multiplier/pp_17 [7]));
 AND2_X1 \u_multiplier/STAGE1/Half_adder_pp_8/_4_  (.A1(\u_multiplier/STAGE1/_179_ ),
    .A2(\u_multiplier/STAGE1/_178_ ),
    .ZN(\u_multiplier/pp_9 [3]));
 XOR2_X2 \u_multiplier/STAGE1/Half_adder_pp_8/_5_  (.A(\u_multiplier/STAGE1/_179_ ),
    .B(\u_multiplier/STAGE1/_178_ ),
    .Z(\u_multiplier/pp_8 [0]));
 AND2_X1 \u_multiplier/STAGE1/_434_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[0]),
    .ZN(\u_multiplier/s_0 ));
 AND2_X1 \u_multiplier/STAGE1/_435_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[1]),
    .ZN(\u_multiplier/s_1 [0]));
 AND2_X1 \u_multiplier/STAGE1/_436_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[1]),
    .ZN(\u_multiplier/s_1 [1]));
 AND2_X1 \u_multiplier/STAGE1/_437_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[2]),
    .ZN(\u_multiplier/s_2 [0]));
 AND2_X1 \u_multiplier/STAGE1/_438_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[1]),
    .ZN(\u_multiplier/s_2 [1]));
 AND2_X1 \u_multiplier/STAGE1/_439_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[2]),
    .ZN(\u_multiplier/s_2 [2]));
 AND2_X1 \u_multiplier/STAGE1/_440_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[3]),
    .ZN(\u_multiplier/s_3 [0]));
 AND2_X1 \u_multiplier/STAGE1/_441_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[2]),
    .ZN(\u_multiplier/s_3 [1]));
 AND2_X1 \u_multiplier/STAGE1/_442_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[2]),
    .ZN(\u_multiplier/s_3 [2]));
 AND2_X1 \u_multiplier/STAGE1/_443_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[3]),
    .ZN(\u_multiplier/s_3 [3]));
 AND2_X1 \u_multiplier/STAGE1/_444_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[4]),
    .ZN(\u_multiplier/pp_4 [0]));
 AND2_X1 \u_multiplier/STAGE1/_445_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[3]),
    .ZN(\u_multiplier/pp_4 [1]));
 AND2_X1 \u_multiplier/STAGE1/_446_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[2]),
    .ZN(\u_multiplier/s_4 [1]));
 AND2_X1 \u_multiplier/STAGE1/_447_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[3]),
    .ZN(\u_multiplier/s_4 [2]));
 AND2_X1 \u_multiplier/STAGE1/_448_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[4]),
    .ZN(\u_multiplier/s_4 [3]));
 AND2_X1 \u_multiplier/STAGE1/_449_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[5]),
    .ZN(\u_multiplier/pp_5 [0]));
 AND2_X1 \u_multiplier/STAGE1/_450_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[4]),
    .ZN(\u_multiplier/pp_5 [1]));
 AND2_X1 \u_multiplier/STAGE1/_451_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[3]),
    .ZN(\u_multiplier/pp_5 [2]));
 AND2_X1 \u_multiplier/STAGE1/_452_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[3]),
    .ZN(\u_multiplier/pp_5 [3]));
 AND2_X1 \u_multiplier/STAGE1/_453_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[4]),
    .ZN(\u_multiplier/s_5 [1]));
 AND2_X1 \u_multiplier/STAGE1/_454_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[5]),
    .ZN(\u_multiplier/s_5 [2]));
 AND2_X1 \u_multiplier/STAGE1/_455_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[6]),
    .ZN(\u_multiplier/pp_6 [0]));
 AND2_X1 \u_multiplier/STAGE1/_456_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[5]),
    .ZN(\u_multiplier/pp_6 [1]));
 AND2_X1 \u_multiplier/STAGE1/_457_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[4]),
    .ZN(\u_multiplier/pp_6 [2]));
 AND2_X1 \u_multiplier/STAGE1/_458_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[3]),
    .ZN(\u_multiplier/pp_6 [3]));
 AND2_X1 \u_multiplier/STAGE1/_459_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[4]),
    .ZN(\u_multiplier/pp_6 [4]));
 AND2_X1 \u_multiplier/STAGE1/_460_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[5]),
    .ZN(\u_multiplier/pp_6 [5]));
 AND2_X1 \u_multiplier/STAGE1/_461_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[6]),
    .ZN(\u_multiplier/s_6 [2]));
 AND2_X1 \u_multiplier/STAGE1/_462_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[7]),
    .ZN(\u_multiplier/pp_7 [0]));
 AND2_X1 \u_multiplier/STAGE1/_463_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[6]),
    .ZN(\u_multiplier/pp_7 [1]));
 AND2_X1 \u_multiplier/STAGE1/_464_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[5]),
    .ZN(\u_multiplier/pp_7 [2]));
 AND2_X1 \u_multiplier/STAGE1/_465_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[4]),
    .ZN(\u_multiplier/pp_7 [3]));
 AND2_X1 \u_multiplier/STAGE1/_466_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[4]),
    .ZN(\u_multiplier/pp_7 [4]));
 AND2_X1 \u_multiplier/STAGE1/_467_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[5]),
    .ZN(\u_multiplier/pp_7 [5]));
 AND2_X1 \u_multiplier/STAGE1/_468_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[6]),
    .ZN(\u_multiplier/pp_7 [6]));
 AND2_X1 \u_multiplier/STAGE1/_469_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[7]),
    .ZN(\u_multiplier/pp_7 [7]));
 AND2_X1 \u_multiplier/STAGE1/_470_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[6]),
    .ZN(\u_multiplier/pp_8 [1]));
 AND2_X1 \u_multiplier/STAGE1/_471_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[5]),
    .ZN(\u_multiplier/pp_8 [2]));
 AND2_X1 \u_multiplier/STAGE1/_472_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[4]),
    .ZN(\u_multiplier/pp_8 [3]));
 AND2_X1 \u_multiplier/STAGE1/_473_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[5]),
    .ZN(\u_multiplier/pp_8 [4]));
 AND2_X1 \u_multiplier/STAGE1/_474_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[6]),
    .ZN(\u_multiplier/pp_8 [5]));
 AND2_X1 \u_multiplier/STAGE1/_475_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[7]),
    .ZN(\u_multiplier/pp_8 [6]));
 AND2_X1 \u_multiplier/STAGE1/_476_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/pp_8 [7]));
 AND2_X1 \u_multiplier/STAGE1/_477_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[5]),
    .ZN(\u_multiplier/pp_9 [1]));
 AND2_X1 \u_multiplier/STAGE1/_478_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[5]),
    .ZN(\u_multiplier/pp_9 [2]));
 AND2_X1 \u_multiplier/STAGE1/_479_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[6]),
    .ZN(\u_multiplier/pp_9 [4]));
 AND2_X1 \u_multiplier/STAGE1/_480_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[7]),
    .ZN(\u_multiplier/pp_9 [5]));
 AND2_X1 \u_multiplier/STAGE1/_481_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/pp_9 [6]));
 AND2_X1 \u_multiplier/STAGE1/_482_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/pp_9 [7]));
 AND2_X1 \u_multiplier/STAGE1/_483_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[6]),
    .ZN(\u_multiplier/pp_10 [2]));
 AND2_X1 \u_multiplier/STAGE1/_484_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[7]),
    .ZN(\u_multiplier/pp_10 [4]));
 AND2_X1 \u_multiplier/STAGE1/_485_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/pp_10 [5]));
 AND2_X1 \u_multiplier/STAGE1/_486_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/pp_10 [6]));
 AND2_X1 \u_multiplier/STAGE1/_487_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/pp_10 [7]));
 AND2_X1 \u_multiplier/STAGE1/_488_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/pp_11 [4]));
 AND2_X1 \u_multiplier/STAGE1/_489_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/pp_11 [5]));
 AND2_X1 \u_multiplier/STAGE1/_490_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/pp_11 [6]));
 AND2_X1 \u_multiplier/STAGE1/_491_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/pp_11 [7]));
 AND2_X1 \u_multiplier/STAGE1/_492_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/pp_12 [5]));
 AND2_X1 \u_multiplier/STAGE1/_493_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/pp_12 [6]));
 AND2_X1 \u_multiplier/STAGE1/_494_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/pp_12 [7]));
 AND2_X1 \u_multiplier/STAGE1/_495_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/pp_13 [5]));
 AND2_X1 \u_multiplier/STAGE1/_496_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/pp_13 [6]));
 AND2_X1 \u_multiplier/STAGE1/_497_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/pp_14 [6]));
 AND2_X1 \u_multiplier/STAGE1/_498_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/pp_18 [7]));
 AND2_X1 \u_multiplier/STAGE1/_499_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/pp_19 [7]));
 AND2_X1 \u_multiplier/STAGE1/_500_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/pp_20 [5]));
 AND2_X1 \u_multiplier/STAGE1/_501_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/pp_20 [6]));
 AND2_X1 \u_multiplier/STAGE1/_502_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/pp_20 [7]));
 AND2_X1 \u_multiplier/STAGE1/_503_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/pp_21 [5]));
 AND2_X1 \u_multiplier/STAGE1/_504_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/pp_21 [6]));
 AND2_X1 \u_multiplier/STAGE1/_505_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/pp_21 [7]));
 AND2_X1 \u_multiplier/STAGE1/_506_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/pp_22 [2]));
 AND2_X1 \u_multiplier/STAGE1/_507_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/pp_22 [3]));
 AND2_X1 \u_multiplier/STAGE1/_508_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/pp_22 [5]));
 AND2_X1 \u_multiplier/STAGE1/_509_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/pp_22 [6]));
 AND2_X1 \u_multiplier/STAGE1/_510_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/pp_22 [7]));
 AND2_X1 \u_multiplier/STAGE1/_511_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/pp_23 [2]));
 AND2_X1 \u_multiplier/STAGE1/_512_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/pp_23 [3]));
 AND2_X1 \u_multiplier/STAGE1/_513_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/pp_23 [5]));
 AND2_X1 \u_multiplier/STAGE1/_514_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/pp_23 [6]));
 AND2_X1 \u_multiplier/STAGE1/_515_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/pp_23 [7]));
 AND2_X1 \u_multiplier/STAGE1/_516_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/pp_24 [1]));
 AND2_X1 \u_multiplier/STAGE1/_517_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/pp_24 [2]));
 AND2_X1 \u_multiplier/STAGE1/_518_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/pp_24 [3]));
 AND2_X1 \u_multiplier/STAGE1/_519_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/pp_24 [4]));
 AND2_X1 \u_multiplier/STAGE1/_520_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/pp_24 [5]));
 AND2_X1 \u_multiplier/STAGE1/_521_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/pp_24 [6]));
 AND2_X1 \u_multiplier/STAGE1/_522_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/pp_24 [7]));
 AND2_X1 \u_multiplier/STAGE1/_523_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/pp_25 [0]));
 AND2_X1 \u_multiplier/STAGE1/_524_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/pp_25 [1]));
 AND2_X1 \u_multiplier/STAGE1/_525_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/pp_25 [2]));
 AND2_X1 \u_multiplier/STAGE1/_526_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/pp_25 [3]));
 AND2_X1 \u_multiplier/STAGE1/_527_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/pp_25 [4]));
 AND2_X1 \u_multiplier/STAGE1/_528_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/pp_25 [5]));
 AND2_X1 \u_multiplier/STAGE1/_529_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/pp_26 [0]));
 AND2_X1 \u_multiplier/STAGE1/_530_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/pp_26 [1]));
 AND2_X1 \u_multiplier/STAGE1/_531_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/pp_26 [2]));
 AND2_X1 \u_multiplier/STAGE1/_532_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/pp_26 [3]));
 AND2_X1 \u_multiplier/STAGE1/_533_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/s_26 [1]));
 AND2_X1 \u_multiplier/STAGE1/_534_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/pp_27 [0]));
 AND2_X1 \u_multiplier/STAGE1/_535_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/pp_27 [1]));
 AND2_X1 \u_multiplier/STAGE1/_536_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/pp_27 [2]));
 AND2_X1 \u_multiplier/STAGE1/_537_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/s_27 [1]));
 AND2_X1 \u_multiplier/STAGE1/_538_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/s_28 [1]));
 AND2_X1 \u_multiplier/STAGE1/_539_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/s_28 [2]));
 AND2_X1 \u_multiplier/STAGE1/_540_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/s_28 [3]));
 AND2_X1 \u_multiplier/STAGE1/_541_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/s_29 [0]));
 AND2_X1 \u_multiplier/STAGE1/_542_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/s_29 [1]));
 AND2_X1 \u_multiplier/STAGE1/_543_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/s_30 ));
 AND2_X1 \u_multiplier/STAGE1/_544_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/STAGE1/_178_ ));
 AND2_X1 \u_multiplier/STAGE1/_545_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[7]),
    .ZN(\u_multiplier/STAGE1/_179_ ));
 AND2_X1 \u_multiplier/STAGE1/_546_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/STAGE1/_180_ ));
 AND2_X1 \u_multiplier/STAGE1/_547_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/STAGE1/_181_ ));
 AND2_X1 \u_multiplier/STAGE1/_548_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[7]),
    .ZN(\u_multiplier/STAGE1/_182_ ));
 AND2_X1 \u_multiplier/STAGE1/_549_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[6]),
    .ZN(\u_multiplier/STAGE1/_183_ ));
 AND2_X1 \u_multiplier/STAGE1/_550_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/STAGE1/_184_ ));
 AND2_X1 \u_multiplier/STAGE1/_551_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/STAGE1/_185_ ));
 AND2_X1 \u_multiplier/STAGE1/_552_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/STAGE1/_186_ ));
 AND2_X1 \u_multiplier/STAGE1/_553_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[7]),
    .ZN(\u_multiplier/STAGE1/_187_ ));
 AND2_X1 \u_multiplier/STAGE1/_554_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[6]),
    .ZN(\u_multiplier/STAGE1/_188_ ));
 AND2_X1 \u_multiplier/STAGE1/_555_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[5]),
    .ZN(\u_multiplier/STAGE1/_189_ ));
 AND2_X1 \u_multiplier/STAGE1/_556_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/STAGE1/_190_ ));
 AND2_X1 \u_multiplier/STAGE1/_557_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/STAGE1/_191_ ));
 AND2_X1 \u_multiplier/STAGE1/_558_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/STAGE1/_192_ ));
 AND2_X1 \u_multiplier/STAGE1/_559_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/STAGE1/_193_ ));
 AND2_X1 \u_multiplier/STAGE1/_560_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[7]),
    .ZN(\u_multiplier/STAGE1/_194_ ));
 AND2_X1 \u_multiplier/STAGE1/_561_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[6]),
    .ZN(\u_multiplier/STAGE1/_195_ ));
 AND2_X1 \u_multiplier/STAGE1/_562_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[6]),
    .ZN(\u_multiplier/STAGE1/_196_ ));
 AND2_X1 \u_multiplier/STAGE1/_563_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[7]),
    .ZN(\u_multiplier/STAGE1/_197_ ));
 AND2_X1 \u_multiplier/STAGE1/_564_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/STAGE1/_198_ ));
 AND2_X1 \u_multiplier/STAGE1/_565_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/STAGE1/_199_ ));
 AND2_X1 \u_multiplier/STAGE1/_566_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/STAGE1/_200_ ));
 AND2_X1 \u_multiplier/STAGE1/_567_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/STAGE1/_201_ ));
 AND2_X1 \u_multiplier/STAGE1/_568_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/STAGE1/_202_ ));
 AND2_X1 \u_multiplier/STAGE1/_569_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[7]),
    .ZN(\u_multiplier/STAGE1/_203_ ));
 AND2_X1 \u_multiplier/STAGE1/_570_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[6]),
    .ZN(\u_multiplier/STAGE1/_204_ ));
 AND2_X1 \u_multiplier/STAGE1/_571_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[7]),
    .ZN(\u_multiplier/STAGE1/_205_ ));
 AND2_X1 \u_multiplier/STAGE1/_572_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/STAGE1/_206_ ));
 AND2_X1 \u_multiplier/STAGE1/_573_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/STAGE1/_207_ ));
 AND2_X1 \u_multiplier/STAGE1/_574_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/STAGE1/_208_ ));
 AND2_X1 \u_multiplier/STAGE1/_575_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/STAGE1/_209_ ));
 AND2_X1 \u_multiplier/STAGE1/_576_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/STAGE1/_210_ ));
 AND2_X1 \u_multiplier/STAGE1/_577_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/STAGE1/_211_ ));
 AND2_X1 \u_multiplier/STAGE1/_578_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/STAGE1/_212_ ));
 AND2_X1 \u_multiplier/STAGE1/_579_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/STAGE1/_213_ ));
 AND2_X1 \u_multiplier/STAGE1/_580_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[7]),
    .ZN(\u_multiplier/STAGE1/_214_ ));
 AND2_X1 \u_multiplier/STAGE1/_581_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[7]),
    .ZN(\u_multiplier/STAGE1/_215_ ));
 AND2_X1 \u_multiplier/STAGE1/_582_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/STAGE1/_216_ ));
 AND2_X1 \u_multiplier/STAGE1/_583_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/STAGE1/_217_ ));
 AND2_X1 \u_multiplier/STAGE1/_584_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/STAGE1/_218_ ));
 AND2_X1 \u_multiplier/STAGE1/_585_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/STAGE1/_219_ ));
 AND2_X1 \u_multiplier/STAGE1/_586_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/STAGE1/_220_ ));
 AND2_X1 \u_multiplier/STAGE1/_587_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/STAGE1/_221_ ));
 AND2_X1 \u_multiplier/STAGE1/_588_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/STAGE1/_222_ ));
 AND2_X1 \u_multiplier/STAGE1/_589_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/STAGE1/_223_ ));
 AND2_X1 \u_multiplier/STAGE1/_590_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/STAGE1/_224_ ));
 AND2_X1 \u_multiplier/STAGE1/_591_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/STAGE1/_225_ ));
 AND2_X1 \u_multiplier/STAGE1/_592_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/STAGE1/_226_ ));
 AND2_X1 \u_multiplier/STAGE1/_593_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[7]),
    .ZN(\u_multiplier/STAGE1/_227_ ));
 AND2_X1 \u_multiplier/STAGE1/_594_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/STAGE1/_228_ ));
 AND2_X1 \u_multiplier/STAGE1/_595_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/STAGE1/_229_ ));
 AND2_X1 \u_multiplier/STAGE1/_596_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/STAGE1/_230_ ));
 AND2_X1 \u_multiplier/STAGE1/_597_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/STAGE1/_231_ ));
 AND2_X1 \u_multiplier/STAGE1/_598_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/STAGE1/_232_ ));
 AND2_X1 \u_multiplier/STAGE1/_599_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/STAGE1/_233_ ));
 AND2_X1 \u_multiplier/STAGE1/_600_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/STAGE1/_234_ ));
 AND2_X1 \u_multiplier/STAGE1/_601_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/STAGE1/_235_ ));
 AND2_X1 \u_multiplier/STAGE1/_602_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/STAGE1/_236_ ));
 AND2_X1 \u_multiplier/STAGE1/_603_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/STAGE1/_237_ ));
 AND2_X1 \u_multiplier/STAGE1/_604_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/STAGE1/_238_ ));
 AND2_X1 \u_multiplier/STAGE1/_605_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/STAGE1/_239_ ));
 AND2_X1 \u_multiplier/STAGE1/_606_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/STAGE1/_240_ ));
 AND2_X1 \u_multiplier/STAGE1/_607_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/STAGE1/_241_ ));
 AND2_X1 \u_multiplier/STAGE1/_608_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/STAGE1/_242_ ));
 AND2_X1 \u_multiplier/STAGE1/_609_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/STAGE1/_243_ ));
 AND2_X1 \u_multiplier/STAGE1/_610_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/STAGE1/_244_ ));
 AND2_X1 \u_multiplier/STAGE1/_611_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/STAGE1/_245_ ));
 AND2_X1 \u_multiplier/STAGE1/_612_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/STAGE1/_246_ ));
 AND2_X1 \u_multiplier/STAGE1/_613_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/STAGE1/_247_ ));
 AND2_X1 \u_multiplier/STAGE1/_614_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/STAGE1/_248_ ));
 AND2_X1 \u_multiplier/STAGE1/_615_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/STAGE1/_249_ ));
 AND2_X1 \u_multiplier/STAGE1/_616_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/STAGE1/_250_ ));
 AND2_X1 \u_multiplier/STAGE1/_617_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/STAGE1/_251_ ));
 AND2_X1 \u_multiplier/STAGE1/_618_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/STAGE1/_252_ ));
 AND2_X1 \u_multiplier/STAGE1/_619_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/STAGE1/_253_ ));
 AND2_X1 \u_multiplier/STAGE1/_620_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/STAGE1/_254_ ));
 AND2_X1 \u_multiplier/STAGE1/_621_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/STAGE1/_255_ ));
 AND2_X1 \u_multiplier/STAGE1/_622_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/STAGE1/_256_ ));
 AND2_X1 \u_multiplier/STAGE1/_623_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/STAGE1/_257_ ));
 AND2_X1 \u_multiplier/STAGE1/_624_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/STAGE1/_258_ ));
 AND2_X1 \u_multiplier/STAGE1/_625_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/STAGE1/_259_ ));
 AND2_X1 \u_multiplier/STAGE1/_626_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/STAGE1/_260_ ));
 AND2_X1 \u_multiplier/STAGE1/_627_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/STAGE1/_261_ ));
 AND2_X1 \u_multiplier/STAGE1/_628_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/STAGE1/_262_ ));
 AND2_X1 \u_multiplier/STAGE1/_629_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/STAGE1/_263_ ));
 AND2_X1 \u_multiplier/STAGE1/_630_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/STAGE1/_264_ ));
 AND2_X1 \u_multiplier/STAGE1/_631_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/STAGE1/_265_ ));
 AND2_X1 \u_multiplier/STAGE1/_632_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/STAGE1/_266_ ));
 AND2_X1 \u_multiplier/STAGE1/_633_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/STAGE1/_267_ ));
 AND2_X1 \u_multiplier/STAGE1/_634_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/STAGE1/_268_ ));
 AND2_X1 \u_multiplier/STAGE1/_635_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/STAGE1/_269_ ));
 AND2_X1 \u_multiplier/STAGE1/_636_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/STAGE1/_270_ ));
 AND2_X1 \u_multiplier/STAGE1/_637_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/STAGE1/_271_ ));
 AND2_X1 \u_multiplier/STAGE1/_638_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/STAGE1/_272_ ));
 AND2_X1 \u_multiplier/STAGE1/_639_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/STAGE1/_273_ ));
 AND2_X1 \u_multiplier/STAGE1/_640_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/STAGE1/_274_ ));
 AND2_X1 \u_multiplier/STAGE1/_641_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/STAGE1/_275_ ));
 AND2_X1 \u_multiplier/STAGE1/_642_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/STAGE1/_276_ ));
 AND2_X1 \u_multiplier/STAGE1/_643_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/STAGE1/_277_ ));
 AND2_X1 \u_multiplier/STAGE1/_644_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/STAGE1/_278_ ));
 AND2_X1 \u_multiplier/STAGE1/_645_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/STAGE1/_279_ ));
 AND2_X1 \u_multiplier/STAGE1/_646_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/STAGE1/_280_ ));
 AND2_X1 \u_multiplier/STAGE1/_647_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/STAGE1/_281_ ));
 AND2_X1 \u_multiplier/STAGE1/_648_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/STAGE1/_282_ ));
 AND2_X1 \u_multiplier/STAGE1/_649_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/STAGE1/_283_ ));
 AND2_X1 \u_multiplier/STAGE1/_650_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/STAGE1/_284_ ));
 AND2_X1 \u_multiplier/STAGE1/_651_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/STAGE1/_285_ ));
 AND2_X1 \u_multiplier/STAGE1/_652_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/STAGE1/_286_ ));
 AND2_X1 \u_multiplier/STAGE1/_653_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/STAGE1/_287_ ));
 AND2_X1 \u_multiplier/STAGE1/_654_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/STAGE1/_288_ ));
 AND2_X1 \u_multiplier/STAGE1/_655_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/STAGE1/_289_ ));
 AND2_X1 \u_multiplier/STAGE1/_656_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/STAGE1/_290_ ));
 AND2_X1 \u_multiplier/STAGE1/_657_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/STAGE1/_291_ ));
 AND2_X1 \u_multiplier/STAGE1/_658_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/STAGE1/_292_ ));
 AND2_X1 \u_multiplier/STAGE1/_659_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/STAGE1/_293_ ));
 AND2_X1 \u_multiplier/STAGE1/_660_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/STAGE1/_294_ ));
 AND2_X1 \u_multiplier/STAGE1/_661_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/STAGE1/_295_ ));
 AND2_X1 \u_multiplier/STAGE1/_662_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/STAGE1/_296_ ));
 AND2_X1 \u_multiplier/STAGE1/_663_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/STAGE1/_297_ ));
 AND2_X1 \u_multiplier/STAGE1/_664_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/STAGE1/_298_ ));
 AND2_X1 \u_multiplier/STAGE1/_665_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/STAGE1/_299_ ));
 AND2_X1 \u_multiplier/STAGE1/_666_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/STAGE1/_300_ ));
 AND2_X1 \u_multiplier/STAGE1/_667_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/STAGE1/_301_ ));
 AND2_X1 \u_multiplier/STAGE1/_668_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/STAGE1/_302_ ));
 AND2_X1 \u_multiplier/STAGE1/_669_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/STAGE1/_303_ ));
 AND2_X1 \u_multiplier/STAGE1/_670_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/STAGE1/_304_ ));
 AND2_X1 \u_multiplier/STAGE1/_671_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/STAGE1/_305_ ));
 AND2_X1 \u_multiplier/STAGE1/_672_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/STAGE1/_306_ ));
 AND2_X1 \u_multiplier/STAGE1/_673_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/STAGE1/_307_ ));
 AND2_X1 \u_multiplier/STAGE1/_674_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/STAGE1/_308_ ));
 AND2_X1 \u_multiplier/STAGE1/_675_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/STAGE1/_309_ ));
 AND2_X1 \u_multiplier/STAGE1/_676_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/STAGE1/_310_ ));
 AND2_X1 \u_multiplier/STAGE1/_677_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/STAGE1/_311_ ));
 AND2_X1 \u_multiplier/STAGE1/_678_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/STAGE1/_312_ ));
 AND2_X1 \u_multiplier/STAGE1/_679_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/STAGE1/_313_ ));
 AND2_X1 \u_multiplier/STAGE1/_680_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/STAGE1/_314_ ));
 AND2_X1 \u_multiplier/STAGE1/_681_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/STAGE1/_315_ ));
 AND2_X1 \u_multiplier/STAGE1/_682_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/STAGE1/_316_ ));
 AND2_X1 \u_multiplier/STAGE1/_683_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/STAGE1/_317_ ));
 AND2_X1 \u_multiplier/STAGE1/_684_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/STAGE1/_318_ ));
 AND2_X1 \u_multiplier/STAGE1/_685_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/STAGE1/_319_ ));
 AND2_X1 \u_multiplier/STAGE1/_686_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/STAGE1/_320_ ));
 AND2_X1 \u_multiplier/STAGE1/_687_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/STAGE1/_321_ ));
 AND2_X1 \u_multiplier/STAGE1/_688_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/STAGE1/_322_ ));
 AND2_X1 \u_multiplier/STAGE1/_689_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/STAGE1/_323_ ));
 NAND3_X1 \u_multiplier/STAGE2/ACCI1_pp_10_1/_21_  (.A1(\u_multiplier/pp_10 [1]),
    .A2(\u_multiplier/pp_10 [0]),
    .A3(\u_multiplier/pp_10 [2]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_10_1/_18_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_10_1/_22_  (.A(\u_multiplier/pp_10 [1]),
    .B(\u_multiplier/pp_10 [0]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_10_1/_19_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_10_1/_23_  (.A(\u_multiplier/pp_10 [2]),
    .B(\u_multiplier/pp_10 [3]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_10_1/_20_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_10_1/_24_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_10_1/_19_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_10_1/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_10_1/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE2/ACCI1_pp_10_1/_25_  (.A(\u_multiplier/STAGE2/ACCI1_pp_10_1/_19_ ),
    .B(\u_multiplier/STAGE2/ACCI1_pp_10_1/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_10_1/_16_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_10_1/_26_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_10_1/_18_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_10_1/_16_ ),
    .ZN(\u_multiplier/s_10 [1]));
 AOI22_X1 \u_multiplier/STAGE2/ACCI1_pp_10_1/_27_  (.A1(\u_multiplier/pp_10 [1]),
    .A2(\u_multiplier/pp_10 [0]),
    .B1(\u_multiplier/pp_10 [2]),
    .B2(\u_multiplier/pp_10 [3]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_10_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_10_1/_28_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_10_1/_15_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_10_1/_17_ ),
    .ZN(\u_multiplier/s_11 [2]));
 NAND3_X1 \u_multiplier/STAGE2/ACCI1_pp_10_2/_21_  (.A1(\u_multiplier/pp_10 [5]),
    .A2(\u_multiplier/pp_10 [4]),
    .A3(\u_multiplier/pp_10 [6]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_10_2/_18_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_10_2/_22_  (.A(\u_multiplier/pp_10 [5]),
    .B(\u_multiplier/pp_10 [4]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_10_2/_19_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_10_2/_23_  (.A(\u_multiplier/pp_10 [6]),
    .B(\u_multiplier/pp_10 [7]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_10_2/_20_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_10_2/_24_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_10_2/_19_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_10_2/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_10_2/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE2/ACCI1_pp_10_2/_25_  (.A(\u_multiplier/STAGE2/ACCI1_pp_10_2/_19_ ),
    .B(\u_multiplier/STAGE2/ACCI1_pp_10_2/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_10_2/_16_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_10_2/_26_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_10_2/_18_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_10_2/_16_ ),
    .ZN(\u_multiplier/s_10 [0]));
 AOI22_X1 \u_multiplier/STAGE2/ACCI1_pp_10_2/_27_  (.A1(\u_multiplier/pp_10 [5]),
    .A2(\u_multiplier/pp_10 [4]),
    .B1(\u_multiplier/pp_10 [6]),
    .B2(\u_multiplier/pp_10 [7]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_10_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_10_2/_28_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_10_2/_15_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_10_2/_17_ ),
    .ZN(\u_multiplier/s_11 [3]));
 NAND3_X1 \u_multiplier/STAGE2/ACCI1_pp_11_1/_21_  (.A1(\u_multiplier/pp_11 [1]),
    .A2(\u_multiplier/pp_11 [0]),
    .A3(\u_multiplier/pp_11 [2]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_11_1/_18_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_11_1/_22_  (.A(\u_multiplier/pp_11 [1]),
    .B(\u_multiplier/pp_11 [0]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_11_1/_19_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_11_1/_23_  (.A(\u_multiplier/pp_11 [2]),
    .B(\u_multiplier/pp_11 [3]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_11_1/_20_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_11_1/_24_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_11_1/_19_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_11_1/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_11_1/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE2/ACCI1_pp_11_1/_25_  (.A(\u_multiplier/STAGE2/ACCI1_pp_11_1/_19_ ),
    .B(\u_multiplier/STAGE2/ACCI1_pp_11_1/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_11_1/_16_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_11_1/_26_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_11_1/_18_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_11_1/_16_ ),
    .ZN(\u_multiplier/s_11 [1]));
 AOI22_X1 \u_multiplier/STAGE2/ACCI1_pp_11_1/_27_  (.A1(\u_multiplier/pp_11 [1]),
    .A2(\u_multiplier/pp_11 [0]),
    .B1(\u_multiplier/pp_11 [2]),
    .B2(\u_multiplier/pp_11 [3]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_11_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_11_1/_28_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_11_1/_15_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_11_1/_17_ ),
    .ZN(\u_multiplier/s_12 [2]));
 NAND3_X1 \u_multiplier/STAGE2/ACCI1_pp_11_2/_21_  (.A1(\u_multiplier/pp_11 [5]),
    .A2(\u_multiplier/pp_11 [4]),
    .A3(\u_multiplier/pp_11 [6]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_11_2/_18_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_11_2/_22_  (.A(\u_multiplier/pp_11 [5]),
    .B(\u_multiplier/pp_11 [4]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_11_2/_19_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_11_2/_23_  (.A(\u_multiplier/pp_11 [6]),
    .B(\u_multiplier/pp_11 [7]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_11_2/_20_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_11_2/_24_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_11_2/_19_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_11_2/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_11_2/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE2/ACCI1_pp_11_2/_25_  (.A(\u_multiplier/STAGE2/ACCI1_pp_11_2/_19_ ),
    .B(\u_multiplier/STAGE2/ACCI1_pp_11_2/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_11_2/_16_ ));
 NAND2_X2 \u_multiplier/STAGE2/ACCI1_pp_11_2/_26_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_11_2/_18_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_11_2/_16_ ),
    .ZN(\u_multiplier/s_11 [0]));
 AOI22_X1 \u_multiplier/STAGE2/ACCI1_pp_11_2/_27_  (.A1(\u_multiplier/pp_11 [5]),
    .A2(\u_multiplier/pp_11 [4]),
    .B1(\u_multiplier/pp_11 [6]),
    .B2(\u_multiplier/pp_11 [7]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_11_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_11_2/_28_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_11_2/_15_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_11_2/_17_ ),
    .ZN(\u_multiplier/s_12 [3]));
 NAND3_X1 \u_multiplier/STAGE2/ACCI1_pp_12_1/_21_  (.A1(\u_multiplier/pp_12 [1]),
    .A2(\u_multiplier/pp_12 [0]),
    .A3(\u_multiplier/pp_12 [2]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_12_1/_18_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_12_1/_22_  (.A(\u_multiplier/pp_12 [1]),
    .B(\u_multiplier/pp_12 [0]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_12_1/_19_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_12_1/_23_  (.A(\u_multiplier/pp_12 [2]),
    .B(\u_multiplier/pp_12 [3]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_12_1/_20_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_12_1/_24_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_12_1/_19_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_12_1/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_12_1/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE2/ACCI1_pp_12_1/_25_  (.A(\u_multiplier/STAGE2/ACCI1_pp_12_1/_19_ ),
    .B(\u_multiplier/STAGE2/ACCI1_pp_12_1/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_12_1/_16_ ));
 NAND2_X2 \u_multiplier/STAGE2/ACCI1_pp_12_1/_26_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_12_1/_18_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_12_1/_16_ ),
    .ZN(\u_multiplier/s_12 [1]));
 AOI22_X1 \u_multiplier/STAGE2/ACCI1_pp_12_1/_27_  (.A1(\u_multiplier/pp_12 [1]),
    .A2(\u_multiplier/pp_12 [0]),
    .B1(\u_multiplier/pp_12 [2]),
    .B2(\u_multiplier/pp_12 [3]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_12_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_12_1/_28_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_12_1/_15_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_12_1/_17_ ),
    .ZN(\u_multiplier/s_13 [2]));
 NAND3_X1 \u_multiplier/STAGE2/ACCI1_pp_12_2/_21_  (.A1(\u_multiplier/pp_12 [5]),
    .A2(\u_multiplier/pp_12 [4]),
    .A3(\u_multiplier/pp_12 [6]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_12_2/_18_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_12_2/_22_  (.A(\u_multiplier/pp_12 [5]),
    .B(\u_multiplier/pp_12 [4]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_12_2/_19_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_12_2/_23_  (.A(\u_multiplier/pp_12 [6]),
    .B(\u_multiplier/pp_12 [7]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_12_2/_20_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_12_2/_24_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_12_2/_19_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_12_2/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_12_2/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE2/ACCI1_pp_12_2/_25_  (.A(\u_multiplier/STAGE2/ACCI1_pp_12_2/_19_ ),
    .B(\u_multiplier/STAGE2/ACCI1_pp_12_2/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_12_2/_16_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_12_2/_26_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_12_2/_18_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_12_2/_16_ ),
    .ZN(\u_multiplier/s_12 [0]));
 AOI22_X1 \u_multiplier/STAGE2/ACCI1_pp_12_2/_27_  (.A1(\u_multiplier/pp_12 [5]),
    .A2(\u_multiplier/pp_12 [4]),
    .B1(\u_multiplier/pp_12 [6]),
    .B2(\u_multiplier/pp_12 [7]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_12_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_12_2/_28_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_12_2/_15_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_12_2/_17_ ),
    .ZN(\u_multiplier/s_13 [3]));
 NAND3_X1 \u_multiplier/STAGE2/ACCI1_pp_13_1/_21_  (.A1(\u_multiplier/pp_13 [1]),
    .A2(\u_multiplier/pp_13 [0]),
    .A3(\u_multiplier/pp_13 [2]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_13_1/_18_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_13_1/_22_  (.A(\u_multiplier/pp_13 [1]),
    .B(\u_multiplier/pp_13 [0]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_13_1/_19_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_13_1/_23_  (.A(\u_multiplier/pp_13 [2]),
    .B(\u_multiplier/pp_13 [3]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_13_1/_20_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_13_1/_24_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_13_1/_19_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_13_1/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_13_1/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE2/ACCI1_pp_13_1/_25_  (.A(\u_multiplier/STAGE2/ACCI1_pp_13_1/_19_ ),
    .B(\u_multiplier/STAGE2/ACCI1_pp_13_1/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_13_1/_16_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_13_1/_26_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_13_1/_18_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_13_1/_16_ ),
    .ZN(\u_multiplier/s_13 [1]));
 AOI22_X2 \u_multiplier/STAGE2/ACCI1_pp_13_1/_27_  (.A1(\u_multiplier/pp_13 [1]),
    .A2(\u_multiplier/pp_13 [0]),
    .B1(\u_multiplier/pp_13 [2]),
    .B2(\u_multiplier/pp_13 [3]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_13_1/_17_ ));
 NAND2_X2 \u_multiplier/STAGE2/ACCI1_pp_13_1/_28_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_13_1/_15_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_13_1/_17_ ),
    .ZN(\u_multiplier/s_14 [2]));
 NAND3_X1 \u_multiplier/STAGE2/ACCI1_pp_13_2/_21_  (.A1(\u_multiplier/pp_13 [5]),
    .A2(\u_multiplier/pp_13 [4]),
    .A3(\u_multiplier/pp_13 [6]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_13_2/_18_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_13_2/_22_  (.A(\u_multiplier/pp_13 [5]),
    .B(\u_multiplier/pp_13 [4]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_13_2/_19_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_13_2/_23_  (.A(\u_multiplier/pp_13 [6]),
    .B(\u_multiplier/pp_13 [7]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_13_2/_20_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_13_2/_24_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_13_2/_19_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_13_2/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_13_2/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE2/ACCI1_pp_13_2/_25_  (.A(\u_multiplier/STAGE2/ACCI1_pp_13_2/_19_ ),
    .B(\u_multiplier/STAGE2/ACCI1_pp_13_2/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_13_2/_16_ ));
 NAND2_X2 \u_multiplier/STAGE2/ACCI1_pp_13_2/_26_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_13_2/_18_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_13_2/_16_ ),
    .ZN(\u_multiplier/s_13 [0]));
 AOI22_X1 \u_multiplier/STAGE2/ACCI1_pp_13_2/_27_  (.A1(\u_multiplier/pp_13 [5]),
    .A2(\u_multiplier/pp_13 [4]),
    .B1(\u_multiplier/pp_13 [6]),
    .B2(\u_multiplier/pp_13 [7]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_13_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_13_2/_28_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_13_2/_15_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_13_2/_17_ ),
    .ZN(\u_multiplier/s_14 [3]));
 NAND3_X1 \u_multiplier/STAGE2/ACCI1_pp_14_1/_21_  (.A1(\u_multiplier/pp_14 [1]),
    .A2(\u_multiplier/pp_14 [0]),
    .A3(\u_multiplier/pp_14 [2]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_14_1/_18_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_14_1/_22_  (.A(\u_multiplier/pp_14 [1]),
    .B(\u_multiplier/pp_14 [0]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_14_1/_19_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_14_1/_23_  (.A(\u_multiplier/pp_14 [2]),
    .B(\u_multiplier/pp_14 [3]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_14_1/_20_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_14_1/_24_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_14_1/_19_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_14_1/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_14_1/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE2/ACCI1_pp_14_1/_25_  (.A(\u_multiplier/STAGE2/ACCI1_pp_14_1/_19_ ),
    .B(\u_multiplier/STAGE2/ACCI1_pp_14_1/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_14_1/_16_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_14_1/_26_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_14_1/_18_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_14_1/_16_ ),
    .ZN(\u_multiplier/s_14 [1]));
 AOI22_X1 \u_multiplier/STAGE2/ACCI1_pp_14_1/_27_  (.A1(\u_multiplier/pp_14 [1]),
    .A2(\u_multiplier/pp_14 [0]),
    .B1(\u_multiplier/pp_14 [2]),
    .B2(\u_multiplier/pp_14 [3]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_14_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_14_1/_28_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_14_1/_15_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_14_1/_17_ ),
    .ZN(\u_multiplier/s_15 [2]));
 NAND3_X1 \u_multiplier/STAGE2/ACCI1_pp_14_2/_21_  (.A1(\u_multiplier/pp_14 [5]),
    .A2(\u_multiplier/pp_14 [4]),
    .A3(\u_multiplier/pp_14 [6]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_14_2/_18_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_14_2/_22_  (.A(\u_multiplier/pp_14 [5]),
    .B(\u_multiplier/pp_14 [4]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_14_2/_19_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_14_2/_23_  (.A(\u_multiplier/pp_14 [6]),
    .B(\u_multiplier/pp_14 [7]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_14_2/_20_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_14_2/_24_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_14_2/_19_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_14_2/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_14_2/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE2/ACCI1_pp_14_2/_25_  (.A(\u_multiplier/STAGE2/ACCI1_pp_14_2/_19_ ),
    .B(\u_multiplier/STAGE2/ACCI1_pp_14_2/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_14_2/_16_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_14_2/_26_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_14_2/_18_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_14_2/_16_ ),
    .ZN(\u_multiplier/s_14 [0]));
 AOI22_X1 \u_multiplier/STAGE2/ACCI1_pp_14_2/_27_  (.A1(\u_multiplier/pp_14 [5]),
    .A2(\u_multiplier/pp_14 [4]),
    .B1(\u_multiplier/pp_14 [6]),
    .B2(\u_multiplier/pp_14 [7]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_14_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_14_2/_28_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_14_2/_15_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_14_2/_17_ ),
    .ZN(\u_multiplier/s_15 [3]));
 NAND3_X1 \u_multiplier/STAGE2/ACCI1_pp_15_1/_21_  (.A1(\u_multiplier/pp_15 [1]),
    .A2(\u_multiplier/pp_15 [0]),
    .A3(\u_multiplier/pp_15 [2]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_15_1/_18_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_15_1/_22_  (.A(\u_multiplier/pp_15 [1]),
    .B(\u_multiplier/pp_15 [0]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_15_1/_19_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_15_1/_23_  (.A(\u_multiplier/pp_15 [2]),
    .B(\u_multiplier/pp_15 [3]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_15_1/_20_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_15_1/_24_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_15_1/_19_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_15_1/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_15_1/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE2/ACCI1_pp_15_1/_25_  (.A(\u_multiplier/STAGE2/ACCI1_pp_15_1/_19_ ),
    .B(\u_multiplier/STAGE2/ACCI1_pp_15_1/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_15_1/_16_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_15_1/_26_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_15_1/_18_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_15_1/_16_ ),
    .ZN(\u_multiplier/s_15 [1]));
 AOI22_X1 \u_multiplier/STAGE2/ACCI1_pp_15_1/_27_  (.A1(\u_multiplier/pp_15 [1]),
    .A2(\u_multiplier/pp_15 [0]),
    .B1(\u_multiplier/pp_15 [2]),
    .B2(\u_multiplier/pp_15 [3]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_15_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_15_1/_28_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_15_1/_15_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_15_1/_17_ ),
    .ZN(\u_multiplier/s_16 [0]));
 NAND3_X1 \u_multiplier/STAGE2/ACCI1_pp_15_2/_21_  (.A1(\u_multiplier/pp_15 [5]),
    .A2(\u_multiplier/pp_15 [4]),
    .A3(\u_multiplier/pp_15 [6]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_15_2/_18_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_15_2/_22_  (.A(\u_multiplier/pp_15 [5]),
    .B(\u_multiplier/pp_15 [4]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_15_2/_19_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_15_2/_23_  (.A(\u_multiplier/pp_15 [6]),
    .B(\u_multiplier/pp_15 [7]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_15_2/_20_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_15_2/_24_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_15_2/_19_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_15_2/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_15_2/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE2/ACCI1_pp_15_2/_25_  (.A(\u_multiplier/STAGE2/ACCI1_pp_15_2/_19_ ),
    .B(\u_multiplier/STAGE2/ACCI1_pp_15_2/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_15_2/_16_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_15_2/_26_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_15_2/_18_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_15_2/_16_ ),
    .ZN(\u_multiplier/s_15 [0]));
 AOI22_X1 \u_multiplier/STAGE2/ACCI1_pp_15_2/_27_  (.A1(\u_multiplier/pp_15 [5]),
    .A2(\u_multiplier/pp_15 [4]),
    .B1(\u_multiplier/pp_15 [6]),
    .B2(\u_multiplier/pp_15 [7]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_15_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_15_2/_28_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_15_2/_15_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_15_2/_17_ ),
    .ZN(\u_multiplier/s_16 [2]));
 NAND3_X1 \u_multiplier/STAGE2/ACCI1_pp_5/_21_  (.A1(\u_multiplier/pp_5 [1]),
    .A2(\u_multiplier/pp_5 [0]),
    .A3(\u_multiplier/pp_5 [2]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_5/_18_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_5/_22_  (.A(\u_multiplier/pp_5 [1]),
    .B(\u_multiplier/pp_5 [0]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_5/_19_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_5/_23_  (.A(\u_multiplier/pp_5 [2]),
    .B(\u_multiplier/pp_5 [3]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_5/_20_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_5/_24_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_5/_19_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_5/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_5/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE2/ACCI1_pp_5/_25_  (.A(\u_multiplier/STAGE2/ACCI1_pp_5/_19_ ),
    .B(\u_multiplier/STAGE2/ACCI1_pp_5/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_5/_16_ ));
 NAND2_X2 \u_multiplier/STAGE2/ACCI1_pp_5/_26_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_5/_18_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_5/_16_ ),
    .ZN(\u_multiplier/s_5 [0]));
 AOI22_X1 \u_multiplier/STAGE2/ACCI1_pp_5/_27_  (.A1(\u_multiplier/pp_5 [1]),
    .A2(\u_multiplier/pp_5 [0]),
    .B1(\u_multiplier/pp_5 [2]),
    .B2(\u_multiplier/pp_5 [3]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_5/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_5/_28_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_5/_15_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_5/_17_ ),
    .ZN(\u_multiplier/s_6 [3]));
 NAND3_X1 \u_multiplier/STAGE2/ACCI1_pp_6/_21_  (.A1(\u_multiplier/pp_6 [1]),
    .A2(\u_multiplier/pp_6 [0]),
    .A3(\u_multiplier/pp_6 [2]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_6/_18_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_6/_22_  (.A(\u_multiplier/pp_6 [1]),
    .B(\u_multiplier/pp_6 [0]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_6/_19_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_6/_23_  (.A(\u_multiplier/pp_6 [2]),
    .B(\u_multiplier/pp_6 [3]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_6/_20_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_6/_24_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_6/_19_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_6/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_6/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE2/ACCI1_pp_6/_25_  (.A(\u_multiplier/STAGE2/ACCI1_pp_6/_19_ ),
    .B(\u_multiplier/STAGE2/ACCI1_pp_6/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_6/_16_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_6/_26_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_6/_18_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_6/_16_ ),
    .ZN(\u_multiplier/s_6 [1]));
 AOI22_X2 \u_multiplier/STAGE2/ACCI1_pp_6/_27_  (.A1(\u_multiplier/pp_6 [1]),
    .A2(\u_multiplier/pp_6 [0]),
    .B1(\u_multiplier/pp_6 [2]),
    .B2(\u_multiplier/pp_6 [3]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_6/_17_ ));
 NAND2_X2 \u_multiplier/STAGE2/ACCI1_pp_6/_28_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_6/_15_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_6/_17_ ),
    .ZN(\u_multiplier/s_7 [2]));
 NAND3_X1 \u_multiplier/STAGE2/ACCI1_pp_7_1/_21_  (.A1(\u_multiplier/pp_7 [1]),
    .A2(\u_multiplier/pp_7 [0]),
    .A3(\u_multiplier/pp_7 [2]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_7_1/_18_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_7_1/_22_  (.A(\u_multiplier/pp_7 [1]),
    .B(\u_multiplier/pp_7 [0]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_7_1/_19_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_7_1/_23_  (.A(\u_multiplier/pp_7 [2]),
    .B(\u_multiplier/pp_7 [3]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_7_1/_20_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_7_1/_24_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_7_1/_19_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_7_1/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_7_1/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE2/ACCI1_pp_7_1/_25_  (.A(\u_multiplier/STAGE2/ACCI1_pp_7_1/_19_ ),
    .B(\u_multiplier/STAGE2/ACCI1_pp_7_1/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_7_1/_16_ ));
 NAND2_X2 \u_multiplier/STAGE2/ACCI1_pp_7_1/_26_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_7_1/_18_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_7_1/_16_ ),
    .ZN(\u_multiplier/s_7 [1]));
 AOI22_X1 \u_multiplier/STAGE2/ACCI1_pp_7_1/_27_  (.A1(\u_multiplier/pp_7 [1]),
    .A2(\u_multiplier/pp_7 [0]),
    .B1(\u_multiplier/pp_7 [2]),
    .B2(\u_multiplier/pp_7 [3]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_7_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_7_1/_28_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_7_1/_15_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_7_1/_17_ ),
    .ZN(\u_multiplier/s_8 [2]));
 NAND3_X1 \u_multiplier/STAGE2/ACCI1_pp_7_2/_21_  (.A1(\u_multiplier/pp_7 [5]),
    .A2(\u_multiplier/pp_7 [4]),
    .A3(\u_multiplier/pp_7 [6]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_7_2/_18_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_7_2/_22_  (.A(\u_multiplier/pp_7 [5]),
    .B(\u_multiplier/pp_7 [4]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_7_2/_19_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_7_2/_23_  (.A(\u_multiplier/pp_7 [6]),
    .B(\u_multiplier/pp_7 [7]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_7_2/_20_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_7_2/_24_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_7_2/_19_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_7_2/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_7_2/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE2/ACCI1_pp_7_2/_25_  (.A(\u_multiplier/STAGE2/ACCI1_pp_7_2/_19_ ),
    .B(\u_multiplier/STAGE2/ACCI1_pp_7_2/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_7_2/_16_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_7_2/_26_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_7_2/_18_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_7_2/_16_ ),
    .ZN(\u_multiplier/s_7 [0]));
 AOI22_X1 \u_multiplier/STAGE2/ACCI1_pp_7_2/_27_  (.A1(\u_multiplier/pp_7 [5]),
    .A2(\u_multiplier/pp_7 [4]),
    .B1(\u_multiplier/pp_7 [6]),
    .B2(\u_multiplier/pp_7 [7]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_7_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_7_2/_28_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_7_2/_15_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_7_2/_17_ ),
    .ZN(\u_multiplier/s_8 [3]));
 NAND3_X1 \u_multiplier/STAGE2/ACCI1_pp_8_1/_21_  (.A1(\u_multiplier/pp_8 [1]),
    .A2(\u_multiplier/pp_8 [0]),
    .A3(\u_multiplier/pp_8 [2]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_8_1/_18_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_8_1/_22_  (.A(\u_multiplier/pp_8 [1]),
    .B(\u_multiplier/pp_8 [0]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_8_1/_19_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_8_1/_23_  (.A(\u_multiplier/pp_8 [2]),
    .B(\u_multiplier/pp_8 [3]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_8_1/_20_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_8_1/_24_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_8_1/_19_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_8_1/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_8_1/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE2/ACCI1_pp_8_1/_25_  (.A(\u_multiplier/STAGE2/ACCI1_pp_8_1/_19_ ),
    .B(\u_multiplier/STAGE2/ACCI1_pp_8_1/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_8_1/_16_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_8_1/_26_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_8_1/_18_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_8_1/_16_ ),
    .ZN(\u_multiplier/s_8 [1]));
 AOI22_X1 \u_multiplier/STAGE2/ACCI1_pp_8_1/_27_  (.A1(\u_multiplier/pp_8 [1]),
    .A2(\u_multiplier/pp_8 [0]),
    .B1(\u_multiplier/pp_8 [2]),
    .B2(\u_multiplier/pp_8 [3]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_8_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_8_1/_28_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_8_1/_15_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_8_1/_17_ ),
    .ZN(\u_multiplier/s_9 [2]));
 NAND3_X1 \u_multiplier/STAGE2/ACCI1_pp_8_2/_21_  (.A1(\u_multiplier/pp_8 [5]),
    .A2(\u_multiplier/pp_8 [4]),
    .A3(\u_multiplier/pp_8 [6]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_8_2/_18_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_8_2/_22_  (.A(\u_multiplier/pp_8 [5]),
    .B(\u_multiplier/pp_8 [4]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_8_2/_19_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_8_2/_23_  (.A(\u_multiplier/pp_8 [6]),
    .B(\u_multiplier/pp_8 [7]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_8_2/_20_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_8_2/_24_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_8_2/_19_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_8_2/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_8_2/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE2/ACCI1_pp_8_2/_25_  (.A(\u_multiplier/STAGE2/ACCI1_pp_8_2/_19_ ),
    .B(\u_multiplier/STAGE2/ACCI1_pp_8_2/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_8_2/_16_ ));
 NAND2_X2 \u_multiplier/STAGE2/ACCI1_pp_8_2/_26_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_8_2/_18_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_8_2/_16_ ),
    .ZN(\u_multiplier/s_8 [0]));
 AOI22_X1 \u_multiplier/STAGE2/ACCI1_pp_8_2/_27_  (.A1(\u_multiplier/pp_8 [5]),
    .A2(\u_multiplier/pp_8 [4]),
    .B1(\u_multiplier/pp_8 [6]),
    .B2(\u_multiplier/pp_8 [7]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_8_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_8_2/_28_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_8_2/_15_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_8_2/_17_ ),
    .ZN(\u_multiplier/s_9 [3]));
 NAND3_X1 \u_multiplier/STAGE2/ACCI1_pp_9_1/_21_  (.A1(\u_multiplier/pp_9 [1]),
    .A2(\u_multiplier/pp_9 [0]),
    .A3(\u_multiplier/pp_9 [2]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_9_1/_18_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_9_1/_22_  (.A(\u_multiplier/pp_9 [1]),
    .B(\u_multiplier/pp_9 [0]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_9_1/_19_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_9_1/_23_  (.A(\u_multiplier/pp_9 [2]),
    .B(\u_multiplier/pp_9 [3]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_9_1/_20_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_9_1/_24_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_9_1/_19_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_9_1/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_9_1/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE2/ACCI1_pp_9_1/_25_  (.A(\u_multiplier/STAGE2/ACCI1_pp_9_1/_19_ ),
    .B(\u_multiplier/STAGE2/ACCI1_pp_9_1/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_9_1/_16_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_9_1/_26_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_9_1/_18_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_9_1/_16_ ),
    .ZN(\u_multiplier/s_9 [1]));
 AOI22_X1 \u_multiplier/STAGE2/ACCI1_pp_9_1/_27_  (.A1(\u_multiplier/pp_9 [1]),
    .A2(\u_multiplier/pp_9 [0]),
    .B1(\u_multiplier/pp_9 [2]),
    .B2(\u_multiplier/pp_9 [3]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_9_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_9_1/_28_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_9_1/_15_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_9_1/_17_ ),
    .ZN(\u_multiplier/s_10 [2]));
 NAND3_X1 \u_multiplier/STAGE2/ACCI1_pp_9_2/_21_  (.A1(\u_multiplier/pp_9 [5]),
    .A2(\u_multiplier/pp_9 [4]),
    .A3(\u_multiplier/pp_9 [6]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_9_2/_18_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_9_2/_22_  (.A(\u_multiplier/pp_9 [5]),
    .B(\u_multiplier/pp_9 [4]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_9_2/_19_ ));
 XOR2_X2 \u_multiplier/STAGE2/ACCI1_pp_9_2/_23_  (.A(\u_multiplier/pp_9 [6]),
    .B(\u_multiplier/pp_9 [7]),
    .Z(\u_multiplier/STAGE2/ACCI1_pp_9_2/_20_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_9_2/_24_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_9_2/_19_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_9_2/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_9_2/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE2/ACCI1_pp_9_2/_25_  (.A(\u_multiplier/STAGE2/ACCI1_pp_9_2/_19_ ),
    .B(\u_multiplier/STAGE2/ACCI1_pp_9_2/_20_ ),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_9_2/_16_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_9_2/_26_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_9_2/_18_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_9_2/_16_ ),
    .ZN(\u_multiplier/s_9 [0]));
 AOI22_X1 \u_multiplier/STAGE2/ACCI1_pp_9_2/_27_  (.A1(\u_multiplier/pp_9 [5]),
    .A2(\u_multiplier/pp_9 [4]),
    .B1(\u_multiplier/pp_9 [6]),
    .B2(\u_multiplier/pp_9 [7]),
    .ZN(\u_multiplier/STAGE2/ACCI1_pp_9_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/ACCI1_pp_9_2/_28_  (.A1(\u_multiplier/STAGE2/ACCI1_pp_9_2/_15_ ),
    .A2(\u_multiplier/STAGE2/ACCI1_pp_9_2/_17_ ),
    .ZN(\u_multiplier/s_10 [3]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_16_1/_18_  (.A(net60),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_16_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_16_1/_19_  (.A1(\u_multiplier/pp_16 [1]),
    .A2(\u_multiplier/pp_16 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_16_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_16_1/_20_  (.A(\u_multiplier/pp_16 [1]),
    .B(\u_multiplier/pp_16 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_16_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_16_1/_21_  (.A1(\u_multiplier/pp_16 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_16_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_16_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_16_1/_22_  (.A(\u_multiplier/pp_16 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_16_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_16_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_16_1/_23_  (.A1(\u_multiplier/pp_16 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_16_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_16_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_16_1/_24_  (.A(\u_multiplier/pp_16 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_16_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_16_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_16_1/_25_  (.A(net61),
    .B(\u_multiplier/STAGE2/E_4_2_pp_16_1/_16_ ),
    .ZN(\u_multiplier/s_16 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_16_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_16_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_16_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_16_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_16_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_16_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_16_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_16_1/_17_ ),
    .ZN(\u_multiplier/s_17 [0]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_16_2/_18_  (.A(net62),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_16_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_16_2/_19_  (.A1(\u_multiplier/pp_16 [5]),
    .A2(\u_multiplier/pp_16 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_16_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_16_2/_20_  (.A(\u_multiplier/pp_16 [5]),
    .B(\u_multiplier/pp_16 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_16_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_16_2/_21_  (.A1(\u_multiplier/pp_16 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_16_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_16_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_16_2/_22_  (.A(\u_multiplier/pp_16 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_16_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_16_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_16_2/_23_  (.A1(\u_multiplier/pp_16 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_16_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_16_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_16_2/_24_  (.A(\u_multiplier/pp_16 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_16_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_16_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_16_2/_25_  (.A(net63),
    .B(\u_multiplier/STAGE2/E_4_2_pp_16_2/_16_ ),
    .ZN(\u_multiplier/s_16 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_16_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_16_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_16_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_16_c4 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_16_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_16_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_16_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_16_2/_17_ ),
    .ZN(\u_multiplier/s_17 [2]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_17_1/_18_  (.A(\u_multiplier/STAGE2/pp_16_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_17_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_17_1/_19_  (.A1(\u_multiplier/pp_17 [1]),
    .A2(\u_multiplier/pp_17 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_17_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_17_1/_20_  (.A(\u_multiplier/pp_17 [1]),
    .B(\u_multiplier/pp_17 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_17_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_17_1/_21_  (.A1(\u_multiplier/pp_17 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_17_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_17_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_17_1/_22_  (.A(\u_multiplier/pp_17 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_17_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_17_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_17_1/_23_  (.A1(\u_multiplier/pp_17 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_17_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_17_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_17_1/_24_  (.A(\u_multiplier/pp_17 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_17_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_17_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_17_1/_25_  (.A(\u_multiplier/STAGE2/pp_16_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_17_1/_16_ ),
    .ZN(\u_multiplier/s_17 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_17_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_17_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_17_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_17_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_17_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_17_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_17_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_17_1/_17_ ),
    .ZN(\u_multiplier/s_18 [0]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_17_2/_18_  (.A(\u_multiplier/STAGE2/pp_16_c4 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_17_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_17_2/_19_  (.A1(\u_multiplier/pp_17 [5]),
    .A2(\u_multiplier/pp_17 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_17_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_17_2/_20_  (.A(\u_multiplier/pp_17 [5]),
    .B(\u_multiplier/pp_17 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_17_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_17_2/_21_  (.A1(\u_multiplier/pp_17 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_17_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_17_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_17_2/_22_  (.A(\u_multiplier/pp_17 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_17_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_17_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_17_2/_23_  (.A1(\u_multiplier/pp_17 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_17_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_17_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_17_2/_24_  (.A(\u_multiplier/pp_17 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_17_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_17_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_17_2/_25_  (.A(\u_multiplier/STAGE2/pp_16_c4 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_17_2/_16_ ),
    .ZN(\u_multiplier/s_17 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_17_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_17_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_17_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_17_c4 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_17_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_17_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_17_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_17_2/_17_ ),
    .ZN(\u_multiplier/s_18 [2]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_18_1/_18_  (.A(\u_multiplier/STAGE2/pp_17_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_18_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_18_1/_19_  (.A1(\u_multiplier/pp_18 [1]),
    .A2(\u_multiplier/pp_18 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_18_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_18_1/_20_  (.A(\u_multiplier/pp_18 [1]),
    .B(\u_multiplier/pp_18 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_18_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_18_1/_21_  (.A1(\u_multiplier/pp_18 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_18_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_18_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_18_1/_22_  (.A(\u_multiplier/pp_18 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_18_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_18_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_18_1/_23_  (.A1(\u_multiplier/pp_18 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_18_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_18_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_18_1/_24_  (.A(\u_multiplier/pp_18 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_18_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_18_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_18_1/_25_  (.A(\u_multiplier/STAGE2/pp_17_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_18_1/_16_ ),
    .ZN(\u_multiplier/s_18 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_18_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_18_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_18_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_18_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_18_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_18_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_18_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_18_1/_17_ ),
    .ZN(\u_multiplier/s_19 [0]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_18_2/_18_  (.A(\u_multiplier/STAGE2/pp_17_c4 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_18_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_18_2/_19_  (.A1(\u_multiplier/pp_18 [5]),
    .A2(\u_multiplier/pp_18 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_18_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_18_2/_20_  (.A(\u_multiplier/pp_18 [5]),
    .B(\u_multiplier/pp_18 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_18_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_18_2/_21_  (.A1(\u_multiplier/pp_18 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_18_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_18_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_18_2/_22_  (.A(\u_multiplier/pp_18 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_18_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_18_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_18_2/_23_  (.A1(\u_multiplier/pp_18 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_18_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_18_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_18_2/_24_  (.A(\u_multiplier/pp_18 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_18_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_18_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_18_2/_25_  (.A(\u_multiplier/STAGE2/pp_17_c4 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_18_2/_16_ ),
    .ZN(\u_multiplier/s_18 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_18_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_18_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_18_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_18_c4 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_18_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_18_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_18_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_18_2/_17_ ),
    .ZN(\u_multiplier/s_19 [2]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_19_1/_18_  (.A(\u_multiplier/STAGE2/pp_18_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_19_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_19_1/_19_  (.A1(\u_multiplier/pp_19 [1]),
    .A2(\u_multiplier/pp_19 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_19_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_19_1/_20_  (.A(\u_multiplier/pp_19 [1]),
    .B(\u_multiplier/pp_19 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_19_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_19_1/_21_  (.A1(\u_multiplier/pp_19 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_19_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_19_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_19_1/_22_  (.A(\u_multiplier/pp_19 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_19_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_19_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_19_1/_23_  (.A1(\u_multiplier/pp_19 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_19_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_19_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_19_1/_24_  (.A(\u_multiplier/pp_19 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_19_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_19_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_19_1/_25_  (.A(\u_multiplier/STAGE2/pp_18_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_19_1/_16_ ),
    .ZN(\u_multiplier/s_19 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_19_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_19_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_19_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_19_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_19_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_19_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_19_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_19_1/_17_ ),
    .ZN(\u_multiplier/s_20 [0]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_19_2/_18_  (.A(\u_multiplier/STAGE2/pp_18_c4 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_19_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_19_2/_19_  (.A1(\u_multiplier/pp_19 [5]),
    .A2(\u_multiplier/pp_19 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_19_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_19_2/_20_  (.A(\u_multiplier/pp_19 [5]),
    .B(\u_multiplier/pp_19 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_19_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_19_2/_21_  (.A1(\u_multiplier/pp_19 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_19_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_19_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_19_2/_22_  (.A(\u_multiplier/pp_19 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_19_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_19_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_19_2/_23_  (.A1(\u_multiplier/pp_19 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_19_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_19_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_19_2/_24_  (.A(\u_multiplier/pp_19 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_19_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_19_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_19_2/_25_  (.A(\u_multiplier/STAGE2/pp_18_c4 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_19_2/_16_ ),
    .ZN(\u_multiplier/s_19 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_19_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_19_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_19_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_19_c4 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_19_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_19_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_19_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_19_2/_17_ ),
    .ZN(\u_multiplier/s_20 [2]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_20_1/_18_  (.A(\u_multiplier/STAGE2/pp_19_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_20_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_20_1/_19_  (.A1(\u_multiplier/pp_20 [1]),
    .A2(\u_multiplier/pp_20 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_20_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_20_1/_20_  (.A(\u_multiplier/pp_20 [1]),
    .B(\u_multiplier/pp_20 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_20_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_20_1/_21_  (.A1(\u_multiplier/pp_20 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_20_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_20_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_20_1/_22_  (.A(\u_multiplier/pp_20 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_20_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_20_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_20_1/_23_  (.A1(\u_multiplier/pp_20 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_20_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_20_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_20_1/_24_  (.A(\u_multiplier/pp_20 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_20_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_20_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_20_1/_25_  (.A(\u_multiplier/STAGE2/pp_19_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_20_1/_16_ ),
    .ZN(\u_multiplier/s_20 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_20_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_20_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_20_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_20_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_20_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_20_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_20_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_20_1/_17_ ),
    .ZN(\u_multiplier/s_21 [0]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_20_2/_18_  (.A(\u_multiplier/STAGE2/pp_19_c4 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_20_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_20_2/_19_  (.A1(\u_multiplier/pp_20 [5]),
    .A2(\u_multiplier/pp_20 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_20_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_20_2/_20_  (.A(\u_multiplier/pp_20 [5]),
    .B(\u_multiplier/pp_20 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_20_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_20_2/_21_  (.A1(\u_multiplier/pp_20 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_20_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_20_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_20_2/_22_  (.A(\u_multiplier/pp_20 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_20_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_20_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_20_2/_23_  (.A1(\u_multiplier/pp_20 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_20_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_20_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_20_2/_24_  (.A(\u_multiplier/pp_20 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_20_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_20_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_20_2/_25_  (.A(\u_multiplier/STAGE2/pp_19_c4 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_20_2/_16_ ),
    .ZN(\u_multiplier/s_20 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_20_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_20_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_20_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_20_c4 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_20_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_20_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_20_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_20_2/_17_ ),
    .ZN(\u_multiplier/s_21 [2]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_21_1/_18_  (.A(\u_multiplier/STAGE2/pp_20_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_21_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_21_1/_19_  (.A1(\u_multiplier/pp_21 [1]),
    .A2(\u_multiplier/pp_21 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_21_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_21_1/_20_  (.A(\u_multiplier/pp_21 [1]),
    .B(\u_multiplier/pp_21 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_21_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_21_1/_21_  (.A1(\u_multiplier/pp_21 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_21_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_21_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_21_1/_22_  (.A(\u_multiplier/pp_21 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_21_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_21_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_21_1/_23_  (.A1(\u_multiplier/pp_21 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_21_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_21_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_21_1/_24_  (.A(\u_multiplier/pp_21 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_21_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_21_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_21_1/_25_  (.A(\u_multiplier/STAGE2/pp_20_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_21_1/_16_ ),
    .ZN(\u_multiplier/s_21 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_21_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_21_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_21_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_21_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_21_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_21_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_21_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_21_1/_17_ ),
    .ZN(\u_multiplier/s_22 [0]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_21_2/_18_  (.A(\u_multiplier/STAGE2/pp_20_c4 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_21_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_21_2/_19_  (.A1(\u_multiplier/pp_21 [5]),
    .A2(\u_multiplier/pp_21 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_21_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_21_2/_20_  (.A(\u_multiplier/pp_21 [5]),
    .B(\u_multiplier/pp_21 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_21_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_21_2/_21_  (.A1(\u_multiplier/pp_21 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_21_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_21_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_21_2/_22_  (.A(\u_multiplier/pp_21 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_21_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_21_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_21_2/_23_  (.A1(\u_multiplier/pp_21 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_21_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_21_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_21_2/_24_  (.A(\u_multiplier/pp_21 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_21_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_21_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_21_2/_25_  (.A(\u_multiplier/STAGE2/pp_20_c4 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_21_2/_16_ ),
    .ZN(\u_multiplier/s_21 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_21_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_21_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_21_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_21_c4 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_21_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_21_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_21_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_21_2/_17_ ),
    .ZN(\u_multiplier/s_22 [2]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_22_1/_18_  (.A(\u_multiplier/STAGE2/pp_21_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_22_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_22_1/_19_  (.A1(\u_multiplier/pp_22 [1]),
    .A2(\u_multiplier/pp_22 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_22_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_22_1/_20_  (.A(\u_multiplier/pp_22 [1]),
    .B(\u_multiplier/pp_22 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_22_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_22_1/_21_  (.A1(\u_multiplier/pp_22 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_22_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_22_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_22_1/_22_  (.A(\u_multiplier/pp_22 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_22_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_22_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_22_1/_23_  (.A1(\u_multiplier/pp_22 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_22_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_22_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_22_1/_24_  (.A(\u_multiplier/pp_22 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_22_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_22_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_22_1/_25_  (.A(\u_multiplier/STAGE2/pp_21_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_22_1/_16_ ),
    .ZN(\u_multiplier/s_22 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_22_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_22_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_22_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_22_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_22_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_22_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_22_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_22_1/_17_ ),
    .ZN(\u_multiplier/s_23 [0]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_22_2/_18_  (.A(\u_multiplier/STAGE2/pp_21_c4 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_22_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_22_2/_19_  (.A1(\u_multiplier/pp_22 [5]),
    .A2(\u_multiplier/pp_22 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_22_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_22_2/_20_  (.A(\u_multiplier/pp_22 [5]),
    .B(\u_multiplier/pp_22 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_22_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_22_2/_21_  (.A1(\u_multiplier/pp_22 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_22_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_22_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_22_2/_22_  (.A(\u_multiplier/pp_22 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_22_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_22_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_22_2/_23_  (.A1(\u_multiplier/pp_22 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_22_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_22_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_22_2/_24_  (.A(\u_multiplier/pp_22 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_22_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_22_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_22_2/_25_  (.A(\u_multiplier/STAGE2/pp_21_c4 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_22_2/_16_ ),
    .ZN(\u_multiplier/s_22 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_22_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_22_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_22_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_22_c4 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_22_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_22_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_22_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_22_2/_17_ ),
    .ZN(\u_multiplier/s_23 [2]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_23_1/_18_  (.A(\u_multiplier/STAGE2/pp_22_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_23_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_23_1/_19_  (.A1(\u_multiplier/pp_23 [1]),
    .A2(\u_multiplier/pp_23 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_23_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_23_1/_20_  (.A(\u_multiplier/pp_23 [1]),
    .B(\u_multiplier/pp_23 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_23_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_23_1/_21_  (.A1(\u_multiplier/pp_23 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_23_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_23_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_23_1/_22_  (.A(\u_multiplier/pp_23 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_23_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_23_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_23_1/_23_  (.A1(\u_multiplier/pp_23 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_23_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_23_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_23_1/_24_  (.A(\u_multiplier/pp_23 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_23_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_23_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_23_1/_25_  (.A(\u_multiplier/STAGE2/pp_22_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_23_1/_16_ ),
    .ZN(\u_multiplier/s_23 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_23_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_23_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_23_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_23_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_23_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_23_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_23_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_23_1/_17_ ),
    .ZN(\u_multiplier/s_24 [0]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_23_2/_18_  (.A(\u_multiplier/STAGE2/pp_22_c4 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_23_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_23_2/_19_  (.A1(\u_multiplier/pp_23 [5]),
    .A2(\u_multiplier/pp_23 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_23_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_23_2/_20_  (.A(\u_multiplier/pp_23 [5]),
    .B(\u_multiplier/pp_23 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_23_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_23_2/_21_  (.A1(\u_multiplier/pp_23 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_23_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_23_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_23_2/_22_  (.A(\u_multiplier/pp_23 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_23_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_23_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_23_2/_23_  (.A1(\u_multiplier/pp_23 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_23_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_23_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_23_2/_24_  (.A(\u_multiplier/pp_23 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_23_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_23_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_23_2/_25_  (.A(\u_multiplier/STAGE2/pp_22_c4 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_23_2/_16_ ),
    .ZN(\u_multiplier/s_23 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_23_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_23_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_23_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_23_c4 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_23_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_23_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_23_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_23_2/_17_ ),
    .ZN(\u_multiplier/s_24 [2]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_24_1/_18_  (.A(\u_multiplier/STAGE2/pp_23_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_24_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_24_1/_19_  (.A1(\u_multiplier/pp_24 [1]),
    .A2(\u_multiplier/pp_24 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_24_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_24_1/_20_  (.A(\u_multiplier/pp_24 [1]),
    .B(\u_multiplier/pp_24 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_24_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_24_1/_21_  (.A1(\u_multiplier/pp_24 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_24_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_24_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_24_1/_22_  (.A(\u_multiplier/pp_24 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_24_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_24_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_24_1/_23_  (.A1(\u_multiplier/pp_24 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_24_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_24_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_24_1/_24_  (.A(\u_multiplier/pp_24 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_24_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_24_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_24_1/_25_  (.A(\u_multiplier/STAGE2/pp_23_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_24_1/_16_ ),
    .ZN(\u_multiplier/s_24 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_24_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_24_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_24_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_24_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_24_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_24_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_24_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_24_1/_17_ ),
    .ZN(\u_multiplier/s_25 [0]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_24_2/_18_  (.A(\u_multiplier/STAGE2/pp_23_c4 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_24_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_24_2/_19_  (.A1(\u_multiplier/pp_24 [5]),
    .A2(\u_multiplier/pp_24 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_24_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_24_2/_20_  (.A(\u_multiplier/pp_24 [5]),
    .B(\u_multiplier/pp_24 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_24_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_24_2/_21_  (.A1(\u_multiplier/pp_24 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_24_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_24_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_24_2/_22_  (.A(\u_multiplier/pp_24 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_24_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_24_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_24_2/_23_  (.A1(\u_multiplier/pp_24 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_24_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_24_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_24_2/_24_  (.A(\u_multiplier/pp_24 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_24_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_24_2/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE2/E_4_2_pp_24_2/_25_  (.A(\u_multiplier/STAGE2/pp_23_c4 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_24_2/_16_ ),
    .ZN(\u_multiplier/s_24 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_24_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_24_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_24_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_24_c4 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_24_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_24_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_24_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_24_2/_17_ ),
    .ZN(\u_multiplier/s_25 [2]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_25_1/_18_  (.A(\u_multiplier/STAGE2/pp_24_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_25_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_25_1/_19_  (.A1(\u_multiplier/pp_25 [1]),
    .A2(\u_multiplier/pp_25 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_25_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_25_1/_20_  (.A(\u_multiplier/pp_25 [1]),
    .B(\u_multiplier/pp_25 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_25_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_25_1/_21_  (.A1(\u_multiplier/pp_25 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_25_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_25_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_25_1/_22_  (.A(\u_multiplier/pp_25 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_25_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_25_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_25_1/_23_  (.A1(\u_multiplier/pp_25 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_25_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_25_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_25_1/_24_  (.A(\u_multiplier/pp_25 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_25_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_25_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_25_1/_25_  (.A(\u_multiplier/STAGE2/pp_24_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_25_1/_16_ ),
    .ZN(\u_multiplier/s_25 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_25_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_25_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_25_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_25_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_25_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_25_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_25_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_25_1/_17_ ),
    .ZN(\u_multiplier/s_26 [0]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_26_1/_18_  (.A(\u_multiplier/STAGE2/pp_25_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_26_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_26_1/_19_  (.A1(\u_multiplier/pp_26 [1]),
    .A2(\u_multiplier/pp_26 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_26_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_26_1/_20_  (.A(\u_multiplier/pp_26 [1]),
    .B(\u_multiplier/pp_26 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_26_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_26_1/_21_  (.A1(\u_multiplier/pp_26 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_26_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_26_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_26_1/_22_  (.A(\u_multiplier/pp_26 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_26_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_26_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_26_1/_23_  (.A1(\u_multiplier/pp_26 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_26_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_26_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_26_1/_24_  (.A(\u_multiplier/pp_26 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_26_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_26_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_26_1/_25_  (.A(\u_multiplier/STAGE2/pp_25_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_26_1/_16_ ),
    .ZN(\u_multiplier/s_26 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_26_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_26_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_26_1/_13_ ),
    .ZN(\u_multiplier/s_27 [2]));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_26_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_26_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_26_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_26_1/_17_ ),
    .ZN(\u_multiplier/s_27 [0]));
 INV_X1 \u_multiplier/STAGE2/Full_adder_pp_25/_12_  (.A(\u_multiplier/STAGE2/pp_24_c4 ),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp_25/_08_ ));
 NAND3_X1 \u_multiplier/STAGE2/Full_adder_pp_25/_13_  (.A1(\u_multiplier/pp_25 [5]),
    .A2(\u_multiplier/pp_25 [4]),
    .A3(\u_multiplier/STAGE2/pp_24_c4 ),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp_25/_09_ ));
 NOR2_X2 \u_multiplier/STAGE2/Full_adder_pp_25/_14_  (.A1(\u_multiplier/pp_25 [5]),
    .A2(\u_multiplier/pp_25 [4]),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp_25/_10_ ));
 AOI21_X1 \u_multiplier/STAGE2/Full_adder_pp_25/_15_  (.A(\u_multiplier/STAGE2/pp_24_c4 ),
    .B1(\u_multiplier/pp_25 [4]),
    .B2(\u_multiplier/pp_25 [5]),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp_25/_11_ ));
 NOR2_X2 \u_multiplier/STAGE2/Full_adder_pp_25/_16_  (.A1(\u_multiplier/STAGE2/Full_adder_pp_25/_10_ ),
    .A2(\u_multiplier/STAGE2/Full_adder_pp_25/_11_ ),
    .ZN(\u_multiplier/s_26 [2]));
 AOI22_X2 \u_multiplier/STAGE2/Full_adder_pp_25/_17_  (.A1(\u_multiplier/STAGE2/Full_adder_pp_25/_08_ ),
    .A2(\u_multiplier/STAGE2/Full_adder_pp_25/_10_ ),
    .B1(\u_multiplier/s_26 [2]),
    .B2(\u_multiplier/STAGE2/Full_adder_pp_25/_09_ ),
    .ZN(\u_multiplier/s_25 [3]));
 INV_X1 \u_multiplier/STAGE2/Full_adder_pp_27/_12_  (.A(\u_multiplier/pp_27 [2]),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp_27/_08_ ));
 NAND3_X2 \u_multiplier/STAGE2/Full_adder_pp_27/_13_  (.A1(\u_multiplier/pp_27 [1]),
    .A2(\u_multiplier/pp_27 [0]),
    .A3(\u_multiplier/pp_27 [2]),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp_27/_09_ ));
 NOR2_X2 \u_multiplier/STAGE2/Full_adder_pp_27/_14_  (.A1(\u_multiplier/pp_27 [1]),
    .A2(\u_multiplier/pp_27 [0]),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp_27/_10_ ));
 AOI21_X1 \u_multiplier/STAGE2/Full_adder_pp_27/_15_  (.A(\u_multiplier/pp_27 [2]),
    .B1(\u_multiplier/pp_27 [0]),
    .B2(\u_multiplier/pp_27 [1]),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp_27/_11_ ));
 NOR2_X2 \u_multiplier/STAGE2/Full_adder_pp_27/_16_  (.A1(\u_multiplier/STAGE2/Full_adder_pp_27/_10_ ),
    .A2(\u_multiplier/STAGE2/Full_adder_pp_27/_11_ ),
    .ZN(\u_multiplier/s_28 [0]));
 AOI22_X4 \u_multiplier/STAGE2/Full_adder_pp_27/_17_  (.A1(\u_multiplier/STAGE2/Full_adder_pp_27/_08_ ),
    .A2(\u_multiplier/STAGE2/Full_adder_pp_27/_10_ ),
    .B1(\u_multiplier/s_28 [0]),
    .B2(\u_multiplier/STAGE2/Full_adder_pp_27/_09_ ),
    .ZN(\u_multiplier/s_27 [3]));
 AND2_X1 \u_multiplier/STAGE2/Half_adder_pp_4/_4_  (.A1(\u_multiplier/pp_4 [1]),
    .A2(\u_multiplier/pp_4 [0]),
    .ZN(\u_multiplier/s_5 [3]));
 XOR2_X2 \u_multiplier/STAGE2/Half_adder_pp_4/_5_  (.A(\u_multiplier/pp_4 [1]),
    .B(\u_multiplier/pp_4 [0]),
    .Z(\u_multiplier/s_4 [0]));
 AND2_X1 \u_multiplier/STAGE2/Half_adder_pp_6/_4_  (.A1(\u_multiplier/pp_6 [5]),
    .A2(\u_multiplier/pp_6 [4]),
    .ZN(\u_multiplier/s_7 [3]));
 XOR2_X2 \u_multiplier/STAGE2/Half_adder_pp_6/_5_  (.A(\u_multiplier/pp_6 [5]),
    .B(\u_multiplier/pp_6 [4]),
    .Z(\u_multiplier/s_6 [0]));
 NAND3_X1 \u_multiplier/STAGE3/ACCI1_pp_10_1/_21_  (.A1(\u_multiplier/s_10 [1]),
    .A2(\u_multiplier/s_10 [0]),
    .A3(\u_multiplier/s_10 [2]),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_10_1/_18_ ));
 XOR2_X2 \u_multiplier/STAGE3/ACCI1_pp_10_1/_22_  (.A(\u_multiplier/s_10 [1]),
    .B(\u_multiplier/s_10 [0]),
    .Z(\u_multiplier/STAGE3/ACCI1_pp_10_1/_19_ ));
 XOR2_X2 \u_multiplier/STAGE3/ACCI1_pp_10_1/_23_  (.A(\u_multiplier/s_10 [2]),
    .B(\u_multiplier/s_10 [3]),
    .Z(\u_multiplier/STAGE3/ACCI1_pp_10_1/_20_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_10_1/_24_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_10_1/_19_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_10_1/_20_ ),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_10_1/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE3/ACCI1_pp_10_1/_25_  (.A(\u_multiplier/STAGE3/ACCI1_pp_10_1/_19_ ),
    .B(\u_multiplier/STAGE3/ACCI1_pp_10_1/_20_ ),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_10_1/_16_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_10_1/_26_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_10_1/_18_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_10_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_10_s ));
 AOI22_X1 \u_multiplier/STAGE3/ACCI1_pp_10_1/_27_  (.A1(\u_multiplier/s_10 [1]),
    .A2(\u_multiplier/s_10 [0]),
    .B1(\u_multiplier/s_10 [2]),
    .B2(\u_multiplier/s_10 [3]),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_10_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_10_1/_28_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_10_1/_15_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_10_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_10_c ));
 NAND3_X1 \u_multiplier/STAGE3/ACCI1_pp_11_1/_21_  (.A1(\u_multiplier/s_11 [1]),
    .A2(\u_multiplier/s_11 [0]),
    .A3(\u_multiplier/s_11 [2]),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_11_1/_18_ ));
 XOR2_X2 \u_multiplier/STAGE3/ACCI1_pp_11_1/_22_  (.A(\u_multiplier/s_11 [1]),
    .B(\u_multiplier/s_11 [0]),
    .Z(\u_multiplier/STAGE3/ACCI1_pp_11_1/_19_ ));
 XOR2_X2 \u_multiplier/STAGE3/ACCI1_pp_11_1/_23_  (.A(\u_multiplier/s_11 [2]),
    .B(\u_multiplier/s_11 [3]),
    .Z(\u_multiplier/STAGE3/ACCI1_pp_11_1/_20_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_11_1/_24_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_11_1/_19_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_11_1/_20_ ),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_11_1/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE3/ACCI1_pp_11_1/_25_  (.A(\u_multiplier/STAGE3/ACCI1_pp_11_1/_19_ ),
    .B(\u_multiplier/STAGE3/ACCI1_pp_11_1/_20_ ),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_11_1/_16_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_11_1/_26_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_11_1/_18_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_11_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_11_s ));
 AOI22_X1 \u_multiplier/STAGE3/ACCI1_pp_11_1/_27_  (.A1(\u_multiplier/s_11 [1]),
    .A2(\u_multiplier/s_11 [0]),
    .B1(\u_multiplier/s_11 [2]),
    .B2(\u_multiplier/s_11 [3]),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_11_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_11_1/_28_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_11_1/_15_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_11_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_11_c ));
 NAND3_X1 \u_multiplier/STAGE3/ACCI1_pp_12_1/_21_  (.A1(\u_multiplier/s_12 [1]),
    .A2(\u_multiplier/s_12 [0]),
    .A3(\u_multiplier/s_12 [2]),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_12_1/_18_ ));
 XOR2_X2 \u_multiplier/STAGE3/ACCI1_pp_12_1/_22_  (.A(\u_multiplier/s_12 [1]),
    .B(\u_multiplier/s_12 [0]),
    .Z(\u_multiplier/STAGE3/ACCI1_pp_12_1/_19_ ));
 XOR2_X2 \u_multiplier/STAGE3/ACCI1_pp_12_1/_23_  (.A(\u_multiplier/s_12 [2]),
    .B(\u_multiplier/s_12 [3]),
    .Z(\u_multiplier/STAGE3/ACCI1_pp_12_1/_20_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_12_1/_24_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_12_1/_19_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_12_1/_20_ ),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_12_1/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE3/ACCI1_pp_12_1/_25_  (.A(\u_multiplier/STAGE3/ACCI1_pp_12_1/_19_ ),
    .B(\u_multiplier/STAGE3/ACCI1_pp_12_1/_20_ ),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_12_1/_16_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_12_1/_26_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_12_1/_18_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_12_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_12_s ));
 AOI22_X1 \u_multiplier/STAGE3/ACCI1_pp_12_1/_27_  (.A1(\u_multiplier/s_12 [1]),
    .A2(\u_multiplier/s_12 [0]),
    .B1(\u_multiplier/s_12 [2]),
    .B2(\u_multiplier/s_12 [3]),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_12_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_12_1/_28_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_12_1/_15_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_12_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_12_c ));
 NAND3_X1 \u_multiplier/STAGE3/ACCI1_pp_13_1/_21_  (.A1(\u_multiplier/s_13 [1]),
    .A2(\u_multiplier/s_13 [0]),
    .A3(\u_multiplier/s_13 [2]),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_13_1/_18_ ));
 XOR2_X2 \u_multiplier/STAGE3/ACCI1_pp_13_1/_22_  (.A(\u_multiplier/s_13 [1]),
    .B(\u_multiplier/s_13 [0]),
    .Z(\u_multiplier/STAGE3/ACCI1_pp_13_1/_19_ ));
 XOR2_X2 \u_multiplier/STAGE3/ACCI1_pp_13_1/_23_  (.A(\u_multiplier/s_13 [2]),
    .B(\u_multiplier/s_13 [3]),
    .Z(\u_multiplier/STAGE3/ACCI1_pp_13_1/_20_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_13_1/_24_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_13_1/_19_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_13_1/_20_ ),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_13_1/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE3/ACCI1_pp_13_1/_25_  (.A(\u_multiplier/STAGE3/ACCI1_pp_13_1/_19_ ),
    .B(\u_multiplier/STAGE3/ACCI1_pp_13_1/_20_ ),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_13_1/_16_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_13_1/_26_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_13_1/_18_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_13_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_13_s ));
 AOI22_X1 \u_multiplier/STAGE3/ACCI1_pp_13_1/_27_  (.A1(\u_multiplier/s_13 [1]),
    .A2(\u_multiplier/s_13 [0]),
    .B1(\u_multiplier/s_13 [2]),
    .B2(\u_multiplier/s_13 [3]),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_13_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_13_1/_28_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_13_1/_15_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_13_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_13_c ));
 NAND3_X1 \u_multiplier/STAGE3/ACCI1_pp_14_1/_21_  (.A1(\u_multiplier/s_14 [1]),
    .A2(\u_multiplier/s_14 [0]),
    .A3(\u_multiplier/s_14 [2]),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_14_1/_18_ ));
 XOR2_X2 \u_multiplier/STAGE3/ACCI1_pp_14_1/_22_  (.A(\u_multiplier/s_14 [1]),
    .B(\u_multiplier/s_14 [0]),
    .Z(\u_multiplier/STAGE3/ACCI1_pp_14_1/_19_ ));
 XOR2_X2 \u_multiplier/STAGE3/ACCI1_pp_14_1/_23_  (.A(\u_multiplier/s_14 [2]),
    .B(\u_multiplier/s_14 [3]),
    .Z(\u_multiplier/STAGE3/ACCI1_pp_14_1/_20_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_14_1/_24_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_14_1/_19_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_14_1/_20_ ),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_14_1/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE3/ACCI1_pp_14_1/_25_  (.A(\u_multiplier/STAGE3/ACCI1_pp_14_1/_19_ ),
    .B(\u_multiplier/STAGE3/ACCI1_pp_14_1/_20_ ),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_14_1/_16_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_14_1/_26_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_14_1/_18_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_14_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_14_s ));
 AOI22_X1 \u_multiplier/STAGE3/ACCI1_pp_14_1/_27_  (.A1(\u_multiplier/s_14 [1]),
    .A2(\u_multiplier/s_14 [0]),
    .B1(\u_multiplier/s_14 [2]),
    .B2(\u_multiplier/s_14 [3]),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_14_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_14_1/_28_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_14_1/_15_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_14_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_14_c ));
 NAND3_X1 \u_multiplier/STAGE3/ACCI1_pp_15_1/_21_  (.A1(\u_multiplier/s_15 [1]),
    .A2(\u_multiplier/s_15 [0]),
    .A3(\u_multiplier/s_15 [2]),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_15_1/_18_ ));
 XOR2_X2 \u_multiplier/STAGE3/ACCI1_pp_15_1/_22_  (.A(\u_multiplier/s_15 [1]),
    .B(\u_multiplier/s_15 [0]),
    .Z(\u_multiplier/STAGE3/ACCI1_pp_15_1/_19_ ));
 XOR2_X2 \u_multiplier/STAGE3/ACCI1_pp_15_1/_23_  (.A(\u_multiplier/s_15 [2]),
    .B(\u_multiplier/s_15 [3]),
    .Z(\u_multiplier/STAGE3/ACCI1_pp_15_1/_20_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_15_1/_24_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_15_1/_19_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_15_1/_20_ ),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_15_1/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE3/ACCI1_pp_15_1/_25_  (.A(\u_multiplier/STAGE3/ACCI1_pp_15_1/_19_ ),
    .B(\u_multiplier/STAGE3/ACCI1_pp_15_1/_20_ ),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_15_1/_16_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_15_1/_26_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_15_1/_18_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_15_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_15_s ));
 AOI22_X1 \u_multiplier/STAGE3/ACCI1_pp_15_1/_27_  (.A1(\u_multiplier/s_15 [1]),
    .A2(\u_multiplier/s_15 [0]),
    .B1(\u_multiplier/s_15 [2]),
    .B2(\u_multiplier/s_15 [3]),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_15_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_15_1/_28_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_15_1/_15_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_15_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_15_c ));
 NAND3_X1 \u_multiplier/STAGE3/ACCI1_pp_3/_21_  (.A1(\u_multiplier/s_3 [1]),
    .A2(\u_multiplier/s_3 [0]),
    .A3(\u_multiplier/s_3 [2]),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_3/_18_ ));
 XOR2_X2 \u_multiplier/STAGE3/ACCI1_pp_3/_22_  (.A(\u_multiplier/s_3 [1]),
    .B(\u_multiplier/s_3 [0]),
    .Z(\u_multiplier/STAGE3/ACCI1_pp_3/_19_ ));
 XOR2_X2 \u_multiplier/STAGE3/ACCI1_pp_3/_23_  (.A(\u_multiplier/s_3 [2]),
    .B(\u_multiplier/s_3 [3]),
    .Z(\u_multiplier/STAGE3/ACCI1_pp_3/_20_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_3/_24_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_3/_19_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_3/_20_ ),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_3/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE3/ACCI1_pp_3/_25_  (.A(\u_multiplier/STAGE3/ACCI1_pp_3/_19_ ),
    .B(\u_multiplier/STAGE3/ACCI1_pp_3/_20_ ),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_3/_16_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_3/_26_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_3/_18_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_3/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_3_s ));
 AOI22_X1 \u_multiplier/STAGE3/ACCI1_pp_3/_27_  (.A1(\u_multiplier/s_3 [1]),
    .A2(\u_multiplier/s_3 [0]),
    .B1(\u_multiplier/s_3 [2]),
    .B2(\u_multiplier/s_3 [3]),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_3/_28_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_3/_15_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_3/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_3_c ));
 NAND3_X1 \u_multiplier/STAGE3/ACCI1_pp_4/_21_  (.A1(\u_multiplier/s_4 [1]),
    .A2(\u_multiplier/s_4 [0]),
    .A3(\u_multiplier/s_4 [2]),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_4/_18_ ));
 XOR2_X2 \u_multiplier/STAGE3/ACCI1_pp_4/_22_  (.A(\u_multiplier/s_4 [1]),
    .B(\u_multiplier/s_4 [0]),
    .Z(\u_multiplier/STAGE3/ACCI1_pp_4/_19_ ));
 XOR2_X2 \u_multiplier/STAGE3/ACCI1_pp_4/_23_  (.A(\u_multiplier/s_4 [2]),
    .B(\u_multiplier/s_4 [3]),
    .Z(\u_multiplier/STAGE3/ACCI1_pp_4/_20_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_4/_24_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_4/_19_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_4/_20_ ),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_4/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE3/ACCI1_pp_4/_25_  (.A(\u_multiplier/STAGE3/ACCI1_pp_4/_19_ ),
    .B(\u_multiplier/STAGE3/ACCI1_pp_4/_20_ ),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_4/_16_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_4/_26_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_4/_18_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_4/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_4_s ));
 AOI22_X1 \u_multiplier/STAGE3/ACCI1_pp_4/_27_  (.A1(\u_multiplier/s_4 [1]),
    .A2(\u_multiplier/s_4 [0]),
    .B1(\u_multiplier/s_4 [2]),
    .B2(\u_multiplier/s_4 [3]),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_4/_28_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_4/_15_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_4/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_4_c ));
 NAND3_X1 \u_multiplier/STAGE3/ACCI1_pp_5/_21_  (.A1(\u_multiplier/s_5 [1]),
    .A2(\u_multiplier/s_5 [0]),
    .A3(\u_multiplier/s_5 [2]),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_5/_18_ ));
 XOR2_X2 \u_multiplier/STAGE3/ACCI1_pp_5/_22_  (.A(\u_multiplier/s_5 [1]),
    .B(\u_multiplier/s_5 [0]),
    .Z(\u_multiplier/STAGE3/ACCI1_pp_5/_19_ ));
 XOR2_X2 \u_multiplier/STAGE3/ACCI1_pp_5/_23_  (.A(\u_multiplier/s_5 [2]),
    .B(\u_multiplier/s_5 [3]),
    .Z(\u_multiplier/STAGE3/ACCI1_pp_5/_20_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_5/_24_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_5/_19_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_5/_20_ ),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_5/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE3/ACCI1_pp_5/_25_  (.A(\u_multiplier/STAGE3/ACCI1_pp_5/_19_ ),
    .B(\u_multiplier/STAGE3/ACCI1_pp_5/_20_ ),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_5/_16_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_5/_26_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_5/_18_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_5/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_5_s ));
 AOI22_X1 \u_multiplier/STAGE3/ACCI1_pp_5/_27_  (.A1(\u_multiplier/s_5 [1]),
    .A2(\u_multiplier/s_5 [0]),
    .B1(\u_multiplier/s_5 [2]),
    .B2(\u_multiplier/s_5 [3]),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_5/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_5/_28_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_5/_15_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_5/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_5_c ));
 NAND3_X1 \u_multiplier/STAGE3/ACCI1_pp_6/_21_  (.A1(\u_multiplier/s_6 [1]),
    .A2(\u_multiplier/s_6 [0]),
    .A3(\u_multiplier/s_6 [2]),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_6/_18_ ));
 XOR2_X2 \u_multiplier/STAGE3/ACCI1_pp_6/_22_  (.A(\u_multiplier/s_6 [1]),
    .B(\u_multiplier/s_6 [0]),
    .Z(\u_multiplier/STAGE3/ACCI1_pp_6/_19_ ));
 XOR2_X2 \u_multiplier/STAGE3/ACCI1_pp_6/_23_  (.A(\u_multiplier/s_6 [2]),
    .B(\u_multiplier/s_6 [3]),
    .Z(\u_multiplier/STAGE3/ACCI1_pp_6/_20_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_6/_24_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_6/_19_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_6/_20_ ),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_6/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE3/ACCI1_pp_6/_25_  (.A(\u_multiplier/STAGE3/ACCI1_pp_6/_19_ ),
    .B(\u_multiplier/STAGE3/ACCI1_pp_6/_20_ ),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_6/_16_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_6/_26_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_6/_18_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_6/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_6_s ));
 AOI22_X1 \u_multiplier/STAGE3/ACCI1_pp_6/_27_  (.A1(\u_multiplier/s_6 [1]),
    .A2(\u_multiplier/s_6 [0]),
    .B1(\u_multiplier/s_6 [2]),
    .B2(\u_multiplier/s_6 [3]),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_6/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_6/_28_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_6/_15_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_6/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_6_c ));
 NAND3_X1 \u_multiplier/STAGE3/ACCI1_pp_7/_21_  (.A1(\u_multiplier/s_7 [1]),
    .A2(\u_multiplier/s_7 [0]),
    .A3(\u_multiplier/s_7 [2]),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_7/_18_ ));
 XOR2_X2 \u_multiplier/STAGE3/ACCI1_pp_7/_22_  (.A(\u_multiplier/s_7 [1]),
    .B(\u_multiplier/s_7 [0]),
    .Z(\u_multiplier/STAGE3/ACCI1_pp_7/_19_ ));
 XOR2_X2 \u_multiplier/STAGE3/ACCI1_pp_7/_23_  (.A(\u_multiplier/s_7 [2]),
    .B(\u_multiplier/s_7 [3]),
    .Z(\u_multiplier/STAGE3/ACCI1_pp_7/_20_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_7/_24_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_7/_19_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_7/_20_ ),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_7/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE3/ACCI1_pp_7/_25_  (.A(\u_multiplier/STAGE3/ACCI1_pp_7/_19_ ),
    .B(\u_multiplier/STAGE3/ACCI1_pp_7/_20_ ),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_7/_16_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_7/_26_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_7/_18_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_7/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_7_s ));
 AOI22_X1 \u_multiplier/STAGE3/ACCI1_pp_7/_27_  (.A1(\u_multiplier/s_7 [1]),
    .A2(\u_multiplier/s_7 [0]),
    .B1(\u_multiplier/s_7 [2]),
    .B2(\u_multiplier/s_7 [3]),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_7/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_7/_28_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_7/_15_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_7/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_7_c ));
 NAND3_X1 \u_multiplier/STAGE3/ACCI1_pp_8/_21_  (.A1(\u_multiplier/s_8 [1]),
    .A2(\u_multiplier/s_8 [0]),
    .A3(\u_multiplier/s_8 [2]),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_8/_18_ ));
 XOR2_X2 \u_multiplier/STAGE3/ACCI1_pp_8/_22_  (.A(\u_multiplier/s_8 [1]),
    .B(\u_multiplier/s_8 [0]),
    .Z(\u_multiplier/STAGE3/ACCI1_pp_8/_19_ ));
 XOR2_X2 \u_multiplier/STAGE3/ACCI1_pp_8/_23_  (.A(\u_multiplier/s_8 [2]),
    .B(\u_multiplier/s_8 [3]),
    .Z(\u_multiplier/STAGE3/ACCI1_pp_8/_20_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_8/_24_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_8/_19_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_8/_20_ ),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_8/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE3/ACCI1_pp_8/_25_  (.A(\u_multiplier/STAGE3/ACCI1_pp_8/_19_ ),
    .B(\u_multiplier/STAGE3/ACCI1_pp_8/_20_ ),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_8/_16_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_8/_26_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_8/_18_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_8/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_8_s ));
 AOI22_X1 \u_multiplier/STAGE3/ACCI1_pp_8/_27_  (.A1(\u_multiplier/s_8 [1]),
    .A2(\u_multiplier/s_8 [0]),
    .B1(\u_multiplier/s_8 [2]),
    .B2(\u_multiplier/s_8 [3]),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_8/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_8/_28_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_8/_15_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_8/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_8_c ));
 NAND3_X1 \u_multiplier/STAGE3/ACCI1_pp_9/_21_  (.A1(\u_multiplier/s_9 [1]),
    .A2(\u_multiplier/s_9 [0]),
    .A3(\u_multiplier/s_9 [2]),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_9/_18_ ));
 XOR2_X2 \u_multiplier/STAGE3/ACCI1_pp_9/_22_  (.A(\u_multiplier/s_9 [1]),
    .B(\u_multiplier/s_9 [0]),
    .Z(\u_multiplier/STAGE3/ACCI1_pp_9/_19_ ));
 XOR2_X2 \u_multiplier/STAGE3/ACCI1_pp_9/_23_  (.A(\u_multiplier/s_9 [2]),
    .B(\u_multiplier/s_9 [3]),
    .Z(\u_multiplier/STAGE3/ACCI1_pp_9/_20_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_9/_24_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_9/_19_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_9/_20_ ),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_9/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE3/ACCI1_pp_9/_25_  (.A(\u_multiplier/STAGE3/ACCI1_pp_9/_19_ ),
    .B(\u_multiplier/STAGE3/ACCI1_pp_9/_20_ ),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_9/_16_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_9/_26_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_9/_18_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_9/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_9_s ));
 AOI22_X1 \u_multiplier/STAGE3/ACCI1_pp_9/_27_  (.A1(\u_multiplier/s_9 [1]),
    .A2(\u_multiplier/s_9 [0]),
    .B1(\u_multiplier/s_9 [2]),
    .B2(\u_multiplier/s_9 [3]),
    .ZN(\u_multiplier/STAGE3/ACCI1_pp_9/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/ACCI1_pp_9/_28_  (.A1(\u_multiplier/STAGE3/ACCI1_pp_9/_15_ ),
    .A2(\u_multiplier/STAGE3/ACCI1_pp_9/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_9_c ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_16_1/_18_  (.A(net64),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_16_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_16_1/_19_  (.A1(\u_multiplier/s_16 [1]),
    .A2(\u_multiplier/s_16 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_16_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_16_1/_20_  (.A(\u_multiplier/s_16 [1]),
    .B(\u_multiplier/s_16 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_16_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_16_1/_21_  (.A1(\u_multiplier/s_16 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_16_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_16_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_16_1/_22_  (.A(\u_multiplier/s_16 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_16_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_16_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_16_1/_23_  (.A1(\u_multiplier/s_16 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_16_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_16_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_16_1/_24_  (.A(\u_multiplier/s_16 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_16_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_16_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_16_1/_25_  (.A(net65),
    .B(\u_multiplier/STAGE3/E_4_2_pp_16_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_16_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_16_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_16_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_16_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_16_c2 ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp_16_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_16_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_16_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_16_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_16_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_17_1/_18_  (.A(\u_multiplier/STAGE3/pp_16_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_17_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_17_1/_19_  (.A1(\u_multiplier/s_17 [1]),
    .A2(\u_multiplier/s_17 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_17_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_17_1/_20_  (.A(\u_multiplier/s_17 [1]),
    .B(\u_multiplier/s_17 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_17_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_17_1/_21_  (.A1(\u_multiplier/s_17 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_17_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_17_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_17_1/_22_  (.A(\u_multiplier/s_17 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_17_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_17_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_17_1/_23_  (.A1(\u_multiplier/s_17 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_17_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_17_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_17_1/_24_  (.A(\u_multiplier/s_17 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_17_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_17_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_17_1/_25_  (.A(\u_multiplier/STAGE3/pp_16_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_17_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_17_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_17_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_17_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_17_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_17_c2 ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp_17_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_17_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_17_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_17_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_17_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_18_1/_18_  (.A(\u_multiplier/STAGE3/pp_17_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_18_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_18_1/_19_  (.A1(\u_multiplier/s_18 [1]),
    .A2(\u_multiplier/s_18 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_18_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_18_1/_20_  (.A(\u_multiplier/s_18 [1]),
    .B(\u_multiplier/s_18 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_18_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_18_1/_21_  (.A1(\u_multiplier/s_18 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_18_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_18_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_18_1/_22_  (.A(\u_multiplier/s_18 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_18_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_18_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_18_1/_23_  (.A1(\u_multiplier/s_18 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_18_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_18_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_18_1/_24_  (.A(\u_multiplier/s_18 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_18_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_18_1/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE3/E_4_2_pp_18_1/_25_  (.A(\u_multiplier/STAGE3/pp_17_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_18_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_18_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_18_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_18_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_18_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_18_c2 ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp_18_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_18_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_18_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_18_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_18_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_19_1/_18_  (.A(\u_multiplier/STAGE3/pp_18_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_19_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_19_1/_19_  (.A1(\u_multiplier/s_19 [1]),
    .A2(\u_multiplier/s_19 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_19_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_19_1/_20_  (.A(\u_multiplier/s_19 [1]),
    .B(\u_multiplier/s_19 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_19_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_19_1/_21_  (.A1(\u_multiplier/s_19 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_19_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_19_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_19_1/_22_  (.A(\u_multiplier/s_19 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_19_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_19_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_19_1/_23_  (.A1(\u_multiplier/s_19 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_19_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_19_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_19_1/_24_  (.A(\u_multiplier/s_19 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_19_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_19_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_19_1/_25_  (.A(\u_multiplier/STAGE3/pp_18_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_19_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_19_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_19_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_19_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_19_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_19_c2 ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp_19_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_19_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_19_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_19_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_19_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_20_1/_18_  (.A(\u_multiplier/STAGE3/pp_19_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_20_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_20_1/_19_  (.A1(\u_multiplier/s_20 [1]),
    .A2(\u_multiplier/s_20 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_20_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_20_1/_20_  (.A(\u_multiplier/s_20 [1]),
    .B(\u_multiplier/s_20 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_20_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_20_1/_21_  (.A1(\u_multiplier/s_20 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_20_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_20_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_20_1/_22_  (.A(\u_multiplier/s_20 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_20_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_20_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_20_1/_23_  (.A1(\u_multiplier/s_20 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_20_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_20_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_20_1/_24_  (.A(\u_multiplier/s_20 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_20_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_20_1/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE3/E_4_2_pp_20_1/_25_  (.A(\u_multiplier/STAGE3/pp_19_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_20_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_20_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_20_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_20_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_20_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_20_c2 ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp_20_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_20_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_20_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_20_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_20_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_21_1/_18_  (.A(\u_multiplier/STAGE3/pp_20_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_21_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_21_1/_19_  (.A1(\u_multiplier/s_21 [1]),
    .A2(\u_multiplier/s_21 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_21_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_21_1/_20_  (.A(\u_multiplier/s_21 [1]),
    .B(\u_multiplier/s_21 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_21_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_21_1/_21_  (.A1(\u_multiplier/s_21 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_21_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_21_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_21_1/_22_  (.A(\u_multiplier/s_21 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_21_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_21_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_21_1/_23_  (.A1(\u_multiplier/s_21 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_21_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_21_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_21_1/_24_  (.A(\u_multiplier/s_21 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_21_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_21_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_21_1/_25_  (.A(\u_multiplier/STAGE3/pp_20_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_21_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_21_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_21_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_21_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_21_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_21_c2 ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp_21_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_21_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_21_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_21_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_21_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_22_1/_18_  (.A(\u_multiplier/STAGE3/pp_21_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_22_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_22_1/_19_  (.A1(\u_multiplier/s_22 [1]),
    .A2(\u_multiplier/s_22 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_22_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_22_1/_20_  (.A(\u_multiplier/s_22 [1]),
    .B(\u_multiplier/s_22 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_22_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_22_1/_21_  (.A1(\u_multiplier/s_22 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_22_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_22_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_22_1/_22_  (.A(\u_multiplier/s_22 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_22_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_22_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_22_1/_23_  (.A1(\u_multiplier/s_22 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_22_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_22_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_22_1/_24_  (.A(\u_multiplier/s_22 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_22_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_22_1/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE3/E_4_2_pp_22_1/_25_  (.A(\u_multiplier/STAGE3/pp_21_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_22_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_22_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_22_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_22_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_22_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_22_c2 ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp_22_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_22_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_22_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_22_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_22_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_23_1/_18_  (.A(\u_multiplier/STAGE3/pp_22_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_23_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_23_1/_19_  (.A1(\u_multiplier/s_23 [1]),
    .A2(\u_multiplier/s_23 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_23_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_23_1/_20_  (.A(\u_multiplier/s_23 [1]),
    .B(\u_multiplier/s_23 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_23_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_23_1/_21_  (.A1(\u_multiplier/s_23 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_23_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_23_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_23_1/_22_  (.A(\u_multiplier/s_23 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_23_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_23_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_23_1/_23_  (.A1(\u_multiplier/s_23 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_23_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_23_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_23_1/_24_  (.A(\u_multiplier/s_23 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_23_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_23_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_23_1/_25_  (.A(\u_multiplier/STAGE3/pp_22_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_23_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_23_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_23_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_23_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_23_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_23_c2 ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp_23_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_23_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_23_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_23_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_23_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_24_1/_18_  (.A(\u_multiplier/STAGE3/pp_23_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_24_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_24_1/_19_  (.A1(\u_multiplier/s_24 [1]),
    .A2(\u_multiplier/s_24 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_24_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_24_1/_20_  (.A(\u_multiplier/s_24 [1]),
    .B(\u_multiplier/s_24 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_24_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_24_1/_21_  (.A1(\u_multiplier/s_24 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_24_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_24_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_24_1/_22_  (.A(\u_multiplier/s_24 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_24_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_24_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_24_1/_23_  (.A1(\u_multiplier/s_24 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_24_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_24_1/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE3/E_4_2_pp_24_1/_24_  (.A(\u_multiplier/s_24 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_24_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_24_1/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE3/E_4_2_pp_24_1/_25_  (.A(\u_multiplier/STAGE3/pp_23_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_24_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_24_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_24_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_24_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_24_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_24_c2 ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp_24_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_24_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_24_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_24_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_24_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_25_1/_18_  (.A(\u_multiplier/STAGE3/pp_24_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_25_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_25_1/_19_  (.A1(\u_multiplier/s_25 [1]),
    .A2(\u_multiplier/s_25 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_25_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_25_1/_20_  (.A(\u_multiplier/s_25 [1]),
    .B(\u_multiplier/s_25 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_25_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_25_1/_21_  (.A1(\u_multiplier/s_25 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_25_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_25_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_25_1/_22_  (.A(\u_multiplier/s_25 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_25_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_25_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_25_1/_23_  (.A1(\u_multiplier/s_25 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_25_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_25_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_25_1/_24_  (.A(\u_multiplier/s_25 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_25_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_25_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_25_1/_25_  (.A(\u_multiplier/STAGE3/pp_24_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_25_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_25_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_25_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_25_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_25_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_25_c2 ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp_25_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_25_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_25_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_25_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_25_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_26_1/_18_  (.A(\u_multiplier/STAGE3/pp_25_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_26_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_26_1/_19_  (.A1(\u_multiplier/s_26 [1]),
    .A2(\u_multiplier/s_26 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_26_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_26_1/_20_  (.A(\u_multiplier/s_26 [1]),
    .B(\u_multiplier/s_26 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_26_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_26_1/_21_  (.A1(\u_multiplier/s_26 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_26_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_26_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_26_1/_22_  (.A(\u_multiplier/s_26 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_26_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_26_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_26_1/_23_  (.A1(\u_multiplier/s_26 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_26_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_26_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_26_1/_24_  (.A(\u_multiplier/s_26 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_26_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_26_1/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE3/E_4_2_pp_26_1/_25_  (.A(\u_multiplier/STAGE3/pp_25_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_26_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_26_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_26_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_26_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_26_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_26_c2 ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp_26_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_26_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_26_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_26_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_26_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_27_1/_18_  (.A(\u_multiplier/STAGE3/pp_26_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_27_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_27_1/_19_  (.A1(\u_multiplier/s_27 [1]),
    .A2(\u_multiplier/s_27 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_27_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_27_1/_20_  (.A(\u_multiplier/s_27 [1]),
    .B(\u_multiplier/s_27 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_27_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_27_1/_21_  (.A1(\u_multiplier/s_27 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_27_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_27_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_27_1/_22_  (.A(\u_multiplier/s_27 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_27_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_27_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_27_1/_23_  (.A1(\u_multiplier/s_27 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_27_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_27_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_27_1/_24_  (.A(\u_multiplier/s_27 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_27_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_27_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_27_1/_25_  (.A(\u_multiplier/STAGE3/pp_26_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_27_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_27_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_27_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_27_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_27_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_27_c2 ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp_27_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_27_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_27_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_27_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_27_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_28_1/_18_  (.A(\u_multiplier/STAGE3/pp_27_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_28_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_28_1/_19_  (.A1(\u_multiplier/s_28 [1]),
    .A2(\u_multiplier/s_28 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_28_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_28_1/_20_  (.A(\u_multiplier/s_28 [1]),
    .B(\u_multiplier/s_28 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_28_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_28_1/_21_  (.A1(\u_multiplier/s_28 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_28_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_28_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_28_1/_22_  (.A(\u_multiplier/s_28 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_28_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_28_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_28_1/_23_  (.A1(\u_multiplier/s_28 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_28_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_28_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_28_1/_24_  (.A(\u_multiplier/s_28 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_28_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_28_1/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE3/E_4_2_pp_28_1/_25_  (.A(\u_multiplier/STAGE3/pp_27_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_28_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_28_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_28_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_28_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_28_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_28_c2 ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp_28_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_28_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_28_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_28_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_28_c1 ));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_40_  (.A1(\u_multiplier/STAGE3/pp_2_c ),
    .A2(\u_multiplier/STAGE3/pp_3_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla1/_25_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_41_  (.A1(\u_multiplier/s_2 [2]),
    .A2(\u_multiplier/STAGE3/pp_2_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla1/_26_ ));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_42_  (.A1(\u_multiplier/s_1 [0]),
    .A2(\u_multiplier/s_1 [1]),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla1/_27_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_43_  (.A1(net66),
    .A2(\u_multiplier/s_0 ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla1/_28_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_44_  (.A1(net67),
    .A2(\u_multiplier/s_0 ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla1/_29_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_45_  (.A(net68),
    .B(\u_multiplier/s_0 ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla1/_30_ ));
 AOI21_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_46_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla1/_28_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla1/_29_ ),
    .B2(net69),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla1/_31_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_47_  (.A1(\u_multiplier/s_1 [0]),
    .A2(\u_multiplier/s_1 [1]),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla1/_32_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_48_  (.A(\u_multiplier/s_1 [0]),
    .B(\u_multiplier/s_1 [1]),
    .Z(\u_multiplier/STAGE3/Final_add/cla1/cla1/_33_ ));
 OAI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla1/_49_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla1/_27_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla1/_31_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/cla1/_32_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla1/_34_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_50_  (.A1(\u_multiplier/s_2 [2]),
    .A2(\u_multiplier/STAGE3/pp_2_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla1/_35_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_51_  (.A(\u_multiplier/s_2 [2]),
    .B(\u_multiplier/STAGE3/pp_2_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla1/_36_ ));
 AOI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla1/_52_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla1/_26_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla1/_34_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/cla1/_35_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla1/_37_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_53_  (.A1(\u_multiplier/STAGE3/pp_2_c ),
    .A2(\u_multiplier/STAGE3/pp_3_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla1/_38_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_54_  (.A(\u_multiplier/STAGE3/pp_2_c ),
    .B(\u_multiplier/STAGE3/pp_3_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla1/cla1/_39_ ));
 OAI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla1/_55_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla1/_25_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla1/_37_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/cla1/_38_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/c1 ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_56_  (.A(net70),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla1/_30_ ),
    .ZN(product[0]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_57_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla1/_31_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla1/_33_ ),
    .ZN(product[1]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_58_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla1/_34_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla1/_36_ ),
    .ZN(product[2]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_59_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla1/_37_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla1/_39_ ),
    .ZN(product[3]));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_40_  (.A1(\u_multiplier/STAGE3/pp_6_c ),
    .A2(\u_multiplier/STAGE3/pp_7_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla2/_25_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_41_  (.A1(\u_multiplier/STAGE3/pp_5_c ),
    .A2(\u_multiplier/STAGE3/pp_6_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla2/_26_ ));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_42_  (.A1(\u_multiplier/STAGE3/pp_4_c ),
    .A2(\u_multiplier/STAGE3/pp_5_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla2/_27_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_43_  (.A1(\u_multiplier/STAGE3/pp_3_c ),
    .A2(\u_multiplier/STAGE3/pp_4_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla2/_28_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_44_  (.A1(\u_multiplier/STAGE3/pp_3_c ),
    .A2(\u_multiplier/STAGE3/pp_4_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla2/_29_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_45_  (.A(\u_multiplier/STAGE3/pp_3_c ),
    .B(\u_multiplier/STAGE3/pp_4_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla2/_30_ ));
 AOI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla2/_46_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla2/_28_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla2/_29_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/c1 ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla2/_31_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_47_  (.A1(\u_multiplier/STAGE3/pp_4_c ),
    .A2(\u_multiplier/STAGE3/pp_5_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla2/_32_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_48_  (.A(\u_multiplier/STAGE3/pp_4_c ),
    .B(\u_multiplier/STAGE3/pp_5_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla1/cla2/_33_ ));
 OAI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla2/_49_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla2/_27_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla2/_31_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/cla2/_32_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla2/_34_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_50_  (.A1(\u_multiplier/STAGE3/pp_5_c ),
    .A2(\u_multiplier/STAGE3/pp_6_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla2/_35_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_51_  (.A(\u_multiplier/STAGE3/pp_5_c ),
    .B(\u_multiplier/STAGE3/pp_6_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla2/_36_ ));
 AOI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla2/_52_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla2/_26_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla2/_34_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/cla2/_35_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla2/_37_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_53_  (.A1(\u_multiplier/STAGE3/pp_6_c ),
    .A2(\u_multiplier/STAGE3/pp_7_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla2/_38_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_54_  (.A(\u_multiplier/STAGE3/pp_6_c ),
    .B(\u_multiplier/STAGE3/pp_7_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla1/cla2/_39_ ));
 OAI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla2/_55_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla2/_25_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla2/_37_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/cla2/_38_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/c2 ));
 XNOR2_X2 \u_multiplier/STAGE3/Final_add/cla1/cla2/_56_  (.A(\u_multiplier/STAGE3/Final_add/cla1/c1 ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla2/_30_ ),
    .ZN(product[4]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_57_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla2/_31_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla2/_33_ ),
    .ZN(product[5]));
 XNOR2_X2 \u_multiplier/STAGE3/Final_add/cla1/cla2/_58_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla2/_34_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla2/_36_ ),
    .ZN(product[6]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_59_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla2/_37_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla2/_39_ ),
    .ZN(product[7]));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_40_  (.A1(\u_multiplier/STAGE3/pp_10_c ),
    .A2(\u_multiplier/STAGE3/pp_11_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla3/_25_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_41_  (.A1(\u_multiplier/STAGE3/pp_9_c ),
    .A2(\u_multiplier/STAGE3/pp_10_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla3/_26_ ));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_42_  (.A1(\u_multiplier/STAGE3/pp_8_c ),
    .A2(\u_multiplier/STAGE3/pp_9_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla3/_27_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_43_  (.A1(\u_multiplier/STAGE3/pp_7_c ),
    .A2(\u_multiplier/STAGE3/pp_8_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla3/_28_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_44_  (.A1(\u_multiplier/STAGE3/pp_7_c ),
    .A2(\u_multiplier/STAGE3/pp_8_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla3/_29_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_45_  (.A(\u_multiplier/STAGE3/pp_7_c ),
    .B(\u_multiplier/STAGE3/pp_8_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla3/_30_ ));
 AOI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla3/_46_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla3/_28_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla3/_29_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/c2 ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla3/_31_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_47_  (.A1(\u_multiplier/STAGE3/pp_8_c ),
    .A2(\u_multiplier/STAGE3/pp_9_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla3/_32_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_48_  (.A(\u_multiplier/STAGE3/pp_8_c ),
    .B(\u_multiplier/STAGE3/pp_9_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla1/cla3/_33_ ));
 OAI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla3/_49_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla3/_27_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla3/_31_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/cla3/_32_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla3/_34_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_50_  (.A1(\u_multiplier/STAGE3/pp_9_c ),
    .A2(\u_multiplier/STAGE3/pp_10_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla3/_35_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_51_  (.A(\u_multiplier/STAGE3/pp_9_c ),
    .B(\u_multiplier/STAGE3/pp_10_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla3/_36_ ));
 AOI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla3/_52_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla3/_26_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla3/_34_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/cla3/_35_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla3/_37_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_53_  (.A1(\u_multiplier/STAGE3/pp_10_c ),
    .A2(\u_multiplier/STAGE3/pp_11_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla3/_38_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_54_  (.A(\u_multiplier/STAGE3/pp_10_c ),
    .B(\u_multiplier/STAGE3/pp_11_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla1/cla3/_39_ ));
 OAI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla3/_55_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla3/_25_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla3/_37_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/cla3/_38_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/c3 ));
 XNOR2_X2 \u_multiplier/STAGE3/Final_add/cla1/cla3/_56_  (.A(\u_multiplier/STAGE3/Final_add/cla1/c2 ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla3/_30_ ),
    .ZN(product[8]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_57_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla3/_31_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla3/_33_ ),
    .ZN(product[9]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_58_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla3/_34_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla3/_36_ ),
    .ZN(product[10]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_59_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla3/_37_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla3/_39_ ),
    .ZN(product[11]));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_40_  (.A1(\u_multiplier/STAGE3/pp_14_c ),
    .A2(\u_multiplier/STAGE3/pp_15_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla4/_25_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_41_  (.A1(\u_multiplier/STAGE3/pp_13_c ),
    .A2(\u_multiplier/STAGE3/pp_14_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla4/_26_ ));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_42_  (.A1(\u_multiplier/STAGE3/pp_12_c ),
    .A2(\u_multiplier/STAGE3/pp_13_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla4/_27_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_43_  (.A1(\u_multiplier/STAGE3/pp_11_c ),
    .A2(\u_multiplier/STAGE3/pp_12_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla4/_28_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_44_  (.A1(\u_multiplier/STAGE3/pp_11_c ),
    .A2(\u_multiplier/STAGE3/pp_12_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla4/_29_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_45_  (.A(\u_multiplier/STAGE3/pp_11_c ),
    .B(\u_multiplier/STAGE3/pp_12_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla4/_30_ ));
 AOI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla4/_46_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla4/_28_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla4/_29_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/c3 ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla4/_31_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_47_  (.A1(\u_multiplier/STAGE3/pp_12_c ),
    .A2(\u_multiplier/STAGE3/pp_13_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla4/_32_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_48_  (.A(\u_multiplier/STAGE3/pp_12_c ),
    .B(\u_multiplier/STAGE3/pp_13_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla1/cla4/_33_ ));
 OAI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla4/_49_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla4/_27_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla4/_31_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/cla4/_32_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla4/_34_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_50_  (.A1(\u_multiplier/STAGE3/pp_13_c ),
    .A2(\u_multiplier/STAGE3/pp_14_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla4/_35_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_51_  (.A(\u_multiplier/STAGE3/pp_13_c ),
    .B(\u_multiplier/STAGE3/pp_14_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla4/_36_ ));
 AOI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla4/_52_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla4/_26_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla4/_34_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/cla4/_35_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla4/_37_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_53_  (.A1(\u_multiplier/STAGE3/pp_14_c ),
    .A2(\u_multiplier/STAGE3/pp_15_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla4/_38_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_54_  (.A(\u_multiplier/STAGE3/pp_14_c ),
    .B(\u_multiplier/STAGE3/pp_15_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla1/cla4/_39_ ));
 OAI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla4/_55_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla4/_25_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla4/_37_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/cla4/_38_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/c1 ));
 XNOR2_X2 \u_multiplier/STAGE3/Final_add/cla1/cla4/_56_  (.A(\u_multiplier/STAGE3/Final_add/cla1/c3 ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla4/_30_ ),
    .ZN(product[12]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_57_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla4/_31_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla4/_33_ ),
    .ZN(product[13]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_58_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla4/_34_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla4/_36_ ),
    .ZN(product[14]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_59_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla4/_37_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla4/_39_ ),
    .ZN(product[15]));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_40_  (.A1(\u_multiplier/STAGE3/pp_18_c1 ),
    .A2(\u_multiplier/STAGE3/pp_19_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla1/_25_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_41_  (.A1(\u_multiplier/STAGE3/pp_17_c1 ),
    .A2(\u_multiplier/STAGE3/pp_18_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla1/_26_ ));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_42_  (.A1(\u_multiplier/STAGE3/pp_16_c1 ),
    .A2(\u_multiplier/STAGE3/pp_17_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla1/_27_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_43_  (.A1(\u_multiplier/STAGE3/pp_15_c ),
    .A2(\u_multiplier/STAGE3/pp_16_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla1/_28_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_44_  (.A1(\u_multiplier/STAGE3/pp_15_c ),
    .A2(\u_multiplier/STAGE3/pp_16_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla1/_29_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_45_  (.A(\u_multiplier/STAGE3/pp_15_c ),
    .B(\u_multiplier/STAGE3/pp_16_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla1/_30_ ));
 AOI21_X2 \u_multiplier/STAGE3/Final_add/cla2/cla1/_46_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla1/_28_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla1/_29_ ),
    .B2(\u_multiplier/STAGE3/Final_add/c1 ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla1/_31_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_47_  (.A1(\u_multiplier/STAGE3/pp_16_c1 ),
    .A2(\u_multiplier/STAGE3/pp_17_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla1/_32_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_48_  (.A(\u_multiplier/STAGE3/pp_16_c1 ),
    .B(\u_multiplier/STAGE3/pp_17_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla2/cla1/_33_ ));
 OAI21_X2 \u_multiplier/STAGE3/Final_add/cla2/cla1/_49_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla1/_27_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla1/_31_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/cla1/_32_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla1/_34_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_50_  (.A1(\u_multiplier/STAGE3/pp_17_c1 ),
    .A2(\u_multiplier/STAGE3/pp_18_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla1/_35_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_51_  (.A(\u_multiplier/STAGE3/pp_17_c1 ),
    .B(\u_multiplier/STAGE3/pp_18_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla1/_36_ ));
 AOI21_X2 \u_multiplier/STAGE3/Final_add/cla2/cla1/_52_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla1/_26_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla1/_34_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/cla1/_35_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla1/_37_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_53_  (.A1(\u_multiplier/STAGE3/pp_18_c1 ),
    .A2(\u_multiplier/STAGE3/pp_19_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla1/_38_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_54_  (.A(\u_multiplier/STAGE3/pp_18_c1 ),
    .B(\u_multiplier/STAGE3/pp_19_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla2/cla1/_39_ ));
 OAI21_X2 \u_multiplier/STAGE3/Final_add/cla2/cla1/_55_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla1/_25_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla1/_37_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/cla1/_38_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/c1 ));
 XNOR2_X2 \u_multiplier/STAGE3/Final_add/cla2/cla1/_56_  (.A(\u_multiplier/STAGE3/Final_add/c1 ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla1/_30_ ),
    .ZN(product[16]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_57_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla1/_31_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla1/_33_ ),
    .ZN(product[17]));
 XNOR2_X2 \u_multiplier/STAGE3/Final_add/cla2/cla1/_58_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla1/_34_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla1/_36_ ),
    .ZN(product[18]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_59_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla1/_37_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla1/_39_ ),
    .ZN(product[19]));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_40_  (.A1(\u_multiplier/STAGE3/pp_22_c1 ),
    .A2(\u_multiplier/STAGE3/pp_23_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla2/_25_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_41_  (.A1(\u_multiplier/STAGE3/pp_21_c1 ),
    .A2(\u_multiplier/STAGE3/pp_22_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla2/_26_ ));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_42_  (.A1(\u_multiplier/STAGE3/pp_20_c1 ),
    .A2(\u_multiplier/STAGE3/pp_21_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla2/_27_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_43_  (.A1(\u_multiplier/STAGE3/pp_19_c1 ),
    .A2(\u_multiplier/STAGE3/pp_20_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla2/_28_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_44_  (.A1(\u_multiplier/STAGE3/pp_19_c1 ),
    .A2(\u_multiplier/STAGE3/pp_20_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla2/_29_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_45_  (.A(\u_multiplier/STAGE3/pp_19_c1 ),
    .B(\u_multiplier/STAGE3/pp_20_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla2/_30_ ));
 AOI21_X2 \u_multiplier/STAGE3/Final_add/cla2/cla2/_46_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla2/_28_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla2/_29_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/c1 ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla2/_31_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_47_  (.A1(\u_multiplier/STAGE3/pp_20_c1 ),
    .A2(\u_multiplier/STAGE3/pp_21_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla2/_32_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_48_  (.A(\u_multiplier/STAGE3/pp_20_c1 ),
    .B(\u_multiplier/STAGE3/pp_21_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla2/cla2/_33_ ));
 OAI21_X2 \u_multiplier/STAGE3/Final_add/cla2/cla2/_49_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla2/_27_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla2/_31_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/cla2/_32_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla2/_34_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_50_  (.A1(\u_multiplier/STAGE3/pp_21_c1 ),
    .A2(\u_multiplier/STAGE3/pp_22_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla2/_35_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_51_  (.A(\u_multiplier/STAGE3/pp_21_c1 ),
    .B(\u_multiplier/STAGE3/pp_22_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla2/_36_ ));
 AOI21_X2 \u_multiplier/STAGE3/Final_add/cla2/cla2/_52_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla2/_26_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla2/_34_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/cla2/_35_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla2/_37_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_53_  (.A1(\u_multiplier/STAGE3/pp_22_c1 ),
    .A2(\u_multiplier/STAGE3/pp_23_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla2/_38_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_54_  (.A(\u_multiplier/STAGE3/pp_22_c1 ),
    .B(\u_multiplier/STAGE3/pp_23_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla2/cla2/_39_ ));
 OAI21_X2 \u_multiplier/STAGE3/Final_add/cla2/cla2/_55_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla2/_25_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla2/_37_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/cla2/_38_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/c2 ));
 XNOR2_X2 \u_multiplier/STAGE3/Final_add/cla2/cla2/_56_  (.A(\u_multiplier/STAGE3/Final_add/cla2/c1 ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla2/_30_ ),
    .ZN(product[20]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_57_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla2/_31_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla2/_33_ ),
    .ZN(product[21]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_58_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla2/_34_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla2/_36_ ),
    .ZN(product[22]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_59_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla2/_37_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla2/_39_ ),
    .ZN(product[23]));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_40_  (.A1(\u_multiplier/STAGE3/pp_26_c1 ),
    .A2(\u_multiplier/STAGE3/pp_27_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla3/_25_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_41_  (.A1(\u_multiplier/STAGE3/pp_25_c1 ),
    .A2(\u_multiplier/STAGE3/pp_26_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla3/_26_ ));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_42_  (.A1(\u_multiplier/STAGE3/pp_24_c1 ),
    .A2(\u_multiplier/STAGE3/pp_25_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla3/_27_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_43_  (.A1(\u_multiplier/STAGE3/pp_23_c1 ),
    .A2(\u_multiplier/STAGE3/pp_24_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla3/_28_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_44_  (.A1(\u_multiplier/STAGE3/pp_23_c1 ),
    .A2(\u_multiplier/STAGE3/pp_24_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla3/_29_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_45_  (.A(\u_multiplier/STAGE3/pp_23_c1 ),
    .B(\u_multiplier/STAGE3/pp_24_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla3/_30_ ));
 AOI21_X2 \u_multiplier/STAGE3/Final_add/cla2/cla3/_46_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla3/_28_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla3/_29_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/c2 ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla3/_31_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_47_  (.A1(\u_multiplier/STAGE3/pp_24_c1 ),
    .A2(\u_multiplier/STAGE3/pp_25_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla3/_32_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_48_  (.A(\u_multiplier/STAGE3/pp_24_c1 ),
    .B(\u_multiplier/STAGE3/pp_25_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla2/cla3/_33_ ));
 OAI21_X2 \u_multiplier/STAGE3/Final_add/cla2/cla3/_49_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla3/_27_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla3/_31_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/cla3/_32_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla3/_34_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_50_  (.A1(\u_multiplier/STAGE3/pp_25_c1 ),
    .A2(\u_multiplier/STAGE3/pp_26_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla3/_35_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_51_  (.A(\u_multiplier/STAGE3/pp_25_c1 ),
    .B(\u_multiplier/STAGE3/pp_26_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla3/_36_ ));
 AOI21_X2 \u_multiplier/STAGE3/Final_add/cla2/cla3/_52_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla3/_26_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla3/_34_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/cla3/_35_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla3/_37_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_53_  (.A1(\u_multiplier/STAGE3/pp_26_c1 ),
    .A2(\u_multiplier/STAGE3/pp_27_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla3/_38_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_54_  (.A(\u_multiplier/STAGE3/pp_26_c1 ),
    .B(\u_multiplier/STAGE3/pp_27_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla2/cla3/_39_ ));
 OAI21_X2 \u_multiplier/STAGE3/Final_add/cla2/cla3/_55_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla3/_25_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla3/_37_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/cla3/_38_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/c3 ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_56_  (.A(\u_multiplier/STAGE3/Final_add/cla2/c2 ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla3/_30_ ),
    .ZN(product[24]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_57_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla3/_31_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla3/_33_ ),
    .ZN(product[25]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_58_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla3/_34_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla3/_36_ ),
    .ZN(product[26]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_59_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla3/_37_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla3/_39_ ),
    .ZN(product[27]));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_40_  (.A1(net71),
    .A2(net72),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla4/_25_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_41_  (.A1(\u_multiplier/STAGE3/pp_29_c ),
    .A2(\u_multiplier/s_30 ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla4/_26_ ));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_42_  (.A1(\u_multiplier/STAGE3/pp_28_c1 ),
    .A2(\u_multiplier/STAGE3/pp_29_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla4/_27_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_43_  (.A1(\u_multiplier/STAGE3/pp_27_c1 ),
    .A2(\u_multiplier/STAGE3/pp_28_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla4/_28_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_44_  (.A1(\u_multiplier/STAGE3/pp_27_c1 ),
    .A2(\u_multiplier/STAGE3/pp_28_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla4/_29_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_45_  (.A(\u_multiplier/STAGE3/pp_27_c1 ),
    .B(\u_multiplier/STAGE3/pp_28_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla4/_30_ ));
 AOI21_X2 \u_multiplier/STAGE3/Final_add/cla2/cla4/_46_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla4/_28_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla4/_29_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/c3 ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla4/_31_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_47_  (.A1(\u_multiplier/STAGE3/pp_28_c1 ),
    .A2(\u_multiplier/STAGE3/pp_29_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla4/_32_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_48_  (.A(\u_multiplier/STAGE3/pp_28_c1 ),
    .B(\u_multiplier/STAGE3/pp_29_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla2/cla4/_33_ ));
 OAI21_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_49_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla4/_27_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla4/_31_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/cla4/_32_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla4/_34_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_50_  (.A1(\u_multiplier/STAGE3/pp_29_c ),
    .A2(\u_multiplier/s_30 ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla4/_35_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_51_  (.A(\u_multiplier/STAGE3/pp_29_c ),
    .B(\u_multiplier/s_30 ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla4/_36_ ));
 AOI21_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_52_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla4/_26_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla4/_34_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/cla4/_35_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla4/_37_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_53_  (.A1(net73),
    .A2(net74),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla4/_38_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_54_  (.A(net75),
    .B(net76),
    .Z(\u_multiplier/STAGE3/Final_add/cla2/cla4/_39_ ));
 OAI21_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_55_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla4/_25_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla4/_37_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/cla4/_38_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/Cout ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_56_  (.A(\u_multiplier/STAGE3/Final_add/cla2/c3 ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla4/_30_ ),
    .ZN(product[28]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_57_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla4/_31_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla4/_33_ ),
    .ZN(product[29]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_58_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla4/_34_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla4/_36_ ),
    .ZN(product[30]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_59_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla4/_37_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla4/_39_ ),
    .ZN(product[31]));
 INV_X1 \u_multiplier/STAGE3/Full_adder_pp_29/_12_  (.A(\u_multiplier/STAGE3/pp_28_c2 ),
    .ZN(\u_multiplier/STAGE3/Full_adder_pp_29/_08_ ));
 NAND3_X1 \u_multiplier/STAGE3/Full_adder_pp_29/_13_  (.A1(\u_multiplier/s_29 [1]),
    .A2(\u_multiplier/s_29 [0]),
    .A3(\u_multiplier/STAGE3/pp_28_c2 ),
    .ZN(\u_multiplier/STAGE3/Full_adder_pp_29/_09_ ));
 NOR2_X2 \u_multiplier/STAGE3/Full_adder_pp_29/_14_  (.A1(\u_multiplier/s_29 [1]),
    .A2(\u_multiplier/s_29 [0]),
    .ZN(\u_multiplier/STAGE3/Full_adder_pp_29/_10_ ));
 AOI21_X1 \u_multiplier/STAGE3/Full_adder_pp_29/_15_  (.A(\u_multiplier/STAGE3/pp_28_c2 ),
    .B1(\u_multiplier/s_29 [0]),
    .B2(\u_multiplier/s_29 [1]),
    .ZN(\u_multiplier/STAGE3/Full_adder_pp_29/_11_ ));
 NOR2_X2 \u_multiplier/STAGE3/Full_adder_pp_29/_16_  (.A1(\u_multiplier/STAGE3/Full_adder_pp_29/_10_ ),
    .A2(\u_multiplier/STAGE3/Full_adder_pp_29/_11_ ),
    .ZN(\u_multiplier/STAGE3/pp_29_c ));
 AOI22_X2 \u_multiplier/STAGE3/Full_adder_pp_29/_17_  (.A1(\u_multiplier/STAGE3/Full_adder_pp_29/_08_ ),
    .A2(\u_multiplier/STAGE3/Full_adder_pp_29/_10_ ),
    .B1(\u_multiplier/STAGE3/pp_29_c ),
    .B2(\u_multiplier/STAGE3/Full_adder_pp_29/_09_ ),
    .ZN(\u_multiplier/STAGE3/pp_29_s ));
 AND2_X1 \u_multiplier/STAGE3/Half_adder_pp_2/_4_  (.A1(\u_multiplier/s_2 [1]),
    .A2(\u_multiplier/s_2 [0]),
    .ZN(\u_multiplier/STAGE3/pp_2_c ));
 XOR2_X2 \u_multiplier/STAGE3/Half_adder_pp_2/_5_  (.A(\u_multiplier/s_2 [1]),
    .B(\u_multiplier/s_2 [0]),
    .Z(\u_multiplier/STAGE3/pp_2_s ));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_2_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_2_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_2_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_2_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_2_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_2_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_2_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_2_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_2_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_2_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_2_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_2_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_2_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_2_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_2_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_2_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_2_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_2_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_2_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_2_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_2_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_2_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_2_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_2_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_2_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_2_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_2_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_2_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_2_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_2_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_2_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_2_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_2_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_2_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_2_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_2_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_2_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_2_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_2_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_2_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_2_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_2_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_2_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_2_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_2_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_2_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_2_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_2_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_2_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_2_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_2_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_2_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_2_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_2_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_2_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_2_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_2_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_2_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_2_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_2_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_2_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_2_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_2_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_2_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_2_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_2_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_2_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_2_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_2_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_2_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_2_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_2_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_2_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_2_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_2_Right_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_2_Right_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_2_Right_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_2_Right_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_2_Right_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_2_Right_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_2_Right_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_2_Right_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_2_Right_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_2_Right_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_2_Right_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_2_Right_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_2_Right_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_2_Right_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_2_Right_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_2_Right_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_2_Right_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_2_Right_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_2_Right_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_2_Right_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_2_Right_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_2_Right_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_2_Right_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_2_Right_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_2_Right_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_2_Right_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_2_Right_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_2_Right_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_2_Right_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_2_Right_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_2_Right_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_1_Left_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_1_Left_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_1_Left_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_1_Left_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_1_Left_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_1_Left_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_1_Left_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_1_Left_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_1_Left_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_1_Left_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_1_Left_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_1_Left_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_1_Left_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_1_Left_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_1_Left_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_1_Left_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_1_Left_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_1_Left_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_1_Left_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_1_Left_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_1_Left_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_1_Left_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_1_Left_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_1_Left_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_1_Left_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_1_Left_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_1_Left_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_1_Left_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_1_Left_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_1_Left_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_1_Left_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_1_Left_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_1_Left_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_1_Left_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_1_Left_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_1_Left_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_1_Left_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_1_Left_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_1_Left_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_1_Left_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_1_Left_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_1_Left_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_1_Left_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_1_Left_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_1_Left_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_1_Left_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_1_Left_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_1_Left_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_1_Left_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_1_Left_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_1_Left_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_1_Left_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_1_Left_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_1_Left_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_1_Left_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_1_Left_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_1_Left_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_1_Left_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_1_Left_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_1_Left_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_1_Left_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_1_Left_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_1_Left_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_1_Left_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_1_Left_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_1_Left_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_1_Left_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_1_Left_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_1_Left_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_1_Left_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_1_Left_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_1_Left_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_1_Left_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_1_Left_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_1_Left_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_1_Left_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_1_Left_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_1_Left_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_1_Left_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_1_Left_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_1_Left_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_1_Left_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_1_Left_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_1_Left_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_1_Left_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_1_Left_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_1_Left_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_1_Left_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_1_Left_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_1_Left_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_1_Left_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_1_Left_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_1_Left_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_1_Left_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_1_Left_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_1_Left_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_1_Left_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_1_Left_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_1_Left_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_1_Left_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_1_Left_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_1_Left_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_1_Left_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_1_Left_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Left_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Left_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Left_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Left_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Left_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Left_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Left_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Left_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Left_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Left_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Left_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Left_265 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Left_266 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Left_267 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Left_268 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Left_269 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Left_270 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Left_271 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Left_272 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Left_273 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Left_274 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_1_Left_275 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_2_Left_276 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_2_Left_277 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_2_Left_278 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_2_Left_279 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_2_Left_280 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_2_Left_281 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_2_Left_282 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_2_Left_283 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_2_Left_284 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_2_Left_285 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_2_Left_286 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_2_Left_287 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_2_Left_288 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_2_Left_289 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_2_Left_290 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_2_Left_291 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_2_Left_292 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_2_Left_293 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_2_Left_294 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_2_Left_295 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_2_Left_296 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_2_Left_297 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_2_Left_298 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_2_Left_299 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_2_Left_300 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_2_Left_301 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_2_Left_302 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_2_Left_303 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_2_Left_304 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_2_Left_305 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_2_Left_306 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_2_Left_307 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_2_Left_308 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_2_Left_309 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_2_Left_310 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_2_Left_311 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_2_Left_312 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_2_Left_313 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_2_Left_314 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_2_Left_315 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_2_Left_316 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_2_Left_317 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_2_Left_318 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_2_Left_319 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_2_Left_320 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_2_Left_321 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_2_Left_322 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_2_Left_323 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_2_Left_324 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_2_Left_325 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_2_Left_326 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_2_Left_327 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_2_Left_328 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_2_Left_329 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_2_Left_330 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_2_Left_331 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_2_Left_332 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_2_Left_333 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_2_Left_334 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_2_Left_335 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_2_Left_336 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_2_Left_337 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_2_Left_338 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_2_Left_339 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_2_Left_340 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_2_Left_341 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_2_Left_342 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_2_Left_343 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_2_Left_344 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_2_Left_345 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_2_Left_346 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_2_Left_347 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_2_Left_348 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_2_Left_349 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_2_Left_350 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_2_Left_351 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_2_Left_352 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_2_Left_353 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_2_Left_354 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_2_Left_355 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_2_Left_356 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_2_Left_357 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_2_Left_358 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_2_Left_359 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_2_Left_360 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_2_Left_361 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_2_Left_362 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_2_Left_363 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_2_Left_364 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_2_Left_365 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_2_Left_366 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_2_Left_367 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_2_Left_368 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_2_Left_369 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_2_Left_370 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_2_Left_371 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_2_Left_372 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_2_Left_373 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_2_Left_374 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_2_Left_375 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_2_Left_376 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_2_Left_377 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_2_Left_378 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_2_Left_379 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_2_Left_380 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_1_Right_381 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_1_Right_382 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_1_Right_383 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_1_Right_384 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_1_Right_385 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_1_Right_386 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_1_Right_387 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_1_Right_388 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_1_Right_389 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_1_Right_390 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_1_Right_391 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_1_Right_392 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_1_Right_393 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_1_Right_394 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_1_Right_395 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_1_Right_396 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_1_Right_397 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_1_Right_398 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_1_Right_399 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_1_Right_400 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_1_Right_401 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_1_Right_402 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_1_Right_403 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_1_Right_404 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_1_Right_405 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_1_Right_406 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_1_Right_407 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_1_Right_408 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_1_Right_409 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_1_Right_410 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_1_Right_411 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_1_Right_412 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_1_Right_413 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_1_Right_414 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_1_Right_415 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_1_Right_416 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_1_Right_417 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_1_Right_418 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_1_Right_419 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_1_Right_420 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_1_Right_421 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_1_Right_422 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_1_Right_423 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_1_Right_424 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_1_Right_425 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_1_Right_426 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_1_Right_427 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_1_Right_428 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_1_Right_429 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_1_Right_430 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_1_Right_431 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_1_Right_432 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_1_Right_433 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_1_Right_434 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_1_Right_435 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_1_Right_436 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_1_Right_437 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_1_Right_438 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_1_Right_439 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_1_Right_440 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_1_Right_441 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_1_Right_442 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_1_Right_443 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_1_Right_444 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_1_Right_445 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_1_Right_446 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_1_Right_447 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_1_Right_448 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_1_Right_449 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_1_Right_450 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_1_Right_451 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_1_Right_452 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_1_Right_453 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_1_Right_454 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_1_Right_455 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_1_Right_456 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_1_Right_457 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_1_Right_458 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_1_Right_459 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_1_Right_460 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_1_Right_461 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_1_Right_462 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_1_Right_463 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_1_Right_464 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_1_Right_465 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_1_Right_466 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_1_Right_467 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_1_Right_468 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_1_Right_469 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_1_Right_470 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_1_Right_471 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_1_Right_472 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_1_Right_473 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_1_Right_474 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_1_Right_475 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_1_Right_476 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_1_Right_477 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_1_Right_478 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_1_Right_479 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_1_Right_480 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_1_Right_481 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_1_Right_482 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_1_Right_483 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_1_Right_484 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_1_Right_485 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_486 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_487 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_488 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_489 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_490 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_491 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_492 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_117_493 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_494 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_495 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_496 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_497 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_498 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_499 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_500 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_501 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_502 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_503 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_137_504 ();
 LOGIC0_X1 \u_multiplier/STAGE2/E_4_2_pp_16_1/_18__60  (.Z(net60));
 LOGIC0_X1 \u_multiplier/STAGE3/E_4_2_pp_16_1/_18__64  (.Z(net64));
 CLKBUF_X1 hold77 (.A(net137),
    .Z(net77));
 BUF_X1 input1 (.A(data_in[0]),
    .Z(net1));
 CLKBUF_X2 input2 (.A(data_in[10]),
    .Z(net2));
 BUF_X1 input3 (.A(data_in[11]),
    .Z(net3));
 CLKBUF_X2 input4 (.A(data_in[12]),
    .Z(net4));
 BUF_X1 input5 (.A(data_in[13]),
    .Z(net5));
 BUF_X2 input6 (.A(data_in[14]),
    .Z(net6));
 BUF_X1 input7 (.A(data_in[15]),
    .Z(net7));
 BUF_X2 input8 (.A(data_in[1]),
    .Z(net8));
 BUF_X1 input9 (.A(data_in[2]),
    .Z(net9));
 BUF_X2 input10 (.A(data_in[3]),
    .Z(net10));
 BUF_X1 input11 (.A(data_in[4]),
    .Z(net11));
 BUF_X1 input12 (.A(data_in[5]),
    .Z(net12));
 BUF_X1 input13 (.A(data_in[6]),
    .Z(net13));
 BUF_X1 input14 (.A(data_in[7]),
    .Z(net14));
 BUF_X2 input15 (.A(data_in[8]),
    .Z(net15));
 BUF_X1 input16 (.A(data_in[9]),
    .Z(net16));
 BUF_X2 input17 (.A(init_enable),
    .Z(net17));
 BUF_X2 input18 (.A(pe_ce),
    .Z(net18));
 BUF_X8 input19 (.A(rst_n),
    .Z(net19));
 BUF_X1 output20 (.A(net20),
    .Z(curr_state[1]));
 BUF_X1 output21 (.A(net21),
    .Z(data_out[0]));
 BUF_X1 output22 (.A(net22),
    .Z(data_out[10]));
 BUF_X1 output23 (.A(net23),
    .Z(data_out[11]));
 BUF_X1 output24 (.A(net24),
    .Z(data_out[12]));
 BUF_X1 output25 (.A(net25),
    .Z(data_out[13]));
 BUF_X1 output26 (.A(net26),
    .Z(data_out[14]));
 BUF_X1 output27 (.A(net27),
    .Z(data_out[15]));
 BUF_X1 output28 (.A(net28),
    .Z(data_out[16]));
 BUF_X1 output29 (.A(net29),
    .Z(data_out[17]));
 BUF_X1 output30 (.A(net30),
    .Z(data_out[18]));
 BUF_X1 output31 (.A(net31),
    .Z(data_out[19]));
 BUF_X1 output32 (.A(net32),
    .Z(data_out[1]));
 BUF_X1 output33 (.A(net33),
    .Z(data_out[20]));
 BUF_X1 output34 (.A(net34),
    .Z(data_out[21]));
 BUF_X1 output35 (.A(net35),
    .Z(data_out[22]));
 BUF_X1 output36 (.A(net36),
    .Z(data_out[23]));
 BUF_X1 output37 (.A(net37),
    .Z(data_out[24]));
 BUF_X1 output38 (.A(net38),
    .Z(data_out[25]));
 BUF_X1 output39 (.A(net39),
    .Z(data_out[26]));
 BUF_X1 output40 (.A(net40),
    .Z(data_out[27]));
 BUF_X1 output41 (.A(net41),
    .Z(data_out[28]));
 BUF_X1 output42 (.A(net42),
    .Z(data_out[29]));
 BUF_X1 output43 (.A(net43),
    .Z(data_out[2]));
 BUF_X1 output44 (.A(net44),
    .Z(data_out[30]));
 BUF_X1 output45 (.A(net45),
    .Z(data_out[31]));
 BUF_X1 output46 (.A(net46),
    .Z(data_out[3]));
 BUF_X1 output47 (.A(net47),
    .Z(data_out[4]));
 BUF_X1 output48 (.A(net48),
    .Z(data_out[5]));
 BUF_X1 output49 (.A(net49),
    .Z(data_out[6]));
 BUF_X1 output50 (.A(net50),
    .Z(data_out[7]));
 BUF_X1 output51 (.A(net51),
    .Z(data_out[8]));
 BUF_X1 output52 (.A(net52),
    .Z(data_out[9]));
 BUF_X1 output53 (.A(net53),
    .Z(valid_reg_out));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_16_1/_18__54  (.Z(net54));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_16_1/_25__55  (.Z(net55));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_16_2/_18__56  (.Z(net56));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_16_2/_25__57  (.Z(net57));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_16_3/_18__58  (.Z(net58));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_16_3/_25__59  (.Z(net59));
 LOGIC0_X1 \u_multiplier/STAGE2/E_4_2_pp_16_1/_25__61  (.Z(net61));
 LOGIC0_X1 \u_multiplier/STAGE2/E_4_2_pp_16_2/_18__62  (.Z(net62));
 LOGIC0_X1 \u_multiplier/STAGE2/E_4_2_pp_16_2/_25__63  (.Z(net63));
 LOGIC0_X1 \u_multiplier/STAGE3/E_4_2_pp_16_1/_25__65  (.Z(net65));
 LOGIC0_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_43__66  (.Z(net66));
 LOGIC0_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_44__67  (.Z(net67));
 LOGIC0_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_45__68  (.Z(net68));
 LOGIC0_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_46__69  (.Z(net69));
 LOGIC0_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_56__70  (.Z(net70));
 LOGIC0_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_40__71  (.Z(net71));
 LOGIC0_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_40__72  (.Z(net72));
 LOGIC0_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_53__73  (.Z(net73));
 LOGIC0_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_53__74  (.Z(net74));
 LOGIC0_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_54__75  (.Z(net75));
 LOGIC0_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_54__76  (.Z(net76));
 CLKBUF_X1 hold78 (.A(_173_),
    .Z(net78));
 CLKBUF_X1 hold79 (.A(net142),
    .Z(net79));
 CLKBUF_X1 hold80 (.A(_192_),
    .Z(net80));
 CLKBUF_X1 hold81 (.A(net93),
    .Z(net81));
 CLKBUF_X1 hold82 (.A(net101),
    .Z(net82));
 CLKBUF_X1 hold83 (.A(net98),
    .Z(net83));
 CLKBUF_X1 hold84 (.A(net108),
    .Z(net84));
 CLKBUF_X1 hold85 (.A(net115),
    .Z(net85));
 CLKBUF_X1 hold86 (.A(net112),
    .Z(net86));
 CLKBUF_X1 hold87 (.A(net126),
    .Z(net87));
 CLKBUF_X1 hold88 (.A(net128),
    .Z(net88));
 CLKBUF_X1 hold89 (.A(net130),
    .Z(net89));
 CLKBUF_X1 hold90 (.A(net123),
    .Z(net90));
 CLKBUF_X1 hold91 (.A(net139),
    .Z(net91));
 CLKBUF_X1 hold92 (.A(net140),
    .Z(net92));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_2_0_0_clk));
 CLKBUF_X3 clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_2_1_0_clk));
 CLKBUF_X3 clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .Z(clknet_2_2_0_clk));
 CLKBUF_X3 clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .Z(clknet_2_3_0_clk));
 CLKBUF_X3 clkbuf_3_0_0_clk (.A(clknet_2_0_0_clk),
    .Z(clknet_3_0_0_clk));
 CLKBUF_X3 clkbuf_3_1_0_clk (.A(clknet_2_0_0_clk),
    .Z(clknet_3_1_0_clk));
 CLKBUF_X3 clkbuf_3_2_0_clk (.A(clknet_2_1_0_clk),
    .Z(clknet_3_2_0_clk));
 CLKBUF_X3 clkbuf_3_3_0_clk (.A(clknet_2_1_0_clk),
    .Z(clknet_3_3_0_clk));
 CLKBUF_X3 clkbuf_3_4_0_clk (.A(clknet_2_2_0_clk),
    .Z(clknet_3_4_0_clk));
 CLKBUF_X3 clkbuf_3_5_0_clk (.A(clknet_2_2_0_clk),
    .Z(clknet_3_5_0_clk));
 CLKBUF_X3 clkbuf_3_6_0_clk (.A(clknet_2_3_0_clk),
    .Z(clknet_3_6_0_clk));
 CLKBUF_X3 clkbuf_3_7_0_clk (.A(clknet_2_3_0_clk),
    .Z(clknet_3_7_0_clk));
 INV_X2 clkload0 (.A(clknet_3_0_0_clk));
 INV_X2 clkload1 (.A(clknet_3_3_0_clk));
 INV_X2 clkload2 (.A(clknet_3_4_0_clk));
 INV_X1 clkload3 (.A(clknet_3_6_0_clk));
 CLKBUF_X1 hold1 (.A(_400_),
    .Z(net93));
 CLKBUF_X1 hold2 (.A(net81),
    .Z(net94));
 CLKBUF_X1 hold3 (.A(_118_),
    .Z(net95));
 CLKBUF_X1 hold4 (.A(_403_),
    .Z(net96));
 CLKBUF_X1 hold5 (.A(_280_),
    .Z(net97));
 CLKBUF_X1 hold6 (.A(_405_),
    .Z(net98));
 CLKBUF_X1 hold7 (.A(net83),
    .Z(net99));
 CLKBUF_X1 hold8 (.A(_171_),
    .Z(net100));
 CLKBUF_X1 hold9 (.A(_406_),
    .Z(net101));
 CLKBUF_X1 hold10 (.A(net82),
    .Z(net102));
 CLKBUF_X1 hold11 (.A(_172_),
    .Z(net103));
 CLKBUF_X1 hold12 (.A(net147),
    .Z(net104));
 CLKBUF_X1 hold13 (.A(curr_state[0]),
    .Z(net105));
 CLKBUF_X1 hold14 (.A(_251_),
    .Z(net106));
 CLKBUF_X1 hold15 (.A(_194_),
    .Z(net107));
 CLKBUF_X1 hold16 (.A(_399_),
    .Z(net108));
 CLKBUF_X1 hold17 (.A(net84),
    .Z(net109));
 CLKBUF_X1 hold18 (.A(_117_),
    .Z(net110));
 CLKBUF_X1 hold19 (.A(net146),
    .Z(net111));
 CLKBUF_X1 hold20 (.A(_401_),
    .Z(net112));
 CLKBUF_X1 hold21 (.A(net86),
    .Z(net113));
 CLKBUF_X1 hold22 (.A(data_in_reg[1]),
    .Z(net114));
 CLKBUF_X1 hold23 (.A(_404_),
    .Z(net115));
 CLKBUF_X1 hold24 (.A(net85),
    .Z(net116));
 CLKBUF_X1 hold25 (.A(_170_),
    .Z(net117));
 CLKBUF_X1 hold26 (.A(data_in_reg[12]),
    .Z(net118));
 CLKBUF_X1 hold27 (.A(data_in_reg[5]),
    .Z(net119));
 CLKBUF_X1 hold28 (.A(data_in_reg[10]),
    .Z(net120));
 CLKBUF_X1 hold29 (.A(data_in_reg[11]),
    .Z(net121));
 CLKBUF_X1 hold30 (.A(data_in_reg[15]),
    .Z(net122));
 CLKBUF_X1 hold31 (.A(_408_),
    .Z(net123));
 CLKBUF_X1 hold32 (.A(net90),
    .Z(net124));
 CLKBUF_X1 hold33 (.A(_174_),
    .Z(net125));
 CLKBUF_X1 hold34 (.A(addr_ptr[4]),
    .Z(net126));
 CLKBUF_X1 hold35 (.A(net87),
    .Z(net127));
 CLKBUF_X1 hold36 (.A(addr_ptr[1]),
    .Z(net128));
 CLKBUF_X1 hold37 (.A(net88),
    .Z(net129));
 CLKBUF_X1 hold38 (.A(addr_ptr[2]),
    .Z(net130));
 CLKBUF_X1 hold39 (.A(data_in_reg[4]),
    .Z(net131));
 CLKBUF_X1 hold40 (.A(_402_),
    .Z(net132));
 CLKBUF_X1 hold41 (.A(_278_),
    .Z(net133));
 CLKBUF_X1 hold42 (.A(data_in_reg[3]),
    .Z(net134));
 CLKBUF_X1 hold43 (.A(data_in_reg[2]),
    .Z(net135));
 CLKBUF_X1 hold44 (.A(data_in_reg[8]),
    .Z(net136));
 CLKBUF_X1 hold45 (.A(_407_),
    .Z(net137));
 CLKBUF_X1 hold46 (.A(data_in_reg[6]),
    .Z(net138));
 CLKBUF_X1 hold47 (.A(addr_ptr[3]),
    .Z(net139));
 CLKBUF_X1 hold48 (.A(addr_ptr[0]),
    .Z(net140));
 CLKBUF_X1 hold49 (.A(curr_state[2]),
    .Z(net141));
 CLKBUF_X1 hold50 (.A(_331_),
    .Z(net142));
 CLKBUF_X1 hold51 (.A(data_in_reg[9]),
    .Z(net143));
 CLKBUF_X1 hold52 (.A(data_in_reg[0]),
    .Z(net144));
 CLKBUF_X1 hold53 (.A(data_in_reg[7]),
    .Z(net145));
 CLKBUF_X1 hold54 (.A(data_in_reg[13]),
    .Z(net146));
 CLKBUF_X1 hold55 (.A(data_in_reg[14]),
    .Z(net147));
 FILLCELL_X4 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_8 ();
 FILLCELL_X16 FILLER_0_40 ();
 FILLCELL_X32 FILLER_0_59 ();
 FILLCELL_X32 FILLER_0_91 ();
 FILLCELL_X8 FILLER_0_123 ();
 FILLCELL_X2 FILLER_0_131 ();
 FILLCELL_X32 FILLER_0_136 ();
 FILLCELL_X32 FILLER_0_168 ();
 FILLCELL_X8 FILLER_0_200 ();
 FILLCELL_X4 FILLER_0_208 ();
 FILLCELL_X2 FILLER_0_212 ();
 FILLCELL_X1 FILLER_0_214 ();
 FILLCELL_X32 FILLER_0_219 ();
 FILLCELL_X32 FILLER_0_251 ();
 FILLCELL_X8 FILLER_0_283 ();
 FILLCELL_X1 FILLER_0_291 ();
 FILLCELL_X32 FILLER_0_295 ();
 FILLCELL_X32 FILLER_0_327 ();
 FILLCELL_X8 FILLER_0_359 ();
 FILLCELL_X4 FILLER_0_367 ();
 FILLCELL_X2 FILLER_0_371 ();
 FILLCELL_X1 FILLER_0_373 ();
 FILLCELL_X32 FILLER_0_377 ();
 FILLCELL_X32 FILLER_0_409 ();
 FILLCELL_X8 FILLER_0_441 ();
 FILLCELL_X2 FILLER_0_449 ();
 FILLCELL_X32 FILLER_0_454 ();
 FILLCELL_X32 FILLER_0_486 ();
 FILLCELL_X8 FILLER_0_518 ();
 FILLCELL_X2 FILLER_0_526 ();
 FILLCELL_X32 FILLER_0_531 ();
 FILLCELL_X32 FILLER_0_563 ();
 FILLCELL_X8 FILLER_0_595 ();
 FILLCELL_X4 FILLER_0_603 ();
 FILLCELL_X2 FILLER_0_607 ();
 FILLCELL_X1 FILLER_0_609 ();
 FILLCELL_X16 FILLER_0_613 ();
 FILLCELL_X2 FILLER_0_629 ();
 FILLCELL_X32 FILLER_0_632 ();
 FILLCELL_X16 FILLER_0_664 ();
 FILLCELL_X4 FILLER_0_680 ();
 FILLCELL_X2 FILLER_0_684 ();
 FILLCELL_X1 FILLER_0_686 ();
 FILLCELL_X32 FILLER_0_691 ();
 FILLCELL_X32 FILLER_0_723 ();
 FILLCELL_X8 FILLER_0_755 ();
 FILLCELL_X4 FILLER_0_763 ();
 FILLCELL_X2 FILLER_0_767 ();
 FILLCELL_X32 FILLER_0_772 ();
 FILLCELL_X32 FILLER_0_804 ();
 FILLCELL_X8 FILLER_0_836 ();
 FILLCELL_X2 FILLER_0_844 ();
 FILLCELL_X16 FILLER_0_849 ();
 FILLCELL_X8 FILLER_0_865 ();
 FILLCELL_X4 FILLER_0_873 ();
 FILLCELL_X2 FILLER_0_877 ();
 FILLCELL_X4 FILLER_0_882 ();
 FILLCELL_X16 FILLER_0_889 ();
 FILLCELL_X4 FILLER_0_905 ();
 FILLCELL_X2 FILLER_0_909 ();
 FILLCELL_X1 FILLER_0_911 ();
 FILLCELL_X4 FILLER_0_916 ();
 FILLCELL_X2 FILLER_0_920 ();
 FILLCELL_X1 FILLER_0_922 ();
 FILLCELL_X32 FILLER_0_926 ();
 FILLCELL_X32 FILLER_0_958 ();
 FILLCELL_X8 FILLER_0_990 ();
 FILLCELL_X4 FILLER_0_998 ();
 FILLCELL_X2 FILLER_0_1002 ();
 FILLCELL_X1 FILLER_0_1004 ();
 FILLCELL_X8 FILLER_0_1008 ();
 FILLCELL_X4 FILLER_0_1016 ();
 FILLCELL_X2 FILLER_0_1020 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X32 FILLER_1_257 ();
 FILLCELL_X32 FILLER_1_289 ();
 FILLCELL_X32 FILLER_1_321 ();
 FILLCELL_X32 FILLER_1_353 ();
 FILLCELL_X32 FILLER_1_385 ();
 FILLCELL_X32 FILLER_1_417 ();
 FILLCELL_X32 FILLER_1_449 ();
 FILLCELL_X32 FILLER_1_481 ();
 FILLCELL_X32 FILLER_1_513 ();
 FILLCELL_X32 FILLER_1_545 ();
 FILLCELL_X32 FILLER_1_577 ();
 FILLCELL_X32 FILLER_1_609 ();
 FILLCELL_X32 FILLER_1_641 ();
 FILLCELL_X32 FILLER_1_673 ();
 FILLCELL_X32 FILLER_1_705 ();
 FILLCELL_X32 FILLER_1_737 ();
 FILLCELL_X32 FILLER_1_769 ();
 FILLCELL_X32 FILLER_1_801 ();
 FILLCELL_X8 FILLER_1_833 ();
 FILLCELL_X4 FILLER_1_841 ();
 FILLCELL_X2 FILLER_1_845 ();
 FILLCELL_X1 FILLER_1_847 ();
 FILLCELL_X4 FILLER_1_855 ();
 FILLCELL_X8 FILLER_1_864 ();
 FILLCELL_X4 FILLER_1_872 ();
 FILLCELL_X4 FILLER_1_885 ();
 FILLCELL_X4 FILLER_1_898 ();
 FILLCELL_X2 FILLER_1_902 ();
 FILLCELL_X4 FILLER_1_910 ();
 FILLCELL_X16 FILLER_1_933 ();
 FILLCELL_X2 FILLER_1_949 ();
 FILLCELL_X1 FILLER_1_951 ();
 FILLCELL_X32 FILLER_1_971 ();
 FILLCELL_X16 FILLER_1_1003 ();
 FILLCELL_X2 FILLER_1_1019 ();
 FILLCELL_X1 FILLER_1_1021 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X32 FILLER_2_289 ();
 FILLCELL_X32 FILLER_2_321 ();
 FILLCELL_X32 FILLER_2_353 ();
 FILLCELL_X32 FILLER_2_385 ();
 FILLCELL_X32 FILLER_2_417 ();
 FILLCELL_X32 FILLER_2_449 ();
 FILLCELL_X32 FILLER_2_481 ();
 FILLCELL_X32 FILLER_2_513 ();
 FILLCELL_X32 FILLER_2_545 ();
 FILLCELL_X32 FILLER_2_577 ();
 FILLCELL_X16 FILLER_2_609 ();
 FILLCELL_X4 FILLER_2_625 ();
 FILLCELL_X2 FILLER_2_629 ();
 FILLCELL_X32 FILLER_2_632 ();
 FILLCELL_X32 FILLER_2_664 ();
 FILLCELL_X32 FILLER_2_696 ();
 FILLCELL_X32 FILLER_2_728 ();
 FILLCELL_X32 FILLER_2_760 ();
 FILLCELL_X32 FILLER_2_792 ();
 FILLCELL_X8 FILLER_2_824 ();
 FILLCELL_X4 FILLER_2_832 ();
 FILLCELL_X2 FILLER_2_836 ();
 FILLCELL_X1 FILLER_2_838 ();
 FILLCELL_X4 FILLER_2_843 ();
 FILLCELL_X4 FILLER_2_864 ();
 FILLCELL_X8 FILLER_2_870 ();
 FILLCELL_X1 FILLER_2_878 ();
 FILLCELL_X4 FILLER_2_889 ();
 FILLCELL_X4 FILLER_2_896 ();
 FILLCELL_X4 FILLER_2_906 ();
 FILLCELL_X4 FILLER_2_917 ();
 FILLCELL_X1 FILLER_2_921 ();
 FILLCELL_X8 FILLER_2_925 ();
 FILLCELL_X4 FILLER_2_933 ();
 FILLCELL_X8 FILLER_2_943 ();
 FILLCELL_X4 FILLER_2_951 ();
 FILLCELL_X4 FILLER_2_959 ();
 FILLCELL_X2 FILLER_2_963 ();
 FILLCELL_X16 FILLER_2_984 ();
 FILLCELL_X8 FILLER_2_1000 ();
 FILLCELL_X4 FILLER_2_1008 ();
 FILLCELL_X2 FILLER_2_1012 ();
 FILLCELL_X1 FILLER_2_1014 ();
 FILLCELL_X4 FILLER_2_1018 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X32 FILLER_3_289 ();
 FILLCELL_X32 FILLER_3_321 ();
 FILLCELL_X32 FILLER_3_353 ();
 FILLCELL_X32 FILLER_3_385 ();
 FILLCELL_X32 FILLER_3_417 ();
 FILLCELL_X32 FILLER_3_449 ();
 FILLCELL_X32 FILLER_3_481 ();
 FILLCELL_X32 FILLER_3_513 ();
 FILLCELL_X32 FILLER_3_545 ();
 FILLCELL_X32 FILLER_3_577 ();
 FILLCELL_X32 FILLER_3_609 ();
 FILLCELL_X32 FILLER_3_641 ();
 FILLCELL_X32 FILLER_3_673 ();
 FILLCELL_X32 FILLER_3_705 ();
 FILLCELL_X32 FILLER_3_737 ();
 FILLCELL_X32 FILLER_3_769 ();
 FILLCELL_X16 FILLER_3_801 ();
 FILLCELL_X8 FILLER_3_817 ();
 FILLCELL_X4 FILLER_3_825 ();
 FILLCELL_X1 FILLER_3_829 ();
 FILLCELL_X8 FILLER_3_833 ();
 FILLCELL_X4 FILLER_3_845 ();
 FILLCELL_X4 FILLER_3_854 ();
 FILLCELL_X8 FILLER_3_862 ();
 FILLCELL_X4 FILLER_3_870 ();
 FILLCELL_X1 FILLER_3_874 ();
 FILLCELL_X4 FILLER_3_879 ();
 FILLCELL_X8 FILLER_3_887 ();
 FILLCELL_X1 FILLER_3_895 ();
 FILLCELL_X4 FILLER_3_899 ();
 FILLCELL_X2 FILLER_3_903 ();
 FILLCELL_X8 FILLER_3_908 ();
 FILLCELL_X4 FILLER_3_920 ();
 FILLCELL_X4 FILLER_3_927 ();
 FILLCELL_X2 FILLER_3_931 ();
 FILLCELL_X1 FILLER_3_933 ();
 FILLCELL_X16 FILLER_3_940 ();
 FILLCELL_X8 FILLER_3_956 ();
 FILLCELL_X1 FILLER_3_964 ();
 FILLCELL_X32 FILLER_3_969 ();
 FILLCELL_X16 FILLER_3_1001 ();
 FILLCELL_X4 FILLER_3_1017 ();
 FILLCELL_X1 FILLER_3_1021 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X32 FILLER_4_289 ();
 FILLCELL_X32 FILLER_4_321 ();
 FILLCELL_X32 FILLER_4_353 ();
 FILLCELL_X32 FILLER_4_385 ();
 FILLCELL_X32 FILLER_4_417 ();
 FILLCELL_X32 FILLER_4_449 ();
 FILLCELL_X32 FILLER_4_481 ();
 FILLCELL_X32 FILLER_4_513 ();
 FILLCELL_X32 FILLER_4_545 ();
 FILLCELL_X32 FILLER_4_577 ();
 FILLCELL_X16 FILLER_4_609 ();
 FILLCELL_X4 FILLER_4_625 ();
 FILLCELL_X2 FILLER_4_629 ();
 FILLCELL_X32 FILLER_4_632 ();
 FILLCELL_X32 FILLER_4_664 ();
 FILLCELL_X32 FILLER_4_696 ();
 FILLCELL_X32 FILLER_4_728 ();
 FILLCELL_X32 FILLER_4_760 ();
 FILLCELL_X16 FILLER_4_792 ();
 FILLCELL_X8 FILLER_4_808 ();
 FILLCELL_X2 FILLER_4_816 ();
 FILLCELL_X1 FILLER_4_818 ();
 FILLCELL_X4 FILLER_4_822 ();
 FILLCELL_X4 FILLER_4_835 ();
 FILLCELL_X4 FILLER_4_842 ();
 FILLCELL_X2 FILLER_4_846 ();
 FILLCELL_X16 FILLER_4_852 ();
 FILLCELL_X4 FILLER_4_872 ();
 FILLCELL_X4 FILLER_4_886 ();
 FILLCELL_X4 FILLER_4_897 ();
 FILLCELL_X2 FILLER_4_901 ();
 FILLCELL_X1 FILLER_4_903 ();
 FILLCELL_X4 FILLER_4_914 ();
 FILLCELL_X8 FILLER_4_928 ();
 FILLCELL_X1 FILLER_4_936 ();
 FILLCELL_X4 FILLER_4_944 ();
 FILLCELL_X8 FILLER_4_952 ();
 FILLCELL_X4 FILLER_4_960 ();
 FILLCELL_X1 FILLER_4_964 ();
 FILLCELL_X4 FILLER_4_971 ();
 FILLCELL_X32 FILLER_4_979 ();
 FILLCELL_X8 FILLER_4_1011 ();
 FILLCELL_X2 FILLER_4_1019 ();
 FILLCELL_X1 FILLER_4_1021 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X32 FILLER_5_257 ();
 FILLCELL_X32 FILLER_5_289 ();
 FILLCELL_X32 FILLER_5_321 ();
 FILLCELL_X32 FILLER_5_353 ();
 FILLCELL_X32 FILLER_5_385 ();
 FILLCELL_X32 FILLER_5_417 ();
 FILLCELL_X32 FILLER_5_449 ();
 FILLCELL_X32 FILLER_5_481 ();
 FILLCELL_X32 FILLER_5_513 ();
 FILLCELL_X32 FILLER_5_545 ();
 FILLCELL_X32 FILLER_5_577 ();
 FILLCELL_X32 FILLER_5_609 ();
 FILLCELL_X32 FILLER_5_641 ();
 FILLCELL_X32 FILLER_5_673 ();
 FILLCELL_X32 FILLER_5_705 ();
 FILLCELL_X32 FILLER_5_737 ();
 FILLCELL_X16 FILLER_5_769 ();
 FILLCELL_X8 FILLER_5_785 ();
 FILLCELL_X2 FILLER_5_793 ();
 FILLCELL_X1 FILLER_5_795 ();
 FILLCELL_X4 FILLER_5_800 ();
 FILLCELL_X4 FILLER_5_808 ();
 FILLCELL_X8 FILLER_5_815 ();
 FILLCELL_X2 FILLER_5_823 ();
 FILLCELL_X1 FILLER_5_825 ();
 FILLCELL_X8 FILLER_5_835 ();
 FILLCELL_X1 FILLER_5_843 ();
 FILLCELL_X4 FILLER_5_850 ();
 FILLCELL_X8 FILLER_5_858 ();
 FILLCELL_X4 FILLER_5_866 ();
 FILLCELL_X1 FILLER_5_870 ();
 FILLCELL_X4 FILLER_5_873 ();
 FILLCELL_X2 FILLER_5_877 ();
 FILLCELL_X4 FILLER_5_886 ();
 FILLCELL_X8 FILLER_5_892 ();
 FILLCELL_X8 FILLER_5_902 ();
 FILLCELL_X2 FILLER_5_910 ();
 FILLCELL_X1 FILLER_5_912 ();
 FILLCELL_X4 FILLER_5_922 ();
 FILLCELL_X4 FILLER_5_929 ();
 FILLCELL_X2 FILLER_5_933 ();
 FILLCELL_X4 FILLER_5_939 ();
 FILLCELL_X4 FILLER_5_953 ();
 FILLCELL_X4 FILLER_5_959 ();
 FILLCELL_X4 FILLER_5_965 ();
 FILLCELL_X4 FILLER_5_975 ();
 FILLCELL_X2 FILLER_5_979 ();
 FILLCELL_X32 FILLER_5_988 ();
 FILLCELL_X2 FILLER_5_1020 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X16 FILLER_6_225 ();
 FILLCELL_X8 FILLER_6_241 ();
 FILLCELL_X4 FILLER_6_249 ();
 FILLCELL_X2 FILLER_6_253 ();
 FILLCELL_X4 FILLER_6_274 ();
 FILLCELL_X32 FILLER_6_282 ();
 FILLCELL_X32 FILLER_6_314 ();
 FILLCELL_X32 FILLER_6_346 ();
 FILLCELL_X32 FILLER_6_378 ();
 FILLCELL_X32 FILLER_6_410 ();
 FILLCELL_X1 FILLER_6_442 ();
 FILLCELL_X4 FILLER_6_447 ();
 FILLCELL_X32 FILLER_6_470 ();
 FILLCELL_X32 FILLER_6_502 ();
 FILLCELL_X32 FILLER_6_534 ();
 FILLCELL_X32 FILLER_6_566 ();
 FILLCELL_X32 FILLER_6_598 ();
 FILLCELL_X1 FILLER_6_630 ();
 FILLCELL_X32 FILLER_6_632 ();
 FILLCELL_X32 FILLER_6_664 ();
 FILLCELL_X32 FILLER_6_696 ();
 FILLCELL_X32 FILLER_6_728 ();
 FILLCELL_X16 FILLER_6_760 ();
 FILLCELL_X8 FILLER_6_776 ();
 FILLCELL_X4 FILLER_6_784 ();
 FILLCELL_X2 FILLER_6_788 ();
 FILLCELL_X1 FILLER_6_790 ();
 FILLCELL_X4 FILLER_6_795 ();
 FILLCELL_X4 FILLER_6_808 ();
 FILLCELL_X4 FILLER_6_821 ();
 FILLCELL_X8 FILLER_6_828 ();
 FILLCELL_X1 FILLER_6_836 ();
 FILLCELL_X4 FILLER_6_847 ();
 FILLCELL_X1 FILLER_6_851 ();
 FILLCELL_X4 FILLER_6_859 ();
 FILLCELL_X4 FILLER_6_869 ();
 FILLCELL_X2 FILLER_6_873 ();
 FILLCELL_X4 FILLER_6_885 ();
 FILLCELL_X16 FILLER_6_892 ();
 FILLCELL_X8 FILLER_6_908 ();
 FILLCELL_X2 FILLER_6_916 ();
 FILLCELL_X4 FILLER_6_927 ();
 FILLCELL_X8 FILLER_6_934 ();
 FILLCELL_X1 FILLER_6_942 ();
 FILLCELL_X4 FILLER_6_949 ();
 FILLCELL_X4 FILLER_6_956 ();
 FILLCELL_X1 FILLER_6_960 ();
 FILLCELL_X8 FILLER_6_968 ();
 FILLCELL_X2 FILLER_6_976 ();
 FILLCELL_X1 FILLER_6_978 ();
 FILLCELL_X4 FILLER_6_989 ();
 FILLCELL_X4 FILLER_6_996 ();
 FILLCELL_X16 FILLER_6_1003 ();
 FILLCELL_X2 FILLER_6_1019 ();
 FILLCELL_X1 FILLER_6_1021 ();
 FILLCELL_X4 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_8 ();
 FILLCELL_X32 FILLER_7_40 ();
 FILLCELL_X32 FILLER_7_72 ();
 FILLCELL_X32 FILLER_7_104 ();
 FILLCELL_X32 FILLER_7_136 ();
 FILLCELL_X32 FILLER_7_168 ();
 FILLCELL_X32 FILLER_7_200 ();
 FILLCELL_X32 FILLER_7_232 ();
 FILLCELL_X32 FILLER_7_264 ();
 FILLCELL_X32 FILLER_7_296 ();
 FILLCELL_X32 FILLER_7_328 ();
 FILLCELL_X32 FILLER_7_360 ();
 FILLCELL_X16 FILLER_7_392 ();
 FILLCELL_X4 FILLER_7_427 ();
 FILLCELL_X2 FILLER_7_431 ();
 FILLCELL_X1 FILLER_7_433 ();
 FILLCELL_X8 FILLER_7_453 ();
 FILLCELL_X2 FILLER_7_461 ();
 FILLCELL_X32 FILLER_7_482 ();
 FILLCELL_X32 FILLER_7_514 ();
 FILLCELL_X32 FILLER_7_546 ();
 FILLCELL_X32 FILLER_7_578 ();
 FILLCELL_X32 FILLER_7_610 ();
 FILLCELL_X32 FILLER_7_642 ();
 FILLCELL_X32 FILLER_7_674 ();
 FILLCELL_X32 FILLER_7_706 ();
 FILLCELL_X32 FILLER_7_738 ();
 FILLCELL_X16 FILLER_7_770 ();
 FILLCELL_X8 FILLER_7_786 ();
 FILLCELL_X2 FILLER_7_794 ();
 FILLCELL_X4 FILLER_7_799 ();
 FILLCELL_X8 FILLER_7_806 ();
 FILLCELL_X2 FILLER_7_814 ();
 FILLCELL_X1 FILLER_7_816 ();
 FILLCELL_X16 FILLER_7_820 ();
 FILLCELL_X8 FILLER_7_836 ();
 FILLCELL_X4 FILLER_7_844 ();
 FILLCELL_X2 FILLER_7_848 ();
 FILLCELL_X1 FILLER_7_850 ();
 FILLCELL_X16 FILLER_7_855 ();
 FILLCELL_X4 FILLER_7_871 ();
 FILLCELL_X4 FILLER_7_884 ();
 FILLCELL_X4 FILLER_7_891 ();
 FILLCELL_X4 FILLER_7_898 ();
 FILLCELL_X1 FILLER_7_902 ();
 FILLCELL_X4 FILLER_7_905 ();
 FILLCELL_X16 FILLER_7_916 ();
 FILLCELL_X8 FILLER_7_942 ();
 FILLCELL_X4 FILLER_7_950 ();
 FILLCELL_X4 FILLER_7_961 ();
 FILLCELL_X4 FILLER_7_974 ();
 FILLCELL_X4 FILLER_7_985 ();
 FILLCELL_X16 FILLER_7_992 ();
 FILLCELL_X8 FILLER_7_1008 ();
 FILLCELL_X4 FILLER_7_1016 ();
 FILLCELL_X2 FILLER_7_1020 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X32 FILLER_8_225 ();
 FILLCELL_X32 FILLER_8_257 ();
 FILLCELL_X32 FILLER_8_289 ();
 FILLCELL_X32 FILLER_8_321 ();
 FILLCELL_X16 FILLER_8_353 ();
 FILLCELL_X8 FILLER_8_369 ();
 FILLCELL_X2 FILLER_8_377 ();
 FILLCELL_X4 FILLER_8_398 ();
 FILLCELL_X2 FILLER_8_402 ();
 FILLCELL_X4 FILLER_8_408 ();
 FILLCELL_X2 FILLER_8_412 ();
 FILLCELL_X8 FILLER_8_418 ();
 FILLCELL_X4 FILLER_8_426 ();
 FILLCELL_X16 FILLER_8_434 ();
 FILLCELL_X4 FILLER_8_450 ();
 FILLCELL_X16 FILLER_8_458 ();
 FILLCELL_X4 FILLER_8_474 ();
 FILLCELL_X2 FILLER_8_478 ();
 FILLCELL_X1 FILLER_8_480 ();
 FILLCELL_X4 FILLER_8_500 ();
 FILLCELL_X2 FILLER_8_504 ();
 FILLCELL_X32 FILLER_8_525 ();
 FILLCELL_X32 FILLER_8_557 ();
 FILLCELL_X32 FILLER_8_589 ();
 FILLCELL_X8 FILLER_8_621 ();
 FILLCELL_X2 FILLER_8_629 ();
 FILLCELL_X32 FILLER_8_632 ();
 FILLCELL_X32 FILLER_8_664 ();
 FILLCELL_X32 FILLER_8_696 ();
 FILLCELL_X32 FILLER_8_728 ();
 FILLCELL_X16 FILLER_8_760 ();
 FILLCELL_X8 FILLER_8_776 ();
 FILLCELL_X4 FILLER_8_788 ();
 FILLCELL_X4 FILLER_8_795 ();
 FILLCELL_X2 FILLER_8_799 ();
 FILLCELL_X4 FILLER_8_804 ();
 FILLCELL_X4 FILLER_8_810 ();
 FILLCELL_X4 FILLER_8_824 ();
 FILLCELL_X4 FILLER_8_835 ();
 FILLCELL_X1 FILLER_8_839 ();
 FILLCELL_X4 FILLER_8_843 ();
 FILLCELL_X4 FILLER_8_857 ();
 FILLCELL_X8 FILLER_8_868 ();
 FILLCELL_X4 FILLER_8_876 ();
 FILLCELL_X2 FILLER_8_880 ();
 FILLCELL_X1 FILLER_8_882 ();
 FILLCELL_X4 FILLER_8_892 ();
 FILLCELL_X2 FILLER_8_896 ();
 FILLCELL_X4 FILLER_8_908 ();
 FILLCELL_X8 FILLER_8_922 ();
 FILLCELL_X4 FILLER_8_930 ();
 FILLCELL_X2 FILLER_8_934 ();
 FILLCELL_X4 FILLER_8_938 ();
 FILLCELL_X8 FILLER_8_952 ();
 FILLCELL_X2 FILLER_8_960 ();
 FILLCELL_X1 FILLER_8_962 ();
 FILLCELL_X8 FILLER_8_973 ();
 FILLCELL_X1 FILLER_8_981 ();
 FILLCELL_X4 FILLER_8_986 ();
 FILLCELL_X16 FILLER_8_999 ();
 FILLCELL_X4 FILLER_8_1015 ();
 FILLCELL_X2 FILLER_8_1019 ();
 FILLCELL_X1 FILLER_8_1021 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X32 FILLER_9_257 ();
 FILLCELL_X32 FILLER_9_289 ();
 FILLCELL_X32 FILLER_9_321 ();
 FILLCELL_X8 FILLER_9_353 ();
 FILLCELL_X2 FILLER_9_361 ();
 FILLCELL_X4 FILLER_9_382 ();
 FILLCELL_X4 FILLER_9_390 ();
 FILLCELL_X2 FILLER_9_394 ();
 FILLCELL_X1 FILLER_9_396 ();
 FILLCELL_X4 FILLER_9_416 ();
 FILLCELL_X2 FILLER_9_420 ();
 FILLCELL_X1 FILLER_9_422 ();
 FILLCELL_X8 FILLER_9_442 ();
 FILLCELL_X4 FILLER_9_450 ();
 FILLCELL_X1 FILLER_9_454 ();
 FILLCELL_X8 FILLER_9_474 ();
 FILLCELL_X2 FILLER_9_482 ();
 FILLCELL_X4 FILLER_9_503 ();
 FILLCELL_X1 FILLER_9_507 ();
 FILLCELL_X8 FILLER_9_527 ();
 FILLCELL_X32 FILLER_9_538 ();
 FILLCELL_X32 FILLER_9_570 ();
 FILLCELL_X32 FILLER_9_602 ();
 FILLCELL_X32 FILLER_9_634 ();
 FILLCELL_X32 FILLER_9_666 ();
 FILLCELL_X32 FILLER_9_698 ();
 FILLCELL_X32 FILLER_9_730 ();
 FILLCELL_X8 FILLER_9_762 ();
 FILLCELL_X4 FILLER_9_770 ();
 FILLCELL_X2 FILLER_9_774 ();
 FILLCELL_X4 FILLER_9_780 ();
 FILLCELL_X4 FILLER_9_793 ();
 FILLCELL_X4 FILLER_9_801 ();
 FILLCELL_X2 FILLER_9_805 ();
 FILLCELL_X1 FILLER_9_807 ();
 FILLCELL_X4 FILLER_9_812 ();
 FILLCELL_X16 FILLER_9_826 ();
 FILLCELL_X8 FILLER_9_842 ();
 FILLCELL_X4 FILLER_9_854 ();
 FILLCELL_X16 FILLER_9_860 ();
 FILLCELL_X1 FILLER_9_876 ();
 FILLCELL_X4 FILLER_9_884 ();
 FILLCELL_X1 FILLER_9_888 ();
 FILLCELL_X16 FILLER_9_892 ();
 FILLCELL_X4 FILLER_9_911 ();
 FILLCELL_X1 FILLER_9_915 ();
 FILLCELL_X4 FILLER_9_925 ();
 FILLCELL_X4 FILLER_9_931 ();
 FILLCELL_X2 FILLER_9_935 ();
 FILLCELL_X8 FILLER_9_941 ();
 FILLCELL_X2 FILLER_9_949 ();
 FILLCELL_X4 FILLER_9_954 ();
 FILLCELL_X4 FILLER_9_961 ();
 FILLCELL_X2 FILLER_9_965 ();
 FILLCELL_X1 FILLER_9_967 ();
 FILLCELL_X4 FILLER_9_971 ();
 FILLCELL_X8 FILLER_9_978 ();
 FILLCELL_X4 FILLER_9_986 ();
 FILLCELL_X2 FILLER_9_990 ();
 FILLCELL_X4 FILLER_9_995 ();
 FILLCELL_X16 FILLER_9_1002 ();
 FILLCELL_X4 FILLER_9_1018 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X32 FILLER_10_257 ();
 FILLCELL_X32 FILLER_10_289 ();
 FILLCELL_X16 FILLER_10_321 ();
 FILLCELL_X8 FILLER_10_337 ();
 FILLCELL_X1 FILLER_10_345 ();
 FILLCELL_X4 FILLER_10_349 ();
 FILLCELL_X2 FILLER_10_353 ();
 FILLCELL_X1 FILLER_10_355 ();
 FILLCELL_X16 FILLER_10_375 ();
 FILLCELL_X8 FILLER_10_410 ();
 FILLCELL_X2 FILLER_10_418 ();
 FILLCELL_X4 FILLER_10_439 ();
 FILLCELL_X1 FILLER_10_443 ();
 FILLCELL_X4 FILLER_10_448 ();
 FILLCELL_X4 FILLER_10_471 ();
 FILLCELL_X32 FILLER_10_479 ();
 FILLCELL_X32 FILLER_10_511 ();
 FILLCELL_X32 FILLER_10_543 ();
 FILLCELL_X16 FILLER_10_575 ();
 FILLCELL_X8 FILLER_10_591 ();
 FILLCELL_X2 FILLER_10_599 ();
 FILLCELL_X16 FILLER_10_604 ();
 FILLCELL_X8 FILLER_10_620 ();
 FILLCELL_X2 FILLER_10_628 ();
 FILLCELL_X1 FILLER_10_630 ();
 FILLCELL_X16 FILLER_10_632 ();
 FILLCELL_X8 FILLER_10_648 ();
 FILLCELL_X4 FILLER_10_656 ();
 FILLCELL_X4 FILLER_10_664 ();
 FILLCELL_X16 FILLER_10_687 ();
 FILLCELL_X8 FILLER_10_703 ();
 FILLCELL_X4 FILLER_10_711 ();
 FILLCELL_X2 FILLER_10_715 ();
 FILLCELL_X4 FILLER_10_720 ();
 FILLCELL_X1 FILLER_10_724 ();
 FILLCELL_X32 FILLER_10_728 ();
 FILLCELL_X16 FILLER_10_760 ();
 FILLCELL_X8 FILLER_10_776 ();
 FILLCELL_X4 FILLER_10_784 ();
 FILLCELL_X2 FILLER_10_788 ();
 FILLCELL_X1 FILLER_10_790 ();
 FILLCELL_X16 FILLER_10_800 ();
 FILLCELL_X2 FILLER_10_816 ();
 FILLCELL_X8 FILLER_10_821 ();
 FILLCELL_X2 FILLER_10_829 ();
 FILLCELL_X1 FILLER_10_831 ();
 FILLCELL_X4 FILLER_10_836 ();
 FILLCELL_X4 FILLER_10_843 ();
 FILLCELL_X4 FILLER_10_857 ();
 FILLCELL_X2 FILLER_10_861 ();
 FILLCELL_X1 FILLER_10_863 ();
 FILLCELL_X4 FILLER_10_868 ();
 FILLCELL_X4 FILLER_10_882 ();
 FILLCELL_X4 FILLER_10_895 ();
 FILLCELL_X4 FILLER_10_902 ();
 FILLCELL_X4 FILLER_10_909 ();
 FILLCELL_X2 FILLER_10_913 ();
 FILLCELL_X4 FILLER_10_918 ();
 FILLCELL_X4 FILLER_10_932 ();
 FILLCELL_X2 FILLER_10_936 ();
 FILLCELL_X1 FILLER_10_938 ();
 FILLCELL_X4 FILLER_10_949 ();
 FILLCELL_X4 FILLER_10_956 ();
 FILLCELL_X2 FILLER_10_960 ();
 FILLCELL_X1 FILLER_10_962 ();
 FILLCELL_X8 FILLER_10_972 ();
 FILLCELL_X2 FILLER_10_980 ();
 FILLCELL_X1 FILLER_10_982 ();
 FILLCELL_X4 FILLER_10_987 ();
 FILLCELL_X4 FILLER_10_1000 ();
 FILLCELL_X8 FILLER_10_1007 ();
 FILLCELL_X4 FILLER_10_1015 ();
 FILLCELL_X2 FILLER_10_1019 ();
 FILLCELL_X1 FILLER_10_1021 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_11_193 ();
 FILLCELL_X32 FILLER_11_225 ();
 FILLCELL_X32 FILLER_11_257 ();
 FILLCELL_X32 FILLER_11_289 ();
 FILLCELL_X16 FILLER_11_321 ();
 FILLCELL_X8 FILLER_11_342 ();
 FILLCELL_X1 FILLER_11_350 ();
 FILLCELL_X4 FILLER_11_354 ();
 FILLCELL_X4 FILLER_11_362 ();
 FILLCELL_X4 FILLER_11_370 ();
 FILLCELL_X8 FILLER_11_377 ();
 FILLCELL_X2 FILLER_11_385 ();
 FILLCELL_X4 FILLER_11_391 ();
 FILLCELL_X8 FILLER_11_399 ();
 FILLCELL_X4 FILLER_11_407 ();
 FILLCELL_X4 FILLER_11_416 ();
 FILLCELL_X16 FILLER_11_424 ();
 FILLCELL_X2 FILLER_11_440 ();
 FILLCELL_X16 FILLER_11_446 ();
 FILLCELL_X4 FILLER_11_465 ();
 FILLCELL_X4 FILLER_11_473 ();
 FILLCELL_X8 FILLER_11_482 ();
 FILLCELL_X1 FILLER_11_490 ();
 FILLCELL_X4 FILLER_11_495 ();
 FILLCELL_X32 FILLER_11_503 ();
 FILLCELL_X32 FILLER_11_535 ();
 FILLCELL_X4 FILLER_11_567 ();
 FILLCELL_X2 FILLER_11_571 ();
 FILLCELL_X1 FILLER_11_573 ();
 FILLCELL_X32 FILLER_11_577 ();
 FILLCELL_X16 FILLER_11_609 ();
 FILLCELL_X4 FILLER_11_625 ();
 FILLCELL_X2 FILLER_11_629 ();
 FILLCELL_X16 FILLER_11_632 ();
 FILLCELL_X1 FILLER_11_648 ();
 FILLCELL_X32 FILLER_11_652 ();
 FILLCELL_X8 FILLER_11_684 ();
 FILLCELL_X2 FILLER_11_692 ();
 FILLCELL_X8 FILLER_11_697 ();
 FILLCELL_X2 FILLER_11_705 ();
 FILLCELL_X4 FILLER_11_711 ();
 FILLCELL_X16 FILLER_11_734 ();
 FILLCELL_X4 FILLER_11_754 ();
 FILLCELL_X16 FILLER_11_777 ();
 FILLCELL_X4 FILLER_11_793 ();
 FILLCELL_X1 FILLER_11_797 ();
 FILLCELL_X4 FILLER_11_802 ();
 FILLCELL_X8 FILLER_11_816 ();
 FILLCELL_X2 FILLER_11_824 ();
 FILLCELL_X4 FILLER_11_830 ();
 FILLCELL_X4 FILLER_11_843 ();
 FILLCELL_X4 FILLER_11_851 ();
 FILLCELL_X8 FILLER_11_858 ();
 FILLCELL_X4 FILLER_11_868 ();
 FILLCELL_X4 FILLER_11_882 ();
 FILLCELL_X4 FILLER_11_889 ();
 FILLCELL_X2 FILLER_11_893 ();
 FILLCELL_X1 FILLER_11_895 ();
 FILLCELL_X4 FILLER_11_905 ();
 FILLCELL_X16 FILLER_11_912 ();
 FILLCELL_X8 FILLER_11_928 ();
 FILLCELL_X2 FILLER_11_936 ();
 FILLCELL_X8 FILLER_11_942 ();
 FILLCELL_X4 FILLER_11_950 ();
 FILLCELL_X2 FILLER_11_954 ();
 FILLCELL_X4 FILLER_11_960 ();
 FILLCELL_X4 FILLER_11_967 ();
 FILLCELL_X4 FILLER_11_974 ();
 FILLCELL_X8 FILLER_11_981 ();
 FILLCELL_X2 FILLER_11_989 ();
 FILLCELL_X8 FILLER_11_1001 ();
 FILLCELL_X8 FILLER_11_1011 ();
 FILLCELL_X2 FILLER_11_1019 ();
 FILLCELL_X1 FILLER_11_1021 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X8 FILLER_12_161 ();
 FILLCELL_X8 FILLER_12_819 ();
 FILLCELL_X4 FILLER_12_827 ();
 FILLCELL_X2 FILLER_12_831 ();
 FILLCELL_X1 FILLER_12_833 ();
 FILLCELL_X4 FILLER_12_837 ();
 FILLCELL_X8 FILLER_12_850 ();
 FILLCELL_X4 FILLER_12_862 ();
 FILLCELL_X16 FILLER_12_869 ();
 FILLCELL_X1 FILLER_12_885 ();
 FILLCELL_X8 FILLER_12_890 ();
 FILLCELL_X4 FILLER_12_902 ();
 FILLCELL_X8 FILLER_12_910 ();
 FILLCELL_X4 FILLER_12_918 ();
 FILLCELL_X4 FILLER_12_931 ();
 FILLCELL_X8 FILLER_12_938 ();
 FILLCELL_X4 FILLER_12_946 ();
 FILLCELL_X2 FILLER_12_950 ();
 FILLCELL_X1 FILLER_12_952 ();
 FILLCELL_X4 FILLER_12_962 ();
 FILLCELL_X4 FILLER_12_975 ();
 FILLCELL_X2 FILLER_12_979 ();
 FILLCELL_X4 FILLER_12_991 ();
 FILLCELL_X2 FILLER_12_995 ();
 FILLCELL_X8 FILLER_12_1007 ();
 FILLCELL_X4 FILLER_12_1018 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X8 FILLER_13_161 ();
 FILLCELL_X4 FILLER_13_819 ();
 FILLCELL_X4 FILLER_13_830 ();
 FILLCELL_X8 FILLER_13_836 ();
 FILLCELL_X4 FILLER_13_844 ();
 FILLCELL_X1 FILLER_13_848 ();
 FILLCELL_X4 FILLER_13_853 ();
 FILLCELL_X4 FILLER_13_866 ();
 FILLCELL_X8 FILLER_13_873 ();
 FILLCELL_X4 FILLER_13_881 ();
 FILLCELL_X2 FILLER_13_885 ();
 FILLCELL_X4 FILLER_13_890 ();
 FILLCELL_X16 FILLER_13_897 ();
 FILLCELL_X2 FILLER_13_913 ();
 FILLCELL_X1 FILLER_13_915 ();
 FILLCELL_X16 FILLER_13_923 ();
 FILLCELL_X8 FILLER_13_939 ();
 FILLCELL_X2 FILLER_13_947 ();
 FILLCELL_X1 FILLER_13_949 ();
 FILLCELL_X4 FILLER_13_954 ();
 FILLCELL_X4 FILLER_13_962 ();
 FILLCELL_X4 FILLER_13_969 ();
 FILLCELL_X2 FILLER_13_973 ();
 FILLCELL_X8 FILLER_13_978 ();
 FILLCELL_X4 FILLER_13_986 ();
 FILLCELL_X1 FILLER_13_990 ();
 FILLCELL_X4 FILLER_13_995 ();
 FILLCELL_X4 FILLER_13_1006 ();
 FILLCELL_X8 FILLER_13_1013 ();
 FILLCELL_X1 FILLER_13_1021 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X8 FILLER_14_161 ();
 FILLCELL_X8 FILLER_14_819 ();
 FILLCELL_X4 FILLER_14_837 ();
 FILLCELL_X4 FILLER_14_844 ();
 FILLCELL_X1 FILLER_14_848 ();
 FILLCELL_X4 FILLER_14_853 ();
 FILLCELL_X16 FILLER_14_866 ();
 FILLCELL_X4 FILLER_14_891 ();
 FILLCELL_X1 FILLER_14_895 ();
 FILLCELL_X8 FILLER_14_899 ();
 FILLCELL_X4 FILLER_14_911 ();
 FILLCELL_X4 FILLER_14_925 ();
 FILLCELL_X4 FILLER_14_938 ();
 FILLCELL_X4 FILLER_14_946 ();
 FILLCELL_X1 FILLER_14_950 ();
 FILLCELL_X16 FILLER_14_954 ();
 FILLCELL_X4 FILLER_14_970 ();
 FILLCELL_X1 FILLER_14_974 ();
 FILLCELL_X4 FILLER_14_977 ();
 FILLCELL_X4 FILLER_14_985 ();
 FILLCELL_X16 FILLER_14_998 ();
 FILLCELL_X8 FILLER_14_1014 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X8 FILLER_15_161 ();
 FILLCELL_X4 FILLER_15_819 ();
 FILLCELL_X2 FILLER_15_823 ();
 FILLCELL_X1 FILLER_15_825 ();
 FILLCELL_X4 FILLER_15_835 ();
 FILLCELL_X4 FILLER_15_842 ();
 FILLCELL_X8 FILLER_15_849 ();
 FILLCELL_X1 FILLER_15_857 ();
 FILLCELL_X4 FILLER_15_861 ();
 FILLCELL_X2 FILLER_15_865 ();
 FILLCELL_X1 FILLER_15_867 ();
 FILLCELL_X8 FILLER_15_871 ();
 FILLCELL_X2 FILLER_15_879 ();
 FILLCELL_X1 FILLER_15_881 ();
 FILLCELL_X4 FILLER_15_885 ();
 FILLCELL_X2 FILLER_15_889 ();
 FILLCELL_X4 FILLER_15_900 ();
 FILLCELL_X4 FILLER_15_914 ();
 FILLCELL_X1 FILLER_15_918 ();
 FILLCELL_X4 FILLER_15_922 ();
 FILLCELL_X4 FILLER_15_930 ();
 FILLCELL_X4 FILLER_15_943 ();
 FILLCELL_X4 FILLER_15_951 ();
 FILLCELL_X1 FILLER_15_955 ();
 FILLCELL_X4 FILLER_15_960 ();
 FILLCELL_X4 FILLER_15_968 ();
 FILLCELL_X8 FILLER_15_976 ();
 FILLCELL_X4 FILLER_15_984 ();
 FILLCELL_X1 FILLER_15_988 ();
 FILLCELL_X4 FILLER_15_992 ();
 FILLCELL_X2 FILLER_15_996 ();
 FILLCELL_X1 FILLER_15_998 ();
 FILLCELL_X4 FILLER_15_1018 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X8 FILLER_16_161 ();
 FILLCELL_X4 FILLER_16_819 ();
 FILLCELL_X2 FILLER_16_823 ();
 FILLCELL_X1 FILLER_16_825 ();
 FILLCELL_X16 FILLER_16_835 ();
 FILLCELL_X4 FILLER_16_851 ();
 FILLCELL_X2 FILLER_16_855 ();
 FILLCELL_X1 FILLER_16_857 ();
 FILLCELL_X4 FILLER_16_862 ();
 FILLCELL_X4 FILLER_16_876 ();
 FILLCELL_X4 FILLER_16_890 ();
 FILLCELL_X8 FILLER_16_901 ();
 FILLCELL_X2 FILLER_16_909 ();
 FILLCELL_X16 FILLER_16_913 ();
 FILLCELL_X4 FILLER_16_929 ();
 FILLCELL_X4 FILLER_16_936 ();
 FILLCELL_X4 FILLER_16_943 ();
 FILLCELL_X2 FILLER_16_947 ();
 FILLCELL_X1 FILLER_16_949 ();
 FILLCELL_X8 FILLER_16_954 ();
 FILLCELL_X4 FILLER_16_969 ();
 FILLCELL_X4 FILLER_16_978 ();
 FILLCELL_X2 FILLER_16_982 ();
 FILLCELL_X1 FILLER_16_984 ();
 FILLCELL_X8 FILLER_16_994 ();
 FILLCELL_X16 FILLER_16_1006 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X8 FILLER_17_161 ();
 FILLCELL_X8 FILLER_17_819 ();
 FILLCELL_X2 FILLER_17_827 ();
 FILLCELL_X4 FILLER_17_839 ();
 FILLCELL_X8 FILLER_17_846 ();
 FILLCELL_X4 FILLER_17_854 ();
 FILLCELL_X2 FILLER_17_858 ();
 FILLCELL_X4 FILLER_17_863 ();
 FILLCELL_X4 FILLER_17_871 ();
 FILLCELL_X4 FILLER_17_885 ();
 FILLCELL_X4 FILLER_17_891 ();
 FILLCELL_X1 FILLER_17_895 ();
 FILLCELL_X4 FILLER_17_899 ();
 FILLCELL_X4 FILLER_17_907 ();
 FILLCELL_X4 FILLER_17_915 ();
 FILLCELL_X4 FILLER_17_922 ();
 FILLCELL_X2 FILLER_17_926 ();
 FILLCELL_X16 FILLER_17_938 ();
 FILLCELL_X2 FILLER_17_954 ();
 FILLCELL_X4 FILLER_17_958 ();
 FILLCELL_X4 FILLER_17_979 ();
 FILLCELL_X4 FILLER_17_987 ();
 FILLCELL_X1 FILLER_17_991 ();
 FILLCELL_X4 FILLER_17_996 ();
 FILLCELL_X4 FILLER_17_1003 ();
 FILLCELL_X8 FILLER_17_1010 ();
 FILLCELL_X4 FILLER_17_1018 ();
 FILLCELL_X4 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_8 ();
 FILLCELL_X32 FILLER_18_40 ();
 FILLCELL_X32 FILLER_18_72 ();
 FILLCELL_X32 FILLER_18_104 ();
 FILLCELL_X32 FILLER_18_136 ();
 FILLCELL_X1 FILLER_18_168 ();
 FILLCELL_X4 FILLER_18_819 ();
 FILLCELL_X16 FILLER_18_827 ();
 FILLCELL_X4 FILLER_18_843 ();
 FILLCELL_X4 FILLER_18_856 ();
 FILLCELL_X4 FILLER_18_863 ();
 FILLCELL_X32 FILLER_18_870 ();
 FILLCELL_X1 FILLER_18_902 ();
 FILLCELL_X4 FILLER_18_912 ();
 FILLCELL_X4 FILLER_18_919 ();
 FILLCELL_X4 FILLER_18_927 ();
 FILLCELL_X1 FILLER_18_931 ();
 FILLCELL_X4 FILLER_18_935 ();
 FILLCELL_X8 FILLER_18_941 ();
 FILLCELL_X2 FILLER_18_949 ();
 FILLCELL_X4 FILLER_18_960 ();
 FILLCELL_X2 FILLER_18_964 ();
 FILLCELL_X16 FILLER_18_971 ();
 FILLCELL_X2 FILLER_18_987 ();
 FILLCELL_X4 FILLER_18_999 ();
 FILLCELL_X8 FILLER_18_1006 ();
 FILLCELL_X4 FILLER_18_1018 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X16 FILLER_19_129 ();
 FILLCELL_X8 FILLER_19_145 ();
 FILLCELL_X2 FILLER_19_153 ();
 FILLCELL_X1 FILLER_19_155 ();
 FILLCELL_X8 FILLER_19_160 ();
 FILLCELL_X1 FILLER_19_168 ();
 FILLCELL_X4 FILLER_19_819 ();
 FILLCELL_X2 FILLER_19_823 ();
 FILLCELL_X4 FILLER_19_829 ();
 FILLCELL_X2 FILLER_19_833 ();
 FILLCELL_X1 FILLER_19_835 ();
 FILLCELL_X4 FILLER_19_843 ();
 FILLCELL_X4 FILLER_19_857 ();
 FILLCELL_X8 FILLER_19_870 ();
 FILLCELL_X2 FILLER_19_878 ();
 FILLCELL_X16 FILLER_19_882 ();
 FILLCELL_X4 FILLER_19_898 ();
 FILLCELL_X2 FILLER_19_902 ();
 FILLCELL_X4 FILLER_19_913 ();
 FILLCELL_X8 FILLER_19_921 ();
 FILLCELL_X4 FILLER_19_939 ();
 FILLCELL_X8 FILLER_19_950 ();
 FILLCELL_X4 FILLER_19_961 ();
 FILLCELL_X16 FILLER_19_968 ();
 FILLCELL_X4 FILLER_19_984 ();
 FILLCELL_X2 FILLER_19_988 ();
 FILLCELL_X1 FILLER_19_990 ();
 FILLCELL_X8 FILLER_19_1000 ();
 FILLCELL_X8 FILLER_19_1014 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X16 FILLER_20_129 ();
 FILLCELL_X1 FILLER_20_145 ();
 FILLCELL_X4 FILLER_20_165 ();
 FILLCELL_X4 FILLER_20_819 ();
 FILLCELL_X4 FILLER_20_827 ();
 FILLCELL_X8 FILLER_20_835 ();
 FILLCELL_X4 FILLER_20_843 ();
 FILLCELL_X2 FILLER_20_847 ();
 FILLCELL_X4 FILLER_20_853 ();
 FILLCELL_X4 FILLER_20_860 ();
 FILLCELL_X2 FILLER_20_864 ();
 FILLCELL_X1 FILLER_20_866 ();
 FILLCELL_X4 FILLER_20_870 ();
 FILLCELL_X4 FILLER_20_884 ();
 FILLCELL_X4 FILLER_20_891 ();
 FILLCELL_X2 FILLER_20_895 ();
 FILLCELL_X4 FILLER_20_904 ();
 FILLCELL_X32 FILLER_20_911 ();
 FILLCELL_X4 FILLER_20_946 ();
 FILLCELL_X4 FILLER_20_959 ();
 FILLCELL_X1 FILLER_20_963 ();
 FILLCELL_X16 FILLER_20_974 ();
 FILLCELL_X2 FILLER_20_990 ();
 FILLCELL_X1 FILLER_20_992 ();
 FILLCELL_X4 FILLER_20_996 ();
 FILLCELL_X4 FILLER_20_1006 ();
 FILLCELL_X4 FILLER_20_1017 ();
 FILLCELL_X1 FILLER_20_1021 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X8 FILLER_21_161 ();
 FILLCELL_X4 FILLER_21_819 ();
 FILLCELL_X16 FILLER_21_842 ();
 FILLCELL_X4 FILLER_21_858 ();
 FILLCELL_X2 FILLER_21_862 ();
 FILLCELL_X4 FILLER_21_867 ();
 FILLCELL_X8 FILLER_21_880 ();
 FILLCELL_X1 FILLER_21_888 ();
 FILLCELL_X4 FILLER_21_899 ();
 FILLCELL_X4 FILLER_21_913 ();
 FILLCELL_X2 FILLER_21_917 ();
 FILLCELL_X1 FILLER_21_919 ();
 FILLCELL_X4 FILLER_21_924 ();
 FILLCELL_X4 FILLER_21_937 ();
 FILLCELL_X4 FILLER_21_944 ();
 FILLCELL_X8 FILLER_21_951 ();
 FILLCELL_X4 FILLER_21_961 ();
 FILLCELL_X4 FILLER_21_972 ();
 FILLCELL_X4 FILLER_21_985 ();
 FILLCELL_X4 FILLER_21_999 ();
 FILLCELL_X2 FILLER_21_1003 ();
 FILLCELL_X1 FILLER_21_1005 ();
 FILLCELL_X4 FILLER_21_1010 ();
 FILLCELL_X4 FILLER_21_1018 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X8 FILLER_22_161 ();
 FILLCELL_X4 FILLER_22_819 ();
 FILLCELL_X4 FILLER_22_832 ();
 FILLCELL_X4 FILLER_22_842 ();
 FILLCELL_X4 FILLER_22_856 ();
 FILLCELL_X4 FILLER_22_862 ();
 FILLCELL_X4 FILLER_22_875 ();
 FILLCELL_X4 FILLER_22_881 ();
 FILLCELL_X4 FILLER_22_888 ();
 FILLCELL_X8 FILLER_22_895 ();
 FILLCELL_X4 FILLER_22_907 ();
 FILLCELL_X4 FILLER_22_914 ();
 FILLCELL_X2 FILLER_22_918 ();
 FILLCELL_X1 FILLER_22_920 ();
 FILLCELL_X4 FILLER_22_925 ();
 FILLCELL_X8 FILLER_22_938 ();
 FILLCELL_X1 FILLER_22_946 ();
 FILLCELL_X8 FILLER_22_957 ();
 FILLCELL_X1 FILLER_22_965 ();
 FILLCELL_X4 FILLER_22_976 ();
 FILLCELL_X4 FILLER_22_983 ();
 FILLCELL_X4 FILLER_22_990 ();
 FILLCELL_X4 FILLER_22_996 ();
 FILLCELL_X4 FILLER_22_1003 ();
 FILLCELL_X8 FILLER_22_1013 ();
 FILLCELL_X1 FILLER_22_1021 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X8 FILLER_23_161 ();
 FILLCELL_X8 FILLER_23_819 ();
 FILLCELL_X2 FILLER_23_827 ();
 FILLCELL_X1 FILLER_23_829 ();
 FILLCELL_X4 FILLER_23_836 ();
 FILLCELL_X4 FILLER_23_847 ();
 FILLCELL_X16 FILLER_23_854 ();
 FILLCELL_X4 FILLER_23_870 ();
 FILLCELL_X1 FILLER_23_874 ();
 FILLCELL_X4 FILLER_23_879 ();
 FILLCELL_X4 FILLER_23_887 ();
 FILLCELL_X8 FILLER_23_894 ();
 FILLCELL_X1 FILLER_23_902 ();
 FILLCELL_X4 FILLER_23_907 ();
 FILLCELL_X8 FILLER_23_915 ();
 FILLCELL_X4 FILLER_23_923 ();
 FILLCELL_X2 FILLER_23_927 ();
 FILLCELL_X1 FILLER_23_929 ();
 FILLCELL_X4 FILLER_23_934 ();
 FILLCELL_X4 FILLER_23_941 ();
 FILLCELL_X2 FILLER_23_945 ();
 FILLCELL_X1 FILLER_23_947 ();
 FILLCELL_X8 FILLER_23_950 ();
 FILLCELL_X2 FILLER_23_958 ();
 FILLCELL_X16 FILLER_23_964 ();
 FILLCELL_X4 FILLER_23_980 ();
 FILLCELL_X4 FILLER_23_986 ();
 FILLCELL_X4 FILLER_23_993 ();
 FILLCELL_X2 FILLER_23_997 ();
 FILLCELL_X4 FILLER_23_1018 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X8 FILLER_24_161 ();
 FILLCELL_X4 FILLER_24_819 ();
 FILLCELL_X2 FILLER_24_823 ();
 FILLCELL_X1 FILLER_24_825 ();
 FILLCELL_X8 FILLER_24_830 ();
 FILLCELL_X4 FILLER_24_841 ();
 FILLCELL_X4 FILLER_24_848 ();
 FILLCELL_X8 FILLER_24_855 ();
 FILLCELL_X4 FILLER_24_863 ();
 FILLCELL_X1 FILLER_24_867 ();
 FILLCELL_X4 FILLER_24_872 ();
 FILLCELL_X4 FILLER_24_885 ();
 FILLCELL_X4 FILLER_24_898 ();
 FILLCELL_X4 FILLER_24_905 ();
 FILLCELL_X4 FILLER_24_918 ();
 FILLCELL_X16 FILLER_24_926 ();
 FILLCELL_X8 FILLER_24_942 ();
 FILLCELL_X4 FILLER_24_957 ();
 FILLCELL_X2 FILLER_24_961 ();
 FILLCELL_X1 FILLER_24_963 ();
 FILLCELL_X4 FILLER_24_973 ();
 FILLCELL_X2 FILLER_24_977 ();
 FILLCELL_X1 FILLER_24_979 ();
 FILLCELL_X4 FILLER_24_984 ();
 FILLCELL_X4 FILLER_24_998 ();
 FILLCELL_X4 FILLER_24_1009 ();
 FILLCELL_X4 FILLER_24_1017 ();
 FILLCELL_X1 FILLER_24_1021 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X8 FILLER_25_161 ();
 FILLCELL_X8 FILLER_25_819 ();
 FILLCELL_X4 FILLER_25_829 ();
 FILLCELL_X4 FILLER_25_836 ();
 FILLCELL_X2 FILLER_25_840 ();
 FILLCELL_X4 FILLER_25_846 ();
 FILLCELL_X16 FILLER_25_860 ();
 FILLCELL_X1 FILLER_25_876 ();
 FILLCELL_X16 FILLER_25_884 ();
 FILLCELL_X4 FILLER_25_900 ();
 FILLCELL_X4 FILLER_25_913 ();
 FILLCELL_X4 FILLER_25_920 ();
 FILLCELL_X8 FILLER_25_928 ();
 FILLCELL_X4 FILLER_25_940 ();
 FILLCELL_X4 FILLER_25_954 ();
 FILLCELL_X4 FILLER_25_967 ();
 FILLCELL_X4 FILLER_25_975 ();
 FILLCELL_X2 FILLER_25_979 ();
 FILLCELL_X1 FILLER_25_981 ();
 FILLCELL_X4 FILLER_25_986 ();
 FILLCELL_X8 FILLER_25_993 ();
 FILLCELL_X4 FILLER_25_1004 ();
 FILLCELL_X8 FILLER_25_1014 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X8 FILLER_26_161 ();
 FILLCELL_X8 FILLER_26_819 ();
 FILLCELL_X1 FILLER_26_827 ();
 FILLCELL_X4 FILLER_26_838 ();
 FILLCELL_X4 FILLER_26_851 ();
 FILLCELL_X2 FILLER_26_855 ();
 FILLCELL_X4 FILLER_26_859 ();
 FILLCELL_X4 FILLER_26_870 ();
 FILLCELL_X2 FILLER_26_874 ();
 FILLCELL_X4 FILLER_26_886 ();
 FILLCELL_X16 FILLER_26_893 ();
 FILLCELL_X8 FILLER_26_909 ();
 FILLCELL_X4 FILLER_26_917 ();
 FILLCELL_X1 FILLER_26_921 ();
 FILLCELL_X4 FILLER_26_926 ();
 FILLCELL_X1 FILLER_26_930 ();
 FILLCELL_X4 FILLER_26_940 ();
 FILLCELL_X2 FILLER_26_944 ();
 FILLCELL_X8 FILLER_26_949 ();
 FILLCELL_X2 FILLER_26_957 ();
 FILLCELL_X8 FILLER_26_962 ();
 FILLCELL_X1 FILLER_26_970 ();
 FILLCELL_X4 FILLER_26_981 ();
 FILLCELL_X4 FILLER_26_994 ();
 FILLCELL_X2 FILLER_26_998 ();
 FILLCELL_X1 FILLER_26_1000 ();
 FILLCELL_X4 FILLER_26_1005 ();
 FILLCELL_X4 FILLER_26_1015 ();
 FILLCELL_X2 FILLER_26_1019 ();
 FILLCELL_X1 FILLER_26_1021 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X8 FILLER_27_161 ();
 FILLCELL_X4 FILLER_27_819 ();
 FILLCELL_X8 FILLER_27_826 ();
 FILLCELL_X8 FILLER_27_837 ();
 FILLCELL_X4 FILLER_27_845 ();
 FILLCELL_X1 FILLER_27_849 ();
 FILLCELL_X8 FILLER_27_857 ();
 FILLCELL_X4 FILLER_27_875 ();
 FILLCELL_X4 FILLER_27_883 ();
 FILLCELL_X2 FILLER_27_887 ();
 FILLCELL_X4 FILLER_27_896 ();
 FILLCELL_X8 FILLER_27_904 ();
 FILLCELL_X4 FILLER_27_912 ();
 FILLCELL_X4 FILLER_27_920 ();
 FILLCELL_X4 FILLER_27_933 ();
 FILLCELL_X8 FILLER_27_940 ();
 FILLCELL_X4 FILLER_27_958 ();
 FILLCELL_X2 FILLER_27_962 ();
 FILLCELL_X4 FILLER_27_967 ();
 FILLCELL_X4 FILLER_27_974 ();
 FILLCELL_X8 FILLER_27_980 ();
 FILLCELL_X2 FILLER_27_988 ();
 FILLCELL_X4 FILLER_27_993 ();
 FILLCELL_X4 FILLER_27_1006 ();
 FILLCELL_X4 FILLER_27_1016 ();
 FILLCELL_X2 FILLER_27_1020 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X8 FILLER_28_161 ();
 FILLCELL_X8 FILLER_28_819 ();
 FILLCELL_X4 FILLER_28_837 ();
 FILLCELL_X4 FILLER_28_850 ();
 FILLCELL_X1 FILLER_28_854 ();
 FILLCELL_X8 FILLER_28_865 ();
 FILLCELL_X1 FILLER_28_873 ();
 FILLCELL_X4 FILLER_28_884 ();
 FILLCELL_X8 FILLER_28_890 ();
 FILLCELL_X4 FILLER_28_908 ();
 FILLCELL_X8 FILLER_28_915 ();
 FILLCELL_X4 FILLER_28_923 ();
 FILLCELL_X4 FILLER_28_930 ();
 FILLCELL_X4 FILLER_28_937 ();
 FILLCELL_X4 FILLER_28_944 ();
 FILLCELL_X4 FILLER_28_950 ();
 FILLCELL_X2 FILLER_28_954 ();
 FILLCELL_X8 FILLER_28_960 ();
 FILLCELL_X1 FILLER_28_968 ();
 FILLCELL_X8 FILLER_28_976 ();
 FILLCELL_X4 FILLER_28_984 ();
 FILLCELL_X1 FILLER_28_988 ();
 FILLCELL_X4 FILLER_28_992 ();
 FILLCELL_X4 FILLER_28_999 ();
 FILLCELL_X4 FILLER_28_1006 ();
 FILLCELL_X4 FILLER_28_1017 ();
 FILLCELL_X1 FILLER_28_1021 ();
 FILLCELL_X4 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_8 ();
 FILLCELL_X32 FILLER_29_40 ();
 FILLCELL_X32 FILLER_29_72 ();
 FILLCELL_X32 FILLER_29_104 ();
 FILLCELL_X32 FILLER_29_136 ();
 FILLCELL_X1 FILLER_29_168 ();
 FILLCELL_X8 FILLER_29_819 ();
 FILLCELL_X2 FILLER_29_827 ();
 FILLCELL_X8 FILLER_29_832 ();
 FILLCELL_X2 FILLER_29_840 ();
 FILLCELL_X1 FILLER_29_842 ();
 FILLCELL_X4 FILLER_29_846 ();
 FILLCELL_X4 FILLER_29_853 ();
 FILLCELL_X8 FILLER_29_859 ();
 FILLCELL_X1 FILLER_29_867 ();
 FILLCELL_X4 FILLER_29_871 ();
 FILLCELL_X1 FILLER_29_875 ();
 FILLCELL_X8 FILLER_29_878 ();
 FILLCELL_X4 FILLER_29_886 ();
 FILLCELL_X1 FILLER_29_890 ();
 FILLCELL_X4 FILLER_29_894 ();
 FILLCELL_X1 FILLER_29_898 ();
 FILLCELL_X4 FILLER_29_903 ();
 FILLCELL_X4 FILLER_29_911 ();
 FILLCELL_X8 FILLER_29_918 ();
 FILLCELL_X8 FILLER_29_929 ();
 FILLCELL_X2 FILLER_29_937 ();
 FILLCELL_X4 FILLER_29_943 ();
 FILLCELL_X8 FILLER_29_954 ();
 FILLCELL_X4 FILLER_29_972 ();
 FILLCELL_X4 FILLER_29_985 ();
 FILLCELL_X4 FILLER_29_998 ();
 FILLCELL_X4 FILLER_29_1008 ();
 FILLCELL_X4 FILLER_29_1015 ();
 FILLCELL_X2 FILLER_29_1019 ();
 FILLCELL_X1 FILLER_29_1021 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X8 FILLER_30_161 ();
 FILLCELL_X4 FILLER_30_819 ();
 FILLCELL_X2 FILLER_30_823 ();
 FILLCELL_X4 FILLER_30_827 ();
 FILLCELL_X4 FILLER_30_834 ();
 FILLCELL_X4 FILLER_30_847 ();
 FILLCELL_X4 FILLER_30_856 ();
 FILLCELL_X4 FILLER_30_863 ();
 FILLCELL_X4 FILLER_30_870 ();
 FILLCELL_X4 FILLER_30_877 ();
 FILLCELL_X4 FILLER_30_884 ();
 FILLCELL_X8 FILLER_30_890 ();
 FILLCELL_X4 FILLER_30_907 ();
 FILLCELL_X4 FILLER_30_913 ();
 FILLCELL_X2 FILLER_30_917 ();
 FILLCELL_X1 FILLER_30_919 ();
 FILLCELL_X4 FILLER_30_924 ();
 FILLCELL_X2 FILLER_30_928 ();
 FILLCELL_X1 FILLER_30_930 ();
 FILLCELL_X4 FILLER_30_940 ();
 FILLCELL_X2 FILLER_30_944 ();
 FILLCELL_X16 FILLER_30_956 ();
 FILLCELL_X2 FILLER_30_972 ();
 FILLCELL_X1 FILLER_30_974 ();
 FILLCELL_X4 FILLER_30_979 ();
 FILLCELL_X4 FILLER_30_986 ();
 FILLCELL_X4 FILLER_30_993 ();
 FILLCELL_X2 FILLER_30_997 ();
 FILLCELL_X4 FILLER_30_1002 ();
 FILLCELL_X4 FILLER_30_1009 ();
 FILLCELL_X4 FILLER_30_1015 ();
 FILLCELL_X2 FILLER_30_1019 ();
 FILLCELL_X1 FILLER_30_1021 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X8 FILLER_31_161 ();
 FILLCELL_X8 FILLER_31_819 ();
 FILLCELL_X2 FILLER_31_827 ();
 FILLCELL_X4 FILLER_31_838 ();
 FILLCELL_X8 FILLER_31_849 ();
 FILLCELL_X4 FILLER_31_860 ();
 FILLCELL_X1 FILLER_31_864 ();
 FILLCELL_X8 FILLER_31_874 ();
 FILLCELL_X1 FILLER_31_882 ();
 FILLCELL_X4 FILLER_31_886 ();
 FILLCELL_X4 FILLER_31_900 ();
 FILLCELL_X8 FILLER_31_907 ();
 FILLCELL_X4 FILLER_31_919 ();
 FILLCELL_X4 FILLER_31_932 ();
 FILLCELL_X4 FILLER_31_940 ();
 FILLCELL_X2 FILLER_31_944 ();
 FILLCELL_X1 FILLER_31_946 ();
 FILLCELL_X32 FILLER_31_950 ();
 FILLCELL_X8 FILLER_31_982 ();
 FILLCELL_X4 FILLER_31_990 ();
 FILLCELL_X2 FILLER_31_994 ();
 FILLCELL_X8 FILLER_31_999 ();
 FILLCELL_X1 FILLER_31_1007 ();
 FILLCELL_X4 FILLER_31_1018 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X8 FILLER_32_161 ();
 FILLCELL_X8 FILLER_32_819 ();
 FILLCELL_X4 FILLER_32_837 ();
 FILLCELL_X4 FILLER_32_848 ();
 FILLCELL_X2 FILLER_32_852 ();
 FILLCELL_X4 FILLER_32_864 ();
 FILLCELL_X4 FILLER_32_877 ();
 FILLCELL_X4 FILLER_32_888 ();
 FILLCELL_X1 FILLER_32_892 ();
 FILLCELL_X4 FILLER_32_902 ();
 FILLCELL_X16 FILLER_32_910 ();
 FILLCELL_X4 FILLER_32_926 ();
 FILLCELL_X8 FILLER_32_933 ();
 FILLCELL_X4 FILLER_32_941 ();
 FILLCELL_X4 FILLER_32_948 ();
 FILLCELL_X4 FILLER_32_961 ();
 FILLCELL_X4 FILLER_32_968 ();
 FILLCELL_X1 FILLER_32_972 ();
 FILLCELL_X8 FILLER_32_977 ();
 FILLCELL_X1 FILLER_32_985 ();
 FILLCELL_X4 FILLER_32_990 ();
 FILLCELL_X1 FILLER_32_994 ();
 FILLCELL_X4 FILLER_32_1005 ();
 FILLCELL_X4 FILLER_32_1016 ();
 FILLCELL_X2 FILLER_32_1020 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X8 FILLER_33_161 ();
 FILLCELL_X8 FILLER_33_819 ();
 FILLCELL_X2 FILLER_33_827 ();
 FILLCELL_X1 FILLER_33_829 ();
 FILLCELL_X4 FILLER_33_833 ();
 FILLCELL_X8 FILLER_33_839 ();
 FILLCELL_X4 FILLER_33_854 ();
 FILLCELL_X8 FILLER_33_860 ();
 FILLCELL_X4 FILLER_33_868 ();
 FILLCELL_X8 FILLER_33_874 ();
 FILLCELL_X4 FILLER_33_892 ();
 FILLCELL_X8 FILLER_33_900 ();
 FILLCELL_X1 FILLER_33_908 ();
 FILLCELL_X8 FILLER_33_928 ();
 FILLCELL_X4 FILLER_33_936 ();
 FILLCELL_X2 FILLER_33_940 ();
 FILLCELL_X1 FILLER_33_942 ();
 FILLCELL_X4 FILLER_33_952 ();
 FILLCELL_X4 FILLER_33_960 ();
 FILLCELL_X2 FILLER_33_964 ();
 FILLCELL_X1 FILLER_33_966 ();
 FILLCELL_X4 FILLER_33_971 ();
 FILLCELL_X4 FILLER_33_984 ();
 FILLCELL_X8 FILLER_33_991 ();
 FILLCELL_X4 FILLER_33_1018 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X8 FILLER_34_161 ();
 FILLCELL_X4 FILLER_34_819 ();
 FILLCELL_X4 FILLER_34_829 ();
 FILLCELL_X4 FILLER_34_835 ();
 FILLCELL_X2 FILLER_34_839 ();
 FILLCELL_X1 FILLER_34_841 ();
 FILLCELL_X4 FILLER_34_844 ();
 FILLCELL_X8 FILLER_34_850 ();
 FILLCELL_X2 FILLER_34_858 ();
 FILLCELL_X1 FILLER_34_860 ();
 FILLCELL_X4 FILLER_34_871 ();
 FILLCELL_X8 FILLER_34_877 ();
 FILLCELL_X4 FILLER_34_885 ();
 FILLCELL_X2 FILLER_34_889 ();
 FILLCELL_X8 FILLER_34_894 ();
 FILLCELL_X1 FILLER_34_902 ();
 FILLCELL_X16 FILLER_34_907 ();
 FILLCELL_X2 FILLER_34_923 ();
 FILLCELL_X4 FILLER_34_929 ();
 FILLCELL_X8 FILLER_34_935 ();
 FILLCELL_X4 FILLER_34_943 ();
 FILLCELL_X2 FILLER_34_947 ();
 FILLCELL_X1 FILLER_34_949 ();
 FILLCELL_X8 FILLER_34_953 ();
 FILLCELL_X2 FILLER_34_961 ();
 FILLCELL_X1 FILLER_34_963 ();
 FILLCELL_X4 FILLER_34_974 ();
 FILLCELL_X4 FILLER_34_982 ();
 FILLCELL_X4 FILLER_34_995 ();
 FILLCELL_X4 FILLER_34_1002 ();
 FILLCELL_X2 FILLER_34_1006 ();
 FILLCELL_X4 FILLER_34_1011 ();
 FILLCELL_X4 FILLER_34_1018 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X16 FILLER_35_129 ();
 FILLCELL_X8 FILLER_35_145 ();
 FILLCELL_X8 FILLER_35_155 ();
 FILLCELL_X4 FILLER_35_163 ();
 FILLCELL_X2 FILLER_35_167 ();
 FILLCELL_X4 FILLER_35_819 ();
 FILLCELL_X4 FILLER_35_826 ();
 FILLCELL_X1 FILLER_35_830 ();
 FILLCELL_X4 FILLER_35_841 ();
 FILLCELL_X8 FILLER_35_855 ();
 FILLCELL_X2 FILLER_35_863 ();
 FILLCELL_X4 FILLER_35_867 ();
 FILLCELL_X4 FILLER_35_878 ();
 FILLCELL_X8 FILLER_35_886 ();
 FILLCELL_X2 FILLER_35_894 ();
 FILLCELL_X4 FILLER_35_900 ();
 FILLCELL_X4 FILLER_35_908 ();
 FILLCELL_X2 FILLER_35_912 ();
 FILLCELL_X1 FILLER_35_914 ();
 FILLCELL_X4 FILLER_35_919 ();
 FILLCELL_X4 FILLER_35_927 ();
 FILLCELL_X8 FILLER_35_948 ();
 FILLCELL_X4 FILLER_35_956 ();
 FILLCELL_X2 FILLER_35_960 ();
 FILLCELL_X1 FILLER_35_962 ();
 FILLCELL_X16 FILLER_35_965 ();
 FILLCELL_X1 FILLER_35_981 ();
 FILLCELL_X8 FILLER_35_985 ();
 FILLCELL_X4 FILLER_35_993 ();
 FILLCELL_X2 FILLER_35_997 ();
 FILLCELL_X1 FILLER_35_999 ();
 FILLCELL_X4 FILLER_35_1002 ();
 FILLCELL_X4 FILLER_35_1010 ();
 FILLCELL_X4 FILLER_35_1018 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X8 FILLER_36_129 ();
 FILLCELL_X2 FILLER_36_137 ();
 FILLCELL_X4 FILLER_36_142 ();
 FILLCELL_X2 FILLER_36_146 ();
 FILLCELL_X4 FILLER_36_165 ();
 FILLCELL_X4 FILLER_36_819 ();
 FILLCELL_X8 FILLER_36_826 ();
 FILLCELL_X4 FILLER_36_834 ();
 FILLCELL_X2 FILLER_36_838 ();
 FILLCELL_X1 FILLER_36_840 ();
 FILLCELL_X4 FILLER_36_844 ();
 FILLCELL_X1 FILLER_36_848 ();
 FILLCELL_X4 FILLER_36_852 ();
 FILLCELL_X4 FILLER_36_859 ();
 FILLCELL_X2 FILLER_36_863 ();
 FILLCELL_X1 FILLER_36_865 ();
 FILLCELL_X4 FILLER_36_876 ();
 FILLCELL_X4 FILLER_36_890 ();
 FILLCELL_X4 FILLER_36_903 ();
 FILLCELL_X8 FILLER_36_916 ();
 FILLCELL_X2 FILLER_36_924 ();
 FILLCELL_X1 FILLER_36_926 ();
 FILLCELL_X4 FILLER_36_934 ();
 FILLCELL_X16 FILLER_36_943 ();
 FILLCELL_X1 FILLER_36_959 ();
 FILLCELL_X4 FILLER_36_970 ();
 FILLCELL_X4 FILLER_36_981 ();
 FILLCELL_X2 FILLER_36_985 ();
 FILLCELL_X4 FILLER_36_991 ();
 FILLCELL_X4 FILLER_36_1004 ();
 FILLCELL_X4 FILLER_36_1018 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X2 FILLER_37_129 ();
 FILLCELL_X1 FILLER_37_131 ();
 FILLCELL_X4 FILLER_37_135 ();
 FILLCELL_X4 FILLER_37_142 ();
 FILLCELL_X8 FILLER_37_149 ();
 FILLCELL_X1 FILLER_37_157 ();
 FILLCELL_X4 FILLER_37_162 ();
 FILLCELL_X2 FILLER_37_166 ();
 FILLCELL_X1 FILLER_37_168 ();
 FILLCELL_X16 FILLER_37_819 ();
 FILLCELL_X1 FILLER_37_835 ();
 FILLCELL_X4 FILLER_37_839 ();
 FILLCELL_X4 FILLER_37_846 ();
 FILLCELL_X1 FILLER_37_850 ();
 FILLCELL_X8 FILLER_37_860 ();
 FILLCELL_X4 FILLER_37_878 ();
 FILLCELL_X8 FILLER_37_885 ();
 FILLCELL_X1 FILLER_37_893 ();
 FILLCELL_X4 FILLER_37_897 ();
 FILLCELL_X4 FILLER_37_905 ();
 FILLCELL_X16 FILLER_37_912 ();
 FILLCELL_X4 FILLER_37_933 ();
 FILLCELL_X8 FILLER_37_941 ();
 FILLCELL_X1 FILLER_37_949 ();
 FILLCELL_X4 FILLER_37_969 ();
 FILLCELL_X4 FILLER_37_976 ();
 FILLCELL_X2 FILLER_37_980 ();
 FILLCELL_X8 FILLER_37_991 ();
 FILLCELL_X4 FILLER_37_1004 ();
 FILLCELL_X4 FILLER_37_1012 ();
 FILLCELL_X4 FILLER_37_1018 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X16 FILLER_38_97 ();
 FILLCELL_X4 FILLER_38_113 ();
 FILLCELL_X2 FILLER_38_117 ();
 FILLCELL_X1 FILLER_38_119 ();
 FILLCELL_X4 FILLER_38_137 ();
 FILLCELL_X4 FILLER_38_144 ();
 FILLCELL_X4 FILLER_38_151 ();
 FILLCELL_X4 FILLER_38_158 ();
 FILLCELL_X4 FILLER_38_165 ();
 FILLCELL_X8 FILLER_38_819 ();
 FILLCELL_X1 FILLER_38_827 ();
 FILLCELL_X4 FILLER_38_834 ();
 FILLCELL_X2 FILLER_38_838 ();
 FILLCELL_X1 FILLER_38_840 ();
 FILLCELL_X4 FILLER_38_850 ();
 FILLCELL_X4 FILLER_38_858 ();
 FILLCELL_X4 FILLER_38_865 ();
 FILLCELL_X2 FILLER_38_869 ();
 FILLCELL_X1 FILLER_38_871 ();
 FILLCELL_X4 FILLER_38_874 ();
 FILLCELL_X4 FILLER_38_881 ();
 FILLCELL_X16 FILLER_38_888 ();
 FILLCELL_X4 FILLER_38_904 ();
 FILLCELL_X4 FILLER_38_912 ();
 FILLCELL_X8 FILLER_38_920 ();
 FILLCELL_X2 FILLER_38_928 ();
 FILLCELL_X8 FILLER_38_934 ();
 FILLCELL_X2 FILLER_38_942 ();
 FILLCELL_X8 FILLER_38_948 ();
 FILLCELL_X4 FILLER_38_960 ();
 FILLCELL_X8 FILLER_38_967 ();
 FILLCELL_X4 FILLER_38_975 ();
 FILLCELL_X4 FILLER_38_982 ();
 FILLCELL_X4 FILLER_38_990 ();
 FILLCELL_X4 FILLER_38_999 ();
 FILLCELL_X8 FILLER_38_1012 ();
 FILLCELL_X2 FILLER_38_1020 ();
 FILLCELL_X4 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_9 ();
 FILLCELL_X32 FILLER_39_41 ();
 FILLCELL_X32 FILLER_39_73 ();
 FILLCELL_X4 FILLER_39_105 ();
 FILLCELL_X2 FILLER_39_109 ();
 FILLCELL_X1 FILLER_39_111 ();
 FILLCELL_X4 FILLER_39_131 ();
 FILLCELL_X4 FILLER_39_140 ();
 FILLCELL_X4 FILLER_39_148 ();
 FILLCELL_X1 FILLER_39_152 ();
 FILLCELL_X4 FILLER_39_162 ();
 FILLCELL_X2 FILLER_39_166 ();
 FILLCELL_X1 FILLER_39_168 ();
 FILLCELL_X4 FILLER_39_819 ();
 FILLCELL_X2 FILLER_39_823 ();
 FILLCELL_X1 FILLER_39_825 ();
 FILLCELL_X4 FILLER_39_836 ();
 FILLCELL_X8 FILLER_39_847 ();
 FILLCELL_X2 FILLER_39_855 ();
 FILLCELL_X4 FILLER_39_866 ();
 FILLCELL_X4 FILLER_39_873 ();
 FILLCELL_X4 FILLER_39_879 ();
 FILLCELL_X4 FILLER_39_892 ();
 FILLCELL_X1 FILLER_39_896 ();
 FILLCELL_X4 FILLER_39_901 ();
 FILLCELL_X4 FILLER_39_910 ();
 FILLCELL_X4 FILLER_39_919 ();
 FILLCELL_X8 FILLER_39_927 ();
 FILLCELL_X1 FILLER_39_935 ();
 FILLCELL_X4 FILLER_39_945 ();
 FILLCELL_X4 FILLER_39_958 ();
 FILLCELL_X4 FILLER_39_966 ();
 FILLCELL_X2 FILLER_39_970 ();
 FILLCELL_X8 FILLER_39_982 ();
 FILLCELL_X4 FILLER_39_993 ();
 FILLCELL_X8 FILLER_39_1001 ();
 FILLCELL_X2 FILLER_39_1009 ();
 FILLCELL_X1 FILLER_39_1011 ();
 FILLCELL_X4 FILLER_39_1015 ();
 FILLCELL_X2 FILLER_39_1019 ();
 FILLCELL_X1 FILLER_39_1021 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X1 FILLER_40_97 ();
 FILLCELL_X4 FILLER_40_101 ();
 FILLCELL_X2 FILLER_40_105 ();
 FILLCELL_X1 FILLER_40_107 ();
 FILLCELL_X4 FILLER_40_112 ();
 FILLCELL_X2 FILLER_40_116 ();
 FILLCELL_X4 FILLER_40_121 ();
 FILLCELL_X4 FILLER_40_128 ();
 FILLCELL_X8 FILLER_40_136 ();
 FILLCELL_X1 FILLER_40_144 ();
 FILLCELL_X4 FILLER_40_164 ();
 FILLCELL_X1 FILLER_40_168 ();
 FILLCELL_X4 FILLER_40_819 ();
 FILLCELL_X1 FILLER_40_823 ();
 FILLCELL_X4 FILLER_40_827 ();
 FILLCELL_X4 FILLER_40_835 ();
 FILLCELL_X1 FILLER_40_839 ();
 FILLCELL_X4 FILLER_40_849 ();
 FILLCELL_X4 FILLER_40_860 ();
 FILLCELL_X8 FILLER_40_874 ();
 FILLCELL_X4 FILLER_40_885 ();
 FILLCELL_X8 FILLER_40_892 ();
 FILLCELL_X1 FILLER_40_900 ();
 FILLCELL_X8 FILLER_40_910 ();
 FILLCELL_X16 FILLER_40_923 ();
 FILLCELL_X4 FILLER_40_942 ();
 FILLCELL_X1 FILLER_40_946 ();
 FILLCELL_X4 FILLER_40_950 ();
 FILLCELL_X1 FILLER_40_954 ();
 FILLCELL_X4 FILLER_40_959 ();
 FILLCELL_X4 FILLER_40_967 ();
 FILLCELL_X4 FILLER_40_974 ();
 FILLCELL_X16 FILLER_40_980 ();
 FILLCELL_X2 FILLER_40_996 ();
 FILLCELL_X1 FILLER_40_998 ();
 FILLCELL_X4 FILLER_40_1018 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X16 FILLER_41_65 ();
 FILLCELL_X8 FILLER_41_81 ();
 FILLCELL_X4 FILLER_41_106 ();
 FILLCELL_X16 FILLER_41_114 ();
 FILLCELL_X2 FILLER_41_130 ();
 FILLCELL_X1 FILLER_41_132 ();
 FILLCELL_X4 FILLER_41_136 ();
 FILLCELL_X4 FILLER_41_143 ();
 FILLCELL_X2 FILLER_41_147 ();
 FILLCELL_X16 FILLER_41_153 ();
 FILLCELL_X8 FILLER_41_819 ();
 FILLCELL_X2 FILLER_41_827 ();
 FILLCELL_X4 FILLER_41_832 ();
 FILLCELL_X4 FILLER_41_846 ();
 FILLCELL_X8 FILLER_41_852 ();
 FILLCELL_X4 FILLER_41_860 ();
 FILLCELL_X4 FILLER_41_866 ();
 FILLCELL_X2 FILLER_41_870 ();
 FILLCELL_X4 FILLER_41_879 ();
 FILLCELL_X1 FILLER_41_883 ();
 FILLCELL_X8 FILLER_41_893 ();
 FILLCELL_X4 FILLER_41_901 ();
 FILLCELL_X1 FILLER_41_905 ();
 FILLCELL_X4 FILLER_41_908 ();
 FILLCELL_X8 FILLER_41_916 ();
 FILLCELL_X1 FILLER_41_924 ();
 FILLCELL_X4 FILLER_41_929 ();
 FILLCELL_X2 FILLER_41_933 ();
 FILLCELL_X8 FILLER_41_939 ();
 FILLCELL_X4 FILLER_41_947 ();
 FILLCELL_X2 FILLER_41_951 ();
 FILLCELL_X8 FILLER_41_959 ();
 FILLCELL_X2 FILLER_41_967 ();
 FILLCELL_X4 FILLER_41_979 ();
 FILLCELL_X4 FILLER_41_990 ();
 FILLCELL_X4 FILLER_41_997 ();
 FILLCELL_X4 FILLER_41_1005 ();
 FILLCELL_X4 FILLER_41_1015 ();
 FILLCELL_X2 FILLER_41_1019 ();
 FILLCELL_X1 FILLER_41_1021 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X8 FILLER_42_65 ();
 FILLCELL_X4 FILLER_42_73 ();
 FILLCELL_X2 FILLER_42_77 ();
 FILLCELL_X4 FILLER_42_82 ();
 FILLCELL_X4 FILLER_42_91 ();
 FILLCELL_X4 FILLER_42_100 ();
 FILLCELL_X4 FILLER_42_109 ();
 FILLCELL_X2 FILLER_42_113 ();
 FILLCELL_X4 FILLER_42_119 ();
 FILLCELL_X4 FILLER_42_125 ();
 FILLCELL_X1 FILLER_42_129 ();
 FILLCELL_X4 FILLER_42_136 ();
 FILLCELL_X4 FILLER_42_143 ();
 FILLCELL_X16 FILLER_42_150 ();
 FILLCELL_X2 FILLER_42_166 ();
 FILLCELL_X1 FILLER_42_168 ();
 FILLCELL_X16 FILLER_42_819 ();
 FILLCELL_X1 FILLER_42_835 ();
 FILLCELL_X4 FILLER_42_840 ();
 FILLCELL_X1 FILLER_42_844 ();
 FILLCELL_X16 FILLER_42_847 ();
 FILLCELL_X8 FILLER_42_873 ();
 FILLCELL_X4 FILLER_42_891 ();
 FILLCELL_X16 FILLER_42_898 ();
 FILLCELL_X8 FILLER_42_914 ();
 FILLCELL_X4 FILLER_42_941 ();
 FILLCELL_X8 FILLER_42_951 ();
 FILLCELL_X2 FILLER_42_959 ();
 FILLCELL_X4 FILLER_42_970 ();
 FILLCELL_X2 FILLER_42_974 ();
 FILLCELL_X1 FILLER_42_976 ();
 FILLCELL_X4 FILLER_42_981 ();
 FILLCELL_X4 FILLER_42_994 ();
 FILLCELL_X2 FILLER_42_998 ();
 FILLCELL_X1 FILLER_42_1000 ();
 FILLCELL_X4 FILLER_42_1005 ();
 FILLCELL_X4 FILLER_42_1015 ();
 FILLCELL_X2 FILLER_42_1019 ();
 FILLCELL_X1 FILLER_42_1021 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X2 FILLER_43_65 ();
 FILLCELL_X4 FILLER_43_70 ();
 FILLCELL_X4 FILLER_43_91 ();
 FILLCELL_X4 FILLER_43_98 ();
 FILLCELL_X4 FILLER_43_109 ();
 FILLCELL_X4 FILLER_43_116 ();
 FILLCELL_X2 FILLER_43_120 ();
 FILLCELL_X4 FILLER_43_139 ();
 FILLCELL_X4 FILLER_43_148 ();
 FILLCELL_X8 FILLER_43_156 ();
 FILLCELL_X4 FILLER_43_164 ();
 FILLCELL_X1 FILLER_43_168 ();
 FILLCELL_X16 FILLER_43_819 ();
 FILLCELL_X4 FILLER_43_837 ();
 FILLCELL_X4 FILLER_43_844 ();
 FILLCELL_X4 FILLER_43_852 ();
 FILLCELL_X8 FILLER_43_859 ();
 FILLCELL_X4 FILLER_43_867 ();
 FILLCELL_X1 FILLER_43_871 ();
 FILLCELL_X8 FILLER_43_882 ();
 FILLCELL_X4 FILLER_43_893 ();
 FILLCELL_X1 FILLER_43_897 ();
 FILLCELL_X4 FILLER_43_903 ();
 FILLCELL_X4 FILLER_43_916 ();
 FILLCELL_X4 FILLER_43_924 ();
 FILLCELL_X8 FILLER_43_932 ();
 FILLCELL_X4 FILLER_43_944 ();
 FILLCELL_X4 FILLER_43_952 ();
 FILLCELL_X4 FILLER_43_960 ();
 FILLCELL_X16 FILLER_43_967 ();
 FILLCELL_X4 FILLER_43_986 ();
 FILLCELL_X4 FILLER_43_999 ();
 FILLCELL_X4 FILLER_43_1006 ();
 FILLCELL_X4 FILLER_43_1017 ();
 FILLCELL_X1 FILLER_43_1021 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X32 FILLER_44_33 ();
 FILLCELL_X1 FILLER_44_65 ();
 FILLCELL_X4 FILLER_44_69 ();
 FILLCELL_X4 FILLER_44_76 ();
 FILLCELL_X4 FILLER_44_83 ();
 FILLCELL_X4 FILLER_44_93 ();
 FILLCELL_X4 FILLER_44_101 ();
 FILLCELL_X8 FILLER_44_109 ();
 FILLCELL_X4 FILLER_44_122 ();
 FILLCELL_X2 FILLER_44_126 ();
 FILLCELL_X1 FILLER_44_128 ();
 FILLCELL_X4 FILLER_44_133 ();
 FILLCELL_X4 FILLER_44_142 ();
 FILLCELL_X4 FILLER_44_165 ();
 FILLCELL_X8 FILLER_44_819 ();
 FILLCELL_X4 FILLER_44_831 ();
 FILLCELL_X4 FILLER_44_840 ();
 FILLCELL_X4 FILLER_44_853 ();
 FILLCELL_X8 FILLER_44_861 ();
 FILLCELL_X4 FILLER_44_869 ();
 FILLCELL_X2 FILLER_44_873 ();
 FILLCELL_X8 FILLER_44_877 ();
 FILLCELL_X2 FILLER_44_885 ();
 FILLCELL_X4 FILLER_44_893 ();
 FILLCELL_X4 FILLER_44_906 ();
 FILLCELL_X4 FILLER_44_914 ();
 FILLCELL_X16 FILLER_44_922 ();
 FILLCELL_X8 FILLER_44_938 ();
 FILLCELL_X1 FILLER_44_946 ();
 FILLCELL_X4 FILLER_44_951 ();
 FILLCELL_X2 FILLER_44_955 ();
 FILLCELL_X16 FILLER_44_966 ();
 FILLCELL_X4 FILLER_44_982 ();
 FILLCELL_X2 FILLER_44_986 ();
 FILLCELL_X1 FILLER_44_988 ();
 FILLCELL_X4 FILLER_44_991 ();
 FILLCELL_X8 FILLER_44_1001 ();
 FILLCELL_X1 FILLER_44_1009 ();
 FILLCELL_X8 FILLER_44_1014 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X32 FILLER_45_33 ();
 FILLCELL_X8 FILLER_45_65 ();
 FILLCELL_X4 FILLER_45_73 ();
 FILLCELL_X2 FILLER_45_77 ();
 FILLCELL_X4 FILLER_45_82 ();
 FILLCELL_X4 FILLER_45_89 ();
 FILLCELL_X4 FILLER_45_97 ();
 FILLCELL_X4 FILLER_45_105 ();
 FILLCELL_X2 FILLER_45_109 ();
 FILLCELL_X1 FILLER_45_111 ();
 FILLCELL_X4 FILLER_45_114 ();
 FILLCELL_X4 FILLER_45_121 ();
 FILLCELL_X4 FILLER_45_129 ();
 FILLCELL_X4 FILLER_45_140 ();
 FILLCELL_X4 FILLER_45_149 ();
 FILLCELL_X4 FILLER_45_156 ();
 FILLCELL_X4 FILLER_45_163 ();
 FILLCELL_X2 FILLER_45_167 ();
 FILLCELL_X4 FILLER_45_819 ();
 FILLCELL_X4 FILLER_45_827 ();
 FILLCELL_X4 FILLER_45_840 ();
 FILLCELL_X4 FILLER_45_850 ();
 FILLCELL_X4 FILLER_45_858 ();
 FILLCELL_X2 FILLER_45_862 ();
 FILLCELL_X1 FILLER_45_864 ();
 FILLCELL_X4 FILLER_45_868 ();
 FILLCELL_X4 FILLER_45_878 ();
 FILLCELL_X8 FILLER_45_884 ();
 FILLCELL_X4 FILLER_45_892 ();
 FILLCELL_X4 FILLER_45_901 ();
 FILLCELL_X8 FILLER_45_909 ();
 FILLCELL_X4 FILLER_45_917 ();
 FILLCELL_X4 FILLER_45_925 ();
 FILLCELL_X8 FILLER_45_934 ();
 FILLCELL_X4 FILLER_45_942 ();
 FILLCELL_X2 FILLER_45_946 ();
 FILLCELL_X1 FILLER_45_948 ();
 FILLCELL_X4 FILLER_45_953 ();
 FILLCELL_X4 FILLER_45_963 ();
 FILLCELL_X4 FILLER_45_970 ();
 FILLCELL_X4 FILLER_45_977 ();
 FILLCELL_X1 FILLER_45_981 ();
 FILLCELL_X4 FILLER_45_985 ();
 FILLCELL_X4 FILLER_45_999 ();
 FILLCELL_X4 FILLER_45_1005 ();
 FILLCELL_X2 FILLER_45_1009 ();
 FILLCELL_X1 FILLER_45_1011 ();
 FILLCELL_X4 FILLER_45_1018 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X32 FILLER_46_33 ();
 FILLCELL_X8 FILLER_46_65 ();
 FILLCELL_X4 FILLER_46_73 ();
 FILLCELL_X4 FILLER_46_80 ();
 FILLCELL_X4 FILLER_46_89 ();
 FILLCELL_X4 FILLER_46_99 ();
 FILLCELL_X4 FILLER_46_108 ();
 FILLCELL_X1 FILLER_46_112 ();
 FILLCELL_X4 FILLER_46_117 ();
 FILLCELL_X4 FILLER_46_123 ();
 FILLCELL_X2 FILLER_46_127 ();
 FILLCELL_X1 FILLER_46_129 ();
 FILLCELL_X4 FILLER_46_133 ();
 FILLCELL_X4 FILLER_46_140 ();
 FILLCELL_X4 FILLER_46_149 ();
 FILLCELL_X2 FILLER_46_153 ();
 FILLCELL_X1 FILLER_46_155 ();
 FILLCELL_X4 FILLER_46_159 ();
 FILLCELL_X4 FILLER_46_165 ();
 FILLCELL_X16 FILLER_46_819 ();
 FILLCELL_X4 FILLER_46_840 ();
 FILLCELL_X8 FILLER_46_854 ();
 FILLCELL_X4 FILLER_46_869 ();
 FILLCELL_X4 FILLER_46_883 ();
 FILLCELL_X8 FILLER_46_890 ();
 FILLCELL_X1 FILLER_46_898 ();
 FILLCELL_X8 FILLER_46_902 ();
 FILLCELL_X1 FILLER_46_910 ();
 FILLCELL_X4 FILLER_46_915 ();
 FILLCELL_X4 FILLER_46_924 ();
 FILLCELL_X4 FILLER_46_937 ();
 FILLCELL_X16 FILLER_46_943 ();
 FILLCELL_X2 FILLER_46_959 ();
 FILLCELL_X4 FILLER_46_967 ();
 FILLCELL_X2 FILLER_46_971 ();
 FILLCELL_X1 FILLER_46_973 ();
 FILLCELL_X4 FILLER_46_976 ();
 FILLCELL_X1 FILLER_46_980 ();
 FILLCELL_X4 FILLER_46_987 ();
 FILLCELL_X2 FILLER_46_991 ();
 FILLCELL_X1 FILLER_46_993 ();
 FILLCELL_X4 FILLER_46_1001 ();
 FILLCELL_X4 FILLER_46_1011 ();
 FILLCELL_X4 FILLER_46_1018 ();
 FILLCELL_X32 FILLER_47_1 ();
 FILLCELL_X32 FILLER_47_33 ();
 FILLCELL_X8 FILLER_47_65 ();
 FILLCELL_X4 FILLER_47_92 ();
 FILLCELL_X1 FILLER_47_96 ();
 FILLCELL_X4 FILLER_47_102 ();
 FILLCELL_X4 FILLER_47_112 ();
 FILLCELL_X1 FILLER_47_116 ();
 FILLCELL_X4 FILLER_47_122 ();
 FILLCELL_X8 FILLER_47_131 ();
 FILLCELL_X2 FILLER_47_139 ();
 FILLCELL_X4 FILLER_47_144 ();
 FILLCELL_X4 FILLER_47_154 ();
 FILLCELL_X2 FILLER_47_158 ();
 FILLCELL_X4 FILLER_47_165 ();
 FILLCELL_X4 FILLER_47_819 ();
 FILLCELL_X16 FILLER_47_826 ();
 FILLCELL_X8 FILLER_47_842 ();
 FILLCELL_X4 FILLER_47_852 ();
 FILLCELL_X8 FILLER_47_859 ();
 FILLCELL_X1 FILLER_47_867 ();
 FILLCELL_X4 FILLER_47_871 ();
 FILLCELL_X4 FILLER_47_879 ();
 FILLCELL_X1 FILLER_47_883 ();
 FILLCELL_X8 FILLER_47_886 ();
 FILLCELL_X4 FILLER_47_897 ();
 FILLCELL_X2 FILLER_47_901 ();
 FILLCELL_X1 FILLER_47_903 ();
 FILLCELL_X8 FILLER_47_908 ();
 FILLCELL_X4 FILLER_47_916 ();
 FILLCELL_X2 FILLER_47_920 ();
 FILLCELL_X4 FILLER_47_926 ();
 FILLCELL_X4 FILLER_47_934 ();
 FILLCELL_X4 FILLER_47_940 ();
 FILLCELL_X2 FILLER_47_944 ();
 FILLCELL_X4 FILLER_47_949 ();
 FILLCELL_X4 FILLER_47_957 ();
 FILLCELL_X2 FILLER_47_961 ();
 FILLCELL_X1 FILLER_47_963 ();
 FILLCELL_X4 FILLER_47_970 ();
 FILLCELL_X4 FILLER_47_977 ();
 FILLCELL_X4 FILLER_47_984 ();
 FILLCELL_X4 FILLER_47_990 ();
 FILLCELL_X4 FILLER_47_997 ();
 FILLCELL_X4 FILLER_47_1018 ();
 FILLCELL_X32 FILLER_48_1 ();
 FILLCELL_X32 FILLER_48_33 ();
 FILLCELL_X8 FILLER_48_65 ();
 FILLCELL_X4 FILLER_48_73 ();
 FILLCELL_X1 FILLER_48_77 ();
 FILLCELL_X4 FILLER_48_81 ();
 FILLCELL_X4 FILLER_48_104 ();
 FILLCELL_X4 FILLER_48_111 ();
 FILLCELL_X4 FILLER_48_134 ();
 FILLCELL_X4 FILLER_48_140 ();
 FILLCELL_X8 FILLER_48_161 ();
 FILLCELL_X8 FILLER_48_819 ();
 FILLCELL_X1 FILLER_48_827 ();
 FILLCELL_X4 FILLER_48_832 ();
 FILLCELL_X2 FILLER_48_836 ();
 FILLCELL_X1 FILLER_48_838 ();
 FILLCELL_X4 FILLER_48_842 ();
 FILLCELL_X4 FILLER_48_849 ();
 FILLCELL_X8 FILLER_48_856 ();
 FILLCELL_X1 FILLER_48_864 ();
 FILLCELL_X4 FILLER_48_874 ();
 FILLCELL_X8 FILLER_48_884 ();
 FILLCELL_X4 FILLER_48_897 ();
 FILLCELL_X4 FILLER_48_910 ();
 FILLCELL_X4 FILLER_48_918 ();
 FILLCELL_X2 FILLER_48_922 ();
 FILLCELL_X1 FILLER_48_924 ();
 FILLCELL_X8 FILLER_48_927 ();
 FILLCELL_X4 FILLER_48_938 ();
 FILLCELL_X16 FILLER_48_944 ();
 FILLCELL_X1 FILLER_48_960 ();
 FILLCELL_X4 FILLER_48_965 ();
 FILLCELL_X4 FILLER_48_972 ();
 FILLCELL_X2 FILLER_48_976 ();
 FILLCELL_X8 FILLER_48_988 ();
 FILLCELL_X1 FILLER_48_996 ();
 FILLCELL_X4 FILLER_48_1000 ();
 FILLCELL_X2 FILLER_48_1004 ();
 FILLCELL_X1 FILLER_48_1006 ();
 FILLCELL_X8 FILLER_48_1014 ();
 FILLCELL_X32 FILLER_49_1 ();
 FILLCELL_X32 FILLER_49_33 ();
 FILLCELL_X16 FILLER_49_65 ();
 FILLCELL_X8 FILLER_49_81 ();
 FILLCELL_X2 FILLER_49_89 ();
 FILLCELL_X4 FILLER_49_94 ();
 FILLCELL_X4 FILLER_49_101 ();
 FILLCELL_X4 FILLER_49_108 ();
 FILLCELL_X4 FILLER_49_115 ();
 FILLCELL_X4 FILLER_49_122 ();
 FILLCELL_X4 FILLER_49_129 ();
 FILLCELL_X8 FILLER_49_139 ();
 FILLCELL_X1 FILLER_49_147 ();
 FILLCELL_X4 FILLER_49_155 ();
 FILLCELL_X2 FILLER_49_159 ();
 FILLCELL_X4 FILLER_49_165 ();
 FILLCELL_X4 FILLER_49_819 ();
 FILLCELL_X4 FILLER_49_827 ();
 FILLCELL_X2 FILLER_49_831 ();
 FILLCELL_X1 FILLER_49_833 ();
 FILLCELL_X4 FILLER_49_843 ();
 FILLCELL_X4 FILLER_49_851 ();
 FILLCELL_X2 FILLER_49_855 ();
 FILLCELL_X4 FILLER_49_866 ();
 FILLCELL_X8 FILLER_49_873 ();
 FILLCELL_X4 FILLER_49_881 ();
 FILLCELL_X2 FILLER_49_885 ();
 FILLCELL_X8 FILLER_49_891 ();
 FILLCELL_X1 FILLER_49_899 ();
 FILLCELL_X16 FILLER_49_904 ();
 FILLCELL_X2 FILLER_49_920 ();
 FILLCELL_X4 FILLER_49_925 ();
 FILLCELL_X4 FILLER_49_933 ();
 FILLCELL_X2 FILLER_49_937 ();
 FILLCELL_X1 FILLER_49_939 ();
 FILLCELL_X4 FILLER_49_949 ();
 FILLCELL_X8 FILLER_49_957 ();
 FILLCELL_X2 FILLER_49_965 ();
 FILLCELL_X1 FILLER_49_967 ();
 FILLCELL_X4 FILLER_49_970 ();
 FILLCELL_X1 FILLER_49_974 ();
 FILLCELL_X4 FILLER_49_977 ();
 FILLCELL_X2 FILLER_49_981 ();
 FILLCELL_X4 FILLER_49_989 ();
 FILLCELL_X1 FILLER_49_993 ();
 FILLCELL_X4 FILLER_49_1001 ();
 FILLCELL_X4 FILLER_49_1009 ();
 FILLCELL_X1 FILLER_49_1013 ();
 FILLCELL_X4 FILLER_49_1018 ();
 FILLCELL_X4 FILLER_50_1 ();
 FILLCELL_X32 FILLER_50_9 ();
 FILLCELL_X32 FILLER_50_41 ();
 FILLCELL_X16 FILLER_50_73 ();
 FILLCELL_X8 FILLER_50_89 ();
 FILLCELL_X2 FILLER_50_97 ();
 FILLCELL_X4 FILLER_50_102 ();
 FILLCELL_X8 FILLER_50_109 ();
 FILLCELL_X1 FILLER_50_117 ();
 FILLCELL_X4 FILLER_50_121 ();
 FILLCELL_X4 FILLER_50_128 ();
 FILLCELL_X8 FILLER_50_137 ();
 FILLCELL_X1 FILLER_50_145 ();
 FILLCELL_X4 FILLER_50_150 ();
 FILLCELL_X8 FILLER_50_159 ();
 FILLCELL_X2 FILLER_50_167 ();
 FILLCELL_X8 FILLER_50_819 ();
 FILLCELL_X4 FILLER_50_832 ();
 FILLCELL_X4 FILLER_50_845 ();
 FILLCELL_X8 FILLER_50_853 ();
 FILLCELL_X4 FILLER_50_861 ();
 FILLCELL_X2 FILLER_50_865 ();
 FILLCELL_X1 FILLER_50_867 ();
 FILLCELL_X4 FILLER_50_871 ();
 FILLCELL_X4 FILLER_50_884 ();
 FILLCELL_X1 FILLER_50_888 ();
 FILLCELL_X4 FILLER_50_895 ();
 FILLCELL_X8 FILLER_50_908 ();
 FILLCELL_X4 FILLER_50_916 ();
 FILLCELL_X1 FILLER_50_920 ();
 FILLCELL_X4 FILLER_50_925 ();
 FILLCELL_X8 FILLER_50_938 ();
 FILLCELL_X4 FILLER_50_946 ();
 FILLCELL_X1 FILLER_50_950 ();
 FILLCELL_X4 FILLER_50_961 ();
 FILLCELL_X4 FILLER_50_972 ();
 FILLCELL_X4 FILLER_50_983 ();
 FILLCELL_X2 FILLER_50_987 ();
 FILLCELL_X4 FILLER_50_991 ();
 FILLCELL_X4 FILLER_50_1005 ();
 FILLCELL_X8 FILLER_50_1013 ();
 FILLCELL_X1 FILLER_50_1021 ();
 FILLCELL_X32 FILLER_51_1 ();
 FILLCELL_X32 FILLER_51_33 ();
 FILLCELL_X32 FILLER_51_65 ();
 FILLCELL_X16 FILLER_51_97 ();
 FILLCELL_X4 FILLER_51_113 ();
 FILLCELL_X4 FILLER_51_119 ();
 FILLCELL_X4 FILLER_51_140 ();
 FILLCELL_X4 FILLER_51_148 ();
 FILLCELL_X2 FILLER_51_152 ();
 FILLCELL_X8 FILLER_51_159 ();
 FILLCELL_X2 FILLER_51_167 ();
 FILLCELL_X4 FILLER_51_819 ();
 FILLCELL_X8 FILLER_51_826 ();
 FILLCELL_X2 FILLER_51_834 ();
 FILLCELL_X4 FILLER_51_842 ();
 FILLCELL_X8 FILLER_51_850 ();
 FILLCELL_X4 FILLER_51_858 ();
 FILLCELL_X1 FILLER_51_862 ();
 FILLCELL_X4 FILLER_51_866 ();
 FILLCELL_X4 FILLER_51_880 ();
 FILLCELL_X1 FILLER_51_884 ();
 FILLCELL_X4 FILLER_51_888 ();
 FILLCELL_X4 FILLER_51_911 ();
 FILLCELL_X8 FILLER_51_919 ();
 FILLCELL_X2 FILLER_51_927 ();
 FILLCELL_X1 FILLER_51_929 ();
 FILLCELL_X16 FILLER_51_933 ();
 FILLCELL_X4 FILLER_51_952 ();
 FILLCELL_X4 FILLER_51_960 ();
 FILLCELL_X16 FILLER_51_974 ();
 FILLCELL_X2 FILLER_51_990 ();
 FILLCELL_X4 FILLER_51_996 ();
 FILLCELL_X4 FILLER_51_1006 ();
 FILLCELL_X4 FILLER_51_1016 ();
 FILLCELL_X2 FILLER_51_1020 ();
 FILLCELL_X32 FILLER_52_1 ();
 FILLCELL_X32 FILLER_52_33 ();
 FILLCELL_X32 FILLER_52_65 ();
 FILLCELL_X16 FILLER_52_97 ();
 FILLCELL_X8 FILLER_52_113 ();
 FILLCELL_X2 FILLER_52_121 ();
 FILLCELL_X1 FILLER_52_123 ();
 FILLCELL_X4 FILLER_52_127 ();
 FILLCELL_X4 FILLER_52_136 ();
 FILLCELL_X4 FILLER_52_145 ();
 FILLCELL_X4 FILLER_52_155 ();
 FILLCELL_X1 FILLER_52_159 ();
 FILLCELL_X4 FILLER_52_165 ();
 FILLCELL_X16 FILLER_52_819 ();
 FILLCELL_X4 FILLER_52_835 ();
 FILLCELL_X16 FILLER_52_842 ();
 FILLCELL_X4 FILLER_52_858 ();
 FILLCELL_X2 FILLER_52_862 ();
 FILLCELL_X1 FILLER_52_864 ();
 FILLCELL_X4 FILLER_52_874 ();
 FILLCELL_X4 FILLER_52_884 ();
 FILLCELL_X8 FILLER_52_892 ();
 FILLCELL_X16 FILLER_52_904 ();
 FILLCELL_X2 FILLER_52_920 ();
 FILLCELL_X1 FILLER_52_922 ();
 FILLCELL_X4 FILLER_52_927 ();
 FILLCELL_X16 FILLER_52_935 ();
 FILLCELL_X1 FILLER_52_951 ();
 FILLCELL_X8 FILLER_52_956 ();
 FILLCELL_X2 FILLER_52_964 ();
 FILLCELL_X4 FILLER_52_969 ();
 FILLCELL_X2 FILLER_52_973 ();
 FILLCELL_X4 FILLER_52_978 ();
 FILLCELL_X8 FILLER_52_986 ();
 FILLCELL_X8 FILLER_52_997 ();
 FILLCELL_X4 FILLER_52_1005 ();
 FILLCELL_X1 FILLER_52_1009 ();
 FILLCELL_X8 FILLER_52_1014 ();
 FILLCELL_X32 FILLER_53_1 ();
 FILLCELL_X32 FILLER_53_33 ();
 FILLCELL_X32 FILLER_53_65 ();
 FILLCELL_X16 FILLER_53_97 ();
 FILLCELL_X8 FILLER_53_113 ();
 FILLCELL_X4 FILLER_53_121 ();
 FILLCELL_X2 FILLER_53_125 ();
 FILLCELL_X4 FILLER_53_130 ();
 FILLCELL_X4 FILLER_53_140 ();
 FILLCELL_X2 FILLER_53_144 ();
 FILLCELL_X1 FILLER_53_146 ();
 FILLCELL_X4 FILLER_53_164 ();
 FILLCELL_X1 FILLER_53_168 ();
 FILLCELL_X16 FILLER_53_819 ();
 FILLCELL_X2 FILLER_53_835 ();
 FILLCELL_X4 FILLER_53_846 ();
 FILLCELL_X16 FILLER_53_853 ();
 FILLCELL_X1 FILLER_53_869 ();
 FILLCELL_X4 FILLER_53_875 ();
 FILLCELL_X8 FILLER_53_882 ();
 FILLCELL_X4 FILLER_53_890 ();
 FILLCELL_X2 FILLER_53_894 ();
 FILLCELL_X1 FILLER_53_896 ();
 FILLCELL_X16 FILLER_53_901 ();
 FILLCELL_X8 FILLER_53_921 ();
 FILLCELL_X4 FILLER_53_934 ();
 FILLCELL_X4 FILLER_53_943 ();
 FILLCELL_X2 FILLER_53_947 ();
 FILLCELL_X1 FILLER_53_949 ();
 FILLCELL_X4 FILLER_53_954 ();
 FILLCELL_X4 FILLER_53_967 ();
 FILLCELL_X2 FILLER_53_971 ();
 FILLCELL_X4 FILLER_53_976 ();
 FILLCELL_X2 FILLER_53_980 ();
 FILLCELL_X1 FILLER_53_982 ();
 FILLCELL_X8 FILLER_53_992 ();
 FILLCELL_X1 FILLER_53_1000 ();
 FILLCELL_X4 FILLER_53_1018 ();
 FILLCELL_X32 FILLER_54_1 ();
 FILLCELL_X32 FILLER_54_33 ();
 FILLCELL_X32 FILLER_54_65 ();
 FILLCELL_X16 FILLER_54_97 ();
 FILLCELL_X8 FILLER_54_113 ();
 FILLCELL_X4 FILLER_54_121 ();
 FILLCELL_X1 FILLER_54_125 ();
 FILLCELL_X4 FILLER_54_145 ();
 FILLCELL_X1 FILLER_54_149 ();
 FILLCELL_X4 FILLER_54_153 ();
 FILLCELL_X4 FILLER_54_162 ();
 FILLCELL_X2 FILLER_54_166 ();
 FILLCELL_X1 FILLER_54_168 ();
 FILLCELL_X8 FILLER_54_819 ();
 FILLCELL_X2 FILLER_54_827 ();
 FILLCELL_X4 FILLER_54_832 ();
 FILLCELL_X4 FILLER_54_845 ();
 FILLCELL_X4 FILLER_54_855 ();
 FILLCELL_X2 FILLER_54_859 ();
 FILLCELL_X4 FILLER_54_865 ();
 FILLCELL_X8 FILLER_54_873 ();
 FILLCELL_X4 FILLER_54_881 ();
 FILLCELL_X2 FILLER_54_885 ();
 FILLCELL_X4 FILLER_54_891 ();
 FILLCELL_X4 FILLER_54_904 ();
 FILLCELL_X8 FILLER_54_912 ();
 FILLCELL_X4 FILLER_54_927 ();
 FILLCELL_X8 FILLER_54_948 ();
 FILLCELL_X1 FILLER_54_956 ();
 FILLCELL_X4 FILLER_54_966 ();
 FILLCELL_X4 FILLER_54_973 ();
 FILLCELL_X4 FILLER_54_986 ();
 FILLCELL_X8 FILLER_54_1000 ();
 FILLCELL_X4 FILLER_54_1008 ();
 FILLCELL_X2 FILLER_54_1012 ();
 FILLCELL_X1 FILLER_54_1014 ();
 FILLCELL_X4 FILLER_54_1018 ();
 FILLCELL_X32 FILLER_55_1 ();
 FILLCELL_X32 FILLER_55_33 ();
 FILLCELL_X32 FILLER_55_65 ();
 FILLCELL_X32 FILLER_55_97 ();
 FILLCELL_X8 FILLER_55_129 ();
 FILLCELL_X2 FILLER_55_137 ();
 FILLCELL_X4 FILLER_55_142 ();
 FILLCELL_X2 FILLER_55_146 ();
 FILLCELL_X8 FILLER_55_151 ();
 FILLCELL_X2 FILLER_55_159 ();
 FILLCELL_X1 FILLER_55_161 ();
 FILLCELL_X4 FILLER_55_165 ();
 FILLCELL_X16 FILLER_55_819 ();
 FILLCELL_X4 FILLER_55_835 ();
 FILLCELL_X4 FILLER_55_844 ();
 FILLCELL_X4 FILLER_55_852 ();
 FILLCELL_X4 FILLER_55_860 ();
 FILLCELL_X2 FILLER_55_864 ();
 FILLCELL_X1 FILLER_55_866 ();
 FILLCELL_X4 FILLER_55_874 ();
 FILLCELL_X2 FILLER_55_878 ();
 FILLCELL_X4 FILLER_55_883 ();
 FILLCELL_X4 FILLER_55_892 ();
 FILLCELL_X4 FILLER_55_905 ();
 FILLCELL_X4 FILLER_55_913 ();
 FILLCELL_X4 FILLER_55_921 ();
 FILLCELL_X2 FILLER_55_925 ();
 FILLCELL_X1 FILLER_55_927 ();
 FILLCELL_X4 FILLER_55_932 ();
 FILLCELL_X16 FILLER_55_938 ();
 FILLCELL_X2 FILLER_55_954 ();
 FILLCELL_X1 FILLER_55_956 ();
 FILLCELL_X4 FILLER_55_961 ();
 FILLCELL_X2 FILLER_55_965 ();
 FILLCELL_X1 FILLER_55_967 ();
 FILLCELL_X4 FILLER_55_972 ();
 FILLCELL_X4 FILLER_55_979 ();
 FILLCELL_X4 FILLER_55_986 ();
 FILLCELL_X1 FILLER_55_990 ();
 FILLCELL_X4 FILLER_55_995 ();
 FILLCELL_X4 FILLER_55_1018 ();
 FILLCELL_X32 FILLER_56_1 ();
 FILLCELL_X32 FILLER_56_33 ();
 FILLCELL_X32 FILLER_56_65 ();
 FILLCELL_X32 FILLER_56_97 ();
 FILLCELL_X32 FILLER_56_129 ();
 FILLCELL_X1 FILLER_56_161 ();
 FILLCELL_X4 FILLER_56_165 ();
 FILLCELL_X4 FILLER_56_819 ();
 FILLCELL_X2 FILLER_56_823 ();
 FILLCELL_X4 FILLER_56_830 ();
 FILLCELL_X8 FILLER_56_838 ();
 FILLCELL_X1 FILLER_56_846 ();
 FILLCELL_X4 FILLER_56_850 ();
 FILLCELL_X2 FILLER_56_854 ();
 FILLCELL_X4 FILLER_56_862 ();
 FILLCELL_X16 FILLER_56_875 ();
 FILLCELL_X4 FILLER_56_891 ();
 FILLCELL_X1 FILLER_56_895 ();
 FILLCELL_X4 FILLER_56_905 ();
 FILLCELL_X8 FILLER_56_912 ();
 FILLCELL_X4 FILLER_56_920 ();
 FILLCELL_X2 FILLER_56_924 ();
 FILLCELL_X8 FILLER_56_930 ();
 FILLCELL_X16 FILLER_56_942 ();
 FILLCELL_X2 FILLER_56_958 ();
 FILLCELL_X4 FILLER_56_964 ();
 FILLCELL_X32 FILLER_56_971 ();
 FILLCELL_X16 FILLER_56_1003 ();
 FILLCELL_X2 FILLER_56_1019 ();
 FILLCELL_X1 FILLER_56_1021 ();
 FILLCELL_X32 FILLER_57_1 ();
 FILLCELL_X32 FILLER_57_33 ();
 FILLCELL_X32 FILLER_57_65 ();
 FILLCELL_X32 FILLER_57_97 ();
 FILLCELL_X4 FILLER_57_129 ();
 FILLCELL_X1 FILLER_57_133 ();
 FILLCELL_X4 FILLER_57_138 ();
 FILLCELL_X8 FILLER_57_161 ();
 FILLCELL_X8 FILLER_57_819 ();
 FILLCELL_X4 FILLER_57_846 ();
 FILLCELL_X1 FILLER_57_850 ();
 FILLCELL_X4 FILLER_57_861 ();
 FILLCELL_X1 FILLER_57_865 ();
 FILLCELL_X4 FILLER_57_871 ();
 FILLCELL_X4 FILLER_57_879 ();
 FILLCELL_X4 FILLER_57_886 ();
 FILLCELL_X4 FILLER_57_893 ();
 FILLCELL_X16 FILLER_57_903 ();
 FILLCELL_X4 FILLER_57_923 ();
 FILLCELL_X4 FILLER_57_936 ();
 FILLCELL_X1 FILLER_57_940 ();
 FILLCELL_X4 FILLER_57_945 ();
 FILLCELL_X2 FILLER_57_949 ();
 FILLCELL_X1 FILLER_57_951 ();
 FILLCELL_X4 FILLER_57_956 ();
 FILLCELL_X4 FILLER_57_969 ();
 FILLCELL_X4 FILLER_57_977 ();
 FILLCELL_X32 FILLER_57_985 ();
 FILLCELL_X4 FILLER_57_1017 ();
 FILLCELL_X1 FILLER_57_1021 ();
 FILLCELL_X32 FILLER_58_1 ();
 FILLCELL_X32 FILLER_58_33 ();
 FILLCELL_X32 FILLER_58_65 ();
 FILLCELL_X32 FILLER_58_97 ();
 FILLCELL_X16 FILLER_58_129 ();
 FILLCELL_X4 FILLER_58_145 ();
 FILLCELL_X2 FILLER_58_149 ();
 FILLCELL_X8 FILLER_58_155 ();
 FILLCELL_X4 FILLER_58_163 ();
 FILLCELL_X2 FILLER_58_167 ();
 FILLCELL_X4 FILLER_58_819 ();
 FILLCELL_X2 FILLER_58_823 ();
 FILLCELL_X4 FILLER_58_830 ();
 FILLCELL_X2 FILLER_58_834 ();
 FILLCELL_X1 FILLER_58_836 ();
 FILLCELL_X16 FILLER_58_840 ();
 FILLCELL_X8 FILLER_58_856 ();
 FILLCELL_X4 FILLER_58_864 ();
 FILLCELL_X16 FILLER_58_874 ();
 FILLCELL_X8 FILLER_58_890 ();
 FILLCELL_X2 FILLER_58_898 ();
 FILLCELL_X4 FILLER_58_905 ();
 FILLCELL_X8 FILLER_58_912 ();
 FILLCELL_X1 FILLER_58_920 ();
 FILLCELL_X4 FILLER_58_926 ();
 FILLCELL_X4 FILLER_58_939 ();
 FILLCELL_X4 FILLER_58_946 ();
 FILLCELL_X4 FILLER_58_955 ();
 FILLCELL_X4 FILLER_58_968 ();
 FILLCELL_X4 FILLER_58_981 ();
 FILLCELL_X1 FILLER_58_985 ();
 FILLCELL_X32 FILLER_58_990 ();
 FILLCELL_X32 FILLER_59_1 ();
 FILLCELL_X32 FILLER_59_33 ();
 FILLCELL_X32 FILLER_59_65 ();
 FILLCELL_X32 FILLER_59_97 ();
 FILLCELL_X8 FILLER_59_129 ();
 FILLCELL_X4 FILLER_59_137 ();
 FILLCELL_X8 FILLER_59_160 ();
 FILLCELL_X1 FILLER_59_168 ();
 FILLCELL_X16 FILLER_59_819 ();
 FILLCELL_X4 FILLER_59_835 ();
 FILLCELL_X4 FILLER_59_845 ();
 FILLCELL_X8 FILLER_59_852 ();
 FILLCELL_X4 FILLER_59_860 ();
 FILLCELL_X2 FILLER_59_864 ();
 FILLCELL_X4 FILLER_59_875 ();
 FILLCELL_X4 FILLER_59_882 ();
 FILLCELL_X2 FILLER_59_886 ();
 FILLCELL_X4 FILLER_59_891 ();
 FILLCELL_X4 FILLER_59_904 ();
 FILLCELL_X4 FILLER_59_917 ();
 FILLCELL_X4 FILLER_59_924 ();
 FILLCELL_X2 FILLER_59_928 ();
 FILLCELL_X1 FILLER_59_930 ();
 FILLCELL_X4 FILLER_59_937 ();
 FILLCELL_X4 FILLER_59_945 ();
 FILLCELL_X2 FILLER_59_949 ();
 FILLCELL_X1 FILLER_59_951 ();
 FILLCELL_X4 FILLER_59_955 ();
 FILLCELL_X4 FILLER_59_965 ();
 FILLCELL_X4 FILLER_59_974 ();
 FILLCELL_X1 FILLER_59_978 ();
 FILLCELL_X16 FILLER_59_998 ();
 FILLCELL_X1 FILLER_59_1014 ();
 FILLCELL_X4 FILLER_59_1018 ();
 FILLCELL_X32 FILLER_60_1 ();
 FILLCELL_X32 FILLER_60_33 ();
 FILLCELL_X32 FILLER_60_65 ();
 FILLCELL_X32 FILLER_60_97 ();
 FILLCELL_X8 FILLER_60_129 ();
 FILLCELL_X4 FILLER_60_137 ();
 FILLCELL_X2 FILLER_60_141 ();
 FILLCELL_X1 FILLER_60_143 ();
 FILLCELL_X4 FILLER_60_148 ();
 FILLCELL_X8 FILLER_60_155 ();
 FILLCELL_X4 FILLER_60_163 ();
 FILLCELL_X2 FILLER_60_167 ();
 FILLCELL_X4 FILLER_60_819 ();
 FILLCELL_X8 FILLER_60_828 ();
 FILLCELL_X1 FILLER_60_836 ();
 FILLCELL_X4 FILLER_60_846 ();
 FILLCELL_X8 FILLER_60_855 ();
 FILLCELL_X4 FILLER_60_863 ();
 FILLCELL_X2 FILLER_60_867 ();
 FILLCELL_X1 FILLER_60_869 ();
 FILLCELL_X4 FILLER_60_873 ();
 FILLCELL_X8 FILLER_60_884 ();
 FILLCELL_X4 FILLER_60_892 ();
 FILLCELL_X2 FILLER_60_896 ();
 FILLCELL_X4 FILLER_60_904 ();
 FILLCELL_X16 FILLER_60_912 ();
 FILLCELL_X8 FILLER_60_928 ();
 FILLCELL_X2 FILLER_60_936 ();
 FILLCELL_X32 FILLER_60_943 ();
 FILLCELL_X4 FILLER_60_975 ();
 FILLCELL_X1 FILLER_60_979 ();
 FILLCELL_X4 FILLER_60_984 ();
 FILLCELL_X4 FILLER_60_992 ();
 FILLCELL_X4 FILLER_60_1000 ();
 FILLCELL_X8 FILLER_60_1013 ();
 FILLCELL_X1 FILLER_60_1021 ();
 FILLCELL_X4 FILLER_61_1 ();
 FILLCELL_X32 FILLER_61_8 ();
 FILLCELL_X32 FILLER_61_40 ();
 FILLCELL_X32 FILLER_61_72 ();
 FILLCELL_X32 FILLER_61_104 ();
 FILLCELL_X4 FILLER_61_136 ();
 FILLCELL_X2 FILLER_61_140 ();
 FILLCELL_X8 FILLER_61_161 ();
 FILLCELL_X4 FILLER_61_819 ();
 FILLCELL_X2 FILLER_61_823 ();
 FILLCELL_X1 FILLER_61_825 ();
 FILLCELL_X4 FILLER_61_830 ();
 FILLCELL_X4 FILLER_61_843 ();
 FILLCELL_X4 FILLER_61_852 ();
 FILLCELL_X4 FILLER_61_860 ();
 FILLCELL_X4 FILLER_61_868 ();
 FILLCELL_X4 FILLER_61_876 ();
 FILLCELL_X2 FILLER_61_880 ();
 FILLCELL_X1 FILLER_61_882 ();
 FILLCELL_X4 FILLER_61_889 ();
 FILLCELL_X8 FILLER_61_899 ();
 FILLCELL_X2 FILLER_61_907 ();
 FILLCELL_X1 FILLER_61_909 ();
 FILLCELL_X8 FILLER_61_929 ();
 FILLCELL_X4 FILLER_61_937 ();
 FILLCELL_X2 FILLER_61_941 ();
 FILLCELL_X4 FILLER_61_952 ();
 FILLCELL_X4 FILLER_61_965 ();
 FILLCELL_X2 FILLER_61_969 ();
 FILLCELL_X8 FILLER_61_975 ();
 FILLCELL_X1 FILLER_61_983 ();
 FILLCELL_X4 FILLER_61_989 ();
 FILLCELL_X4 FILLER_61_1002 ();
 FILLCELL_X4 FILLER_61_1015 ();
 FILLCELL_X2 FILLER_61_1019 ();
 FILLCELL_X1 FILLER_61_1021 ();
 FILLCELL_X32 FILLER_62_1 ();
 FILLCELL_X32 FILLER_62_33 ();
 FILLCELL_X32 FILLER_62_65 ();
 FILLCELL_X32 FILLER_62_97 ();
 FILLCELL_X16 FILLER_62_129 ();
 FILLCELL_X1 FILLER_62_145 ();
 FILLCELL_X8 FILLER_62_150 ();
 FILLCELL_X4 FILLER_62_158 ();
 FILLCELL_X4 FILLER_62_165 ();
 FILLCELL_X8 FILLER_62_819 ();
 FILLCELL_X4 FILLER_62_827 ();
 FILLCELL_X2 FILLER_62_831 ();
 FILLCELL_X4 FILLER_62_837 ();
 FILLCELL_X16 FILLER_62_845 ();
 FILLCELL_X4 FILLER_62_870 ();
 FILLCELL_X4 FILLER_62_878 ();
 FILLCELL_X4 FILLER_62_885 ();
 FILLCELL_X2 FILLER_62_889 ();
 FILLCELL_X8 FILLER_62_894 ();
 FILLCELL_X4 FILLER_62_906 ();
 FILLCELL_X8 FILLER_62_913 ();
 FILLCELL_X4 FILLER_62_921 ();
 FILLCELL_X2 FILLER_62_925 ();
 FILLCELL_X4 FILLER_62_931 ();
 FILLCELL_X4 FILLER_62_938 ();
 FILLCELL_X4 FILLER_62_951 ();
 FILLCELL_X4 FILLER_62_961 ();
 FILLCELL_X16 FILLER_62_969 ();
 FILLCELL_X4 FILLER_62_985 ();
 FILLCELL_X2 FILLER_62_989 ();
 FILLCELL_X4 FILLER_62_994 ();
 FILLCELL_X4 FILLER_62_1002 ();
 FILLCELL_X8 FILLER_62_1012 ();
 FILLCELL_X2 FILLER_62_1020 ();
 FILLCELL_X32 FILLER_63_1 ();
 FILLCELL_X32 FILLER_63_33 ();
 FILLCELL_X32 FILLER_63_65 ();
 FILLCELL_X32 FILLER_63_97 ();
 FILLCELL_X8 FILLER_63_129 ();
 FILLCELL_X4 FILLER_63_137 ();
 FILLCELL_X2 FILLER_63_141 ();
 FILLCELL_X4 FILLER_63_162 ();
 FILLCELL_X2 FILLER_63_166 ();
 FILLCELL_X1 FILLER_63_168 ();
 FILLCELL_X16 FILLER_63_819 ();
 FILLCELL_X16 FILLER_63_839 ();
 FILLCELL_X1 FILLER_63_855 ();
 FILLCELL_X4 FILLER_63_859 ();
 FILLCELL_X8 FILLER_63_869 ();
 FILLCELL_X1 FILLER_63_877 ();
 FILLCELL_X4 FILLER_63_882 ();
 FILLCELL_X4 FILLER_63_889 ();
 FILLCELL_X2 FILLER_63_893 ();
 FILLCELL_X1 FILLER_63_895 ();
 FILLCELL_X8 FILLER_63_905 ();
 FILLCELL_X4 FILLER_63_913 ();
 FILLCELL_X2 FILLER_63_917 ();
 FILLCELL_X4 FILLER_63_923 ();
 FILLCELL_X4 FILLER_63_934 ();
 FILLCELL_X4 FILLER_63_944 ();
 FILLCELL_X4 FILLER_63_953 ();
 FILLCELL_X4 FILLER_63_963 ();
 FILLCELL_X1 FILLER_63_967 ();
 FILLCELL_X4 FILLER_63_972 ();
 FILLCELL_X4 FILLER_63_980 ();
 FILLCELL_X1 FILLER_63_984 ();
 FILLCELL_X16 FILLER_63_991 ();
 FILLCELL_X8 FILLER_63_1007 ();
 FILLCELL_X4 FILLER_63_1015 ();
 FILLCELL_X2 FILLER_63_1019 ();
 FILLCELL_X1 FILLER_63_1021 ();
 FILLCELL_X32 FILLER_64_1 ();
 FILLCELL_X32 FILLER_64_33 ();
 FILLCELL_X32 FILLER_64_65 ();
 FILLCELL_X32 FILLER_64_97 ();
 FILLCELL_X16 FILLER_64_129 ();
 FILLCELL_X8 FILLER_64_145 ();
 FILLCELL_X4 FILLER_64_156 ();
 FILLCELL_X2 FILLER_64_160 ();
 FILLCELL_X4 FILLER_64_165 ();
 FILLCELL_X32 FILLER_64_819 ();
 FILLCELL_X4 FILLER_64_851 ();
 FILLCELL_X4 FILLER_64_864 ();
 FILLCELL_X8 FILLER_64_877 ();
 FILLCELL_X1 FILLER_64_885 ();
 FILLCELL_X4 FILLER_64_891 ();
 FILLCELL_X4 FILLER_64_904 ();
 FILLCELL_X4 FILLER_64_914 ();
 FILLCELL_X32 FILLER_64_921 ();
 FILLCELL_X4 FILLER_64_957 ();
 FILLCELL_X4 FILLER_64_964 ();
 FILLCELL_X4 FILLER_64_973 ();
 FILLCELL_X4 FILLER_64_986 ();
 FILLCELL_X8 FILLER_64_999 ();
 FILLCELL_X8 FILLER_64_1011 ();
 FILLCELL_X2 FILLER_64_1019 ();
 FILLCELL_X1 FILLER_64_1021 ();
 FILLCELL_X32 FILLER_65_1 ();
 FILLCELL_X32 FILLER_65_33 ();
 FILLCELL_X32 FILLER_65_65 ();
 FILLCELL_X32 FILLER_65_97 ();
 FILLCELL_X32 FILLER_65_129 ();
 FILLCELL_X1 FILLER_65_161 ();
 FILLCELL_X4 FILLER_65_165 ();
 FILLCELL_X4 FILLER_65_819 ();
 FILLCELL_X2 FILLER_65_823 ();
 FILLCELL_X1 FILLER_65_825 ();
 FILLCELL_X4 FILLER_65_830 ();
 FILLCELL_X4 FILLER_65_843 ();
 FILLCELL_X8 FILLER_65_850 ();
 FILLCELL_X4 FILLER_65_863 ();
 FILLCELL_X8 FILLER_65_871 ();
 FILLCELL_X8 FILLER_65_883 ();
 FILLCELL_X4 FILLER_65_891 ();
 FILLCELL_X1 FILLER_65_895 ();
 FILLCELL_X4 FILLER_65_899 ();
 FILLCELL_X16 FILLER_65_907 ();
 FILLCELL_X4 FILLER_65_923 ();
 FILLCELL_X2 FILLER_65_927 ();
 FILLCELL_X16 FILLER_65_934 ();
 FILLCELL_X1 FILLER_65_950 ();
 FILLCELL_X4 FILLER_65_956 ();
 FILLCELL_X8 FILLER_65_963 ();
 FILLCELL_X2 FILLER_65_971 ();
 FILLCELL_X1 FILLER_65_973 ();
 FILLCELL_X8 FILLER_65_977 ();
 FILLCELL_X8 FILLER_65_989 ();
 FILLCELL_X2 FILLER_65_997 ();
 FILLCELL_X4 FILLER_65_1018 ();
 FILLCELL_X32 FILLER_66_1 ();
 FILLCELL_X32 FILLER_66_33 ();
 FILLCELL_X32 FILLER_66_65 ();
 FILLCELL_X32 FILLER_66_97 ();
 FILLCELL_X32 FILLER_66_129 ();
 FILLCELL_X8 FILLER_66_161 ();
 FILLCELL_X8 FILLER_66_819 ();
 FILLCELL_X1 FILLER_66_827 ();
 FILLCELL_X4 FILLER_66_831 ();
 FILLCELL_X4 FILLER_66_844 ();
 FILLCELL_X4 FILLER_66_854 ();
 FILLCELL_X8 FILLER_66_861 ();
 FILLCELL_X2 FILLER_66_869 ();
 FILLCELL_X8 FILLER_66_874 ();
 FILLCELL_X1 FILLER_66_882 ();
 FILLCELL_X4 FILLER_66_888 ();
 FILLCELL_X4 FILLER_66_895 ();
 FILLCELL_X8 FILLER_66_902 ();
 FILLCELL_X1 FILLER_66_910 ();
 FILLCELL_X4 FILLER_66_915 ();
 FILLCELL_X4 FILLER_66_928 ();
 FILLCELL_X4 FILLER_66_936 ();
 FILLCELL_X4 FILLER_66_943 ();
 FILLCELL_X2 FILLER_66_947 ();
 FILLCELL_X1 FILLER_66_949 ();
 FILLCELL_X4 FILLER_66_959 ();
 FILLCELL_X4 FILLER_66_972 ();
 FILLCELL_X4 FILLER_66_979 ();
 FILLCELL_X2 FILLER_66_983 ();
 FILLCELL_X1 FILLER_66_985 ();
 FILLCELL_X4 FILLER_66_990 ();
 FILLCELL_X4 FILLER_66_997 ();
 FILLCELL_X8 FILLER_66_1004 ();
 FILLCELL_X2 FILLER_66_1012 ();
 FILLCELL_X1 FILLER_66_1014 ();
 FILLCELL_X4 FILLER_66_1018 ();
 FILLCELL_X32 FILLER_67_1 ();
 FILLCELL_X32 FILLER_67_33 ();
 FILLCELL_X32 FILLER_67_65 ();
 FILLCELL_X32 FILLER_67_97 ();
 FILLCELL_X32 FILLER_67_129 ();
 FILLCELL_X8 FILLER_67_161 ();
 FILLCELL_X8 FILLER_67_819 ();
 FILLCELL_X1 FILLER_67_827 ();
 FILLCELL_X4 FILLER_67_832 ();
 FILLCELL_X4 FILLER_67_841 ();
 FILLCELL_X16 FILLER_67_849 ();
 FILLCELL_X4 FILLER_67_865 ();
 FILLCELL_X2 FILLER_67_869 ();
 FILLCELL_X4 FILLER_67_875 ();
 FILLCELL_X4 FILLER_67_888 ();
 FILLCELL_X4 FILLER_67_898 ();
 FILLCELL_X4 FILLER_67_907 ();
 FILLCELL_X2 FILLER_67_911 ();
 FILLCELL_X4 FILLER_67_917 ();
 FILLCELL_X4 FILLER_67_930 ();
 FILLCELL_X4 FILLER_67_940 ();
 FILLCELL_X1 FILLER_67_944 ();
 FILLCELL_X4 FILLER_67_948 ();
 FILLCELL_X2 FILLER_67_952 ();
 FILLCELL_X4 FILLER_67_960 ();
 FILLCELL_X4 FILLER_67_968 ();
 FILLCELL_X1 FILLER_67_972 ();
 FILLCELL_X8 FILLER_67_979 ();
 FILLCELL_X2 FILLER_67_987 ();
 FILLCELL_X4 FILLER_67_993 ();
 FILLCELL_X2 FILLER_67_997 ();
 FILLCELL_X4 FILLER_67_1018 ();
 FILLCELL_X32 FILLER_68_1 ();
 FILLCELL_X32 FILLER_68_33 ();
 FILLCELL_X32 FILLER_68_65 ();
 FILLCELL_X32 FILLER_68_97 ();
 FILLCELL_X16 FILLER_68_129 ();
 FILLCELL_X8 FILLER_68_145 ();
 FILLCELL_X4 FILLER_68_153 ();
 FILLCELL_X2 FILLER_68_157 ();
 FILLCELL_X1 FILLER_68_159 ();
 FILLCELL_X4 FILLER_68_163 ();
 FILLCELL_X2 FILLER_68_167 ();
 FILLCELL_X8 FILLER_68_819 ();
 FILLCELL_X4 FILLER_68_827 ();
 FILLCELL_X2 FILLER_68_831 ();
 FILLCELL_X4 FILLER_68_837 ();
 FILLCELL_X8 FILLER_68_845 ();
 FILLCELL_X4 FILLER_68_853 ();
 FILLCELL_X2 FILLER_68_857 ();
 FILLCELL_X1 FILLER_68_859 ();
 FILLCELL_X4 FILLER_68_865 ();
 FILLCELL_X8 FILLER_68_872 ();
 FILLCELL_X4 FILLER_68_880 ();
 FILLCELL_X8 FILLER_68_893 ();
 FILLCELL_X4 FILLER_68_905 ();
 FILLCELL_X8 FILLER_68_913 ();
 FILLCELL_X4 FILLER_68_930 ();
 FILLCELL_X4 FILLER_68_938 ();
 FILLCELL_X4 FILLER_68_945 ();
 FILLCELL_X2 FILLER_68_949 ();
 FILLCELL_X4 FILLER_68_954 ();
 FILLCELL_X2 FILLER_68_958 ();
 FILLCELL_X4 FILLER_68_963 ();
 FILLCELL_X4 FILLER_68_974 ();
 FILLCELL_X4 FILLER_68_984 ();
 FILLCELL_X4 FILLER_68_991 ();
 FILLCELL_X2 FILLER_68_995 ();
 FILLCELL_X4 FILLER_68_1006 ();
 FILLCELL_X8 FILLER_68_1013 ();
 FILLCELL_X1 FILLER_68_1021 ();
 FILLCELL_X32 FILLER_69_1 ();
 FILLCELL_X32 FILLER_69_33 ();
 FILLCELL_X32 FILLER_69_65 ();
 FILLCELL_X32 FILLER_69_97 ();
 FILLCELL_X32 FILLER_69_129 ();
 FILLCELL_X8 FILLER_69_161 ();
 FILLCELL_X16 FILLER_69_819 ();
 FILLCELL_X8 FILLER_69_835 ();
 FILLCELL_X2 FILLER_69_843 ();
 FILLCELL_X4 FILLER_69_849 ();
 FILLCELL_X1 FILLER_69_853 ();
 FILLCELL_X4 FILLER_69_863 ();
 FILLCELL_X4 FILLER_69_873 ();
 FILLCELL_X8 FILLER_69_880 ();
 FILLCELL_X4 FILLER_69_888 ();
 FILLCELL_X2 FILLER_69_892 ();
 FILLCELL_X1 FILLER_69_894 ();
 FILLCELL_X8 FILLER_69_899 ();
 FILLCELL_X4 FILLER_69_916 ();
 FILLCELL_X8 FILLER_69_924 ();
 FILLCELL_X4 FILLER_69_932 ();
 FILLCELL_X4 FILLER_69_941 ();
 FILLCELL_X4 FILLER_69_950 ();
 FILLCELL_X8 FILLER_69_958 ();
 FILLCELL_X4 FILLER_69_966 ();
 FILLCELL_X8 FILLER_69_973 ();
 FILLCELL_X4 FILLER_69_981 ();
 FILLCELL_X2 FILLER_69_985 ();
 FILLCELL_X1 FILLER_69_987 ();
 FILLCELL_X4 FILLER_69_993 ();
 FILLCELL_X4 FILLER_69_1006 ();
 FILLCELL_X4 FILLER_69_1016 ();
 FILLCELL_X2 FILLER_69_1020 ();
 FILLCELL_X32 FILLER_70_1 ();
 FILLCELL_X32 FILLER_70_33 ();
 FILLCELL_X32 FILLER_70_65 ();
 FILLCELL_X32 FILLER_70_97 ();
 FILLCELL_X32 FILLER_70_129 ();
 FILLCELL_X8 FILLER_70_161 ();
 FILLCELL_X8 FILLER_70_819 ();
 FILLCELL_X4 FILLER_70_827 ();
 FILLCELL_X2 FILLER_70_831 ();
 FILLCELL_X4 FILLER_70_837 ();
 FILLCELL_X4 FILLER_70_845 ();
 FILLCELL_X4 FILLER_70_858 ();
 FILLCELL_X4 FILLER_70_871 ();
 FILLCELL_X2 FILLER_70_875 ();
 FILLCELL_X1 FILLER_70_877 ();
 FILLCELL_X4 FILLER_70_882 ();
 FILLCELL_X4 FILLER_70_889 ();
 FILLCELL_X32 FILLER_70_896 ();
 FILLCELL_X8 FILLER_70_928 ();
 FILLCELL_X4 FILLER_70_945 ();
 FILLCELL_X4 FILLER_70_955 ();
 FILLCELL_X8 FILLER_70_964 ();
 FILLCELL_X4 FILLER_70_972 ();
 FILLCELL_X1 FILLER_70_976 ();
 FILLCELL_X4 FILLER_70_981 ();
 FILLCELL_X2 FILLER_70_985 ();
 FILLCELL_X4 FILLER_70_990 ();
 FILLCELL_X4 FILLER_70_998 ();
 FILLCELL_X4 FILLER_70_1005 ();
 FILLCELL_X2 FILLER_70_1009 ();
 FILLCELL_X1 FILLER_70_1011 ();
 FILLCELL_X4 FILLER_70_1018 ();
 FILLCELL_X4 FILLER_71_1 ();
 FILLCELL_X32 FILLER_71_8 ();
 FILLCELL_X32 FILLER_71_40 ();
 FILLCELL_X32 FILLER_71_72 ();
 FILLCELL_X32 FILLER_71_104 ();
 FILLCELL_X16 FILLER_71_136 ();
 FILLCELL_X4 FILLER_71_156 ();
 FILLCELL_X2 FILLER_71_160 ();
 FILLCELL_X4 FILLER_71_165 ();
 FILLCELL_X16 FILLER_71_819 ();
 FILLCELL_X8 FILLER_71_835 ();
 FILLCELL_X4 FILLER_71_843 ();
 FILLCELL_X4 FILLER_71_851 ();
 FILLCELL_X8 FILLER_71_859 ();
 FILLCELL_X4 FILLER_71_867 ();
 FILLCELL_X4 FILLER_71_875 ();
 FILLCELL_X4 FILLER_71_888 ();
 FILLCELL_X8 FILLER_71_897 ();
 FILLCELL_X4 FILLER_71_905 ();
 FILLCELL_X16 FILLER_71_913 ();
 FILLCELL_X2 FILLER_71_929 ();
 FILLCELL_X1 FILLER_71_931 ();
 FILLCELL_X4 FILLER_71_934 ();
 FILLCELL_X8 FILLER_71_947 ();
 FILLCELL_X4 FILLER_71_961 ();
 FILLCELL_X4 FILLER_71_968 ();
 FILLCELL_X2 FILLER_71_972 ();
 FILLCELL_X1 FILLER_71_974 ();
 FILLCELL_X4 FILLER_71_980 ();
 FILLCELL_X8 FILLER_71_993 ();
 FILLCELL_X8 FILLER_71_1010 ();
 FILLCELL_X4 FILLER_71_1018 ();
 FILLCELL_X32 FILLER_72_1 ();
 FILLCELL_X32 FILLER_72_33 ();
 FILLCELL_X32 FILLER_72_65 ();
 FILLCELL_X32 FILLER_72_97 ();
 FILLCELL_X8 FILLER_72_129 ();
 FILLCELL_X4 FILLER_72_137 ();
 FILLCELL_X2 FILLER_72_141 ();
 FILLCELL_X4 FILLER_72_162 ();
 FILLCELL_X2 FILLER_72_166 ();
 FILLCELL_X1 FILLER_72_168 ();
 FILLCELL_X16 FILLER_72_819 ();
 FILLCELL_X16 FILLER_72_839 ();
 FILLCELL_X8 FILLER_72_855 ();
 FILLCELL_X4 FILLER_72_863 ();
 FILLCELL_X2 FILLER_72_867 ();
 FILLCELL_X8 FILLER_72_873 ();
 FILLCELL_X4 FILLER_72_890 ();
 FILLCELL_X4 FILLER_72_900 ();
 FILLCELL_X2 FILLER_72_904 ();
 FILLCELL_X1 FILLER_72_906 ();
 FILLCELL_X4 FILLER_72_911 ();
 FILLCELL_X1 FILLER_72_915 ();
 FILLCELL_X4 FILLER_72_925 ();
 FILLCELL_X4 FILLER_72_932 ();
 FILLCELL_X4 FILLER_72_939 ();
 FILLCELL_X8 FILLER_72_953 ();
 FILLCELL_X1 FILLER_72_961 ();
 FILLCELL_X4 FILLER_72_969 ();
 FILLCELL_X8 FILLER_72_977 ();
 FILLCELL_X4 FILLER_72_994 ();
 FILLCELL_X1 FILLER_72_998 ();
 FILLCELL_X4 FILLER_72_1018 ();
 FILLCELL_X32 FILLER_73_1 ();
 FILLCELL_X32 FILLER_73_33 ();
 FILLCELL_X32 FILLER_73_65 ();
 FILLCELL_X32 FILLER_73_97 ();
 FILLCELL_X16 FILLER_73_129 ();
 FILLCELL_X8 FILLER_73_145 ();
 FILLCELL_X2 FILLER_73_153 ();
 FILLCELL_X4 FILLER_73_158 ();
 FILLCELL_X4 FILLER_73_165 ();
 FILLCELL_X4 FILLER_73_819 ();
 FILLCELL_X2 FILLER_73_823 ();
 FILLCELL_X1 FILLER_73_825 ();
 FILLCELL_X4 FILLER_73_830 ();
 FILLCELL_X4 FILLER_73_843 ();
 FILLCELL_X16 FILLER_73_851 ();
 FILLCELL_X8 FILLER_73_867 ();
 FILLCELL_X4 FILLER_73_875 ();
 FILLCELL_X8 FILLER_73_883 ();
 FILLCELL_X1 FILLER_73_891 ();
 FILLCELL_X4 FILLER_73_897 ();
 FILLCELL_X8 FILLER_73_905 ();
 FILLCELL_X4 FILLER_73_922 ();
 FILLCELL_X4 FILLER_73_932 ();
 FILLCELL_X8 FILLER_73_941 ();
 FILLCELL_X4 FILLER_73_949 ();
 FILLCELL_X2 FILLER_73_953 ();
 FILLCELL_X1 FILLER_73_955 ();
 FILLCELL_X16 FILLER_73_960 ();
 FILLCELL_X4 FILLER_73_980 ();
 FILLCELL_X8 FILLER_73_988 ();
 FILLCELL_X1 FILLER_73_996 ();
 FILLCELL_X4 FILLER_73_1001 ();
 FILLCELL_X8 FILLER_73_1008 ();
 FILLCELL_X4 FILLER_73_1016 ();
 FILLCELL_X2 FILLER_73_1020 ();
 FILLCELL_X32 FILLER_74_1 ();
 FILLCELL_X32 FILLER_74_33 ();
 FILLCELL_X32 FILLER_74_65 ();
 FILLCELL_X32 FILLER_74_97 ();
 FILLCELL_X32 FILLER_74_129 ();
 FILLCELL_X8 FILLER_74_161 ();
 FILLCELL_X8 FILLER_74_819 ();
 FILLCELL_X4 FILLER_74_832 ();
 FILLCELL_X4 FILLER_74_845 ();
 FILLCELL_X8 FILLER_74_853 ();
 FILLCELL_X4 FILLER_74_865 ();
 FILLCELL_X8 FILLER_74_873 ();
 FILLCELL_X4 FILLER_74_881 ();
 FILLCELL_X4 FILLER_74_889 ();
 FILLCELL_X2 FILLER_74_893 ();
 FILLCELL_X1 FILLER_74_895 ();
 FILLCELL_X4 FILLER_74_900 ();
 FILLCELL_X2 FILLER_74_904 ();
 FILLCELL_X1 FILLER_74_906 ();
 FILLCELL_X4 FILLER_74_911 ();
 FILLCELL_X4 FILLER_74_920 ();
 FILLCELL_X8 FILLER_74_928 ();
 FILLCELL_X4 FILLER_74_936 ();
 FILLCELL_X2 FILLER_74_940 ();
 FILLCELL_X4 FILLER_74_945 ();
 FILLCELL_X2 FILLER_74_949 ();
 FILLCELL_X1 FILLER_74_951 ();
 FILLCELL_X4 FILLER_74_957 ();
 FILLCELL_X8 FILLER_74_964 ();
 FILLCELL_X2 FILLER_74_972 ();
 FILLCELL_X1 FILLER_74_974 ();
 FILLCELL_X8 FILLER_74_979 ();
 FILLCELL_X4 FILLER_74_987 ();
 FILLCELL_X4 FILLER_74_994 ();
 FILLCELL_X2 FILLER_74_998 ();
 FILLCELL_X1 FILLER_74_1000 ();
 FILLCELL_X4 FILLER_74_1007 ();
 FILLCELL_X8 FILLER_74_1014 ();
 FILLCELL_X32 FILLER_75_1 ();
 FILLCELL_X32 FILLER_75_33 ();
 FILLCELL_X32 FILLER_75_65 ();
 FILLCELL_X32 FILLER_75_97 ();
 FILLCELL_X32 FILLER_75_129 ();
 FILLCELL_X8 FILLER_75_161 ();
 FILLCELL_X4 FILLER_75_819 ();
 FILLCELL_X8 FILLER_75_827 ();
 FILLCELL_X2 FILLER_75_835 ();
 FILLCELL_X4 FILLER_75_843 ();
 FILLCELL_X4 FILLER_75_850 ();
 FILLCELL_X4 FILLER_75_858 ();
 FILLCELL_X4 FILLER_75_871 ();
 FILLCELL_X32 FILLER_75_879 ();
 FILLCELL_X2 FILLER_75_911 ();
 FILLCELL_X16 FILLER_75_918 ();
 FILLCELL_X2 FILLER_75_934 ();
 FILLCELL_X1 FILLER_75_936 ();
 FILLCELL_X4 FILLER_75_940 ();
 FILLCELL_X1 FILLER_75_944 ();
 FILLCELL_X4 FILLER_75_951 ();
 FILLCELL_X4 FILLER_75_964 ();
 FILLCELL_X8 FILLER_75_972 ();
 FILLCELL_X4 FILLER_75_980 ();
 FILLCELL_X2 FILLER_75_984 ();
 FILLCELL_X4 FILLER_75_990 ();
 FILLCELL_X4 FILLER_75_1003 ();
 FILLCELL_X4 FILLER_75_1016 ();
 FILLCELL_X2 FILLER_75_1020 ();
 FILLCELL_X32 FILLER_76_1 ();
 FILLCELL_X32 FILLER_76_33 ();
 FILLCELL_X32 FILLER_76_65 ();
 FILLCELL_X32 FILLER_76_97 ();
 FILLCELL_X32 FILLER_76_129 ();
 FILLCELL_X8 FILLER_76_161 ();
 FILLCELL_X16 FILLER_76_819 ();
 FILLCELL_X1 FILLER_76_835 ();
 FILLCELL_X8 FILLER_76_839 ();
 FILLCELL_X2 FILLER_76_847 ();
 FILLCELL_X1 FILLER_76_849 ();
 FILLCELL_X4 FILLER_76_853 ();
 FILLCELL_X8 FILLER_76_860 ();
 FILLCELL_X2 FILLER_76_868 ();
 FILLCELL_X1 FILLER_76_870 ();
 FILLCELL_X8 FILLER_76_888 ();
 FILLCELL_X4 FILLER_76_896 ();
 FILLCELL_X4 FILLER_76_909 ();
 FILLCELL_X4 FILLER_76_917 ();
 FILLCELL_X4 FILLER_76_924 ();
 FILLCELL_X4 FILLER_76_934 ();
 FILLCELL_X4 FILLER_76_945 ();
 FILLCELL_X2 FILLER_76_949 ();
 FILLCELL_X4 FILLER_76_960 ();
 FILLCELL_X4 FILLER_76_967 ();
 FILLCELL_X2 FILLER_76_971 ();
 FILLCELL_X8 FILLER_76_977 ();
 FILLCELL_X2 FILLER_76_985 ();
 FILLCELL_X1 FILLER_76_987 ();
 FILLCELL_X4 FILLER_76_991 ();
 FILLCELL_X4 FILLER_76_1000 ();
 FILLCELL_X4 FILLER_76_1007 ();
 FILLCELL_X8 FILLER_76_1014 ();
 FILLCELL_X32 FILLER_77_1 ();
 FILLCELL_X32 FILLER_77_33 ();
 FILLCELL_X32 FILLER_77_65 ();
 FILLCELL_X32 FILLER_77_97 ();
 FILLCELL_X32 FILLER_77_129 ();
 FILLCELL_X8 FILLER_77_161 ();
 FILLCELL_X16 FILLER_77_819 ();
 FILLCELL_X8 FILLER_77_835 ();
 FILLCELL_X2 FILLER_77_843 ();
 FILLCELL_X4 FILLER_77_848 ();
 FILLCELL_X2 FILLER_77_852 ();
 FILLCELL_X1 FILLER_77_854 ();
 FILLCELL_X4 FILLER_77_861 ();
 FILLCELL_X4 FILLER_77_871 ();
 FILLCELL_X4 FILLER_77_879 ();
 FILLCELL_X2 FILLER_77_883 ();
 FILLCELL_X4 FILLER_77_889 ();
 FILLCELL_X4 FILLER_77_898 ();
 FILLCELL_X8 FILLER_77_911 ();
 FILLCELL_X4 FILLER_77_938 ();
 FILLCELL_X4 FILLER_77_948 ();
 FILLCELL_X8 FILLER_77_955 ();
 FILLCELL_X4 FILLER_77_963 ();
 FILLCELL_X8 FILLER_77_971 ();
 FILLCELL_X2 FILLER_77_979 ();
 FILLCELL_X4 FILLER_77_986 ();
 FILLCELL_X4 FILLER_77_994 ();
 FILLCELL_X1 FILLER_77_998 ();
 FILLCELL_X4 FILLER_77_1018 ();
 FILLCELL_X32 FILLER_78_1 ();
 FILLCELL_X32 FILLER_78_33 ();
 FILLCELL_X32 FILLER_78_65 ();
 FILLCELL_X32 FILLER_78_97 ();
 FILLCELL_X32 FILLER_78_129 ();
 FILLCELL_X8 FILLER_78_161 ();
 FILLCELL_X8 FILLER_78_819 ();
 FILLCELL_X4 FILLER_78_827 ();
 FILLCELL_X1 FILLER_78_831 ();
 FILLCELL_X4 FILLER_78_838 ();
 FILLCELL_X4 FILLER_78_846 ();
 FILLCELL_X8 FILLER_78_857 ();
 FILLCELL_X2 FILLER_78_865 ();
 FILLCELL_X1 FILLER_78_867 ();
 FILLCELL_X4 FILLER_78_875 ();
 FILLCELL_X4 FILLER_78_885 ();
 FILLCELL_X4 FILLER_78_893 ();
 FILLCELL_X4 FILLER_78_901 ();
 FILLCELL_X2 FILLER_78_905 ();
 FILLCELL_X1 FILLER_78_907 ();
 FILLCELL_X4 FILLER_78_914 ();
 FILLCELL_X4 FILLER_78_922 ();
 FILLCELL_X1 FILLER_78_926 ();
 FILLCELL_X16 FILLER_78_931 ();
 FILLCELL_X1 FILLER_78_947 ();
 FILLCELL_X4 FILLER_78_952 ();
 FILLCELL_X4 FILLER_78_960 ();
 FILLCELL_X4 FILLER_78_968 ();
 FILLCELL_X4 FILLER_78_976 ();
 FILLCELL_X4 FILLER_78_989 ();
 FILLCELL_X4 FILLER_78_1002 ();
 FILLCELL_X4 FILLER_78_1010 ();
 FILLCELL_X1 FILLER_78_1014 ();
 FILLCELL_X4 FILLER_78_1018 ();
 FILLCELL_X32 FILLER_79_1 ();
 FILLCELL_X32 FILLER_79_33 ();
 FILLCELL_X32 FILLER_79_65 ();
 FILLCELL_X32 FILLER_79_97 ();
 FILLCELL_X16 FILLER_79_129 ();
 FILLCELL_X4 FILLER_79_145 ();
 FILLCELL_X2 FILLER_79_149 ();
 FILLCELL_X8 FILLER_79_155 ();
 FILLCELL_X4 FILLER_79_163 ();
 FILLCELL_X2 FILLER_79_167 ();
 FILLCELL_X8 FILLER_79_819 ();
 FILLCELL_X2 FILLER_79_827 ();
 FILLCELL_X1 FILLER_79_829 ();
 FILLCELL_X4 FILLER_79_840 ();
 FILLCELL_X8 FILLER_79_851 ();
 FILLCELL_X1 FILLER_79_859 ();
 FILLCELL_X4 FILLER_79_866 ();
 FILLCELL_X4 FILLER_79_874 ();
 FILLCELL_X32 FILLER_79_882 ();
 FILLCELL_X2 FILLER_79_914 ();
 FILLCELL_X4 FILLER_79_919 ();
 FILLCELL_X8 FILLER_79_926 ();
 FILLCELL_X4 FILLER_79_934 ();
 FILLCELL_X8 FILLER_79_941 ();
 FILLCELL_X4 FILLER_79_949 ();
 FILLCELL_X2 FILLER_79_953 ();
 FILLCELL_X1 FILLER_79_955 ();
 FILLCELL_X8 FILLER_79_965 ();
 FILLCELL_X2 FILLER_79_973 ();
 FILLCELL_X1 FILLER_79_975 ();
 FILLCELL_X4 FILLER_79_979 ();
 FILLCELL_X8 FILLER_79_989 ();
 FILLCELL_X2 FILLER_79_997 ();
 FILLCELL_X4 FILLER_79_1018 ();
 FILLCELL_X32 FILLER_80_1 ();
 FILLCELL_X32 FILLER_80_33 ();
 FILLCELL_X32 FILLER_80_65 ();
 FILLCELL_X32 FILLER_80_97 ();
 FILLCELL_X8 FILLER_80_129 ();
 FILLCELL_X4 FILLER_80_137 ();
 FILLCELL_X1 FILLER_80_141 ();
 FILLCELL_X8 FILLER_80_161 ();
 FILLCELL_X16 FILLER_80_819 ();
 FILLCELL_X2 FILLER_80_835 ();
 FILLCELL_X32 FILLER_80_841 ();
 FILLCELL_X16 FILLER_80_873 ();
 FILLCELL_X1 FILLER_80_889 ();
 FILLCELL_X4 FILLER_80_899 ();
 FILLCELL_X8 FILLER_80_906 ();
 FILLCELL_X4 FILLER_80_914 ();
 FILLCELL_X2 FILLER_80_918 ();
 FILLCELL_X4 FILLER_80_923 ();
 FILLCELL_X8 FILLER_80_936 ();
 FILLCELL_X8 FILLER_80_948 ();
 FILLCELL_X2 FILLER_80_956 ();
 FILLCELL_X4 FILLER_80_967 ();
 FILLCELL_X16 FILLER_80_974 ();
 FILLCELL_X4 FILLER_80_990 ();
 FILLCELL_X1 FILLER_80_994 ();
 FILLCELL_X16 FILLER_80_999 ();
 FILLCELL_X4 FILLER_80_1015 ();
 FILLCELL_X2 FILLER_80_1019 ();
 FILLCELL_X1 FILLER_80_1021 ();
 FILLCELL_X32 FILLER_81_1 ();
 FILLCELL_X32 FILLER_81_33 ();
 FILLCELL_X32 FILLER_81_65 ();
 FILLCELL_X32 FILLER_81_97 ();
 FILLCELL_X32 FILLER_81_129 ();
 FILLCELL_X8 FILLER_81_161 ();
 FILLCELL_X8 FILLER_81_819 ();
 FILLCELL_X4 FILLER_81_827 ();
 FILLCELL_X4 FILLER_81_834 ();
 FILLCELL_X4 FILLER_81_844 ();
 FILLCELL_X4 FILLER_81_852 ();
 FILLCELL_X1 FILLER_81_856 ();
 FILLCELL_X4 FILLER_81_863 ();
 FILLCELL_X4 FILLER_81_873 ();
 FILLCELL_X2 FILLER_81_877 ();
 FILLCELL_X8 FILLER_81_883 ();
 FILLCELL_X4 FILLER_81_900 ();
 FILLCELL_X4 FILLER_81_910 ();
 FILLCELL_X4 FILLER_81_917 ();
 FILLCELL_X2 FILLER_81_921 ();
 FILLCELL_X4 FILLER_81_932 ();
 FILLCELL_X4 FILLER_81_942 ();
 FILLCELL_X2 FILLER_81_946 ();
 FILLCELL_X1 FILLER_81_948 ();
 FILLCELL_X4 FILLER_81_955 ();
 FILLCELL_X4 FILLER_81_968 ();
 FILLCELL_X8 FILLER_81_976 ();
 FILLCELL_X32 FILLER_81_988 ();
 FILLCELL_X2 FILLER_81_1020 ();
 FILLCELL_X4 FILLER_82_1 ();
 FILLCELL_X32 FILLER_82_8 ();
 FILLCELL_X32 FILLER_82_40 ();
 FILLCELL_X32 FILLER_82_72 ();
 FILLCELL_X32 FILLER_82_104 ();
 FILLCELL_X32 FILLER_82_136 ();
 FILLCELL_X1 FILLER_82_168 ();
 FILLCELL_X8 FILLER_82_819 ();
 FILLCELL_X4 FILLER_82_827 ();
 FILLCELL_X2 FILLER_82_831 ();
 FILLCELL_X1 FILLER_82_833 ();
 FILLCELL_X4 FILLER_82_843 ();
 FILLCELL_X4 FILLER_82_856 ();
 FILLCELL_X2 FILLER_82_860 ();
 FILLCELL_X4 FILLER_82_869 ();
 FILLCELL_X8 FILLER_82_876 ();
 FILLCELL_X4 FILLER_82_888 ();
 FILLCELL_X4 FILLER_82_897 ();
 FILLCELL_X4 FILLER_82_905 ();
 FILLCELL_X4 FILLER_82_912 ();
 FILLCELL_X2 FILLER_82_916 ();
 FILLCELL_X1 FILLER_82_918 ();
 FILLCELL_X4 FILLER_82_922 ();
 FILLCELL_X4 FILLER_82_931 ();
 FILLCELL_X8 FILLER_82_939 ();
 FILLCELL_X4 FILLER_82_947 ();
 FILLCELL_X1 FILLER_82_951 ();
 FILLCELL_X4 FILLER_82_955 ();
 FILLCELL_X4 FILLER_82_964 ();
 FILLCELL_X4 FILLER_82_971 ();
 FILLCELL_X4 FILLER_82_978 ();
 FILLCELL_X4 FILLER_82_986 ();
 FILLCELL_X4 FILLER_82_994 ();
 FILLCELL_X16 FILLER_82_1002 ();
 FILLCELL_X4 FILLER_82_1018 ();
 FILLCELL_X32 FILLER_83_1 ();
 FILLCELL_X32 FILLER_83_33 ();
 FILLCELL_X32 FILLER_83_65 ();
 FILLCELL_X32 FILLER_83_97 ();
 FILLCELL_X32 FILLER_83_129 ();
 FILLCELL_X1 FILLER_83_161 ();
 FILLCELL_X4 FILLER_83_165 ();
 FILLCELL_X4 FILLER_83_819 ();
 FILLCELL_X2 FILLER_83_823 ();
 FILLCELL_X8 FILLER_83_829 ();
 FILLCELL_X2 FILLER_83_837 ();
 FILLCELL_X4 FILLER_83_844 ();
 FILLCELL_X4 FILLER_83_851 ();
 FILLCELL_X1 FILLER_83_855 ();
 FILLCELL_X4 FILLER_83_859 ();
 FILLCELL_X16 FILLER_83_866 ();
 FILLCELL_X4 FILLER_83_882 ();
 FILLCELL_X16 FILLER_83_890 ();
 FILLCELL_X4 FILLER_83_906 ();
 FILLCELL_X2 FILLER_83_910 ();
 FILLCELL_X1 FILLER_83_912 ();
 FILLCELL_X8 FILLER_83_917 ();
 FILLCELL_X4 FILLER_83_932 ();
 FILLCELL_X16 FILLER_83_940 ();
 FILLCELL_X8 FILLER_83_956 ();
 FILLCELL_X4 FILLER_83_964 ();
 FILLCELL_X4 FILLER_83_972 ();
 FILLCELL_X4 FILLER_83_981 ();
 FILLCELL_X4 FILLER_83_994 ();
 FILLCELL_X4 FILLER_83_1007 ();
 FILLCELL_X4 FILLER_83_1015 ();
 FILLCELL_X2 FILLER_83_1019 ();
 FILLCELL_X1 FILLER_83_1021 ();
 FILLCELL_X32 FILLER_84_1 ();
 FILLCELL_X32 FILLER_84_33 ();
 FILLCELL_X32 FILLER_84_65 ();
 FILLCELL_X32 FILLER_84_97 ();
 FILLCELL_X32 FILLER_84_129 ();
 FILLCELL_X8 FILLER_84_161 ();
 FILLCELL_X8 FILLER_84_819 ();
 FILLCELL_X4 FILLER_84_827 ();
 FILLCELL_X4 FILLER_84_835 ();
 FILLCELL_X8 FILLER_84_843 ();
 FILLCELL_X2 FILLER_84_851 ();
 FILLCELL_X4 FILLER_84_856 ();
 FILLCELL_X4 FILLER_84_864 ();
 FILLCELL_X4 FILLER_84_874 ();
 FILLCELL_X8 FILLER_84_882 ();
 FILLCELL_X2 FILLER_84_890 ();
 FILLCELL_X1 FILLER_84_892 ();
 FILLCELL_X4 FILLER_84_897 ();
 FILLCELL_X4 FILLER_84_907 ();
 FILLCELL_X4 FILLER_84_914 ();
 FILLCELL_X2 FILLER_84_918 ();
 FILLCELL_X4 FILLER_84_926 ();
 FILLCELL_X1 FILLER_84_930 ();
 FILLCELL_X4 FILLER_84_934 ();
 FILLCELL_X1 FILLER_84_938 ();
 FILLCELL_X4 FILLER_84_942 ();
 FILLCELL_X1 FILLER_84_946 ();
 FILLCELL_X4 FILLER_84_951 ();
 FILLCELL_X4 FILLER_84_958 ();
 FILLCELL_X1 FILLER_84_962 ();
 FILLCELL_X8 FILLER_84_967 ();
 FILLCELL_X4 FILLER_84_975 ();
 FILLCELL_X4 FILLER_84_984 ();
 FILLCELL_X4 FILLER_84_994 ();
 FILLCELL_X1 FILLER_84_998 ();
 FILLCELL_X4 FILLER_84_1018 ();
 FILLCELL_X32 FILLER_85_1 ();
 FILLCELL_X32 FILLER_85_33 ();
 FILLCELL_X32 FILLER_85_65 ();
 FILLCELL_X32 FILLER_85_97 ();
 FILLCELL_X32 FILLER_85_129 ();
 FILLCELL_X8 FILLER_85_161 ();
 FILLCELL_X8 FILLER_85_819 ();
 FILLCELL_X4 FILLER_85_827 ();
 FILLCELL_X8 FILLER_85_835 ();
 FILLCELL_X4 FILLER_85_843 ();
 FILLCELL_X8 FILLER_85_856 ();
 FILLCELL_X2 FILLER_85_864 ();
 FILLCELL_X4 FILLER_85_875 ();
 FILLCELL_X4 FILLER_85_888 ();
 FILLCELL_X1 FILLER_85_892 ();
 FILLCELL_X4 FILLER_85_902 ();
 FILLCELL_X4 FILLER_85_915 ();
 FILLCELL_X2 FILLER_85_919 ();
 FILLCELL_X4 FILLER_85_927 ();
 FILLCELL_X1 FILLER_85_931 ();
 FILLCELL_X4 FILLER_85_937 ();
 FILLCELL_X4 FILLER_85_947 ();
 FILLCELL_X4 FILLER_85_960 ();
 FILLCELL_X2 FILLER_85_964 ();
 FILLCELL_X16 FILLER_85_968 ();
 FILLCELL_X8 FILLER_85_984 ();
 FILLCELL_X4 FILLER_85_992 ();
 FILLCELL_X16 FILLER_85_999 ();
 FILLCELL_X4 FILLER_85_1015 ();
 FILLCELL_X2 FILLER_85_1019 ();
 FILLCELL_X1 FILLER_85_1021 ();
 FILLCELL_X32 FILLER_86_1 ();
 FILLCELL_X32 FILLER_86_33 ();
 FILLCELL_X32 FILLER_86_65 ();
 FILLCELL_X32 FILLER_86_97 ();
 FILLCELL_X32 FILLER_86_129 ();
 FILLCELL_X8 FILLER_86_161 ();
 FILLCELL_X16 FILLER_86_819 ();
 FILLCELL_X4 FILLER_86_835 ();
 FILLCELL_X1 FILLER_86_839 ();
 FILLCELL_X4 FILLER_86_843 ();
 FILLCELL_X2 FILLER_86_847 ();
 FILLCELL_X1 FILLER_86_849 ();
 FILLCELL_X4 FILLER_86_854 ();
 FILLCELL_X4 FILLER_86_862 ();
 FILLCELL_X2 FILLER_86_866 ();
 FILLCELL_X1 FILLER_86_868 ();
 FILLCELL_X4 FILLER_86_874 ();
 FILLCELL_X4 FILLER_86_882 ();
 FILLCELL_X2 FILLER_86_886 ();
 FILLCELL_X4 FILLER_86_891 ();
 FILLCELL_X2 FILLER_86_895 ();
 FILLCELL_X1 FILLER_86_897 ();
 FILLCELL_X4 FILLER_86_903 ();
 FILLCELL_X4 FILLER_86_911 ();
 FILLCELL_X8 FILLER_86_918 ();
 FILLCELL_X4 FILLER_86_926 ();
 FILLCELL_X1 FILLER_86_930 ();
 FILLCELL_X4 FILLER_86_935 ();
 FILLCELL_X4 FILLER_86_948 ();
 FILLCELL_X4 FILLER_86_956 ();
 FILLCELL_X1 FILLER_86_960 ();
 FILLCELL_X4 FILLER_86_980 ();
 FILLCELL_X4 FILLER_86_987 ();
 FILLCELL_X4 FILLER_86_994 ();
 FILLCELL_X2 FILLER_86_998 ();
 FILLCELL_X1 FILLER_86_1000 ();
 FILLCELL_X4 FILLER_86_1018 ();
 FILLCELL_X32 FILLER_87_1 ();
 FILLCELL_X32 FILLER_87_33 ();
 FILLCELL_X32 FILLER_87_65 ();
 FILLCELL_X32 FILLER_87_97 ();
 FILLCELL_X32 FILLER_87_129 ();
 FILLCELL_X8 FILLER_87_161 ();
 FILLCELL_X4 FILLER_87_819 ();
 FILLCELL_X2 FILLER_87_823 ();
 FILLCELL_X4 FILLER_87_829 ();
 FILLCELL_X4 FILLER_87_842 ();
 FILLCELL_X4 FILLER_87_851 ();
 FILLCELL_X4 FILLER_87_858 ();
 FILLCELL_X4 FILLER_87_866 ();
 FILLCELL_X16 FILLER_87_873 ();
 FILLCELL_X8 FILLER_87_889 ();
 FILLCELL_X4 FILLER_87_897 ();
 FILLCELL_X4 FILLER_87_905 ();
 FILLCELL_X2 FILLER_87_909 ();
 FILLCELL_X8 FILLER_87_914 ();
 FILLCELL_X2 FILLER_87_922 ();
 FILLCELL_X16 FILLER_87_928 ();
 FILLCELL_X4 FILLER_87_944 ();
 FILLCELL_X2 FILLER_87_948 ();
 FILLCELL_X8 FILLER_87_952 ();
 FILLCELL_X4 FILLER_87_960 ();
 FILLCELL_X2 FILLER_87_964 ();
 FILLCELL_X4 FILLER_87_968 ();
 FILLCELL_X4 FILLER_87_976 ();
 FILLCELL_X4 FILLER_87_987 ();
 FILLCELL_X4 FILLER_87_997 ();
 FILLCELL_X8 FILLER_87_1005 ();
 FILLCELL_X2 FILLER_87_1013 ();
 FILLCELL_X4 FILLER_87_1018 ();
 FILLCELL_X32 FILLER_88_1 ();
 FILLCELL_X32 FILLER_88_33 ();
 FILLCELL_X32 FILLER_88_65 ();
 FILLCELL_X32 FILLER_88_97 ();
 FILLCELL_X32 FILLER_88_129 ();
 FILLCELL_X8 FILLER_88_161 ();
 FILLCELL_X4 FILLER_88_819 ();
 FILLCELL_X2 FILLER_88_823 ();
 FILLCELL_X1 FILLER_88_825 ();
 FILLCELL_X4 FILLER_88_830 ();
 FILLCELL_X4 FILLER_88_843 ();
 FILLCELL_X16 FILLER_88_851 ();
 FILLCELL_X8 FILLER_88_867 ();
 FILLCELL_X4 FILLER_88_875 ();
 FILLCELL_X8 FILLER_88_882 ();
 FILLCELL_X4 FILLER_88_899 ();
 FILLCELL_X8 FILLER_88_907 ();
 FILLCELL_X8 FILLER_88_919 ();
 FILLCELL_X1 FILLER_88_927 ();
 FILLCELL_X4 FILLER_88_933 ();
 FILLCELL_X4 FILLER_88_941 ();
 FILLCELL_X4 FILLER_88_947 ();
 FILLCELL_X4 FILLER_88_953 ();
 FILLCELL_X2 FILLER_88_957 ();
 FILLCELL_X1 FILLER_88_959 ();
 FILLCELL_X4 FILLER_88_964 ();
 FILLCELL_X4 FILLER_88_972 ();
 FILLCELL_X2 FILLER_88_976 ();
 FILLCELL_X1 FILLER_88_978 ();
 FILLCELL_X4 FILLER_88_983 ();
 FILLCELL_X16 FILLER_88_993 ();
 FILLCELL_X8 FILLER_88_1009 ();
 FILLCELL_X4 FILLER_88_1017 ();
 FILLCELL_X1 FILLER_88_1021 ();
 FILLCELL_X32 FILLER_89_1 ();
 FILLCELL_X32 FILLER_89_33 ();
 FILLCELL_X32 FILLER_89_65 ();
 FILLCELL_X32 FILLER_89_97 ();
 FILLCELL_X32 FILLER_89_129 ();
 FILLCELL_X8 FILLER_89_161 ();
 FILLCELL_X8 FILLER_89_819 ();
 FILLCELL_X2 FILLER_89_827 ();
 FILLCELL_X4 FILLER_89_833 ();
 FILLCELL_X16 FILLER_89_843 ();
 FILLCELL_X2 FILLER_89_859 ();
 FILLCELL_X4 FILLER_89_866 ();
 FILLCELL_X4 FILLER_89_879 ();
 FILLCELL_X8 FILLER_89_886 ();
 FILLCELL_X2 FILLER_89_894 ();
 FILLCELL_X4 FILLER_89_900 ();
 FILLCELL_X4 FILLER_89_908 ();
 FILLCELL_X4 FILLER_89_916 ();
 FILLCELL_X1 FILLER_89_920 ();
 FILLCELL_X4 FILLER_89_940 ();
 FILLCELL_X8 FILLER_89_948 ();
 FILLCELL_X4 FILLER_89_960 ();
 FILLCELL_X4 FILLER_89_970 ();
 FILLCELL_X32 FILLER_89_978 ();
 FILLCELL_X8 FILLER_89_1010 ();
 FILLCELL_X4 FILLER_89_1018 ();
 FILLCELL_X32 FILLER_90_1 ();
 FILLCELL_X32 FILLER_90_33 ();
 FILLCELL_X32 FILLER_90_65 ();
 FILLCELL_X32 FILLER_90_97 ();
 FILLCELL_X32 FILLER_90_129 ();
 FILLCELL_X8 FILLER_90_161 ();
 FILLCELL_X8 FILLER_90_819 ();
 FILLCELL_X4 FILLER_90_827 ();
 FILLCELL_X2 FILLER_90_831 ();
 FILLCELL_X1 FILLER_90_833 ();
 FILLCELL_X4 FILLER_90_838 ();
 FILLCELL_X2 FILLER_90_842 ();
 FILLCELL_X4 FILLER_90_849 ();
 FILLCELL_X4 FILLER_90_857 ();
 FILLCELL_X2 FILLER_90_861 ();
 FILLCELL_X4 FILLER_90_872 ();
 FILLCELL_X16 FILLER_90_882 ();
 FILLCELL_X1 FILLER_90_898 ();
 FILLCELL_X16 FILLER_90_903 ();
 FILLCELL_X8 FILLER_90_919 ();
 FILLCELL_X2 FILLER_90_927 ();
 FILLCELL_X1 FILLER_90_929 ();
 FILLCELL_X4 FILLER_90_934 ();
 FILLCELL_X4 FILLER_90_942 ();
 FILLCELL_X4 FILLER_90_950 ();
 FILLCELL_X8 FILLER_90_958 ();
 FILLCELL_X4 FILLER_90_966 ();
 FILLCELL_X1 FILLER_90_970 ();
 FILLCELL_X8 FILLER_90_977 ();
 FILLCELL_X2 FILLER_90_985 ();
 FILLCELL_X16 FILLER_90_1004 ();
 FILLCELL_X2 FILLER_90_1020 ();
 FILLCELL_X32 FILLER_91_1 ();
 FILLCELL_X32 FILLER_91_33 ();
 FILLCELL_X32 FILLER_91_65 ();
 FILLCELL_X32 FILLER_91_97 ();
 FILLCELL_X32 FILLER_91_129 ();
 FILLCELL_X8 FILLER_91_161 ();
 FILLCELL_X4 FILLER_91_819 ();
 FILLCELL_X2 FILLER_91_823 ();
 FILLCELL_X1 FILLER_91_825 ();
 FILLCELL_X4 FILLER_91_830 ();
 FILLCELL_X4 FILLER_91_838 ();
 FILLCELL_X4 FILLER_91_846 ();
 FILLCELL_X4 FILLER_91_853 ();
 FILLCELL_X4 FILLER_91_861 ();
 FILLCELL_X4 FILLER_91_869 ();
 FILLCELL_X8 FILLER_91_877 ();
 FILLCELL_X2 FILLER_91_885 ();
 FILLCELL_X4 FILLER_91_892 ();
 FILLCELL_X8 FILLER_91_905 ();
 FILLCELL_X4 FILLER_91_913 ();
 FILLCELL_X4 FILLER_91_921 ();
 FILLCELL_X4 FILLER_91_931 ();
 FILLCELL_X8 FILLER_91_944 ();
 FILLCELL_X4 FILLER_91_952 ();
 FILLCELL_X4 FILLER_91_960 ();
 FILLCELL_X4 FILLER_91_968 ();
 FILLCELL_X4 FILLER_91_976 ();
 FILLCELL_X1 FILLER_91_980 ();
 FILLCELL_X32 FILLER_91_985 ();
 FILLCELL_X4 FILLER_91_1017 ();
 FILLCELL_X1 FILLER_91_1021 ();
 FILLCELL_X32 FILLER_92_1 ();
 FILLCELL_X32 FILLER_92_33 ();
 FILLCELL_X32 FILLER_92_65 ();
 FILLCELL_X32 FILLER_92_97 ();
 FILLCELL_X32 FILLER_92_129 ();
 FILLCELL_X8 FILLER_92_161 ();
 FILLCELL_X16 FILLER_92_819 ();
 FILLCELL_X1 FILLER_92_835 ();
 FILLCELL_X4 FILLER_92_841 ();
 FILLCELL_X8 FILLER_92_849 ();
 FILLCELL_X4 FILLER_92_861 ();
 FILLCELL_X2 FILLER_92_865 ();
 FILLCELL_X4 FILLER_92_872 ();
 FILLCELL_X1 FILLER_92_876 ();
 FILLCELL_X8 FILLER_92_880 ();
 FILLCELL_X4 FILLER_92_894 ();
 FILLCELL_X4 FILLER_92_907 ();
 FILLCELL_X8 FILLER_92_914 ();
 FILLCELL_X1 FILLER_92_922 ();
 FILLCELL_X4 FILLER_92_926 ();
 FILLCELL_X4 FILLER_92_939 ();
 FILLCELL_X4 FILLER_92_948 ();
 FILLCELL_X4 FILLER_92_956 ();
 FILLCELL_X32 FILLER_92_969 ();
 FILLCELL_X16 FILLER_92_1001 ();
 FILLCELL_X4 FILLER_92_1017 ();
 FILLCELL_X1 FILLER_92_1021 ();
 FILLCELL_X4 FILLER_93_1 ();
 FILLCELL_X32 FILLER_93_8 ();
 FILLCELL_X32 FILLER_93_40 ();
 FILLCELL_X32 FILLER_93_72 ();
 FILLCELL_X32 FILLER_93_104 ();
 FILLCELL_X32 FILLER_93_136 ();
 FILLCELL_X1 FILLER_93_168 ();
 FILLCELL_X8 FILLER_93_819 ();
 FILLCELL_X4 FILLER_93_827 ();
 FILLCELL_X2 FILLER_93_831 ();
 FILLCELL_X4 FILLER_93_842 ();
 FILLCELL_X8 FILLER_93_855 ();
 FILLCELL_X4 FILLER_93_872 ();
 FILLCELL_X4 FILLER_93_885 ();
 FILLCELL_X4 FILLER_93_892 ();
 FILLCELL_X2 FILLER_93_896 ();
 FILLCELL_X1 FILLER_93_898 ();
 FILLCELL_X4 FILLER_93_903 ();
 FILLCELL_X4 FILLER_93_910 ();
 FILLCELL_X4 FILLER_93_918 ();
 FILLCELL_X4 FILLER_93_931 ();
 FILLCELL_X16 FILLER_93_938 ();
 FILLCELL_X4 FILLER_93_954 ();
 FILLCELL_X2 FILLER_93_958 ();
 FILLCELL_X1 FILLER_93_960 ();
 FILLCELL_X32 FILLER_93_970 ();
 FILLCELL_X16 FILLER_93_1002 ();
 FILLCELL_X4 FILLER_93_1018 ();
 FILLCELL_X32 FILLER_94_1 ();
 FILLCELL_X32 FILLER_94_33 ();
 FILLCELL_X32 FILLER_94_65 ();
 FILLCELL_X32 FILLER_94_97 ();
 FILLCELL_X32 FILLER_94_129 ();
 FILLCELL_X8 FILLER_94_161 ();
 FILLCELL_X8 FILLER_94_819 ();
 FILLCELL_X4 FILLER_94_827 ();
 FILLCELL_X4 FILLER_94_834 ();
 FILLCELL_X4 FILLER_94_844 ();
 FILLCELL_X8 FILLER_94_853 ();
 FILLCELL_X4 FILLER_94_861 ();
 FILLCELL_X4 FILLER_94_871 ();
 FILLCELL_X16 FILLER_94_878 ();
 FILLCELL_X2 FILLER_94_894 ();
 FILLCELL_X16 FILLER_94_901 ();
 FILLCELL_X4 FILLER_94_917 ();
 FILLCELL_X16 FILLER_94_924 ();
 FILLCELL_X8 FILLER_94_940 ();
 FILLCELL_X4 FILLER_94_948 ();
 FILLCELL_X4 FILLER_94_957 ();
 FILLCELL_X4 FILLER_94_970 ();
 FILLCELL_X32 FILLER_94_978 ();
 FILLCELL_X8 FILLER_94_1010 ();
 FILLCELL_X4 FILLER_94_1018 ();
 FILLCELL_X32 FILLER_95_1 ();
 FILLCELL_X32 FILLER_95_33 ();
 FILLCELL_X32 FILLER_95_65 ();
 FILLCELL_X32 FILLER_95_97 ();
 FILLCELL_X32 FILLER_95_129 ();
 FILLCELL_X8 FILLER_95_161 ();
 FILLCELL_X32 FILLER_95_819 ();
 FILLCELL_X16 FILLER_95_851 ();
 FILLCELL_X2 FILLER_95_867 ();
 FILLCELL_X4 FILLER_95_872 ();
 FILLCELL_X1 FILLER_95_876 ();
 FILLCELL_X8 FILLER_95_880 ();
 FILLCELL_X4 FILLER_95_888 ();
 FILLCELL_X4 FILLER_95_901 ();
 FILLCELL_X8 FILLER_95_914 ();
 FILLCELL_X4 FILLER_95_927 ();
 FILLCELL_X4 FILLER_95_940 ();
 FILLCELL_X4 FILLER_95_948 ();
 FILLCELL_X4 FILLER_95_955 ();
 FILLCELL_X4 FILLER_95_965 ();
 FILLCELL_X16 FILLER_95_972 ();
 FILLCELL_X8 FILLER_95_988 ();
 FILLCELL_X4 FILLER_95_996 ();
 FILLCELL_X1 FILLER_95_1000 ();
 FILLCELL_X4 FILLER_95_1018 ();
 FILLCELL_X32 FILLER_96_1 ();
 FILLCELL_X32 FILLER_96_33 ();
 FILLCELL_X32 FILLER_96_65 ();
 FILLCELL_X32 FILLER_96_97 ();
 FILLCELL_X32 FILLER_96_129 ();
 FILLCELL_X8 FILLER_96_161 ();
 FILLCELL_X32 FILLER_96_819 ();
 FILLCELL_X4 FILLER_96_851 ();
 FILLCELL_X2 FILLER_96_855 ();
 FILLCELL_X1 FILLER_96_857 ();
 FILLCELL_X4 FILLER_96_864 ();
 FILLCELL_X8 FILLER_96_872 ();
 FILLCELL_X4 FILLER_96_880 ();
 FILLCELL_X2 FILLER_96_884 ();
 FILLCELL_X1 FILLER_96_886 ();
 FILLCELL_X4 FILLER_96_890 ();
 FILLCELL_X4 FILLER_96_900 ();
 FILLCELL_X4 FILLER_96_908 ();
 FILLCELL_X8 FILLER_96_915 ();
 FILLCELL_X1 FILLER_96_923 ();
 FILLCELL_X4 FILLER_96_930 ();
 FILLCELL_X32 FILLER_96_943 ();
 FILLCELL_X32 FILLER_96_975 ();
 FILLCELL_X8 FILLER_96_1007 ();
 FILLCELL_X4 FILLER_96_1015 ();
 FILLCELL_X2 FILLER_96_1019 ();
 FILLCELL_X1 FILLER_96_1021 ();
 FILLCELL_X32 FILLER_97_1 ();
 FILLCELL_X32 FILLER_97_33 ();
 FILLCELL_X32 FILLER_97_65 ();
 FILLCELL_X32 FILLER_97_97 ();
 FILLCELL_X32 FILLER_97_129 ();
 FILLCELL_X8 FILLER_97_161 ();
 FILLCELL_X32 FILLER_97_819 ();
 FILLCELL_X2 FILLER_97_851 ();
 FILLCELL_X4 FILLER_97_863 ();
 FILLCELL_X4 FILLER_97_874 ();
 FILLCELL_X1 FILLER_97_878 ();
 FILLCELL_X8 FILLER_97_883 ();
 FILLCELL_X4 FILLER_97_891 ();
 FILLCELL_X8 FILLER_97_898 ();
 FILLCELL_X1 FILLER_97_906 ();
 FILLCELL_X4 FILLER_97_913 ();
 FILLCELL_X4 FILLER_97_920 ();
 FILLCELL_X4 FILLER_97_927 ();
 FILLCELL_X1 FILLER_97_931 ();
 FILLCELL_X4 FILLER_97_935 ();
 FILLCELL_X32 FILLER_97_942 ();
 FILLCELL_X32 FILLER_97_974 ();
 FILLCELL_X16 FILLER_97_1006 ();
 FILLCELL_X32 FILLER_98_1 ();
 FILLCELL_X32 FILLER_98_33 ();
 FILLCELL_X32 FILLER_98_65 ();
 FILLCELL_X32 FILLER_98_97 ();
 FILLCELL_X16 FILLER_98_129 ();
 FILLCELL_X8 FILLER_98_145 ();
 FILLCELL_X4 FILLER_98_153 ();
 FILLCELL_X2 FILLER_98_157 ();
 FILLCELL_X1 FILLER_98_159 ();
 FILLCELL_X4 FILLER_98_164 ();
 FILLCELL_X1 FILLER_98_168 ();
 FILLCELL_X32 FILLER_98_819 ();
 FILLCELL_X8 FILLER_98_851 ();
 FILLCELL_X2 FILLER_98_859 ();
 FILLCELL_X1 FILLER_98_861 ();
 FILLCELL_X4 FILLER_98_866 ();
 FILLCELL_X2 FILLER_98_870 ();
 FILLCELL_X1 FILLER_98_872 ();
 FILLCELL_X8 FILLER_98_877 ();
 FILLCELL_X2 FILLER_98_885 ();
 FILLCELL_X1 FILLER_98_887 ();
 FILLCELL_X4 FILLER_98_895 ();
 FILLCELL_X8 FILLER_98_905 ();
 FILLCELL_X2 FILLER_98_913 ();
 FILLCELL_X4 FILLER_98_922 ();
 FILLCELL_X32 FILLER_98_929 ();
 FILLCELL_X32 FILLER_98_961 ();
 FILLCELL_X16 FILLER_98_993 ();
 FILLCELL_X4 FILLER_98_1009 ();
 FILLCELL_X2 FILLER_98_1013 ();
 FILLCELL_X4 FILLER_98_1018 ();
 FILLCELL_X32 FILLER_99_1 ();
 FILLCELL_X32 FILLER_99_33 ();
 FILLCELL_X32 FILLER_99_65 ();
 FILLCELL_X32 FILLER_99_97 ();
 FILLCELL_X16 FILLER_99_129 ();
 FILLCELL_X2 FILLER_99_145 ();
 FILLCELL_X1 FILLER_99_147 ();
 FILLCELL_X4 FILLER_99_165 ();
 FILLCELL_X32 FILLER_99_819 ();
 FILLCELL_X16 FILLER_99_851 ();
 FILLCELL_X4 FILLER_99_867 ();
 FILLCELL_X1 FILLER_99_871 ();
 FILLCELL_X4 FILLER_99_878 ();
 FILLCELL_X2 FILLER_99_882 ();
 FILLCELL_X1 FILLER_99_884 ();
 FILLCELL_X4 FILLER_99_892 ();
 FILLCELL_X4 FILLER_99_902 ();
 FILLCELL_X8 FILLER_99_909 ();
 FILLCELL_X32 FILLER_99_923 ();
 FILLCELL_X32 FILLER_99_955 ();
 FILLCELL_X32 FILLER_99_987 ();
 FILLCELL_X2 FILLER_99_1019 ();
 FILLCELL_X1 FILLER_99_1021 ();
 FILLCELL_X32 FILLER_100_1 ();
 FILLCELL_X32 FILLER_100_33 ();
 FILLCELL_X32 FILLER_100_65 ();
 FILLCELL_X32 FILLER_100_97 ();
 FILLCELL_X32 FILLER_100_129 ();
 FILLCELL_X8 FILLER_100_161 ();
 FILLCELL_X32 FILLER_100_819 ();
 FILLCELL_X16 FILLER_100_851 ();
 FILLCELL_X4 FILLER_100_867 ();
 FILLCELL_X16 FILLER_100_881 ();
 FILLCELL_X2 FILLER_100_897 ();
 FILLCELL_X16 FILLER_100_903 ();
 FILLCELL_X1 FILLER_100_919 ();
 FILLCELL_X4 FILLER_100_924 ();
 FILLCELL_X32 FILLER_100_947 ();
 FILLCELL_X32 FILLER_100_979 ();
 FILLCELL_X8 FILLER_100_1011 ();
 FILLCELL_X2 FILLER_100_1019 ();
 FILLCELL_X1 FILLER_100_1021 ();
 FILLCELL_X32 FILLER_101_1 ();
 FILLCELL_X32 FILLER_101_33 ();
 FILLCELL_X32 FILLER_101_65 ();
 FILLCELL_X32 FILLER_101_97 ();
 FILLCELL_X32 FILLER_101_129 ();
 FILLCELL_X8 FILLER_101_161 ();
 FILLCELL_X32 FILLER_101_819 ();
 FILLCELL_X32 FILLER_101_851 ();
 FILLCELL_X16 FILLER_101_883 ();
 FILLCELL_X1 FILLER_101_899 ();
 FILLCELL_X32 FILLER_101_917 ();
 FILLCELL_X32 FILLER_101_949 ();
 FILLCELL_X32 FILLER_101_981 ();
 FILLCELL_X8 FILLER_101_1013 ();
 FILLCELL_X1 FILLER_101_1021 ();
 FILLCELL_X32 FILLER_102_1 ();
 FILLCELL_X32 FILLER_102_33 ();
 FILLCELL_X32 FILLER_102_65 ();
 FILLCELL_X32 FILLER_102_97 ();
 FILLCELL_X32 FILLER_102_129 ();
 FILLCELL_X8 FILLER_102_161 ();
 FILLCELL_X32 FILLER_102_819 ();
 FILLCELL_X32 FILLER_102_851 ();
 FILLCELL_X32 FILLER_102_883 ();
 FILLCELL_X32 FILLER_102_915 ();
 FILLCELL_X32 FILLER_102_947 ();
 FILLCELL_X32 FILLER_102_979 ();
 FILLCELL_X8 FILLER_102_1011 ();
 FILLCELL_X2 FILLER_102_1019 ();
 FILLCELL_X1 FILLER_102_1021 ();
 FILLCELL_X32 FILLER_103_1 ();
 FILLCELL_X32 FILLER_103_33 ();
 FILLCELL_X32 FILLER_103_65 ();
 FILLCELL_X32 FILLER_103_97 ();
 FILLCELL_X32 FILLER_103_129 ();
 FILLCELL_X8 FILLER_103_161 ();
 FILLCELL_X32 FILLER_103_819 ();
 FILLCELL_X32 FILLER_103_851 ();
 FILLCELL_X32 FILLER_103_883 ();
 FILLCELL_X32 FILLER_103_915 ();
 FILLCELL_X32 FILLER_103_947 ();
 FILLCELL_X32 FILLER_103_979 ();
 FILLCELL_X8 FILLER_103_1011 ();
 FILLCELL_X2 FILLER_103_1019 ();
 FILLCELL_X1 FILLER_103_1021 ();
 FILLCELL_X32 FILLER_104_1 ();
 FILLCELL_X32 FILLER_104_33 ();
 FILLCELL_X32 FILLER_104_65 ();
 FILLCELL_X32 FILLER_104_97 ();
 FILLCELL_X32 FILLER_104_129 ();
 FILLCELL_X8 FILLER_104_161 ();
 FILLCELL_X32 FILLER_104_819 ();
 FILLCELL_X32 FILLER_104_851 ();
 FILLCELL_X32 FILLER_104_883 ();
 FILLCELL_X32 FILLER_104_915 ();
 FILLCELL_X32 FILLER_104_947 ();
 FILLCELL_X32 FILLER_104_979 ();
 FILLCELL_X8 FILLER_104_1011 ();
 FILLCELL_X2 FILLER_104_1019 ();
 FILLCELL_X1 FILLER_104_1021 ();
 FILLCELL_X32 FILLER_105_1 ();
 FILLCELL_X32 FILLER_105_33 ();
 FILLCELL_X32 FILLER_105_65 ();
 FILLCELL_X32 FILLER_105_97 ();
 FILLCELL_X32 FILLER_105_129 ();
 FILLCELL_X8 FILLER_105_161 ();
 FILLCELL_X32 FILLER_105_819 ();
 FILLCELL_X32 FILLER_105_851 ();
 FILLCELL_X32 FILLER_105_883 ();
 FILLCELL_X32 FILLER_105_915 ();
 FILLCELL_X32 FILLER_105_947 ();
 FILLCELL_X32 FILLER_105_979 ();
 FILLCELL_X8 FILLER_105_1011 ();
 FILLCELL_X2 FILLER_105_1019 ();
 FILLCELL_X1 FILLER_105_1021 ();
 FILLCELL_X32 FILLER_106_1 ();
 FILLCELL_X32 FILLER_106_33 ();
 FILLCELL_X32 FILLER_106_65 ();
 FILLCELL_X32 FILLER_106_97 ();
 FILLCELL_X32 FILLER_106_129 ();
 FILLCELL_X8 FILLER_106_161 ();
 FILLCELL_X32 FILLER_106_819 ();
 FILLCELL_X32 FILLER_106_851 ();
 FILLCELL_X32 FILLER_106_883 ();
 FILLCELL_X32 FILLER_106_915 ();
 FILLCELL_X32 FILLER_106_947 ();
 FILLCELL_X32 FILLER_106_979 ();
 FILLCELL_X8 FILLER_106_1011 ();
 FILLCELL_X2 FILLER_106_1019 ();
 FILLCELL_X1 FILLER_106_1021 ();
 FILLCELL_X32 FILLER_107_1 ();
 FILLCELL_X32 FILLER_107_33 ();
 FILLCELL_X32 FILLER_107_65 ();
 FILLCELL_X32 FILLER_107_97 ();
 FILLCELL_X32 FILLER_107_129 ();
 FILLCELL_X8 FILLER_107_161 ();
 FILLCELL_X32 FILLER_107_819 ();
 FILLCELL_X32 FILLER_107_851 ();
 FILLCELL_X32 FILLER_107_883 ();
 FILLCELL_X32 FILLER_107_915 ();
 FILLCELL_X32 FILLER_107_947 ();
 FILLCELL_X32 FILLER_107_979 ();
 FILLCELL_X8 FILLER_107_1011 ();
 FILLCELL_X2 FILLER_107_1019 ();
 FILLCELL_X1 FILLER_107_1021 ();
 FILLCELL_X32 FILLER_108_1 ();
 FILLCELL_X32 FILLER_108_33 ();
 FILLCELL_X32 FILLER_108_65 ();
 FILLCELL_X32 FILLER_108_97 ();
 FILLCELL_X32 FILLER_108_129 ();
 FILLCELL_X8 FILLER_108_161 ();
 FILLCELL_X32 FILLER_108_819 ();
 FILLCELL_X32 FILLER_108_851 ();
 FILLCELL_X32 FILLER_108_883 ();
 FILLCELL_X32 FILLER_108_915 ();
 FILLCELL_X32 FILLER_108_947 ();
 FILLCELL_X32 FILLER_108_979 ();
 FILLCELL_X8 FILLER_108_1011 ();
 FILLCELL_X2 FILLER_108_1019 ();
 FILLCELL_X1 FILLER_108_1021 ();
 FILLCELL_X32 FILLER_109_1 ();
 FILLCELL_X32 FILLER_109_33 ();
 FILLCELL_X32 FILLER_109_65 ();
 FILLCELL_X32 FILLER_109_97 ();
 FILLCELL_X32 FILLER_109_129 ();
 FILLCELL_X8 FILLER_109_161 ();
 FILLCELL_X32 FILLER_109_819 ();
 FILLCELL_X32 FILLER_109_851 ();
 FILLCELL_X32 FILLER_109_883 ();
 FILLCELL_X32 FILLER_109_915 ();
 FILLCELL_X32 FILLER_109_947 ();
 FILLCELL_X32 FILLER_109_979 ();
 FILLCELL_X4 FILLER_109_1011 ();
 FILLCELL_X4 FILLER_109_1018 ();
 FILLCELL_X32 FILLER_110_1 ();
 FILLCELL_X32 FILLER_110_33 ();
 FILLCELL_X32 FILLER_110_65 ();
 FILLCELL_X32 FILLER_110_97 ();
 FILLCELL_X32 FILLER_110_129 ();
 FILLCELL_X8 FILLER_110_161 ();
 FILLCELL_X32 FILLER_110_819 ();
 FILLCELL_X32 FILLER_110_851 ();
 FILLCELL_X32 FILLER_110_883 ();
 FILLCELL_X32 FILLER_110_915 ();
 FILLCELL_X32 FILLER_110_947 ();
 FILLCELL_X32 FILLER_110_979 ();
 FILLCELL_X8 FILLER_110_1011 ();
 FILLCELL_X2 FILLER_110_1019 ();
 FILLCELL_X1 FILLER_110_1021 ();
 FILLCELL_X32 FILLER_111_1 ();
 FILLCELL_X32 FILLER_111_33 ();
 FILLCELL_X32 FILLER_111_65 ();
 FILLCELL_X32 FILLER_111_97 ();
 FILLCELL_X32 FILLER_111_129 ();
 FILLCELL_X8 FILLER_111_161 ();
 FILLCELL_X32 FILLER_111_819 ();
 FILLCELL_X32 FILLER_111_851 ();
 FILLCELL_X32 FILLER_111_883 ();
 FILLCELL_X32 FILLER_111_915 ();
 FILLCELL_X32 FILLER_111_947 ();
 FILLCELL_X32 FILLER_111_979 ();
 FILLCELL_X8 FILLER_111_1011 ();
 FILLCELL_X2 FILLER_111_1019 ();
 FILLCELL_X1 FILLER_111_1021 ();
 FILLCELL_X32 FILLER_112_1 ();
 FILLCELL_X32 FILLER_112_33 ();
 FILLCELL_X32 FILLER_112_65 ();
 FILLCELL_X32 FILLER_112_97 ();
 FILLCELL_X32 FILLER_112_129 ();
 FILLCELL_X8 FILLER_112_161 ();
 FILLCELL_X32 FILLER_112_819 ();
 FILLCELL_X32 FILLER_112_851 ();
 FILLCELL_X32 FILLER_112_883 ();
 FILLCELL_X32 FILLER_112_915 ();
 FILLCELL_X32 FILLER_112_947 ();
 FILLCELL_X32 FILLER_112_979 ();
 FILLCELL_X8 FILLER_112_1011 ();
 FILLCELL_X2 FILLER_112_1019 ();
 FILLCELL_X1 FILLER_112_1021 ();
 FILLCELL_X32 FILLER_113_1 ();
 FILLCELL_X32 FILLER_113_33 ();
 FILLCELL_X32 FILLER_113_65 ();
 FILLCELL_X32 FILLER_113_97 ();
 FILLCELL_X32 FILLER_113_129 ();
 FILLCELL_X8 FILLER_113_161 ();
 FILLCELL_X32 FILLER_113_819 ();
 FILLCELL_X32 FILLER_113_851 ();
 FILLCELL_X32 FILLER_113_883 ();
 FILLCELL_X32 FILLER_113_915 ();
 FILLCELL_X32 FILLER_113_947 ();
 FILLCELL_X32 FILLER_113_979 ();
 FILLCELL_X8 FILLER_113_1011 ();
 FILLCELL_X2 FILLER_113_1019 ();
 FILLCELL_X1 FILLER_113_1021 ();
 FILLCELL_X4 FILLER_114_1 ();
 FILLCELL_X32 FILLER_114_8 ();
 FILLCELL_X32 FILLER_114_40 ();
 FILLCELL_X32 FILLER_114_72 ();
 FILLCELL_X32 FILLER_114_104 ();
 FILLCELL_X32 FILLER_114_136 ();
 FILLCELL_X1 FILLER_114_168 ();
 FILLCELL_X32 FILLER_114_819 ();
 FILLCELL_X32 FILLER_114_851 ();
 FILLCELL_X32 FILLER_114_883 ();
 FILLCELL_X32 FILLER_114_915 ();
 FILLCELL_X32 FILLER_114_947 ();
 FILLCELL_X32 FILLER_114_979 ();
 FILLCELL_X8 FILLER_114_1011 ();
 FILLCELL_X2 FILLER_114_1019 ();
 FILLCELL_X1 FILLER_114_1021 ();
 FILLCELL_X32 FILLER_115_1 ();
 FILLCELL_X32 FILLER_115_33 ();
 FILLCELL_X32 FILLER_115_65 ();
 FILLCELL_X32 FILLER_115_97 ();
 FILLCELL_X32 FILLER_115_129 ();
 FILLCELL_X8 FILLER_115_161 ();
 FILLCELL_X32 FILLER_115_819 ();
 FILLCELL_X32 FILLER_115_851 ();
 FILLCELL_X32 FILLER_115_883 ();
 FILLCELL_X32 FILLER_115_915 ();
 FILLCELL_X32 FILLER_115_947 ();
 FILLCELL_X32 FILLER_115_979 ();
 FILLCELL_X8 FILLER_115_1011 ();
 FILLCELL_X2 FILLER_115_1019 ();
 FILLCELL_X1 FILLER_115_1021 ();
 FILLCELL_X32 FILLER_116_1 ();
 FILLCELL_X32 FILLER_116_33 ();
 FILLCELL_X32 FILLER_116_65 ();
 FILLCELL_X32 FILLER_116_97 ();
 FILLCELL_X32 FILLER_116_129 ();
 FILLCELL_X8 FILLER_116_161 ();
 FILLCELL_X32 FILLER_116_819 ();
 FILLCELL_X32 FILLER_116_851 ();
 FILLCELL_X32 FILLER_116_883 ();
 FILLCELL_X32 FILLER_116_915 ();
 FILLCELL_X32 FILLER_116_947 ();
 FILLCELL_X32 FILLER_116_979 ();
 FILLCELL_X8 FILLER_116_1011 ();
 FILLCELL_X2 FILLER_116_1019 ();
 FILLCELL_X1 FILLER_116_1021 ();
 FILLCELL_X32 FILLER_117_1 ();
 FILLCELL_X32 FILLER_117_33 ();
 FILLCELL_X32 FILLER_117_65 ();
 FILLCELL_X32 FILLER_117_97 ();
 FILLCELL_X32 FILLER_117_129 ();
 FILLCELL_X32 FILLER_117_161 ();
 FILLCELL_X32 FILLER_117_193 ();
 FILLCELL_X32 FILLER_117_225 ();
 FILLCELL_X32 FILLER_117_257 ();
 FILLCELL_X32 FILLER_117_289 ();
 FILLCELL_X32 FILLER_117_321 ();
 FILLCELL_X32 FILLER_117_353 ();
 FILLCELL_X32 FILLER_117_385 ();
 FILLCELL_X32 FILLER_117_417 ();
 FILLCELL_X32 FILLER_117_449 ();
 FILLCELL_X32 FILLER_117_481 ();
 FILLCELL_X32 FILLER_117_513 ();
 FILLCELL_X32 FILLER_117_545 ();
 FILLCELL_X32 FILLER_117_577 ();
 FILLCELL_X16 FILLER_117_609 ();
 FILLCELL_X4 FILLER_117_625 ();
 FILLCELL_X2 FILLER_117_629 ();
 FILLCELL_X8 FILLER_117_632 ();
 FILLCELL_X1 FILLER_117_640 ();
 FILLCELL_X4 FILLER_117_660 ();
 FILLCELL_X32 FILLER_117_668 ();
 FILLCELL_X32 FILLER_117_700 ();
 FILLCELL_X32 FILLER_117_732 ();
 FILLCELL_X32 FILLER_117_764 ();
 FILLCELL_X32 FILLER_117_796 ();
 FILLCELL_X32 FILLER_117_828 ();
 FILLCELL_X32 FILLER_117_860 ();
 FILLCELL_X32 FILLER_117_892 ();
 FILLCELL_X32 FILLER_117_924 ();
 FILLCELL_X32 FILLER_117_956 ();
 FILLCELL_X32 FILLER_117_988 ();
 FILLCELL_X2 FILLER_117_1020 ();
 FILLCELL_X32 FILLER_118_1 ();
 FILLCELL_X32 FILLER_118_33 ();
 FILLCELL_X32 FILLER_118_65 ();
 FILLCELL_X32 FILLER_118_97 ();
 FILLCELL_X32 FILLER_118_129 ();
 FILLCELL_X32 FILLER_118_161 ();
 FILLCELL_X32 FILLER_118_193 ();
 FILLCELL_X32 FILLER_118_225 ();
 FILLCELL_X32 FILLER_118_257 ();
 FILLCELL_X32 FILLER_118_289 ();
 FILLCELL_X32 FILLER_118_321 ();
 FILLCELL_X32 FILLER_118_353 ();
 FILLCELL_X32 FILLER_118_385 ();
 FILLCELL_X32 FILLER_118_417 ();
 FILLCELL_X32 FILLER_118_449 ();
 FILLCELL_X32 FILLER_118_481 ();
 FILLCELL_X32 FILLER_118_513 ();
 FILLCELL_X32 FILLER_118_545 ();
 FILLCELL_X32 FILLER_118_577 ();
 FILLCELL_X16 FILLER_118_609 ();
 FILLCELL_X4 FILLER_118_625 ();
 FILLCELL_X2 FILLER_118_629 ();
 FILLCELL_X32 FILLER_118_632 ();
 FILLCELL_X32 FILLER_118_664 ();
 FILLCELL_X32 FILLER_118_696 ();
 FILLCELL_X32 FILLER_118_728 ();
 FILLCELL_X32 FILLER_118_760 ();
 FILLCELL_X32 FILLER_118_792 ();
 FILLCELL_X32 FILLER_118_824 ();
 FILLCELL_X32 FILLER_118_856 ();
 FILLCELL_X32 FILLER_118_888 ();
 FILLCELL_X32 FILLER_118_920 ();
 FILLCELL_X32 FILLER_118_952 ();
 FILLCELL_X32 FILLER_118_984 ();
 FILLCELL_X4 FILLER_118_1016 ();
 FILLCELL_X2 FILLER_118_1020 ();
 FILLCELL_X32 FILLER_119_1 ();
 FILLCELL_X32 FILLER_119_33 ();
 FILLCELL_X32 FILLER_119_65 ();
 FILLCELL_X32 FILLER_119_97 ();
 FILLCELL_X32 FILLER_119_129 ();
 FILLCELL_X32 FILLER_119_161 ();
 FILLCELL_X32 FILLER_119_193 ();
 FILLCELL_X32 FILLER_119_225 ();
 FILLCELL_X32 FILLER_119_257 ();
 FILLCELL_X32 FILLER_119_289 ();
 FILLCELL_X32 FILLER_119_321 ();
 FILLCELL_X32 FILLER_119_353 ();
 FILLCELL_X32 FILLER_119_385 ();
 FILLCELL_X32 FILLER_119_417 ();
 FILLCELL_X32 FILLER_119_449 ();
 FILLCELL_X32 FILLER_119_481 ();
 FILLCELL_X32 FILLER_119_513 ();
 FILLCELL_X32 FILLER_119_545 ();
 FILLCELL_X32 FILLER_119_577 ();
 FILLCELL_X32 FILLER_119_609 ();
 FILLCELL_X32 FILLER_119_641 ();
 FILLCELL_X32 FILLER_119_673 ();
 FILLCELL_X32 FILLER_119_705 ();
 FILLCELL_X32 FILLER_119_737 ();
 FILLCELL_X32 FILLER_119_769 ();
 FILLCELL_X32 FILLER_119_801 ();
 FILLCELL_X32 FILLER_119_833 ();
 FILLCELL_X32 FILLER_119_865 ();
 FILLCELL_X32 FILLER_119_897 ();
 FILLCELL_X32 FILLER_119_929 ();
 FILLCELL_X32 FILLER_119_961 ();
 FILLCELL_X16 FILLER_119_993 ();
 FILLCELL_X8 FILLER_119_1009 ();
 FILLCELL_X4 FILLER_119_1017 ();
 FILLCELL_X1 FILLER_119_1021 ();
 FILLCELL_X32 FILLER_120_1 ();
 FILLCELL_X32 FILLER_120_33 ();
 FILLCELL_X32 FILLER_120_65 ();
 FILLCELL_X32 FILLER_120_97 ();
 FILLCELL_X32 FILLER_120_129 ();
 FILLCELL_X32 FILLER_120_161 ();
 FILLCELL_X32 FILLER_120_193 ();
 FILLCELL_X32 FILLER_120_225 ();
 FILLCELL_X32 FILLER_120_257 ();
 FILLCELL_X32 FILLER_120_289 ();
 FILLCELL_X32 FILLER_120_321 ();
 FILLCELL_X32 FILLER_120_353 ();
 FILLCELL_X32 FILLER_120_385 ();
 FILLCELL_X32 FILLER_120_417 ();
 FILLCELL_X32 FILLER_120_449 ();
 FILLCELL_X32 FILLER_120_481 ();
 FILLCELL_X32 FILLER_120_513 ();
 FILLCELL_X32 FILLER_120_545 ();
 FILLCELL_X32 FILLER_120_577 ();
 FILLCELL_X16 FILLER_120_609 ();
 FILLCELL_X4 FILLER_120_625 ();
 FILLCELL_X2 FILLER_120_629 ();
 FILLCELL_X32 FILLER_120_632 ();
 FILLCELL_X32 FILLER_120_664 ();
 FILLCELL_X32 FILLER_120_696 ();
 FILLCELL_X32 FILLER_120_728 ();
 FILLCELL_X32 FILLER_120_760 ();
 FILLCELL_X32 FILLER_120_792 ();
 FILLCELL_X32 FILLER_120_824 ();
 FILLCELL_X32 FILLER_120_856 ();
 FILLCELL_X32 FILLER_120_888 ();
 FILLCELL_X32 FILLER_120_920 ();
 FILLCELL_X32 FILLER_120_952 ();
 FILLCELL_X16 FILLER_120_984 ();
 FILLCELL_X8 FILLER_120_1000 ();
 FILLCELL_X4 FILLER_120_1008 ();
 FILLCELL_X2 FILLER_120_1012 ();
 FILLCELL_X1 FILLER_120_1014 ();
 FILLCELL_X4 FILLER_120_1018 ();
 FILLCELL_X32 FILLER_121_1 ();
 FILLCELL_X32 FILLER_121_33 ();
 FILLCELL_X32 FILLER_121_65 ();
 FILLCELL_X32 FILLER_121_97 ();
 FILLCELL_X32 FILLER_121_129 ();
 FILLCELL_X32 FILLER_121_161 ();
 FILLCELL_X32 FILLER_121_193 ();
 FILLCELL_X32 FILLER_121_225 ();
 FILLCELL_X32 FILLER_121_257 ();
 FILLCELL_X32 FILLER_121_289 ();
 FILLCELL_X32 FILLER_121_321 ();
 FILLCELL_X32 FILLER_121_353 ();
 FILLCELL_X32 FILLER_121_385 ();
 FILLCELL_X32 FILLER_121_417 ();
 FILLCELL_X32 FILLER_121_449 ();
 FILLCELL_X32 FILLER_121_481 ();
 FILLCELL_X32 FILLER_121_513 ();
 FILLCELL_X32 FILLER_121_545 ();
 FILLCELL_X32 FILLER_121_577 ();
 FILLCELL_X32 FILLER_121_609 ();
 FILLCELL_X32 FILLER_121_641 ();
 FILLCELL_X32 FILLER_121_673 ();
 FILLCELL_X32 FILLER_121_705 ();
 FILLCELL_X32 FILLER_121_737 ();
 FILLCELL_X32 FILLER_121_769 ();
 FILLCELL_X32 FILLER_121_801 ();
 FILLCELL_X32 FILLER_121_833 ();
 FILLCELL_X32 FILLER_121_865 ();
 FILLCELL_X32 FILLER_121_897 ();
 FILLCELL_X32 FILLER_121_929 ();
 FILLCELL_X32 FILLER_121_961 ();
 FILLCELL_X16 FILLER_121_993 ();
 FILLCELL_X8 FILLER_121_1009 ();
 FILLCELL_X4 FILLER_121_1017 ();
 FILLCELL_X1 FILLER_121_1021 ();
 FILLCELL_X32 FILLER_122_1 ();
 FILLCELL_X32 FILLER_122_33 ();
 FILLCELL_X32 FILLER_122_65 ();
 FILLCELL_X32 FILLER_122_97 ();
 FILLCELL_X32 FILLER_122_129 ();
 FILLCELL_X32 FILLER_122_161 ();
 FILLCELL_X32 FILLER_122_193 ();
 FILLCELL_X32 FILLER_122_225 ();
 FILLCELL_X32 FILLER_122_257 ();
 FILLCELL_X32 FILLER_122_289 ();
 FILLCELL_X32 FILLER_122_321 ();
 FILLCELL_X32 FILLER_122_353 ();
 FILLCELL_X32 FILLER_122_385 ();
 FILLCELL_X32 FILLER_122_417 ();
 FILLCELL_X32 FILLER_122_449 ();
 FILLCELL_X32 FILLER_122_481 ();
 FILLCELL_X32 FILLER_122_513 ();
 FILLCELL_X32 FILLER_122_545 ();
 FILLCELL_X32 FILLER_122_577 ();
 FILLCELL_X16 FILLER_122_609 ();
 FILLCELL_X4 FILLER_122_625 ();
 FILLCELL_X2 FILLER_122_629 ();
 FILLCELL_X32 FILLER_122_632 ();
 FILLCELL_X32 FILLER_122_664 ();
 FILLCELL_X32 FILLER_122_696 ();
 FILLCELL_X32 FILLER_122_728 ();
 FILLCELL_X32 FILLER_122_760 ();
 FILLCELL_X32 FILLER_122_792 ();
 FILLCELL_X32 FILLER_122_824 ();
 FILLCELL_X32 FILLER_122_856 ();
 FILLCELL_X32 FILLER_122_888 ();
 FILLCELL_X32 FILLER_122_920 ();
 FILLCELL_X32 FILLER_122_952 ();
 FILLCELL_X32 FILLER_122_984 ();
 FILLCELL_X4 FILLER_122_1016 ();
 FILLCELL_X2 FILLER_122_1020 ();
 FILLCELL_X32 FILLER_123_1 ();
 FILLCELL_X32 FILLER_123_33 ();
 FILLCELL_X32 FILLER_123_65 ();
 FILLCELL_X32 FILLER_123_97 ();
 FILLCELL_X32 FILLER_123_129 ();
 FILLCELL_X32 FILLER_123_161 ();
 FILLCELL_X32 FILLER_123_193 ();
 FILLCELL_X32 FILLER_123_225 ();
 FILLCELL_X32 FILLER_123_257 ();
 FILLCELL_X32 FILLER_123_289 ();
 FILLCELL_X32 FILLER_123_321 ();
 FILLCELL_X32 FILLER_123_353 ();
 FILLCELL_X32 FILLER_123_385 ();
 FILLCELL_X32 FILLER_123_417 ();
 FILLCELL_X32 FILLER_123_449 ();
 FILLCELL_X32 FILLER_123_481 ();
 FILLCELL_X32 FILLER_123_513 ();
 FILLCELL_X32 FILLER_123_545 ();
 FILLCELL_X32 FILLER_123_577 ();
 FILLCELL_X32 FILLER_123_609 ();
 FILLCELL_X32 FILLER_123_641 ();
 FILLCELL_X32 FILLER_123_673 ();
 FILLCELL_X32 FILLER_123_705 ();
 FILLCELL_X32 FILLER_123_737 ();
 FILLCELL_X32 FILLER_123_769 ();
 FILLCELL_X32 FILLER_123_801 ();
 FILLCELL_X32 FILLER_123_833 ();
 FILLCELL_X32 FILLER_123_865 ();
 FILLCELL_X32 FILLER_123_897 ();
 FILLCELL_X32 FILLER_123_929 ();
 FILLCELL_X32 FILLER_123_961 ();
 FILLCELL_X16 FILLER_123_993 ();
 FILLCELL_X8 FILLER_123_1009 ();
 FILLCELL_X4 FILLER_123_1017 ();
 FILLCELL_X1 FILLER_123_1021 ();
 FILLCELL_X32 FILLER_124_1 ();
 FILLCELL_X32 FILLER_124_33 ();
 FILLCELL_X32 FILLER_124_65 ();
 FILLCELL_X32 FILLER_124_97 ();
 FILLCELL_X32 FILLER_124_129 ();
 FILLCELL_X32 FILLER_124_161 ();
 FILLCELL_X32 FILLER_124_193 ();
 FILLCELL_X32 FILLER_124_225 ();
 FILLCELL_X32 FILLER_124_257 ();
 FILLCELL_X32 FILLER_124_289 ();
 FILLCELL_X32 FILLER_124_321 ();
 FILLCELL_X32 FILLER_124_353 ();
 FILLCELL_X32 FILLER_124_385 ();
 FILLCELL_X32 FILLER_124_417 ();
 FILLCELL_X32 FILLER_124_449 ();
 FILLCELL_X32 FILLER_124_481 ();
 FILLCELL_X32 FILLER_124_513 ();
 FILLCELL_X32 FILLER_124_545 ();
 FILLCELL_X32 FILLER_124_577 ();
 FILLCELL_X16 FILLER_124_609 ();
 FILLCELL_X4 FILLER_124_625 ();
 FILLCELL_X2 FILLER_124_629 ();
 FILLCELL_X32 FILLER_124_632 ();
 FILLCELL_X32 FILLER_124_664 ();
 FILLCELL_X32 FILLER_124_696 ();
 FILLCELL_X32 FILLER_124_728 ();
 FILLCELL_X32 FILLER_124_760 ();
 FILLCELL_X32 FILLER_124_792 ();
 FILLCELL_X32 FILLER_124_824 ();
 FILLCELL_X32 FILLER_124_856 ();
 FILLCELL_X32 FILLER_124_888 ();
 FILLCELL_X32 FILLER_124_920 ();
 FILLCELL_X32 FILLER_124_952 ();
 FILLCELL_X32 FILLER_124_984 ();
 FILLCELL_X4 FILLER_124_1016 ();
 FILLCELL_X2 FILLER_124_1020 ();
 FILLCELL_X4 FILLER_125_1 ();
 FILLCELL_X32 FILLER_125_18 ();
 FILLCELL_X32 FILLER_125_50 ();
 FILLCELL_X32 FILLER_125_82 ();
 FILLCELL_X32 FILLER_125_114 ();
 FILLCELL_X32 FILLER_125_146 ();
 FILLCELL_X32 FILLER_125_178 ();
 FILLCELL_X32 FILLER_125_210 ();
 FILLCELL_X32 FILLER_125_242 ();
 FILLCELL_X32 FILLER_125_274 ();
 FILLCELL_X32 FILLER_125_306 ();
 FILLCELL_X32 FILLER_125_338 ();
 FILLCELL_X32 FILLER_125_370 ();
 FILLCELL_X32 FILLER_125_402 ();
 FILLCELL_X32 FILLER_125_434 ();
 FILLCELL_X32 FILLER_125_466 ();
 FILLCELL_X32 FILLER_125_498 ();
 FILLCELL_X32 FILLER_125_530 ();
 FILLCELL_X32 FILLER_125_562 ();
 FILLCELL_X32 FILLER_125_594 ();
 FILLCELL_X32 FILLER_125_626 ();
 FILLCELL_X32 FILLER_125_658 ();
 FILLCELL_X32 FILLER_125_690 ();
 FILLCELL_X32 FILLER_125_722 ();
 FILLCELL_X32 FILLER_125_754 ();
 FILLCELL_X32 FILLER_125_786 ();
 FILLCELL_X32 FILLER_125_818 ();
 FILLCELL_X32 FILLER_125_850 ();
 FILLCELL_X32 FILLER_125_882 ();
 FILLCELL_X32 FILLER_125_914 ();
 FILLCELL_X32 FILLER_125_946 ();
 FILLCELL_X32 FILLER_125_978 ();
 FILLCELL_X8 FILLER_125_1010 ();
 FILLCELL_X4 FILLER_125_1018 ();
 FILLCELL_X32 FILLER_126_1 ();
 FILLCELL_X32 FILLER_126_33 ();
 FILLCELL_X32 FILLER_126_65 ();
 FILLCELL_X32 FILLER_126_97 ();
 FILLCELL_X32 FILLER_126_129 ();
 FILLCELL_X32 FILLER_126_161 ();
 FILLCELL_X32 FILLER_126_193 ();
 FILLCELL_X32 FILLER_126_225 ();
 FILLCELL_X32 FILLER_126_257 ();
 FILLCELL_X32 FILLER_126_289 ();
 FILLCELL_X32 FILLER_126_321 ();
 FILLCELL_X32 FILLER_126_353 ();
 FILLCELL_X32 FILLER_126_385 ();
 FILLCELL_X32 FILLER_126_417 ();
 FILLCELL_X32 FILLER_126_449 ();
 FILLCELL_X32 FILLER_126_481 ();
 FILLCELL_X32 FILLER_126_513 ();
 FILLCELL_X32 FILLER_126_545 ();
 FILLCELL_X32 FILLER_126_577 ();
 FILLCELL_X16 FILLER_126_609 ();
 FILLCELL_X4 FILLER_126_625 ();
 FILLCELL_X2 FILLER_126_629 ();
 FILLCELL_X32 FILLER_126_632 ();
 FILLCELL_X32 FILLER_126_664 ();
 FILLCELL_X32 FILLER_126_696 ();
 FILLCELL_X32 FILLER_126_728 ();
 FILLCELL_X32 FILLER_126_760 ();
 FILLCELL_X32 FILLER_126_792 ();
 FILLCELL_X32 FILLER_126_824 ();
 FILLCELL_X32 FILLER_126_856 ();
 FILLCELL_X32 FILLER_126_888 ();
 FILLCELL_X32 FILLER_126_920 ();
 FILLCELL_X32 FILLER_126_952 ();
 FILLCELL_X32 FILLER_126_984 ();
 FILLCELL_X4 FILLER_126_1016 ();
 FILLCELL_X2 FILLER_126_1020 ();
 FILLCELL_X32 FILLER_127_1 ();
 FILLCELL_X32 FILLER_127_33 ();
 FILLCELL_X32 FILLER_127_65 ();
 FILLCELL_X32 FILLER_127_97 ();
 FILLCELL_X32 FILLER_127_129 ();
 FILLCELL_X32 FILLER_127_161 ();
 FILLCELL_X32 FILLER_127_193 ();
 FILLCELL_X32 FILLER_127_225 ();
 FILLCELL_X32 FILLER_127_257 ();
 FILLCELL_X32 FILLER_127_289 ();
 FILLCELL_X32 FILLER_127_321 ();
 FILLCELL_X32 FILLER_127_353 ();
 FILLCELL_X32 FILLER_127_385 ();
 FILLCELL_X32 FILLER_127_417 ();
 FILLCELL_X32 FILLER_127_449 ();
 FILLCELL_X32 FILLER_127_481 ();
 FILLCELL_X32 FILLER_127_513 ();
 FILLCELL_X32 FILLER_127_545 ();
 FILLCELL_X32 FILLER_127_577 ();
 FILLCELL_X32 FILLER_127_609 ();
 FILLCELL_X32 FILLER_127_641 ();
 FILLCELL_X32 FILLER_127_673 ();
 FILLCELL_X32 FILLER_127_705 ();
 FILLCELL_X32 FILLER_127_737 ();
 FILLCELL_X32 FILLER_127_769 ();
 FILLCELL_X32 FILLER_127_801 ();
 FILLCELL_X32 FILLER_127_833 ();
 FILLCELL_X32 FILLER_127_865 ();
 FILLCELL_X32 FILLER_127_897 ();
 FILLCELL_X32 FILLER_127_929 ();
 FILLCELL_X32 FILLER_127_961 ();
 FILLCELL_X16 FILLER_127_993 ();
 FILLCELL_X8 FILLER_127_1009 ();
 FILLCELL_X4 FILLER_127_1017 ();
 FILLCELL_X1 FILLER_127_1021 ();
 FILLCELL_X32 FILLER_128_1 ();
 FILLCELL_X32 FILLER_128_33 ();
 FILLCELL_X32 FILLER_128_65 ();
 FILLCELL_X32 FILLER_128_97 ();
 FILLCELL_X32 FILLER_128_129 ();
 FILLCELL_X32 FILLER_128_161 ();
 FILLCELL_X32 FILLER_128_193 ();
 FILLCELL_X32 FILLER_128_225 ();
 FILLCELL_X32 FILLER_128_257 ();
 FILLCELL_X32 FILLER_128_289 ();
 FILLCELL_X32 FILLER_128_321 ();
 FILLCELL_X32 FILLER_128_353 ();
 FILLCELL_X32 FILLER_128_385 ();
 FILLCELL_X32 FILLER_128_417 ();
 FILLCELL_X32 FILLER_128_449 ();
 FILLCELL_X32 FILLER_128_481 ();
 FILLCELL_X32 FILLER_128_513 ();
 FILLCELL_X32 FILLER_128_545 ();
 FILLCELL_X32 FILLER_128_577 ();
 FILLCELL_X16 FILLER_128_609 ();
 FILLCELL_X4 FILLER_128_625 ();
 FILLCELL_X2 FILLER_128_629 ();
 FILLCELL_X32 FILLER_128_632 ();
 FILLCELL_X32 FILLER_128_664 ();
 FILLCELL_X32 FILLER_128_696 ();
 FILLCELL_X32 FILLER_128_728 ();
 FILLCELL_X32 FILLER_128_760 ();
 FILLCELL_X32 FILLER_128_792 ();
 FILLCELL_X32 FILLER_128_824 ();
 FILLCELL_X32 FILLER_128_856 ();
 FILLCELL_X32 FILLER_128_888 ();
 FILLCELL_X32 FILLER_128_920 ();
 FILLCELL_X32 FILLER_128_952 ();
 FILLCELL_X32 FILLER_128_984 ();
 FILLCELL_X4 FILLER_128_1016 ();
 FILLCELL_X2 FILLER_128_1020 ();
 FILLCELL_X32 FILLER_129_1 ();
 FILLCELL_X32 FILLER_129_33 ();
 FILLCELL_X32 FILLER_129_65 ();
 FILLCELL_X32 FILLER_129_97 ();
 FILLCELL_X32 FILLER_129_129 ();
 FILLCELL_X32 FILLER_129_161 ();
 FILLCELL_X32 FILLER_129_193 ();
 FILLCELL_X32 FILLER_129_225 ();
 FILLCELL_X32 FILLER_129_257 ();
 FILLCELL_X32 FILLER_129_289 ();
 FILLCELL_X32 FILLER_129_321 ();
 FILLCELL_X32 FILLER_129_353 ();
 FILLCELL_X32 FILLER_129_385 ();
 FILLCELL_X32 FILLER_129_417 ();
 FILLCELL_X32 FILLER_129_449 ();
 FILLCELL_X32 FILLER_129_481 ();
 FILLCELL_X32 FILLER_129_513 ();
 FILLCELL_X32 FILLER_129_545 ();
 FILLCELL_X32 FILLER_129_577 ();
 FILLCELL_X32 FILLER_129_609 ();
 FILLCELL_X32 FILLER_129_641 ();
 FILLCELL_X32 FILLER_129_673 ();
 FILLCELL_X32 FILLER_129_705 ();
 FILLCELL_X32 FILLER_129_737 ();
 FILLCELL_X32 FILLER_129_769 ();
 FILLCELL_X32 FILLER_129_801 ();
 FILLCELL_X32 FILLER_129_833 ();
 FILLCELL_X32 FILLER_129_865 ();
 FILLCELL_X32 FILLER_129_897 ();
 FILLCELL_X32 FILLER_129_929 ();
 FILLCELL_X32 FILLER_129_961 ();
 FILLCELL_X16 FILLER_129_993 ();
 FILLCELL_X8 FILLER_129_1009 ();
 FILLCELL_X4 FILLER_129_1017 ();
 FILLCELL_X1 FILLER_129_1021 ();
 FILLCELL_X32 FILLER_130_1 ();
 FILLCELL_X32 FILLER_130_33 ();
 FILLCELL_X32 FILLER_130_65 ();
 FILLCELL_X32 FILLER_130_97 ();
 FILLCELL_X32 FILLER_130_129 ();
 FILLCELL_X32 FILLER_130_161 ();
 FILLCELL_X32 FILLER_130_193 ();
 FILLCELL_X32 FILLER_130_225 ();
 FILLCELL_X32 FILLER_130_257 ();
 FILLCELL_X32 FILLER_130_289 ();
 FILLCELL_X32 FILLER_130_321 ();
 FILLCELL_X32 FILLER_130_353 ();
 FILLCELL_X32 FILLER_130_385 ();
 FILLCELL_X32 FILLER_130_417 ();
 FILLCELL_X32 FILLER_130_449 ();
 FILLCELL_X32 FILLER_130_481 ();
 FILLCELL_X32 FILLER_130_513 ();
 FILLCELL_X32 FILLER_130_545 ();
 FILLCELL_X32 FILLER_130_577 ();
 FILLCELL_X16 FILLER_130_609 ();
 FILLCELL_X4 FILLER_130_625 ();
 FILLCELL_X2 FILLER_130_629 ();
 FILLCELL_X32 FILLER_130_632 ();
 FILLCELL_X32 FILLER_130_664 ();
 FILLCELL_X32 FILLER_130_696 ();
 FILLCELL_X32 FILLER_130_728 ();
 FILLCELL_X32 FILLER_130_760 ();
 FILLCELL_X32 FILLER_130_792 ();
 FILLCELL_X32 FILLER_130_824 ();
 FILLCELL_X32 FILLER_130_856 ();
 FILLCELL_X32 FILLER_130_888 ();
 FILLCELL_X32 FILLER_130_920 ();
 FILLCELL_X32 FILLER_130_952 ();
 FILLCELL_X16 FILLER_130_984 ();
 FILLCELL_X8 FILLER_130_1000 ();
 FILLCELL_X4 FILLER_130_1008 ();
 FILLCELL_X2 FILLER_130_1012 ();
 FILLCELL_X1 FILLER_130_1014 ();
 FILLCELL_X4 FILLER_130_1018 ();
 FILLCELL_X32 FILLER_131_1 ();
 FILLCELL_X32 FILLER_131_33 ();
 FILLCELL_X32 FILLER_131_65 ();
 FILLCELL_X32 FILLER_131_97 ();
 FILLCELL_X32 FILLER_131_129 ();
 FILLCELL_X32 FILLER_131_161 ();
 FILLCELL_X32 FILLER_131_193 ();
 FILLCELL_X32 FILLER_131_225 ();
 FILLCELL_X32 FILLER_131_257 ();
 FILLCELL_X32 FILLER_131_289 ();
 FILLCELL_X32 FILLER_131_321 ();
 FILLCELL_X32 FILLER_131_353 ();
 FILLCELL_X32 FILLER_131_385 ();
 FILLCELL_X32 FILLER_131_417 ();
 FILLCELL_X32 FILLER_131_449 ();
 FILLCELL_X32 FILLER_131_481 ();
 FILLCELL_X32 FILLER_131_513 ();
 FILLCELL_X32 FILLER_131_545 ();
 FILLCELL_X32 FILLER_131_577 ();
 FILLCELL_X32 FILLER_131_609 ();
 FILLCELL_X32 FILLER_131_641 ();
 FILLCELL_X32 FILLER_131_673 ();
 FILLCELL_X32 FILLER_131_705 ();
 FILLCELL_X32 FILLER_131_737 ();
 FILLCELL_X32 FILLER_131_769 ();
 FILLCELL_X32 FILLER_131_801 ();
 FILLCELL_X32 FILLER_131_833 ();
 FILLCELL_X32 FILLER_131_865 ();
 FILLCELL_X32 FILLER_131_897 ();
 FILLCELL_X32 FILLER_131_929 ();
 FILLCELL_X32 FILLER_131_961 ();
 FILLCELL_X16 FILLER_131_993 ();
 FILLCELL_X8 FILLER_131_1009 ();
 FILLCELL_X4 FILLER_131_1017 ();
 FILLCELL_X1 FILLER_131_1021 ();
 FILLCELL_X32 FILLER_132_1 ();
 FILLCELL_X32 FILLER_132_33 ();
 FILLCELL_X32 FILLER_132_65 ();
 FILLCELL_X32 FILLER_132_97 ();
 FILLCELL_X32 FILLER_132_129 ();
 FILLCELL_X32 FILLER_132_161 ();
 FILLCELL_X32 FILLER_132_193 ();
 FILLCELL_X32 FILLER_132_225 ();
 FILLCELL_X32 FILLER_132_257 ();
 FILLCELL_X32 FILLER_132_289 ();
 FILLCELL_X32 FILLER_132_321 ();
 FILLCELL_X32 FILLER_132_353 ();
 FILLCELL_X32 FILLER_132_385 ();
 FILLCELL_X32 FILLER_132_417 ();
 FILLCELL_X32 FILLER_132_449 ();
 FILLCELL_X32 FILLER_132_481 ();
 FILLCELL_X32 FILLER_132_513 ();
 FILLCELL_X32 FILLER_132_545 ();
 FILLCELL_X32 FILLER_132_577 ();
 FILLCELL_X16 FILLER_132_609 ();
 FILLCELL_X4 FILLER_132_625 ();
 FILLCELL_X2 FILLER_132_629 ();
 FILLCELL_X32 FILLER_132_632 ();
 FILLCELL_X32 FILLER_132_664 ();
 FILLCELL_X32 FILLER_132_696 ();
 FILLCELL_X32 FILLER_132_728 ();
 FILLCELL_X32 FILLER_132_760 ();
 FILLCELL_X32 FILLER_132_792 ();
 FILLCELL_X32 FILLER_132_824 ();
 FILLCELL_X32 FILLER_132_856 ();
 FILLCELL_X32 FILLER_132_888 ();
 FILLCELL_X32 FILLER_132_920 ();
 FILLCELL_X32 FILLER_132_952 ();
 FILLCELL_X32 FILLER_132_984 ();
 FILLCELL_X4 FILLER_132_1016 ();
 FILLCELL_X2 FILLER_132_1020 ();
 FILLCELL_X32 FILLER_133_1 ();
 FILLCELL_X32 FILLER_133_33 ();
 FILLCELL_X32 FILLER_133_65 ();
 FILLCELL_X32 FILLER_133_97 ();
 FILLCELL_X32 FILLER_133_129 ();
 FILLCELL_X32 FILLER_133_161 ();
 FILLCELL_X32 FILLER_133_193 ();
 FILLCELL_X32 FILLER_133_225 ();
 FILLCELL_X32 FILLER_133_257 ();
 FILLCELL_X32 FILLER_133_289 ();
 FILLCELL_X32 FILLER_133_321 ();
 FILLCELL_X32 FILLER_133_353 ();
 FILLCELL_X32 FILLER_133_385 ();
 FILLCELL_X32 FILLER_133_417 ();
 FILLCELL_X32 FILLER_133_449 ();
 FILLCELL_X32 FILLER_133_481 ();
 FILLCELL_X32 FILLER_133_513 ();
 FILLCELL_X32 FILLER_133_545 ();
 FILLCELL_X32 FILLER_133_577 ();
 FILLCELL_X32 FILLER_133_609 ();
 FILLCELL_X32 FILLER_133_641 ();
 FILLCELL_X32 FILLER_133_673 ();
 FILLCELL_X32 FILLER_133_705 ();
 FILLCELL_X32 FILLER_133_737 ();
 FILLCELL_X32 FILLER_133_769 ();
 FILLCELL_X32 FILLER_133_801 ();
 FILLCELL_X32 FILLER_133_833 ();
 FILLCELL_X32 FILLER_133_865 ();
 FILLCELL_X32 FILLER_133_897 ();
 FILLCELL_X32 FILLER_133_929 ();
 FILLCELL_X32 FILLER_133_961 ();
 FILLCELL_X16 FILLER_133_993 ();
 FILLCELL_X8 FILLER_133_1009 ();
 FILLCELL_X4 FILLER_133_1017 ();
 FILLCELL_X1 FILLER_133_1021 ();
 FILLCELL_X32 FILLER_134_1 ();
 FILLCELL_X32 FILLER_134_33 ();
 FILLCELL_X32 FILLER_134_65 ();
 FILLCELL_X32 FILLER_134_97 ();
 FILLCELL_X32 FILLER_134_129 ();
 FILLCELL_X32 FILLER_134_161 ();
 FILLCELL_X32 FILLER_134_193 ();
 FILLCELL_X32 FILLER_134_225 ();
 FILLCELL_X32 FILLER_134_257 ();
 FILLCELL_X32 FILLER_134_289 ();
 FILLCELL_X32 FILLER_134_321 ();
 FILLCELL_X32 FILLER_134_353 ();
 FILLCELL_X32 FILLER_134_385 ();
 FILLCELL_X32 FILLER_134_417 ();
 FILLCELL_X32 FILLER_134_449 ();
 FILLCELL_X32 FILLER_134_481 ();
 FILLCELL_X32 FILLER_134_513 ();
 FILLCELL_X32 FILLER_134_545 ();
 FILLCELL_X32 FILLER_134_577 ();
 FILLCELL_X16 FILLER_134_609 ();
 FILLCELL_X4 FILLER_134_625 ();
 FILLCELL_X2 FILLER_134_629 ();
 FILLCELL_X32 FILLER_134_632 ();
 FILLCELL_X32 FILLER_134_664 ();
 FILLCELL_X32 FILLER_134_696 ();
 FILLCELL_X32 FILLER_134_728 ();
 FILLCELL_X32 FILLER_134_760 ();
 FILLCELL_X32 FILLER_134_792 ();
 FILLCELL_X32 FILLER_134_824 ();
 FILLCELL_X32 FILLER_134_856 ();
 FILLCELL_X32 FILLER_134_888 ();
 FILLCELL_X32 FILLER_134_920 ();
 FILLCELL_X32 FILLER_134_952 ();
 FILLCELL_X32 FILLER_134_984 ();
 FILLCELL_X4 FILLER_134_1016 ();
 FILLCELL_X2 FILLER_134_1020 ();
 FILLCELL_X32 FILLER_135_1 ();
 FILLCELL_X32 FILLER_135_33 ();
 FILLCELL_X32 FILLER_135_65 ();
 FILLCELL_X32 FILLER_135_97 ();
 FILLCELL_X32 FILLER_135_129 ();
 FILLCELL_X32 FILLER_135_161 ();
 FILLCELL_X32 FILLER_135_193 ();
 FILLCELL_X32 FILLER_135_225 ();
 FILLCELL_X32 FILLER_135_257 ();
 FILLCELL_X32 FILLER_135_289 ();
 FILLCELL_X32 FILLER_135_321 ();
 FILLCELL_X32 FILLER_135_353 ();
 FILLCELL_X32 FILLER_135_385 ();
 FILLCELL_X32 FILLER_135_417 ();
 FILLCELL_X32 FILLER_135_449 ();
 FILLCELL_X32 FILLER_135_481 ();
 FILLCELL_X32 FILLER_135_513 ();
 FILLCELL_X32 FILLER_135_545 ();
 FILLCELL_X32 FILLER_135_577 ();
 FILLCELL_X32 FILLER_135_609 ();
 FILLCELL_X32 FILLER_135_641 ();
 FILLCELL_X32 FILLER_135_673 ();
 FILLCELL_X32 FILLER_135_705 ();
 FILLCELL_X32 FILLER_135_737 ();
 FILLCELL_X32 FILLER_135_769 ();
 FILLCELL_X32 FILLER_135_801 ();
 FILLCELL_X32 FILLER_135_833 ();
 FILLCELL_X32 FILLER_135_865 ();
 FILLCELL_X32 FILLER_135_897 ();
 FILLCELL_X32 FILLER_135_929 ();
 FILLCELL_X32 FILLER_135_961 ();
 FILLCELL_X16 FILLER_135_993 ();
 FILLCELL_X8 FILLER_135_1009 ();
 FILLCELL_X4 FILLER_135_1017 ();
 FILLCELL_X1 FILLER_135_1021 ();
 FILLCELL_X4 FILLER_136_1 ();
 FILLCELL_X32 FILLER_136_9 ();
 FILLCELL_X32 FILLER_136_41 ();
 FILLCELL_X32 FILLER_136_73 ();
 FILLCELL_X32 FILLER_136_105 ();
 FILLCELL_X32 FILLER_136_137 ();
 FILLCELL_X32 FILLER_136_169 ();
 FILLCELL_X32 FILLER_136_201 ();
 FILLCELL_X32 FILLER_136_233 ();
 FILLCELL_X32 FILLER_136_265 ();
 FILLCELL_X32 FILLER_136_297 ();
 FILLCELL_X32 FILLER_136_329 ();
 FILLCELL_X32 FILLER_136_361 ();
 FILLCELL_X32 FILLER_136_393 ();
 FILLCELL_X32 FILLER_136_425 ();
 FILLCELL_X32 FILLER_136_457 ();
 FILLCELL_X32 FILLER_136_489 ();
 FILLCELL_X32 FILLER_136_521 ();
 FILLCELL_X32 FILLER_136_553 ();
 FILLCELL_X32 FILLER_136_585 ();
 FILLCELL_X8 FILLER_136_617 ();
 FILLCELL_X4 FILLER_136_625 ();
 FILLCELL_X2 FILLER_136_629 ();
 FILLCELL_X32 FILLER_136_632 ();
 FILLCELL_X32 FILLER_136_664 ();
 FILLCELL_X32 FILLER_136_696 ();
 FILLCELL_X32 FILLER_136_728 ();
 FILLCELL_X32 FILLER_136_760 ();
 FILLCELL_X32 FILLER_136_792 ();
 FILLCELL_X32 FILLER_136_824 ();
 FILLCELL_X32 FILLER_136_856 ();
 FILLCELL_X32 FILLER_136_888 ();
 FILLCELL_X32 FILLER_136_920 ();
 FILLCELL_X32 FILLER_136_952 ();
 FILLCELL_X32 FILLER_136_984 ();
 FILLCELL_X4 FILLER_136_1016 ();
 FILLCELL_X2 FILLER_136_1020 ();
 FILLCELL_X8 FILLER_137_1 ();
 FILLCELL_X4 FILLER_137_9 ();
 FILLCELL_X2 FILLER_137_13 ();
 FILLCELL_X32 FILLER_137_19 ();
 FILLCELL_X32 FILLER_137_51 ();
 FILLCELL_X8 FILLER_137_83 ();
 FILLCELL_X4 FILLER_137_91 ();
 FILLCELL_X2 FILLER_137_95 ();
 FILLCELL_X32 FILLER_137_100 ();
 FILLCELL_X32 FILLER_137_132 ();
 FILLCELL_X8 FILLER_137_164 ();
 FILLCELL_X2 FILLER_137_172 ();
 FILLCELL_X32 FILLER_137_177 ();
 FILLCELL_X32 FILLER_137_209 ();
 FILLCELL_X8 FILLER_137_241 ();
 FILLCELL_X2 FILLER_137_249 ();
 FILLCELL_X32 FILLER_137_254 ();
 FILLCELL_X32 FILLER_137_286 ();
 FILLCELL_X8 FILLER_137_318 ();
 FILLCELL_X4 FILLER_137_326 ();
 FILLCELL_X2 FILLER_137_330 ();
 FILLCELL_X1 FILLER_137_332 ();
 FILLCELL_X32 FILLER_137_336 ();
 FILLCELL_X32 FILLER_137_368 ();
 FILLCELL_X8 FILLER_137_400 ();
 FILLCELL_X2 FILLER_137_408 ();
 FILLCELL_X32 FILLER_137_413 ();
 FILLCELL_X32 FILLER_137_445 ();
 FILLCELL_X8 FILLER_137_477 ();
 FILLCELL_X4 FILLER_137_485 ();
 FILLCELL_X2 FILLER_137_489 ();
 FILLCELL_X1 FILLER_137_491 ();
 FILLCELL_X32 FILLER_137_495 ();
 FILLCELL_X32 FILLER_137_527 ();
 FILLCELL_X8 FILLER_137_559 ();
 FILLCELL_X2 FILLER_137_567 ();
 FILLCELL_X32 FILLER_137_572 ();
 FILLCELL_X16 FILLER_137_604 ();
 FILLCELL_X8 FILLER_137_620 ();
 FILLCELL_X2 FILLER_137_628 ();
 FILLCELL_X1 FILLER_137_630 ();
 FILLCELL_X8 FILLER_137_632 ();
 FILLCELL_X4 FILLER_137_640 ();
 FILLCELL_X2 FILLER_137_644 ();
 FILLCELL_X32 FILLER_137_650 ();
 FILLCELL_X32 FILLER_137_682 ();
 FILLCELL_X8 FILLER_137_714 ();
 FILLCELL_X4 FILLER_137_722 ();
 FILLCELL_X2 FILLER_137_726 ();
 FILLCELL_X32 FILLER_137_731 ();
 FILLCELL_X32 FILLER_137_763 ();
 FILLCELL_X8 FILLER_137_795 ();
 FILLCELL_X2 FILLER_137_803 ();
 FILLCELL_X32 FILLER_137_809 ();
 FILLCELL_X32 FILLER_137_841 ();
 FILLCELL_X8 FILLER_137_873 ();
 FILLCELL_X4 FILLER_137_881 ();
 FILLCELL_X2 FILLER_137_885 ();
 FILLCELL_X32 FILLER_137_890 ();
 FILLCELL_X32 FILLER_137_922 ();
 FILLCELL_X8 FILLER_137_954 ();
 FILLCELL_X2 FILLER_137_962 ();
 FILLCELL_X32 FILLER_137_967 ();
 FILLCELL_X16 FILLER_137_999 ();
 FILLCELL_X4 FILLER_137_1018 ();
 assign init_done = curr_state[1];
 assign valid_out = valid_reg_out;
endmodule
