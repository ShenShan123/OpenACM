module TAPCELL_X1 ();
endmodule

module FILL_X1 ();
endmodule