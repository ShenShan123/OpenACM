* 标准单元SPICE库



.SUBCKT NAND2_X1 A1 A2 ZN VDD VSS 
*.PININFO A1:I A2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(A1 * A2)
M_i_1 net_0 A2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 ZN A1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 ZN A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_2 VDD A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

.SUBCKT XNOR2_X1 A B ZN VDD VSS 
*.PININFO A:I B:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(A ^ B)
M_i_0 net_001 A net_000 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_5 VSS B net_001 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_11 net_002 net_000 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_17 ZN A net_002 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_23 net_002 B ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_29 net_000 A VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_36 VDD B net_000 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_42 ZN net_000 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_48 net_003 A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_53 VDD B net_003 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

.SUBCKT AOI22_X1 A1 A2 B1 B2 ZN VDD VSS 
*.PININFO A1:I A2:I B1:I B2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!((A1 * A2) + (B1 * B2))
M_i_3 net_1 B2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 ZN B1 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 net_0 A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1 VSS A2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_7 VDD B2 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6 net_2 B1 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4 ZN A1 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5 net_2 A2 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

.SUBCKT NAND3_X1 A1 A2 A3 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I ZN:O VDD:P VSS:G 
*.EQN ZN=!((A1 * A2) * A3)
M_i_2 net_1 A3 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1 net_0 A2 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 ZN A1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5 ZN A3 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4 VDD A2 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3 ZN A1 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

.SUBCKT XOR2_X1 A B Z VDD VSS 
*.PININFO A:I B:I Z:O VDD:P VSS:G 
*.EQN Z=(A ^ B)
M_i_0 net_000 A VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_7 VSS B net_000 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_13 Z net_000 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_19 net_001 A Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_24 VSS B net_001 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_30 net_002 A net_000 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_35 VDD B net_002 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_41 net_003 net_000 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_47 Z A net_003 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_53 net_003 B Z VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

.SUBCKT INV_X1 A ZN VDD VSS 
*.PININFO A:I ZN:O VDD:P VSS:G 
*.EQN ZN=!A
M_i_0 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

.SUBCKT OAI21_X1 A B1 B2 ZN VDD VSS 
*.PININFO A:I B1:I B2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(A * (B1 + B2))
M_i_1 ZN B2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 net_0 B1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 VSS A net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4 net_1 B2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3 ZN B1 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

.SUBCKT OR2_X1 A1 A2 ZN VDD VSS 
*.PININFO A1:I A2:I ZN:O VDD:P VSS:G 
*.EQN ZN=(A1 + A2)
M_i_2 ZN_neg A1 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_3 VSS A2 ZN_neg VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4 net_0 A1 ZN_neg VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_5 VDD A2 net_0 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

.SUBCKT AOI21_X1 A B1 B2 ZN VDD VSS 
*.PININFO A:I B1:I B2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(A + (B1 * B2))
M_i_1 net_0 B2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 ZN B1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4 ZN B2 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3 net_1 B1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5 VDD A net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS

.SUBCKT NOR2_X1 A1 A2 ZN VDD VSS 
*.PININFO A1:I A2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(A1 + A2)
M_i_1 ZN A2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 VSS A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 net_0 A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_2 ZN A1 net_0 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

.SUBCKT NOR3_X1 A1 A2 A3 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I ZN:O VDD:P VSS:G 
*.EQN ZN=!((A1 + A2) + A3)
M_i_2 ZN A3 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1 VSS A2 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 ZN A1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5 net_1 A3 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4 net_0 A2 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3 ZN A1 net_0 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

.SUBCKT AND2_X1 A1 A2 ZN VDD VSS 
*.PININFO A1:I A2:I ZN:O VDD:P VSS:G 
*.EQN ZN=(A1 * A2)
M_i_2 net_0 A1 ZN_neg VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_3 VSS A2 net_0 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4 ZN_neg A1 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_5 VDD A2 ZN_neg VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

.SUBCKT OAI22_X1 A1 A2 B1 B2 ZN VDD VSS 
*.PININFO A1:I A2:I B1:I B2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!((A1 + A2) * (B1 + B2))
M_i_3 VSS B2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 net_0 B1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 ZN A1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1 net_0 A2 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_7 net_2 B2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6 ZN B1 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4 net_1 A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5 VDD A2 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

.SUBCKT OR3_X1 A1 A2 A3 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I ZN:O VDD:P VSS:G 
*.EQN ZN=((A1 + A2) + A3)
M_i_2 VSS A1 ZN_neg VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_3 ZN_neg A2 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_4 VSS A3 ZN_neg VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5 net_0 A1 ZN_neg VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_6 net_1 A2 net_0 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_7 VDD A3 net_1 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

.SUBCKT BUF_X1 A Z VDD VSS 
*.PININFO A:I Z:O VDD:P VSS:G 
*.EQN Z=A
M_i_2 VSS A Z_neg VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_0 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 VDD A Z_neg VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_1 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS

.SUBCKT AND3_X1 A1 A2 A3 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I ZN:O VDD:P VSS:G 
*.EQN ZN=((A1 * A2) * A3)
M_i_2 net_0 A1 ZN_neg VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_3 net_1 A2 net_0 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_4 VSS A3 net_1 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5 VDD A1 ZN_neg VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_6 ZN_neg A2 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_7 VDD A3 ZN_neg VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

.SUBCKT MUX2_X1 A B S Z VDD VSS 
*.PININFO A:I B:I S:I Z:O VDD:P VSS:G 
*.EQN Z=((S * B) + (A * !S))
M_i_10 VSS S x1 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_4 net_1 A VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_5 Z_neg x1 net_1 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_2 Z_neg S net_0 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_3 net_0 B VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_0 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_11 VDD S x1 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_8 VDD A net_2 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_6 net_2 S Z_neg VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_9 net_3 x1 Z_neg VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_7 VDD B net_3 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_1 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

.SUBCKT NAND4_X1 A1 A2 A3 A4 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I A4:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(((A1 * A2) * A3) * A4)
M_i_3 net_2 A4 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 net_1 A3 net_2 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1 net_0 A2 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 ZN A1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_7 ZN A4 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6 VDD A3 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5 ZN A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4 VDD A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

.SUBCKT DFFR_X1 D RN CK Q QN VDD VSS 
*.PININFO D:I RN:I CK:I Q:O QN:O VDD:P VSS:G 
M_i_0 VSS CK net_000 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_7 net_001 net_000 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_13 net_002 D VSS VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_18 net_003 net_000 net_002 VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_24 net_004 net_001 net_003 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_28 net_005 net_006 net_004 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_32 VSS RN net_005 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_38 VSS net_003 net_006 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_45 net_007 net_003 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_49 net_008 net_001 net_007 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_55 net_009 net_000 net_008 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_59 VSS net_011 net_009 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_65 net_010 RN VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_70 net_011 net_008 net_010 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_76 VSS net_008 QN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_83 Q net_011 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_89 VDD CK net_000 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_96 net_001 net_000 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_103 net_012 D VDD VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_108 net_003 net_001 net_012 VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_114 net_013 net_000 net_003 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_119 VDD net_006 net_013 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_125 net_013 RN VDD VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_136 VDD net_003 net_006 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_143 net_015 net_003 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_147 net_008 net_000 net_015 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_153 net_016 net_001 net_008 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_159 VDD net_011 net_016 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_165 net_011 RN VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_172 VDD net_008 net_011 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_180 VDD net_008 QN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_187 Q net_011 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 