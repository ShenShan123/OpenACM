module sram_multiplier_system (clk,
    init_done,
    init_enable,
    pe_ce,
    rst_n,
    valid_out,
    data_in,
    data_out);
 input clk;
 output init_done;
 input init_enable;
 input pe_ce;
 input rst_n;
 output valid_out;
 input [7:0] data_in;
 output [15:0] data_out;

 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire \u_multiplier/_0345_ ;
 wire \u_multiplier/_0346_ ;
 wire \u_multiplier/_0347_ ;
 wire \u_multiplier/_0348_ ;
 wire \u_multiplier/_0349_ ;
 wire \u_multiplier/_0350_ ;
 wire \u_multiplier/_0351_ ;
 wire \u_multiplier/_0352_ ;
 wire \u_multiplier/_0353_ ;
 wire \u_multiplier/_0354_ ;
 wire \u_multiplier/_0355_ ;
 wire \u_multiplier/_0392_ ;
 wire \u_multiplier/_0393_ ;
 wire \u_multiplier/_0394_ ;
 wire \u_multiplier/_0395_ ;
 wire \u_multiplier/_0396_ ;
 wire \u_multiplier/_0397_ ;
 wire \u_multiplier/_0398_ ;
 wire \u_multiplier/_0399_ ;
 wire \u_multiplier/_0400_ ;
 wire \u_multiplier/_0401_ ;
 wire \u_multiplier/_0402_ ;
 wire \u_multiplier/_0403_ ;
 wire \u_multiplier/_0404_ ;
 wire \u_multiplier/_0405_ ;
 wire \u_multiplier/_0406_ ;
 wire \u_multiplier/_0407_ ;
 wire \u_multiplier/_0408_ ;
 wire \u_multiplier/_0409_ ;
 wire \u_multiplier/_0410_ ;
 wire \u_multiplier/_0411_ ;
 wire \u_multiplier/_0412_ ;
 wire \u_multiplier/_0413_ ;
 wire \u_multiplier/_0414_ ;
 wire \u_multiplier/_0415_ ;
 wire \u_multiplier/_0416_ ;
 wire \u_multiplier/_0417_ ;
 wire \u_multiplier/_0418_ ;
 wire \u_multiplier/_0419_ ;
 wire \u_multiplier/_0420_ ;
 wire \u_multiplier/_0421_ ;
 wire \u_multiplier/_0422_ ;
 wire \u_multiplier/_0423_ ;
 wire \u_multiplier/_0424_ ;
 wire \u_multiplier/_0425_ ;
 wire \u_multiplier/_0426_ ;
 wire \u_multiplier/_0427_ ;
 wire \u_multiplier/_0428_ ;
 wire \u_multiplier/_0429_ ;
 wire \u_multiplier/_0430_ ;
 wire \u_multiplier/_0431_ ;
 wire \u_multiplier/_0432_ ;
 wire \u_multiplier/_0433_ ;
 wire \u_multiplier/_0434_ ;
 wire \u_multiplier/_0435_ ;
 wire \u_multiplier/_0436_ ;
 wire \u_multiplier/_0437_ ;
 wire \u_multiplier/_0438_ ;
 wire \u_multiplier/_0439_ ;
 wire \u_multiplier/_0440_ ;
 wire \u_multiplier/_0441_ ;
 wire \u_multiplier/_0442_ ;
 wire \u_multiplier/_0443_ ;
 wire \u_multiplier/_0444_ ;
 wire \u_multiplier/_0445_ ;
 wire \u_multiplier/_0446_ ;
 wire \u_multiplier/_0447_ ;
 wire \u_multiplier/_0448_ ;
 wire \u_multiplier/_0449_ ;
 wire \u_multiplier/_0450_ ;
 wire \u_multiplier/_0451_ ;
 wire \u_multiplier/_0452_ ;
 wire \u_multiplier/_0453_ ;
 wire \u_multiplier/_0454_ ;
 wire \u_multiplier/_0455_ ;
 wire \u_multiplier/_0456_ ;
 wire \u_multiplier/_0457_ ;
 wire \u_multiplier/_0458_ ;
 wire \u_multiplier/_0459_ ;
 wire \u_multiplier/_0460_ ;
 wire \u_multiplier/_0461_ ;
 wire \u_multiplier/_0462_ ;
 wire \u_multiplier/_0463_ ;
 wire \u_multiplier/_0464_ ;
 wire \u_multiplier/_0465_ ;
 wire \u_multiplier/_0466_ ;
 wire \u_multiplier/_0467_ ;
 wire \u_multiplier/_0468_ ;
 wire \u_multiplier/_0469_ ;
 wire \u_multiplier/_0470_ ;
 wire \u_multiplier/_0471_ ;
 wire \u_multiplier/_0472_ ;
 wire \u_multiplier/_0473_ ;
 wire \u_multiplier/_0474_ ;
 wire \u_multiplier/_0475_ ;
 wire \u_multiplier/_0476_ ;
 wire \u_multiplier/_0477_ ;
 wire \u_multiplier/_0478_ ;
 wire \u_multiplier/_0479_ ;
 wire \u_multiplier/_0480_ ;
 wire \u_multiplier/_0481_ ;
 wire \u_multiplier/_0482_ ;
 wire \u_multiplier/_0483_ ;
 wire \u_multiplier/_0484_ ;
 wire \u_multiplier/_0485_ ;
 wire \u_multiplier/_0486_ ;
 wire \u_multiplier/_0487_ ;
 wire \u_multiplier/_0488_ ;
 wire \u_multiplier/_0489_ ;
 wire \u_multiplier/_0490_ ;
 wire \u_multiplier/_0491_ ;
 wire \u_multiplier/_0492_ ;
 wire \u_multiplier/_0493_ ;
 wire \u_multiplier/_0494_ ;
 wire \u_multiplier/_0495_ ;
 wire \u_multiplier/_0496_ ;
 wire \u_multiplier/_0497_ ;
 wire \u_multiplier/_0498_ ;
 wire \u_multiplier/_0499_ ;
 wire \u_multiplier/_0500_ ;
 wire \u_multiplier/_0501_ ;
 wire \u_multiplier/_0502_ ;
 wire \u_multiplier/_0503_ ;
 wire \u_multiplier/_0504_ ;
 wire \u_multiplier/_0505_ ;
 wire \u_multiplier/_0506_ ;
 wire \u_multiplier/_0507_ ;
 wire \u_multiplier/_0508_ ;
 wire \u_multiplier/_0509_ ;
 wire \u_multiplier/_0510_ ;
 wire \u_multiplier/_0511_ ;
 wire \u_multiplier/_0512_ ;
 wire \u_multiplier/_0513_ ;
 wire \u_multiplier/_0514_ ;
 wire \u_multiplier/_0515_ ;
 wire \u_multiplier/_0516_ ;
 wire \u_multiplier/_0517_ ;
 wire \u_multiplier/_0518_ ;
 wire \u_multiplier/_0519_ ;
 wire \u_multiplier/_0520_ ;
 wire \u_multiplier/_0521_ ;
 wire \u_multiplier/_0522_ ;
 wire \u_multiplier/_0523_ ;
 wire \u_multiplier/_0524_ ;
 wire \u_multiplier/_0525_ ;
 wire \u_multiplier/_0526_ ;
 wire \u_multiplier/_0527_ ;
 wire \u_multiplier/_0528_ ;
 wire \u_multiplier/_0529_ ;
 wire \u_multiplier/_0530_ ;
 wire \u_multiplier/_0531_ ;
 wire \u_multiplier/_0532_ ;
 wire \u_multiplier/_0533_ ;
 wire \u_multiplier/_0534_ ;
 wire \u_multiplier/_0535_ ;
 wire \u_multiplier/_0536_ ;
 wire \u_multiplier/_0537_ ;
 wire \u_multiplier/_0538_ ;
 wire \u_multiplier/_0539_ ;
 wire \u_multiplier/_0540_ ;
 wire \u_multiplier/_0541_ ;
 wire \u_multiplier/_0542_ ;
 wire \u_multiplier/_0543_ ;
 wire \u_multiplier/_0544_ ;
 wire \u_multiplier/_0545_ ;
 wire \u_multiplier/_0546_ ;
 wire \u_multiplier/_0547_ ;
 wire \u_multiplier/_0548_ ;
 wire \u_multiplier/_0549_ ;
 wire \u_multiplier/_0550_ ;
 wire \u_multiplier/_0551_ ;
 wire \u_multiplier/_0552_ ;
 wire \u_multiplier/_0553_ ;
 wire \u_multiplier/_0554_ ;
 wire \u_multiplier/_0555_ ;
 wire \u_multiplier/_0556_ ;
 wire \u_multiplier/_0557_ ;
 wire \u_multiplier/_0558_ ;
 wire \u_multiplier/_0559_ ;
 wire \u_multiplier/_0560_ ;
 wire \u_multiplier/_0561_ ;
 wire \u_multiplier/_0562_ ;
 wire \u_multiplier/_0563_ ;
 wire \u_multiplier/_0564_ ;
 wire \u_multiplier/_0565_ ;
 wire \u_multiplier/_0566_ ;
 wire \u_multiplier/_0567_ ;
 wire \u_multiplier/_0568_ ;
 wire \u_multiplier/_0569_ ;
 wire \u_multiplier/_0570_ ;
 wire \u_multiplier/_0571_ ;
 wire \u_multiplier/_0572_ ;
 wire \u_multiplier/_0573_ ;
 wire \u_multiplier/_0574_ ;
 wire \u_multiplier/_0575_ ;
 wire \u_multiplier/_0576_ ;
 wire \u_multiplier/_0577_ ;
 wire \u_multiplier/_0578_ ;
 wire \u_multiplier/_0579_ ;
 wire \u_multiplier/_0580_ ;
 wire \u_multiplier/_0581_ ;
 wire \u_multiplier/_0582_ ;
 wire \u_multiplier/_0583_ ;
 wire \u_multiplier/_0584_ ;
 wire \u_multiplier/_0585_ ;
 wire \u_multiplier/_0586_ ;
 wire \u_multiplier/_0587_ ;
 wire \u_multiplier/_0588_ ;
 wire \u_multiplier/_0589_ ;
 wire \u_multiplier/_0590_ ;
 wire \u_multiplier/_0591_ ;
 wire \u_multiplier/_0592_ ;
 wire \u_multiplier/_0593_ ;
 wire \u_multiplier/_0594_ ;
 wire \u_multiplier/_0595_ ;
 wire \u_multiplier/_0596_ ;
 wire \u_multiplier/_0597_ ;
 wire \u_multiplier/_0598_ ;
 wire \u_multiplier/_0599_ ;
 wire \u_multiplier/_0600_ ;
 wire \u_multiplier/_0601_ ;
 wire \u_multiplier/_0602_ ;
 wire \u_multiplier/_0603_ ;
 wire \u_multiplier/_0604_ ;
 wire \u_multiplier/_0605_ ;
 wire \u_multiplier/_0606_ ;
 wire \u_multiplier/_0607_ ;
 wire \u_multiplier/_0608_ ;
 wire \u_multiplier/_0609_ ;
 wire \u_multiplier/_0610_ ;
 wire \u_multiplier/_0611_ ;
 wire \u_multiplier/_0612_ ;
 wire \u_multiplier/_0613_ ;
 wire \u_multiplier/_0614_ ;
 wire \u_multiplier/_0615_ ;
 wire \u_multiplier/_0616_ ;
 wire \u_multiplier/_0617_ ;
 wire \u_multiplier/_0618_ ;
 wire \u_multiplier/_0619_ ;
 wire \u_multiplier/_0620_ ;
 wire \u_multiplier/_0621_ ;
 wire \u_multiplier/_0622_ ;
 wire \u_multiplier/_0623_ ;
 wire \u_multiplier/_0624_ ;
 wire \u_multiplier/_0625_ ;
 wire \u_multiplier/_0626_ ;
 wire \u_multiplier/_0627_ ;
 wire \u_multiplier/_0628_ ;
 wire \u_multiplier/_0629_ ;
 wire \u_multiplier/_0630_ ;
 wire \u_multiplier/_0631_ ;
 wire \u_multiplier/_0632_ ;
 wire \u_multiplier/_0633_ ;
 wire \u_multiplier/_0634_ ;
 wire \u_multiplier/_0635_ ;
 wire \u_multiplier/_0636_ ;
 wire \u_multiplier/_0637_ ;
 wire \u_multiplier/_0638_ ;
 wire \u_multiplier/_0639_ ;
 wire \u_multiplier/_0640_ ;
 wire \u_multiplier/_0641_ ;
 wire \u_multiplier/_0642_ ;
 wire \u_multiplier/_0643_ ;
 wire \u_multiplier/_0644_ ;
 wire \u_multiplier/_0645_ ;
 wire \u_multiplier/_0646_ ;
 wire \u_multiplier/_0647_ ;
 wire \u_multiplier/_0648_ ;
 wire \u_multiplier/_0649_ ;
 wire \u_multiplier/_0650_ ;
 wire \u_multiplier/_0651_ ;
 wire \u_multiplier/_0652_ ;
 wire \u_multiplier/_0653_ ;
 wire \u_multiplier/_0654_ ;
 wire \u_multiplier/_0655_ ;
 wire \u_multiplier/_0656_ ;
 wire \u_multiplier/_0657_ ;
 wire \u_multiplier/_0658_ ;
 wire \u_multiplier/_0659_ ;
 wire \u_multiplier/_0660_ ;
 wire \u_multiplier/_0661_ ;
 wire \u_multiplier/_0662_ ;
 wire \u_multiplier/_0663_ ;
 wire \u_multiplier/_0664_ ;
 wire \u_multiplier/_0665_ ;
 wire \u_multiplier/_0666_ ;
 wire \u_multiplier/_0667_ ;
 wire \u_multiplier/_0668_ ;
 wire \u_multiplier/_0669_ ;
 wire \u_multiplier/_0670_ ;
 wire \u_multiplier/_0671_ ;
 wire \u_multiplier/_0672_ ;
 wire \u_multiplier/_0673_ ;
 wire \u_multiplier/_0674_ ;
 wire \u_multiplier/_0675_ ;
 wire \u_multiplier/_0676_ ;
 wire \u_multiplier/_0677_ ;
 wire \u_multiplier/_0678_ ;
 wire \u_multiplier/_0679_ ;
 wire \u_multiplier/_0680_ ;
 wire \u_multiplier/_0681_ ;
 wire \u_multiplier/_0682_ ;
 wire \u_multiplier/_0683_ ;
 wire \u_multiplier/_0684_ ;
 wire \u_multiplier/_0685_ ;
 wire \u_multiplier/_0686_ ;
 wire \u_multiplier/_0687_ ;
 wire \u_multiplier/_0688_ ;
 wire \u_multiplier/_0689_ ;
 wire \u_multiplier/_0690_ ;
 wire \u_multiplier/_0691_ ;
 wire \u_multiplier/_0692_ ;
 wire \u_multiplier/_0693_ ;
 wire \u_multiplier/_0694_ ;
 wire \u_multiplier/_0695_ ;
 wire \u_multiplier/_0696_ ;
 wire \u_multiplier/_0697_ ;
 wire \u_multiplier/_0698_ ;
 wire \u_multiplier/_0699_ ;
 wire \u_multiplier/_0700_ ;
 wire \u_multiplier/_0701_ ;
 wire \u_multiplier/_0702_ ;
 wire \u_multiplier/_0703_ ;
 wire \u_multiplier/_0704_ ;
 wire \u_multiplier/_0705_ ;
 wire \u_multiplier/_0706_ ;
 wire \u_multiplier/_0707_ ;
 wire \u_multiplier/_0708_ ;
 wire \u_multiplier/_0709_ ;
 wire \u_multiplier/_0710_ ;
 wire \u_multiplier/_0711_ ;
 wire \u_multiplier/_0712_ ;
 wire \u_multiplier/_0713_ ;
 wire \u_multiplier/_0714_ ;
 wire \u_multiplier/_0715_ ;
 wire \u_multiplier/_0716_ ;
 wire \u_multiplier/_0717_ ;
 wire \u_multiplier/_0718_ ;
 wire \u_multiplier/_0719_ ;
 wire \u_multiplier/_0720_ ;
 wire \u_multiplier/_0721_ ;
 wire \u_multiplier/_0722_ ;
 wire \u_multiplier/_0723_ ;
 wire net30;
 wire \u_multiplier/zero_x ;
 wire \u_multiplier/zero_y ;
 wire \u_multiplier/LODx/_12_ ;
 wire \u_multiplier/LODx/_13_ ;
 wire \u_multiplier/LODx/Middle/_3_ ;
 wire \u_multiplier/LODx/lod2_0/_09_ ;
 wire \u_multiplier/LODx/lod2_0/_10_ ;
 wire \u_multiplier/LODx/lod2_0/_11_ ;
 wire \u_multiplier/LODx/lod2_1/_09_ ;
 wire \u_multiplier/LODx/lod2_1/_10_ ;
 wire \u_multiplier/LODx/lod2_1/_11_ ;
 wire \u_multiplier/LODy/_12_ ;
 wire \u_multiplier/LODy/_13_ ;
 wire \u_multiplier/LODy/Middle/_3_ ;
 wire \u_multiplier/LODy/lod2_0/_09_ ;
 wire \u_multiplier/LODy/lod2_0/_10_ ;
 wire \u_multiplier/LODy/lod2_0/_11_ ;
 wire \u_multiplier/LODy/lod2_1/_09_ ;
 wire \u_multiplier/LODy/lod2_1/_10_ ;
 wire \u_multiplier/LODy/lod2_1/_11_ ;
 wire \u_multiplier/NOD/_11_ ;
 wire \u_multiplier/NOD/_12_ ;
 wire \u_multiplier/NOD/_13_ ;
 wire net31;
 wire \u_multiplier/NOD/nod_basic_unit15/_5_ ;
 wire \u_multiplier/NOD/nod_cels[2].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[2].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[2].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[2].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[3].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[3].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[3].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[3].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[4].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[4].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[4].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[4].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[5].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[5].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[5].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[5].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/dec/_34_ ;
 wire \u_multiplier/dec/_35_ ;
 wire \u_multiplier/dec/_36_ ;
 wire \u_multiplier/dec/_37_ ;
 wire \u_multiplier/dec/_38_ ;
 wire \u_multiplier/dec/_39_ ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire valid_reg_out;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire [3:0] addr_ptr;
 wire [2:0] curr_state;
 wire [7:0] data_in_reg;
 wire [3:0] init_count;
 wire [15:0] product;
 wire [7:0] sram_rdata;
 wire [7:0] sram_rdata_reg;
 wire [2:0] \u_multiplier/K ;
 wire [1:0] \u_multiplier/LODx/select ;
 wire [7:0] \u_multiplier/LODx/z ;
 wire [1:0] \u_multiplier/LODy/select ;
 wire [7:0] \u_multiplier/LODy/z ;
 wire [4:0] \u_multiplier/NOD/t_in ;
 wire [7:0] \u_multiplier/NOD_Q1 ;
 wire [2:0] \u_multiplier/code_x ;
 wire [2:0] \u_multiplier/code_y ;
 wire [15:0] \u_multiplier/dec_out ;
 wire [7:0] \u_multiplier/kx ;
 wire [7:0] \u_multiplier/ky ;

 INV_X2 _281_ (.A(net11),
    .ZN(_165_));
 INV_X4 _282_ (.A(net10),
    .ZN(_134_));
 INV_X1 _283_ (.A(init_count[2]),
    .ZN(_166_));
 INV_X1 _284_ (.A(addr_ptr[0]),
    .ZN(_167_));
 INV_X1 _285_ (.A(addr_ptr[3]),
    .ZN(_168_));
 NAND2_X2 _286_ (.A1(net11),
    .A2(net82),
    .ZN(_135_));
 NAND2_X1 _287_ (.A1(init_count[3]),
    .A2(init_count[2]),
    .ZN(_169_));
 NAND2_X1 _288_ (.A1(init_count[1]),
    .A2(init_count[0]),
    .ZN(_170_));
 NAND4_X4 _289_ (.A1(init_count[1]),
    .A2(init_count[0]),
    .A3(init_count[3]),
    .A4(init_count[2]),
    .ZN(_171_));
 NOR2_X1 _290_ (.A1(_134_),
    .A2(_171_),
    .ZN(_172_));
 NAND3_X1 _291_ (.A1(net11),
    .A2(net10),
    .A3(net9),
    .ZN(_173_));
 OAI22_X1 _292_ (.A1(_135_),
    .A2(_172_),
    .B1(_173_),
    .B2(net57),
    .ZN(_133_));
 OR2_X1 _293_ (.A1(_165_),
    .A2(net85),
    .ZN(_174_));
 AND2_X1 _294_ (.A1(_173_),
    .A2(_174_),
    .ZN(_131_));
 AND2_X4 _295_ (.A1(net11),
    .A2(net12),
    .ZN(_130_));
 NOR3_X1 _296_ (.A1(_134_),
    .A2(_135_),
    .A3(_171_),
    .ZN(_175_));
 OR2_X1 _297_ (.A1(_130_),
    .A2(_175_),
    .ZN(_132_));
 AND2_X1 _298_ (.A1(net11),
    .A2(sram_rdata[0]),
    .ZN(_122_));
 AND2_X1 _299_ (.A1(net11),
    .A2(sram_rdata[1]),
    .ZN(_123_));
 AND2_X1 _300_ (.A1(net11),
    .A2(sram_rdata[2]),
    .ZN(_124_));
 AND2_X1 _301_ (.A1(net11),
    .A2(sram_rdata[3]),
    .ZN(_125_));
 AND2_X1 _302_ (.A1(net11),
    .A2(sram_rdata[4]),
    .ZN(_126_));
 AND2_X1 _303_ (.A1(net11),
    .A2(sram_rdata[5]),
    .ZN(_127_));
 AND2_X1 _304_ (.A1(net11),
    .A2(sram_rdata[6]),
    .ZN(_128_));
 AND2_X1 _305_ (.A1(net11),
    .A2(sram_rdata[7]),
    .ZN(_129_));
 AND2_X1 _306_ (.A1(product[0]),
    .A2(_130_),
    .ZN(_102_));
 AND2_X1 _307_ (.A1(product[1]),
    .A2(_130_),
    .ZN(_109_));
 AND2_X1 _308_ (.A1(product[2]),
    .A2(_130_),
    .ZN(_110_));
 AND2_X1 _309_ (.A1(product[3]),
    .A2(_130_),
    .ZN(_111_));
 AND2_X1 _310_ (.A1(product[4]),
    .A2(_130_),
    .ZN(_112_));
 AND2_X1 _311_ (.A1(product[5]),
    .A2(_130_),
    .ZN(_113_));
 AND2_X1 _312_ (.A1(product[6]),
    .A2(_130_),
    .ZN(_114_));
 AND2_X1 _313_ (.A1(product[7]),
    .A2(_130_),
    .ZN(_115_));
 AND2_X1 _314_ (.A1(product[8]),
    .A2(_130_),
    .ZN(_116_));
 AND2_X1 _315_ (.A1(product[9]),
    .A2(_130_),
    .ZN(_117_));
 AND2_X1 _316_ (.A1(product[10]),
    .A2(_130_),
    .ZN(_103_));
 AND2_X1 _317_ (.A1(product[11]),
    .A2(_130_),
    .ZN(_104_));
 AND2_X1 _318_ (.A1(product[12]),
    .A2(_130_),
    .ZN(_105_));
 AND2_X1 _319_ (.A1(product[13]),
    .A2(_130_),
    .ZN(_106_));
 AND2_X1 _320_ (.A1(product[14]),
    .A2(_130_),
    .ZN(_107_));
 AND2_X1 _321_ (.A1(product[15]),
    .A2(_130_),
    .ZN(_108_));
 AND2_X1 _322_ (.A1(net11),
    .A2(net1),
    .ZN(_094_));
 AND2_X1 _323_ (.A1(net11),
    .A2(net2),
    .ZN(_095_));
 AND2_X1 _324_ (.A1(net11),
    .A2(net3),
    .ZN(_096_));
 AND2_X1 _325_ (.A1(net11),
    .A2(net4),
    .ZN(_097_));
 AND2_X1 _326_ (.A1(net11),
    .A2(net5),
    .ZN(_098_));
 AND2_X1 _327_ (.A1(net11),
    .A2(net6),
    .ZN(_099_));
 AND2_X1 _328_ (.A1(net11),
    .A2(net7),
    .ZN(_100_));
 AND2_X1 _329_ (.A1(net11),
    .A2(net8),
    .ZN(_101_));
 OAI21_X1 _330_ (.A(init_count[0]),
    .B1(_269_),
    .B2(_169_),
    .ZN(_176_));
 AOI221_X2 _331_ (.A(_134_),
    .B1(init_count[0]),
    .B2(net12),
    .C1(_176_),
    .C2(curr_state[2]),
    .ZN(_177_));
 AOI211_X1 _332_ (.A(_165_),
    .B(_177_),
    .C1(net61),
    .C2(_134_),
    .ZN(_118_));
 NAND3_X1 _333_ (.A1(init_count[1]),
    .A2(init_count[0]),
    .A3(_169_),
    .ZN(_178_));
 AOI21_X1 _334_ (.A(_134_),
    .B1(init_count[1]),
    .B2(net12),
    .ZN(_179_));
 OAI211_X1 _335_ (.A(curr_state[2]),
    .B(_178_),
    .C1(init_count[1]),
    .C2(init_count[0]),
    .ZN(_180_));
 AOI221_X1 _336_ (.A(_165_),
    .B1(_134_),
    .B2(net79),
    .C1(_179_),
    .C2(_180_),
    .ZN(_119_));
 OR2_X1 _337_ (.A1(init_count[3]),
    .A2(_166_),
    .ZN(_181_));
 NAND2_X1 _338_ (.A1(_166_),
    .A2(_170_),
    .ZN(_182_));
 OAI211_X1 _339_ (.A(curr_state[2]),
    .B(_182_),
    .C1(_181_),
    .C2(_170_),
    .ZN(_183_));
 AOI21_X1 _340_ (.A(_134_),
    .B1(init_count[2]),
    .B2(net12),
    .ZN(_184_));
 AOI221_X1 _341_ (.A(_165_),
    .B1(_134_),
    .B2(net72),
    .C1(_183_),
    .C2(_184_),
    .ZN(_120_));
 NAND2_X1 _342_ (.A1(init_count[3]),
    .A2(net12),
    .ZN(_185_));
 OAI21_X1 _343_ (.A(net76),
    .B1(_170_),
    .B2(net71),
    .ZN(_186_));
 OAI21_X1 _344_ (.A(_186_),
    .B1(curr_state[2]),
    .B2(_134_),
    .ZN(_187_));
 AOI221_X1 _345_ (.A(_165_),
    .B1(_134_),
    .B2(net39),
    .C1(_185_),
    .C2(_187_),
    .ZN(_121_));
 NAND3_X1 _346_ (.A1(curr_state[2]),
    .A2(net63),
    .A3(_171_),
    .ZN(_188_));
 AOI21_X1 _347_ (.A(_134_),
    .B1(net12),
    .B2(_167_),
    .ZN(_189_));
 AOI221_X1 _348_ (.A(_165_),
    .B1(_134_),
    .B2(net40),
    .C1(net64),
    .C2(_189_),
    .ZN(_090_));
 AOI21_X2 _349_ (.A(net12),
    .B1(_171_),
    .B2(curr_state[2]),
    .ZN(_190_));
 NAND2_X1 _350_ (.A1(addr_ptr[0]),
    .A2(addr_ptr[1]),
    .ZN(_191_));
 XNOR2_X1 _351_ (.A(addr_ptr[0]),
    .B(addr_ptr[1]),
    .ZN(_192_));
 OAI21_X1 _352_ (.A(net10),
    .B1(_190_),
    .B2(_192_),
    .ZN(_193_));
 AOI21_X1 _353_ (.A(_165_),
    .B1(_134_),
    .B2(net47),
    .ZN(_194_));
 AND2_X1 _354_ (.A1(_193_),
    .A2(net48),
    .ZN(_091_));
 XOR2_X1 _355_ (.A(addr_ptr[2]),
    .B(_191_),
    .Z(_195_));
 OAI21_X1 _356_ (.A(net10),
    .B1(_190_),
    .B2(_195_),
    .ZN(_196_));
 AOI21_X1 _357_ (.A(_165_),
    .B1(_134_),
    .B2(net49),
    .ZN(_197_));
 AND2_X1 _358_ (.A1(_196_),
    .A2(net50),
    .ZN(_092_));
 AOI21_X1 _359_ (.A(_168_),
    .B1(_171_),
    .B2(curr_state[2]),
    .ZN(_198_));
 NAND4_X1 _360_ (.A1(net10),
    .A2(addr_ptr[0]),
    .A3(addr_ptr[1]),
    .A4(addr_ptr[2]),
    .ZN(_199_));
 OR2_X1 _361_ (.A1(_198_),
    .A2(_199_),
    .ZN(_200_));
 OAI21_X1 _362_ (.A(net11),
    .B1(net53),
    .B2(_199_),
    .ZN(_201_));
 AOI221_X1 _363_ (.A(net54),
    .B1(_200_),
    .B2(net34),
    .C1(net10),
    .C2(_190_),
    .ZN(_093_));
 DFF_X1 _364_ (.D(_102_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net13),
    .QN(_228_));
 DFF_X1 _365_ (.D(_109_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net20),
    .QN(_229_));
 DFF_X1 _366_ (.D(_110_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net21),
    .QN(_230_));
 DFF_X1 _367_ (.D(_111_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net22),
    .QN(_231_));
 DFF_X1 _368_ (.D(_112_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net23),
    .QN(_232_));
 DFF_X2 _369_ (.D(_113_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net24),
    .QN(_233_));
 DFF_X1 _370_ (.D(_114_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net25),
    .QN(_234_));
 DFF_X1 _371_ (.D(_115_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net26),
    .QN(_235_));
 DFF_X1 _372_ (.D(_116_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net27),
    .QN(_236_));
 DFF_X2 _373_ (.D(_117_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net28),
    .QN(_237_));
 DFF_X1 _374_ (.D(_103_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net14),
    .QN(_238_));
 DFF_X1 _375_ (.D(_104_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net15),
    .QN(_239_));
 DFF_X1 _376_ (.D(_105_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net16),
    .QN(_240_));
 DFF_X1 _377_ (.D(_106_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net17),
    .QN(_241_));
 DFF_X1 _378_ (.D(_107_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net18),
    .QN(_242_));
 DFF_X1 _379_ (.D(_108_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net19),
    .QN(_243_));
 DFF_X1 _380_ (.D(_131_),
    .CK(clknet_2_1__leaf_clk),
    .Q(curr_state[0]),
    .QN(_244_));
 DFF_X2 _381_ (.D(_132_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net12),
    .QN(_245_));
 DFF_X2 _382_ (.D(net58),
    .CK(clknet_2_1__leaf_clk),
    .Q(curr_state[2]),
    .QN(_246_));
 DFF_X2 _383_ (.D(_094_),
    .CK(clknet_2_0__leaf_clk),
    .Q(data_in_reg[0]),
    .QN(_247_));
 DFF_X2 _384_ (.D(_095_),
    .CK(clknet_2_2__leaf_clk),
    .Q(data_in_reg[1]),
    .QN(_248_));
 DFF_X2 _385_ (.D(_096_),
    .CK(clknet_2_2__leaf_clk),
    .Q(data_in_reg[2]),
    .QN(_249_));
 DFF_X2 _386_ (.D(_097_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\u_multiplier/LODx/z [3]),
    .QN(_250_));
 DFF_X2 _387_ (.D(_098_),
    .CK(clknet_2_2__leaf_clk),
    .Q(data_in_reg[4]),
    .QN(_251_));
 DFF_X2 _388_ (.D(_099_),
    .CK(clknet_2_2__leaf_clk),
    .Q(data_in_reg[5]),
    .QN(_252_));
 DFF_X2 _389_ (.D(_100_),
    .CK(clknet_2_0__leaf_clk),
    .Q(data_in_reg[6]),
    .QN(_253_));
 DFF_X2 _390_ (.D(_101_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\u_multiplier/LODx/z [7]),
    .QN(_254_));
 DFF_X2 _391_ (.D(_122_),
    .CK(clknet_2_0__leaf_clk),
    .Q(sram_rdata_reg[0]),
    .QN(_255_));
 DFF_X2 _392_ (.D(_123_),
    .CK(clknet_2_0__leaf_clk),
    .Q(sram_rdata_reg[1]),
    .QN(_256_));
 DFF_X2 _393_ (.D(_124_),
    .CK(clknet_2_0__leaf_clk),
    .Q(sram_rdata_reg[2]),
    .QN(_257_));
 DFF_X2 _394_ (.D(_125_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\u_multiplier/LODy/z [3]),
    .QN(_258_));
 DFF_X2 _395_ (.D(_126_),
    .CK(clknet_2_2__leaf_clk),
    .Q(sram_rdata_reg[4]),
    .QN(_259_));
 DFF_X2 _396_ (.D(_127_),
    .CK(clknet_2_2__leaf_clk),
    .Q(sram_rdata_reg[5]),
    .QN(_260_));
 DFF_X2 _397_ (.D(_128_),
    .CK(clknet_2_2__leaf_clk),
    .Q(sram_rdata_reg[6]),
    .QN(_261_));
 DFF_X2 _398_ (.D(_129_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\u_multiplier/LODy/z [7]),
    .QN(_262_));
 DFF_X1 _399_ (.D(_130_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net29),
    .QN(_263_));
 DFF_X2 _400_ (.D(_090_),
    .CK(clknet_2_1__leaf_clk),
    .Q(addr_ptr[0]),
    .QN(_264_));
 DFF_X1 _401_ (.D(_091_),
    .CK(clknet_2_1__leaf_clk),
    .Q(addr_ptr[1]),
    .QN(_265_));
 DFF_X1 _402_ (.D(_092_),
    .CK(clknet_2_1__leaf_clk),
    .Q(addr_ptr[2]),
    .QN(_266_));
 DFF_X1 _403_ (.D(net55),
    .CK(clknet_2_1__leaf_clk),
    .Q(addr_ptr[3]),
    .QN(_267_));
 DFF_X2 _404_ (.D(net62),
    .CK(clknet_2_1__leaf_clk),
    .Q(init_count[0]),
    .QN(_268_));
 DFF_X2 _405_ (.D(net80),
    .CK(clknet_2_1__leaf_clk),
    .Q(init_count[1]),
    .QN(_269_));
 DFF_X2 _406_ (.D(net73),
    .CK(clknet_2_1__leaf_clk),
    .Q(init_count[2]),
    .QN(_270_));
 DFF_X2 _407_ (.D(net77),
    .CK(clknet_2_1__leaf_clk),
    .Q(init_count[3]),
    .QN(_271_));
 SRAM_6T_CORE_16x8_MC_TB sram_inst (.ce_in(_134_),
    .we_in(_135_),
    .clk(clknet_2_0__leaf_clk),
    .addr_in({net68,
    net70,
    net66,
    net75}),
    .rd_out({sram_rdata[7],
    sram_rdata[6],
    sram_rdata[5],
    sram_rdata[4],
    sram_rdata[3],
    sram_rdata[2],
    sram_rdata[1],
    sram_rdata[0]}),
    .wd_in({net42,
    net59,
    net43,
    net44,
    net52,
    net51,
    net46,
    net45}));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_0/_09_  (.A1(\u_multiplier/LODx/z [1]),
    .A2(\u_multiplier/LODx/select [0]),
    .ZN(\u_multiplier/kx [1]));
 AND2_X1 \u_multiplier/LODx/Inst_MUX214_0/_10_  (.A1(\u_multiplier/LODx/select [0]),
    .A2(\u_multiplier/LODx/z [0]),
    .ZN(\u_multiplier/kx [0]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_0/_11_  (.A1(\u_multiplier/LODx/select [0]),
    .A2(\u_multiplier/LODx/z [3]),
    .ZN(\u_multiplier/kx [3]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_0/_12_  (.A1(\u_multiplier/LODx/select [0]),
    .A2(\u_multiplier/LODx/z [2]),
    .ZN(\u_multiplier/kx [2]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_1/_09_  (.A1(\u_multiplier/LODx/z [5]),
    .A2(\u_multiplier/LODx/select [1]),
    .ZN(\u_multiplier/kx [5]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_1/_10_  (.A1(\u_multiplier/LODx/select [1]),
    .A2(\u_multiplier/LODx/z [4]),
    .ZN(\u_multiplier/kx [4]));
 AND2_X1 \u_multiplier/LODx/Inst_MUX214_1/_11_  (.A1(\u_multiplier/LODx/select [1]),
    .A2(\u_multiplier/LODx/z [7]),
    .ZN(\u_multiplier/kx [7]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_1/_12_  (.A1(\u_multiplier/LODx/select [1]),
    .A2(\u_multiplier/LODx/z [6]),
    .ZN(\u_multiplier/kx [6]));
 INV_X1 \u_multiplier/LODx/Middle/_4_  (.A(\u_multiplier/LODx/_12_ ),
    .ZN(\u_multiplier/LODx/Middle/_3_ ));
 NOR2_X1 \u_multiplier/LODx/Middle/_5_  (.A1(\u_multiplier/LODx/Middle/_3_ ),
    .A2(\u_multiplier/LODx/select [1]),
    .ZN(\u_multiplier/LODx/select [0]));
 OR4_X1 \u_multiplier/LODx/_15_  (.A1(data_in_reg[2]),
    .A2(\u_multiplier/LODx/z [3]),
    .A3(data_in_reg[0]),
    .A4(data_in_reg[1]),
    .ZN(\u_multiplier/LODx/_12_ ));
 OR4_X2 \u_multiplier/LODx/_16_  (.A1(data_in_reg[6]),
    .A2(\u_multiplier/LODx/z [7]),
    .A3(data_in_reg[4]),
    .A4(data_in_reg[5]),
    .ZN(\u_multiplier/LODx/select [1]));
 NOR2_X2 \u_multiplier/LODx/_17_  (.A1(\u_multiplier/LODx/_12_ ),
    .A2(\u_multiplier/LODx/select [1]),
    .ZN(\u_multiplier/zero_x ));
 INV_X1 \u_multiplier/LODx/lod2_0/_12_  (.A(data_in_reg[2]),
    .ZN(\u_multiplier/LODx/lod2_0/_10_ ));
 INV_X1 \u_multiplier/LODx/lod2_0/_13_  (.A(data_in_reg[1]),
    .ZN(\u_multiplier/LODx/lod2_0/_11_ ));
 INV_X1 \u_multiplier/LODx/lod2_0/_14_  (.A(data_in_reg[0]),
    .ZN(\u_multiplier/LODx/lod2_0/_09_ ));
 NOR2_X1 \u_multiplier/LODx/lod2_0/_15_  (.A1(\u_multiplier/LODx/lod2_0/_10_ ),
    .A2(\u_multiplier/LODx/z [3]),
    .ZN(\u_multiplier/LODx/z [2]));
 NOR3_X1 \u_multiplier/LODx/lod2_0/_16_  (.A1(data_in_reg[2]),
    .A2(\u_multiplier/LODx/z [3]),
    .A3(\u_multiplier/LODx/lod2_0/_11_ ),
    .ZN(\u_multiplier/LODx/z [1]));
 NOR4_X1 \u_multiplier/LODx/lod2_0/_17_  (.A1(data_in_reg[2]),
    .A2(\u_multiplier/LODx/z [3]),
    .A3(data_in_reg[1]),
    .A4(\u_multiplier/LODx/lod2_0/_09_ ),
    .ZN(\u_multiplier/LODx/z [0]));
 INV_X1 \u_multiplier/LODx/lod2_1/_12_  (.A(data_in_reg[6]),
    .ZN(\u_multiplier/LODx/lod2_1/_10_ ));
 INV_X1 \u_multiplier/LODx/lod2_1/_13_  (.A(data_in_reg[5]),
    .ZN(\u_multiplier/LODx/lod2_1/_11_ ));
 INV_X1 \u_multiplier/LODx/lod2_1/_14_  (.A(data_in_reg[4]),
    .ZN(\u_multiplier/LODx/lod2_1/_09_ ));
 NOR2_X1 \u_multiplier/LODx/lod2_1/_15_  (.A1(\u_multiplier/LODx/lod2_1/_10_ ),
    .A2(\u_multiplier/LODx/z [7]),
    .ZN(\u_multiplier/LODx/z [6]));
 NOR3_X1 \u_multiplier/LODx/lod2_1/_16_  (.A1(data_in_reg[6]),
    .A2(\u_multiplier/LODx/z [7]),
    .A3(\u_multiplier/LODx/lod2_1/_11_ ),
    .ZN(\u_multiplier/LODx/z [5]));
 NOR4_X1 \u_multiplier/LODx/lod2_1/_17_  (.A1(data_in_reg[6]),
    .A2(\u_multiplier/LODx/z [7]),
    .A3(data_in_reg[5]),
    .A4(\u_multiplier/LODx/lod2_1/_09_ ),
    .ZN(\u_multiplier/LODx/z [4]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_0/_09_  (.A1(\u_multiplier/LODy/z [1]),
    .A2(\u_multiplier/LODy/select [0]),
    .ZN(\u_multiplier/ky [1]));
 AND2_X1 \u_multiplier/LODy/Inst_MUX214_0/_10_  (.A1(\u_multiplier/LODy/select [0]),
    .A2(\u_multiplier/LODy/z [0]),
    .ZN(\u_multiplier/ky [0]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_0/_11_  (.A1(\u_multiplier/LODy/select [0]),
    .A2(\u_multiplier/LODy/z [3]),
    .ZN(\u_multiplier/ky [3]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_0/_12_  (.A1(\u_multiplier/LODy/select [0]),
    .A2(\u_multiplier/LODy/z [2]),
    .ZN(\u_multiplier/ky [2]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_1/_09_  (.A1(\u_multiplier/LODy/z [5]),
    .A2(\u_multiplier/LODy/select [1]),
    .ZN(\u_multiplier/ky [5]));
 AND2_X1 \u_multiplier/LODy/Inst_MUX214_1/_10_  (.A1(\u_multiplier/LODy/select [1]),
    .A2(\u_multiplier/LODy/z [4]),
    .ZN(\u_multiplier/ky [4]));
 AND2_X1 \u_multiplier/LODy/Inst_MUX214_1/_11_  (.A1(\u_multiplier/LODy/select [1]),
    .A2(\u_multiplier/LODy/z [7]),
    .ZN(\u_multiplier/ky [7]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_1/_12_  (.A1(\u_multiplier/LODy/select [1]),
    .A2(\u_multiplier/LODy/z [6]),
    .ZN(\u_multiplier/ky [6]));
 INV_X1 \u_multiplier/LODy/Middle/_4_  (.A(\u_multiplier/LODy/_12_ ),
    .ZN(\u_multiplier/LODy/Middle/_3_ ));
 NOR2_X1 \u_multiplier/LODy/Middle/_5_  (.A1(\u_multiplier/LODy/Middle/_3_ ),
    .A2(\u_multiplier/LODy/select [1]),
    .ZN(\u_multiplier/LODy/select [0]));
 OR4_X1 \u_multiplier/LODy/_15_  (.A1(sram_rdata_reg[2]),
    .A2(\u_multiplier/LODy/z [3]),
    .A3(sram_rdata_reg[0]),
    .A4(sram_rdata_reg[1]),
    .ZN(\u_multiplier/LODy/_12_ ));
 OR4_X2 \u_multiplier/LODy/_16_  (.A1(sram_rdata_reg[6]),
    .A2(\u_multiplier/LODy/z [7]),
    .A3(sram_rdata_reg[4]),
    .A4(sram_rdata_reg[5]),
    .ZN(\u_multiplier/LODy/select [1]));
 NOR2_X2 \u_multiplier/LODy/_17_  (.A1(\u_multiplier/LODy/_12_ ),
    .A2(\u_multiplier/LODy/select [1]),
    .ZN(\u_multiplier/zero_y ));
 INV_X1 \u_multiplier/LODy/lod2_0/_12_  (.A(sram_rdata_reg[2]),
    .ZN(\u_multiplier/LODy/lod2_0/_10_ ));
 INV_X1 \u_multiplier/LODy/lod2_0/_13_  (.A(sram_rdata_reg[1]),
    .ZN(\u_multiplier/LODy/lod2_0/_11_ ));
 INV_X1 \u_multiplier/LODy/lod2_0/_14_  (.A(sram_rdata_reg[0]),
    .ZN(\u_multiplier/LODy/lod2_0/_09_ ));
 NOR2_X1 \u_multiplier/LODy/lod2_0/_15_  (.A1(\u_multiplier/LODy/lod2_0/_10_ ),
    .A2(\u_multiplier/LODy/z [3]),
    .ZN(\u_multiplier/LODy/z [2]));
 NOR3_X1 \u_multiplier/LODy/lod2_0/_16_  (.A1(sram_rdata_reg[2]),
    .A2(\u_multiplier/LODy/z [3]),
    .A3(\u_multiplier/LODy/lod2_0/_11_ ),
    .ZN(\u_multiplier/LODy/z [1]));
 NOR4_X1 \u_multiplier/LODy/lod2_0/_17_  (.A1(sram_rdata_reg[2]),
    .A2(\u_multiplier/LODy/z [3]),
    .A3(sram_rdata_reg[1]),
    .A4(\u_multiplier/LODy/lod2_0/_09_ ),
    .ZN(\u_multiplier/LODy/z [0]));
 INV_X1 \u_multiplier/LODy/lod2_1/_12_  (.A(sram_rdata_reg[6]),
    .ZN(\u_multiplier/LODy/lod2_1/_10_ ));
 INV_X1 \u_multiplier/LODy/lod2_1/_13_  (.A(sram_rdata_reg[5]),
    .ZN(\u_multiplier/LODy/lod2_1/_11_ ));
 INV_X1 \u_multiplier/LODy/lod2_1/_14_  (.A(sram_rdata_reg[4]),
    .ZN(\u_multiplier/LODy/lod2_1/_09_ ));
 NOR2_X1 \u_multiplier/LODy/lod2_1/_15_  (.A1(\u_multiplier/LODy/lod2_1/_10_ ),
    .A2(\u_multiplier/LODy/z [7]),
    .ZN(\u_multiplier/LODy/z [6]));
 NOR3_X1 \u_multiplier/LODy/lod2_1/_16_  (.A1(sram_rdata_reg[6]),
    .A2(\u_multiplier/LODy/z [7]),
    .A3(\u_multiplier/LODy/lod2_1/_11_ ),
    .ZN(\u_multiplier/LODy/z [5]));
 NOR4_X1 \u_multiplier/LODy/lod2_1/_17_  (.A1(sram_rdata_reg[6]),
    .A2(\u_multiplier/LODy/z [7]),
    .A3(sram_rdata_reg[5]),
    .A4(\u_multiplier/LODy/lod2_1/_09_ ),
    .ZN(\u_multiplier/LODy/z [4]));
 INV_X1 \u_multiplier/NOD/_15_  (.A(\u_multiplier/NOD/t_in [1]),
    .ZN(\u_multiplier/NOD/_11_ ));
 INV_X1 \u_multiplier/NOD/_16_  (.A(\u_multiplier/_0346_ ),
    .ZN(\u_multiplier/NOD/_12_ ));
 INV_X1 \u_multiplier/NOD/_17_  (.A(\u_multiplier/_0345_ ),
    .ZN(\u_multiplier/NOD/_13_ ));
 AND2_X1 \u_multiplier/NOD/_18_  (.A1(\u_multiplier/_0350_ ),
    .A2(\u_multiplier/_0351_ ),
    .ZN(\u_multiplier/NOD_Q1 [7]));
 NOR4_X2 \u_multiplier/NOD/_19_  (.A1(\u_multiplier/_0347_ ),
    .A2(\u_multiplier/NOD/_11_ ),
    .A3(\u_multiplier/NOD/_12_ ),
    .A4(\u_multiplier/_0345_ ),
    .ZN(\u_multiplier/NOD_Q1 [1]));
 NOR4_X1 \u_multiplier/NOD/_20_  (.A1(\u_multiplier/_0347_ ),
    .A2(\u_multiplier/NOD/_11_ ),
    .A3(\u_multiplier/_0346_ ),
    .A4(\u_multiplier/NOD/_13_ ),
    .ZN(\u_multiplier/NOD_Q1 [0]));
 AOI21_X1 \u_multiplier/NOD/nod_basic_unit15/_7_  (.A(\u_multiplier/_0351_ ),
    .B1(\u_multiplier/_0349_ ),
    .B2(\u_multiplier/_0350_ ),
    .ZN(\u_multiplier/NOD/nod_basic_unit15/_5_ ));
 AOI21_X2 \u_multiplier/NOD/nod_basic_unit15/_8_  (.A(\u_multiplier/NOD/nod_basic_unit15/_5_ ),
    .B1(\u_multiplier/_0351_ ),
    .B2(\u_multiplier/_0350_ ),
    .ZN(\u_multiplier/NOD_Q1 [6]));
 INV_X1 \u_multiplier/NOD/nod_cels[2].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [2]),
    .ZN(\u_multiplier/NOD/nod_cels[2].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[2].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[2].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[2].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[2].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[2].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0348_ ),
    .ZN(\u_multiplier/NOD/t_in [1]));
 NOR3_X1 \u_multiplier/NOD/nod_cels[2].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[2].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0348_ ),
    .A3(\u_multiplier/NOD/nod_cels[2].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [2]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[2].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_0347_ ),
    .B1(\u_multiplier/_0345_ ),
    .B2(\u_multiplier/_0346_ ),
    .ZN(\u_multiplier/NOD/nod_cels[2].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[2].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[2].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_0347_ ),
    .B2(\u_multiplier/_0346_ ),
    .ZN(\u_multiplier/NOD/nod_cels[2].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[3].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [3]),
    .ZN(\u_multiplier/NOD/nod_cels[3].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[3].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[3].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[3].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[3].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[3].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0349_ ),
    .ZN(\u_multiplier/NOD/t_in [2]));
 NOR3_X2 \u_multiplier/NOD/nod_cels[3].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[3].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0349_ ),
    .A3(\u_multiplier/NOD/nod_cels[3].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [3]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[3].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_0348_ ),
    .B1(\u_multiplier/_0346_ ),
    .B2(\u_multiplier/_0347_ ),
    .ZN(\u_multiplier/NOD/nod_cels[3].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[3].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[3].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_0348_ ),
    .B2(\u_multiplier/_0347_ ),
    .ZN(\u_multiplier/NOD/nod_cels[3].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[4].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [4]),
    .ZN(\u_multiplier/NOD/nod_cels[4].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[4].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[4].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[4].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[4].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[4].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0350_ ),
    .ZN(\u_multiplier/NOD/t_in [3]));
 NOR3_X1 \u_multiplier/NOD/nod_cels[4].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[4].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0350_ ),
    .A3(\u_multiplier/NOD/nod_cels[4].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [4]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[4].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_0349_ ),
    .B1(\u_multiplier/_0347_ ),
    .B2(\u_multiplier/_0348_ ),
    .ZN(\u_multiplier/NOD/nod_cels[4].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[4].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[4].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_0349_ ),
    .B2(\u_multiplier/_0348_ ),
    .ZN(\u_multiplier/NOD/nod_cels[4].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[5].Nod_bits/_07_  (.A(net30),
    .ZN(\u_multiplier/NOD/nod_cels[5].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[5].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[5].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[5].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[5].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[5].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0351_ ),
    .ZN(\u_multiplier/NOD/t_in [4]));
 NOR3_X2 \u_multiplier/NOD/nod_cels[5].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[5].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0351_ ),
    .A3(\u_multiplier/NOD/nod_cels[5].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [5]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[5].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_0350_ ),
    .B1(\u_multiplier/_0348_ ),
    .B2(\u_multiplier/_0349_ ),
    .ZN(\u_multiplier/NOD/nod_cels[5].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[5].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[5].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_0350_ ),
    .B2(\u_multiplier/_0349_ ),
    .ZN(\u_multiplier/NOD/nod_cels[5].Nod_bits/tmp1 ));
 OR4_X4 \u_multiplier/PE/code0/_7_  (.A1(\u_multiplier/NOD_Q1 [5]),
    .A2(\u_multiplier/NOD_Q1 [1]),
    .A3(\u_multiplier/NOD_Q1 [7]),
    .A4(\u_multiplier/NOD_Q1 [3]),
    .ZN(\u_multiplier/K [0]));
 OR4_X4 \u_multiplier/PE/code1/_7_  (.A1(\u_multiplier/NOD_Q1 [6]),
    .A2(\u_multiplier/NOD_Q1 [2]),
    .A3(\u_multiplier/NOD_Q1 [7]),
    .A4(\u_multiplier/NOD_Q1 [3]),
    .ZN(\u_multiplier/K [1]));
 OR4_X4 \u_multiplier/PE/code2/_7_  (.A1(\u_multiplier/NOD_Q1 [6]),
    .A2(\u_multiplier/NOD_Q1 [4]),
    .A3(\u_multiplier/NOD_Q1 [7]),
    .A4(\u_multiplier/NOD_Q1 [5]),
    .ZN(\u_multiplier/K [2]));
 OR4_X4 \u_multiplier/PEx/code0/_7_  (.A1(\u_multiplier/kx [5]),
    .A2(\u_multiplier/kx [1]),
    .A3(\u_multiplier/kx [7]),
    .A4(\u_multiplier/kx [3]),
    .ZN(\u_multiplier/code_x [0]));
 OR4_X4 \u_multiplier/PEx/code1/_7_  (.A1(\u_multiplier/kx [6]),
    .A2(\u_multiplier/kx [2]),
    .A3(\u_multiplier/kx [7]),
    .A4(\u_multiplier/kx [3]),
    .ZN(\u_multiplier/code_x [1]));
 OR4_X4 \u_multiplier/PEx/code2/_7_  (.A1(\u_multiplier/kx [6]),
    .A2(\u_multiplier/kx [4]),
    .A3(\u_multiplier/kx [7]),
    .A4(\u_multiplier/kx [5]),
    .ZN(\u_multiplier/code_x [2]));
 OR4_X4 \u_multiplier/PEy/code0/_7_  (.A1(\u_multiplier/ky [5]),
    .A2(\u_multiplier/ky [1]),
    .A3(\u_multiplier/ky [7]),
    .A4(\u_multiplier/ky [3]),
    .ZN(\u_multiplier/code_y [0]));
 OR4_X4 \u_multiplier/PEy/code1/_7_  (.A1(\u_multiplier/ky [6]),
    .A2(\u_multiplier/ky [2]),
    .A3(\u_multiplier/ky [7]),
    .A4(\u_multiplier/ky [3]),
    .ZN(\u_multiplier/code_y [1]));
 OR4_X4 \u_multiplier/PEy/code2/_7_  (.A1(\u_multiplier/ky [6]),
    .A2(\u_multiplier/ky [4]),
    .A3(\u_multiplier/ky [7]),
    .A4(\u_multiplier/ky [5]),
    .ZN(\u_multiplier/code_y [2]));
 INV_X1 \u_multiplier/_0756_  (.A(\u_multiplier/code_y [2]),
    .ZN(\u_multiplier/_0707_ ));
 INV_X1 \u_multiplier/_0757_  (.A(\u_multiplier/code_x [2]),
    .ZN(\u_multiplier/_0708_ ));
 INV_X2 \u_multiplier/_0758_  (.A(\u_multiplier/K [0]),
    .ZN(\u_multiplier/_0709_ ));
 INV_X2 \u_multiplier/_0759_  (.A(\u_multiplier/K [1]),
    .ZN(\u_multiplier/_0710_ ));
 INV_X4 \u_multiplier/_0760_  (.A(\u_multiplier/K [2]),
    .ZN(\u_multiplier/_0711_ ));
 INV_X1 \u_multiplier/_0761_  (.A(\u_multiplier/dec_out [12]),
    .ZN(\u_multiplier/_0712_ ));
 INV_X1 \u_multiplier/_0762_  (.A(\u_multiplier/dec_out [15]),
    .ZN(\u_multiplier/_0713_ ));
 XNOR2_X2 \u_multiplier/_0763_  (.A(\u_multiplier/ky [0]),
    .B(sram_rdata_reg[0]),
    .ZN(\u_multiplier/_0714_ ));
 XOR2_X2 \u_multiplier/_0764_  (.A(\u_multiplier/ky [0]),
    .B(sram_rdata_reg[0]),
    .Z(\u_multiplier/_0715_ ));
 XOR2_X2 \u_multiplier/_0765_  (.A(\u_multiplier/kx [6]),
    .B(data_in_reg[6]),
    .Z(\u_multiplier/_0716_ ));
 XNOR2_X2 \u_multiplier/_0766_  (.A(\u_multiplier/kx [6]),
    .B(data_in_reg[6]),
    .ZN(\u_multiplier/_0717_ ));
 XOR2_X2 \u_multiplier/_0767_  (.A(\u_multiplier/ky [6]),
    .B(sram_rdata_reg[6]),
    .Z(\u_multiplier/_0718_ ));
 XNOR2_X2 \u_multiplier/_0768_  (.A(\u_multiplier/ky [6]),
    .B(sram_rdata_reg[6]),
    .ZN(\u_multiplier/_0719_ ));
 NOR2_X2 \u_multiplier/_0769_  (.A1(\u_multiplier/_0716_ ),
    .A2(\u_multiplier/_0719_ ),
    .ZN(\u_multiplier/_0720_ ));
 XOR2_X2 \u_multiplier/_0770_  (.A(\u_multiplier/ky [1]),
    .B(sram_rdata_reg[1]),
    .Z(\u_multiplier/_0721_ ));
 XNOR2_X2 \u_multiplier/_0771_  (.A(\u_multiplier/ky [1]),
    .B(sram_rdata_reg[1]),
    .ZN(\u_multiplier/_0722_ ));
 XNOR2_X2 \u_multiplier/_0772_  (.A(\u_multiplier/kx [1]),
    .B(data_in_reg[1]),
    .ZN(\u_multiplier/_0723_ ));
 XOR2_X2 \u_multiplier/_0773_  (.A(\u_multiplier/kx [1]),
    .B(data_in_reg[1]),
    .Z(\u_multiplier/_0392_ ));
 XNOR2_X2 \u_multiplier/_0774_  (.A(\u_multiplier/kx [0]),
    .B(data_in_reg[0]),
    .ZN(\u_multiplier/_0393_ ));
 XOR2_X2 \u_multiplier/_0775_  (.A(\u_multiplier/kx [0]),
    .B(data_in_reg[0]),
    .Z(\u_multiplier/_0394_ ));
 AOI211_X1 \u_multiplier/_0776_  (.A(\u_multiplier/_0715_ ),
    .B(\u_multiplier/_0393_ ),
    .C1(\u_multiplier/_0723_ ),
    .C2(\u_multiplier/_0721_ ),
    .ZN(\u_multiplier/_0395_ ));
 OAI211_X1 \u_multiplier/_0777_  (.A(\u_multiplier/_0714_ ),
    .B(\u_multiplier/_0394_ ),
    .C1(\u_multiplier/_0392_ ),
    .C2(\u_multiplier/_0722_ ),
    .ZN(\u_multiplier/_0396_ ));
 XOR2_X2 \u_multiplier/_0778_  (.A(\u_multiplier/ky [2]),
    .B(sram_rdata_reg[2]),
    .Z(\u_multiplier/_0397_ ));
 XNOR2_X2 \u_multiplier/_0779_  (.A(\u_multiplier/ky [2]),
    .B(sram_rdata_reg[2]),
    .ZN(\u_multiplier/_0398_ ));
 XNOR2_X2 \u_multiplier/_0780_  (.A(\u_multiplier/kx [2]),
    .B(data_in_reg[2]),
    .ZN(\u_multiplier/_0399_ ));
 XOR2_X2 \u_multiplier/_0781_  (.A(\u_multiplier/kx [2]),
    .B(data_in_reg[2]),
    .Z(\u_multiplier/_0400_ ));
 AOI22_X1 \u_multiplier/_0782_  (.A1(\u_multiplier/_0722_ ),
    .A2(\u_multiplier/_0392_ ),
    .B1(\u_multiplier/_0398_ ),
    .B2(\u_multiplier/_0400_ ),
    .ZN(\u_multiplier/_0401_ ));
 OAI22_X1 \u_multiplier/_0783_  (.A1(\u_multiplier/_0721_ ),
    .A2(\u_multiplier/_0723_ ),
    .B1(\u_multiplier/_0397_ ),
    .B2(\u_multiplier/_0399_ ),
    .ZN(\u_multiplier/_0402_ ));
 XOR2_X2 \u_multiplier/_0784_  (.A(\u_multiplier/ky [3]),
    .B(\u_multiplier/LODy/z [3]),
    .Z(\u_multiplier/_0403_ ));
 XNOR2_X2 \u_multiplier/_0785_  (.A(\u_multiplier/kx [3]),
    .B(\u_multiplier/LODx/z [3]),
    .ZN(\u_multiplier/_0404_ ));
 XOR2_X2 \u_multiplier/_0786_  (.A(\u_multiplier/kx [3]),
    .B(\u_multiplier/LODx/z [3]),
    .Z(\u_multiplier/_0405_ ));
 AOI22_X1 \u_multiplier/_0787_  (.A1(\u_multiplier/_0397_ ),
    .A2(\u_multiplier/_0399_ ),
    .B1(\u_multiplier/_0403_ ),
    .B2(\u_multiplier/_0404_ ),
    .ZN(\u_multiplier/_0406_ ));
 AOI222_X2 \u_multiplier/_0788_  (.A1(\u_multiplier/_0397_ ),
    .A2(\u_multiplier/_0399_ ),
    .B1(\u_multiplier/_0403_ ),
    .B2(\u_multiplier/_0404_ ),
    .C1(\u_multiplier/_0401_ ),
    .C2(\u_multiplier/_0396_ ),
    .ZN(\u_multiplier/_0407_ ));
 OAI21_X1 \u_multiplier/_0789_  (.A(\u_multiplier/_0406_ ),
    .B1(\u_multiplier/_0402_ ),
    .B2(\u_multiplier/_0395_ ),
    .ZN(\u_multiplier/_0408_ ));
 XOR2_X2 \u_multiplier/_0790_  (.A(\u_multiplier/ky [4]),
    .B(sram_rdata_reg[4]),
    .Z(\u_multiplier/_0409_ ));
 XNOR2_X2 \u_multiplier/_0791_  (.A(\u_multiplier/kx [4]),
    .B(data_in_reg[4]),
    .ZN(\u_multiplier/_0410_ ));
 XOR2_X2 \u_multiplier/_0792_  (.A(\u_multiplier/kx [4]),
    .B(data_in_reg[4]),
    .Z(\u_multiplier/_0411_ ));
 OAI22_X2 \u_multiplier/_0793_  (.A1(\u_multiplier/_0403_ ),
    .A2(\u_multiplier/_0404_ ),
    .B1(\u_multiplier/_0409_ ),
    .B2(\u_multiplier/_0410_ ),
    .ZN(\u_multiplier/_0412_ ));
 INV_X1 \u_multiplier/_0794_  (.A(\u_multiplier/_0412_ ),
    .ZN(\u_multiplier/_0413_ ));
 XOR2_X2 \u_multiplier/_0795_  (.A(\u_multiplier/kx [5]),
    .B(data_in_reg[5]),
    .Z(\u_multiplier/_0414_ ));
 XNOR2_X2 \u_multiplier/_0796_  (.A(\u_multiplier/ky [5]),
    .B(sram_rdata_reg[5]),
    .ZN(\u_multiplier/_0415_ ));
 XOR2_X2 \u_multiplier/_0797_  (.A(\u_multiplier/ky [5]),
    .B(sram_rdata_reg[5]),
    .Z(\u_multiplier/_0416_ ));
 NOR2_X1 \u_multiplier/_0798_  (.A1(\u_multiplier/_0414_ ),
    .A2(\u_multiplier/_0415_ ),
    .ZN(\u_multiplier/_0417_ ));
 NAND2_X1 \u_multiplier/_0799_  (.A1(\u_multiplier/_0409_ ),
    .A2(\u_multiplier/_0410_ ),
    .ZN(\u_multiplier/_0418_ ));
 AOI221_X2 \u_multiplier/_0800_  (.A(\u_multiplier/_0417_ ),
    .B1(\u_multiplier/_0410_ ),
    .B2(\u_multiplier/_0409_ ),
    .C1(\u_multiplier/_0408_ ),
    .C2(\u_multiplier/_0413_ ),
    .ZN(\u_multiplier/_0419_ ));
 OAI221_X2 \u_multiplier/_0801_  (.A(\u_multiplier/_0418_ ),
    .B1(\u_multiplier/_0415_ ),
    .B2(\u_multiplier/_0414_ ),
    .C1(\u_multiplier/_0407_ ),
    .C2(\u_multiplier/_0412_ ),
    .ZN(\u_multiplier/_0420_ ));
 NAND2_X1 \u_multiplier/_0802_  (.A1(\u_multiplier/_0414_ ),
    .A2(\u_multiplier/_0415_ ),
    .ZN(\u_multiplier/_0421_ ));
 AOI22_X4 \u_multiplier/_0803_  (.A1(\u_multiplier/_0716_ ),
    .A2(\u_multiplier/_0719_ ),
    .B1(\u_multiplier/_0414_ ),
    .B2(\u_multiplier/_0415_ ),
    .ZN(\u_multiplier/_0422_ ));
 OAI21_X2 \u_multiplier/_0804_  (.A(\u_multiplier/_0421_ ),
    .B1(\u_multiplier/_0718_ ),
    .B2(\u_multiplier/_0717_ ),
    .ZN(\u_multiplier/_0423_ ));
 AOI21_X4 \u_multiplier/_0805_  (.A(\u_multiplier/_0720_ ),
    .B1(\u_multiplier/_0420_ ),
    .B2(\u_multiplier/_0422_ ),
    .ZN(\u_multiplier/_0424_ ));
 OAI22_X4 \u_multiplier/_0806_  (.A1(\u_multiplier/_0716_ ),
    .A2(\u_multiplier/_0719_ ),
    .B1(\u_multiplier/_0419_ ),
    .B2(\u_multiplier/_0423_ ),
    .ZN(\u_multiplier/_0425_ ));
 MUX2_X1 \u_multiplier/_0807_  (.A(\u_multiplier/_0715_ ),
    .B(\u_multiplier/_0394_ ),
    .S(\u_multiplier/_0424_ ),
    .Z(\u_multiplier/_0345_ ));
 MUX2_X2 \u_multiplier/_0808_  (.A(\u_multiplier/_0721_ ),
    .B(\u_multiplier/_0392_ ),
    .S(\u_multiplier/_0424_ ),
    .Z(\u_multiplier/_0346_ ));
 MUX2_X2 \u_multiplier/_0809_  (.A(\u_multiplier/_0397_ ),
    .B(\u_multiplier/_0400_ ),
    .S(\u_multiplier/_0424_ ),
    .Z(\u_multiplier/_0347_ ));
 MUX2_X2 \u_multiplier/_0810_  (.A(\u_multiplier/_0403_ ),
    .B(\u_multiplier/_0405_ ),
    .S(\u_multiplier/_0424_ ),
    .Z(\u_multiplier/_0348_ ));
 MUX2_X2 \u_multiplier/_0811_  (.A(\u_multiplier/_0409_ ),
    .B(\u_multiplier/_0411_ ),
    .S(\u_multiplier/_0424_ ),
    .Z(\u_multiplier/_0349_ ));
 MUX2_X2 \u_multiplier/_0812_  (.A(\u_multiplier/_0414_ ),
    .B(\u_multiplier/_0416_ ),
    .S(\u_multiplier/_0425_ ),
    .Z(\u_multiplier/_0350_ ));
 NAND2_X2 \u_multiplier/_0813_  (.A1(\u_multiplier/_0717_ ),
    .A2(\u_multiplier/_0719_ ),
    .ZN(\u_multiplier/_0351_ ));
 MUX2_X2 \u_multiplier/_0814_  (.A(\u_multiplier/_0714_ ),
    .B(\u_multiplier/_0393_ ),
    .S(\u_multiplier/_0425_ ),
    .Z(\u_multiplier/_0426_ ));
 NOR3_X1 \u_multiplier/_0815_  (.A1(\u_multiplier/K [0]),
    .A2(\u_multiplier/K [1]),
    .A3(\u_multiplier/_0426_ ),
    .ZN(\u_multiplier/_0427_ ));
 NOR4_X2 \u_multiplier/_0816_  (.A1(\u_multiplier/K [0]),
    .A2(\u_multiplier/K [1]),
    .A3(\u_multiplier/K [2]),
    .A4(\u_multiplier/_0426_ ),
    .ZN(\u_multiplier/_0428_ ));
 NOR2_X1 \u_multiplier/_0817_  (.A1(\u_multiplier/code_x [0]),
    .A2(\u_multiplier/_0714_ ),
    .ZN(\u_multiplier/_0429_ ));
 NOR3_X1 \u_multiplier/_0818_  (.A1(\u_multiplier/code_x [0]),
    .A2(\u_multiplier/code_x [1]),
    .A3(\u_multiplier/_0714_ ),
    .ZN(\u_multiplier/_0430_ ));
 AND2_X1 \u_multiplier/_0819_  (.A1(\u_multiplier/_0708_ ),
    .A2(\u_multiplier/_0430_ ),
    .ZN(\u_multiplier/_0431_ ));
 NOR2_X1 \u_multiplier/_0820_  (.A1(\u_multiplier/code_y [0]),
    .A2(\u_multiplier/_0393_ ),
    .ZN(\u_multiplier/_0432_ ));
 OR3_X1 \u_multiplier/_0821_  (.A1(\u_multiplier/code_y [0]),
    .A2(\u_multiplier/code_y [1]),
    .A3(\u_multiplier/_0393_ ),
    .ZN(\u_multiplier/_0433_ ));
 NOR2_X1 \u_multiplier/_0822_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_0433_ ),
    .ZN(\u_multiplier/_0434_ ));
 NAND2_X1 \u_multiplier/_0823_  (.A1(\u_multiplier/_0431_ ),
    .A2(\u_multiplier/_0434_ ),
    .ZN(\u_multiplier/_0435_ ));
 XOR2_X1 \u_multiplier/_0824_  (.A(\u_multiplier/_0431_ ),
    .B(\u_multiplier/_0434_ ),
    .Z(\u_multiplier/_0436_ ));
 OR3_X1 \u_multiplier/_0825_  (.A1(\u_multiplier/dec_out [0]),
    .A2(\u_multiplier/_0428_ ),
    .A3(\u_multiplier/_0436_ ),
    .ZN(\u_multiplier/_0437_ ));
 OAI21_X1 \u_multiplier/_0826_  (.A(\u_multiplier/_0436_ ),
    .B1(\u_multiplier/_0428_ ),
    .B2(\u_multiplier/dec_out [0]),
    .ZN(\u_multiplier/_0438_ ));
 NOR2_X4 \u_multiplier/_0827_  (.A1(\u_multiplier/zero_y ),
    .A2(\u_multiplier/zero_x ),
    .ZN(\u_multiplier/_0439_ ));
 OR2_X2 \u_multiplier/_0828_  (.A1(\u_multiplier/zero_y ),
    .A2(\u_multiplier/zero_x ),
    .ZN(\u_multiplier/_0440_ ));
 AND3_X1 \u_multiplier/_0829_  (.A1(\u_multiplier/_0437_ ),
    .A2(\u_multiplier/_0438_ ),
    .A3(\u_multiplier/_0439_ ),
    .ZN(product[0]));
 NAND2_X1 \u_multiplier/_0830_  (.A1(\u_multiplier/_0435_ ),
    .A2(\u_multiplier/_0438_ ),
    .ZN(\u_multiplier/_0441_ ));
 AOI211_X2 \u_multiplier/_0831_  (.A(\u_multiplier/_0720_ ),
    .B(\u_multiplier/_0722_ ),
    .C1(\u_multiplier/_0420_ ),
    .C2(\u_multiplier/_0422_ ),
    .ZN(\u_multiplier/_0442_ ));
 AOI211_X2 \u_multiplier/_0832_  (.A(\u_multiplier/K [0]),
    .B(\u_multiplier/_0442_ ),
    .C1(\u_multiplier/_0425_ ),
    .C2(\u_multiplier/_0392_ ),
    .ZN(\u_multiplier/_0443_ ));
 AOI21_X1 \u_multiplier/_0833_  (.A(\u_multiplier/_0443_ ),
    .B1(\u_multiplier/_0426_ ),
    .B2(\u_multiplier/K [0]),
    .ZN(\u_multiplier/_0444_ ));
 AOI211_X2 \u_multiplier/_0834_  (.A(\u_multiplier/K [1]),
    .B(\u_multiplier/_0443_ ),
    .C1(\u_multiplier/_0426_ ),
    .C2(\u_multiplier/K [0]),
    .ZN(\u_multiplier/_0445_ ));
 AOI21_X4 \u_multiplier/_0835_  (.A(\u_multiplier/dec_out [1]),
    .B1(\u_multiplier/_0445_ ),
    .B2(\u_multiplier/_0711_ ),
    .ZN(\u_multiplier/_0446_ ));
 MUX2_X1 \u_multiplier/_0836_  (.A(\u_multiplier/_0722_ ),
    .B(\u_multiplier/_0714_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_0447_ ));
 OR2_X1 \u_multiplier/_0837_  (.A1(\u_multiplier/code_x [1]),
    .A2(\u_multiplier/_0447_ ),
    .ZN(\u_multiplier/_0448_ ));
 MUX2_X1 \u_multiplier/_0838_  (.A(\u_multiplier/_0723_ ),
    .B(\u_multiplier/_0393_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_0449_ ));
 OR2_X1 \u_multiplier/_0839_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_0449_ ),
    .ZN(\u_multiplier/_0450_ ));
 OAI22_X1 \u_multiplier/_0840_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_0448_ ),
    .B1(\u_multiplier/_0450_ ),
    .B2(\u_multiplier/code_y [2]),
    .ZN(\u_multiplier/_0451_ ));
 OR4_X1 \u_multiplier/_0841_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/code_x [2]),
    .A3(\u_multiplier/_0448_ ),
    .A4(\u_multiplier/_0450_ ),
    .ZN(\u_multiplier/_0452_ ));
 NAND2_X1 \u_multiplier/_0842_  (.A1(\u_multiplier/_0451_ ),
    .A2(\u_multiplier/_0452_ ),
    .ZN(\u_multiplier/_0453_ ));
 XOR2_X2 \u_multiplier/_0843_  (.A(\u_multiplier/_0446_ ),
    .B(\u_multiplier/_0453_ ),
    .Z(\u_multiplier/_0454_ ));
 NAND2_X2 \u_multiplier/_0844_  (.A1(\u_multiplier/_0441_ ),
    .A2(\u_multiplier/_0454_ ),
    .ZN(\u_multiplier/_0455_ ));
 OAI21_X1 \u_multiplier/_0845_  (.A(\u_multiplier/_0439_ ),
    .B1(\u_multiplier/_0441_ ),
    .B2(\u_multiplier/_0454_ ),
    .ZN(\u_multiplier/_0456_ ));
 AOI21_X1 \u_multiplier/_0846_  (.A(\u_multiplier/_0456_ ),
    .B1(\u_multiplier/_0454_ ),
    .B2(\u_multiplier/_0441_ ),
    .ZN(product[1]));
 OAI21_X2 \u_multiplier/_0847_  (.A(\u_multiplier/_0452_ ),
    .B1(\u_multiplier/_0453_ ),
    .B2(\u_multiplier/_0446_ ),
    .ZN(\u_multiplier/_0457_ ));
 AOI211_X2 \u_multiplier/_0848_  (.A(\u_multiplier/_0720_ ),
    .B(\u_multiplier/_0398_ ),
    .C1(\u_multiplier/_0420_ ),
    .C2(\u_multiplier/_0422_ ),
    .ZN(\u_multiplier/_0458_ ));
 MUX2_X1 \u_multiplier/_0849_  (.A(\u_multiplier/_0397_ ),
    .B(\u_multiplier/_0400_ ),
    .S(\u_multiplier/_0425_ ),
    .Z(\u_multiplier/_0459_ ));
 AOI211_X2 \u_multiplier/_0850_  (.A(\u_multiplier/_0709_ ),
    .B(\u_multiplier/_0442_ ),
    .C1(\u_multiplier/_0425_ ),
    .C2(\u_multiplier/_0392_ ),
    .ZN(\u_multiplier/_0460_ ));
 AOI211_X2 \u_multiplier/_0851_  (.A(\u_multiplier/K [0]),
    .B(\u_multiplier/_0458_ ),
    .C1(\u_multiplier/_0425_ ),
    .C2(\u_multiplier/_0400_ ),
    .ZN(\u_multiplier/_0461_ ));
 OAI21_X1 \u_multiplier/_0852_  (.A(\u_multiplier/K [1]),
    .B1(\u_multiplier/_0426_ ),
    .B2(\u_multiplier/K [0]),
    .ZN(\u_multiplier/_0462_ ));
 OAI21_X1 \u_multiplier/_0853_  (.A(\u_multiplier/_0710_ ),
    .B1(\u_multiplier/_0460_ ),
    .B2(\u_multiplier/_0461_ ),
    .ZN(\u_multiplier/_0463_ ));
 AND3_X1 \u_multiplier/_0854_  (.A1(\u_multiplier/_0711_ ),
    .A2(\u_multiplier/_0462_ ),
    .A3(\u_multiplier/_0463_ ),
    .ZN(\u_multiplier/_0464_ ));
 MUX2_X1 \u_multiplier/_0855_  (.A(\u_multiplier/_0398_ ),
    .B(\u_multiplier/_0722_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_0465_ ));
 NOR2_X1 \u_multiplier/_0856_  (.A1(\u_multiplier/code_x [1]),
    .A2(\u_multiplier/_0465_ ),
    .ZN(\u_multiplier/_0466_ ));
 AOI21_X2 \u_multiplier/_0857_  (.A(\u_multiplier/_0466_ ),
    .B1(\u_multiplier/_0429_ ),
    .B2(\u_multiplier/code_x [1]),
    .ZN(\u_multiplier/_0467_ ));
 NOR2_X1 \u_multiplier/_0858_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_0467_ ),
    .ZN(\u_multiplier/_0468_ ));
 MUX2_X1 \u_multiplier/_0859_  (.A(\u_multiplier/_0399_ ),
    .B(\u_multiplier/_0723_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_0469_ ));
 NOR2_X1 \u_multiplier/_0860_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_0469_ ),
    .ZN(\u_multiplier/_0470_ ));
 AOI21_X2 \u_multiplier/_0861_  (.A(\u_multiplier/_0470_ ),
    .B1(\u_multiplier/_0432_ ),
    .B2(\u_multiplier/code_y [1]),
    .ZN(\u_multiplier/_0471_ ));
 NOR2_X1 \u_multiplier/_0862_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_0471_ ),
    .ZN(\u_multiplier/_0472_ ));
 NAND2_X1 \u_multiplier/_0863_  (.A1(\u_multiplier/_0468_ ),
    .A2(\u_multiplier/_0472_ ),
    .ZN(\u_multiplier/_0473_ ));
 XOR2_X2 \u_multiplier/_0864_  (.A(\u_multiplier/_0468_ ),
    .B(\u_multiplier/_0472_ ),
    .Z(\u_multiplier/_0474_ ));
 OAI21_X2 \u_multiplier/_0865_  (.A(\u_multiplier/_0474_ ),
    .B1(\u_multiplier/_0464_ ),
    .B2(\u_multiplier/dec_out [2]),
    .ZN(\u_multiplier/_0475_ ));
 OR3_X1 \u_multiplier/_0866_  (.A1(\u_multiplier/dec_out [2]),
    .A2(\u_multiplier/_0464_ ),
    .A3(\u_multiplier/_0474_ ),
    .ZN(\u_multiplier/_0476_ ));
 AND2_X1 \u_multiplier/_0867_  (.A1(\u_multiplier/_0475_ ),
    .A2(\u_multiplier/_0476_ ),
    .ZN(\u_multiplier/_0477_ ));
 NAND3_X1 \u_multiplier/_0868_  (.A1(\u_multiplier/_0457_ ),
    .A2(\u_multiplier/_0475_ ),
    .A3(\u_multiplier/_0476_ ),
    .ZN(\u_multiplier/_0478_ ));
 AOI21_X1 \u_multiplier/_0869_  (.A(\u_multiplier/_0457_ ),
    .B1(\u_multiplier/_0475_ ),
    .B2(\u_multiplier/_0476_ ),
    .ZN(\u_multiplier/_0479_ ));
 XNOR2_X1 \u_multiplier/_0870_  (.A(\u_multiplier/_0457_ ),
    .B(\u_multiplier/_0477_ ),
    .ZN(\u_multiplier/_0480_ ));
 OAI21_X1 \u_multiplier/_0871_  (.A(\u_multiplier/_0439_ ),
    .B1(\u_multiplier/_0455_ ),
    .B2(\u_multiplier/_0480_ ),
    .ZN(\u_multiplier/_0481_ ));
 AOI21_X2 \u_multiplier/_0872_  (.A(\u_multiplier/_0481_ ),
    .B1(\u_multiplier/_0480_ ),
    .B2(\u_multiplier/_0455_ ),
    .ZN(product[2]));
 OAI21_X2 \u_multiplier/_0873_  (.A(\u_multiplier/_0478_ ),
    .B1(\u_multiplier/_0479_ ),
    .B2(\u_multiplier/_0455_ ),
    .ZN(\u_multiplier/_0482_ ));
 NAND2_X1 \u_multiplier/_0874_  (.A1(\u_multiplier/_0473_ ),
    .A2(\u_multiplier/_0475_ ),
    .ZN(\u_multiplier/_0483_ ));
 MUX2_X1 \u_multiplier/_0875_  (.A(\u_multiplier/_0403_ ),
    .B(\u_multiplier/_0405_ ),
    .S(\u_multiplier/_0425_ ),
    .Z(\u_multiplier/_0484_ ));
 MUX2_X1 \u_multiplier/_0876_  (.A(\u_multiplier/_0459_ ),
    .B(\u_multiplier/_0484_ ),
    .S(\u_multiplier/_0709_ ),
    .Z(\u_multiplier/_0485_ ));
 MUX2_X1 \u_multiplier/_0877_  (.A(\u_multiplier/_0444_ ),
    .B(\u_multiplier/_0485_ ),
    .S(\u_multiplier/_0710_ ),
    .Z(\u_multiplier/_0486_ ));
 AOI21_X2 \u_multiplier/_0878_  (.A(\u_multiplier/dec_out [3]),
    .B1(\u_multiplier/_0486_ ),
    .B2(\u_multiplier/_0711_ ),
    .ZN(\u_multiplier/_0487_ ));
 MUX2_X1 \u_multiplier/_0879_  (.A(\u_multiplier/_0403_ ),
    .B(\u_multiplier/_0397_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_0488_ ));
 NAND2_X1 \u_multiplier/_0880_  (.A1(\u_multiplier/code_x [1]),
    .A2(\u_multiplier/_0447_ ),
    .ZN(\u_multiplier/_0489_ ));
 OAI21_X2 \u_multiplier/_0881_  (.A(\u_multiplier/_0489_ ),
    .B1(\u_multiplier/_0488_ ),
    .B2(\u_multiplier/code_x [1]),
    .ZN(\u_multiplier/_0490_ ));
 NOR2_X2 \u_multiplier/_0882_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_0490_ ),
    .ZN(\u_multiplier/_0491_ ));
 MUX2_X1 \u_multiplier/_0883_  (.A(\u_multiplier/_0404_ ),
    .B(\u_multiplier/_0399_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_0492_ ));
 MUX2_X1 \u_multiplier/_0884_  (.A(\u_multiplier/_0492_ ),
    .B(\u_multiplier/_0449_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_0493_ ));
 NOR2_X2 \u_multiplier/_0885_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_0493_ ),
    .ZN(\u_multiplier/_0494_ ));
 XNOR2_X2 \u_multiplier/_0886_  (.A(\u_multiplier/_0491_ ),
    .B(\u_multiplier/_0494_ ),
    .ZN(\u_multiplier/_0495_ ));
 NOR2_X1 \u_multiplier/_0887_  (.A1(\u_multiplier/_0487_ ),
    .A2(\u_multiplier/_0495_ ),
    .ZN(\u_multiplier/_0496_ ));
 XOR2_X2 \u_multiplier/_0888_  (.A(\u_multiplier/_0487_ ),
    .B(\u_multiplier/_0495_ ),
    .Z(\u_multiplier/_0497_ ));
 AND2_X1 \u_multiplier/_0889_  (.A1(\u_multiplier/_0483_ ),
    .A2(\u_multiplier/_0497_ ),
    .ZN(\u_multiplier/_0498_ ));
 XOR2_X2 \u_multiplier/_0890_  (.A(\u_multiplier/_0483_ ),
    .B(\u_multiplier/_0497_ ),
    .Z(\u_multiplier/_0499_ ));
 NAND2_X1 \u_multiplier/_0891_  (.A1(\u_multiplier/_0482_ ),
    .A2(\u_multiplier/_0499_ ),
    .ZN(\u_multiplier/_0500_ ));
 OR2_X1 \u_multiplier/_0892_  (.A1(\u_multiplier/_0482_ ),
    .A2(\u_multiplier/_0499_ ),
    .ZN(\u_multiplier/_0501_ ));
 NAND3_X1 \u_multiplier/_0893_  (.A1(\u_multiplier/_0439_ ),
    .A2(\u_multiplier/_0500_ ),
    .A3(\u_multiplier/_0501_ ),
    .ZN(\u_multiplier/_0502_ ));
 INV_X1 \u_multiplier/_0894_  (.A(\u_multiplier/_0502_ ),
    .ZN(product[3]));
 AOI21_X2 \u_multiplier/_0895_  (.A(\u_multiplier/_0498_ ),
    .B1(\u_multiplier/_0499_ ),
    .B2(\u_multiplier/_0482_ ),
    .ZN(\u_multiplier/_0503_ ));
 AOI21_X2 \u_multiplier/_0896_  (.A(\u_multiplier/_0496_ ),
    .B1(\u_multiplier/_0494_ ),
    .B2(\u_multiplier/_0491_ ),
    .ZN(\u_multiplier/_0504_ ));
 MUX2_X1 \u_multiplier/_0897_  (.A(\u_multiplier/_0409_ ),
    .B(\u_multiplier/_0411_ ),
    .S(\u_multiplier/_0425_ ),
    .Z(\u_multiplier/_0505_ ));
 MUX2_X1 \u_multiplier/_0898_  (.A(\u_multiplier/_0484_ ),
    .B(\u_multiplier/_0505_ ),
    .S(\u_multiplier/_0709_ ),
    .Z(\u_multiplier/_0506_ ));
 NAND2_X1 \u_multiplier/_0899_  (.A1(\u_multiplier/_0710_ ),
    .A2(\u_multiplier/_0506_ ),
    .ZN(\u_multiplier/_0507_ ));
 OR3_X1 \u_multiplier/_0900_  (.A1(\u_multiplier/_0710_ ),
    .A2(\u_multiplier/_0460_ ),
    .A3(\u_multiplier/_0461_ ),
    .ZN(\u_multiplier/_0508_ ));
 AND2_X1 \u_multiplier/_0901_  (.A1(\u_multiplier/_0507_ ),
    .A2(\u_multiplier/_0508_ ),
    .ZN(\u_multiplier/_0509_ ));
 AOI21_X1 \u_multiplier/_0902_  (.A(\u_multiplier/dec_out [4]),
    .B1(\u_multiplier/_0427_ ),
    .B2(\u_multiplier/K [2]),
    .ZN(\u_multiplier/_0510_ ));
 OAI21_X2 \u_multiplier/_0903_  (.A(\u_multiplier/_0510_ ),
    .B1(\u_multiplier/_0509_ ),
    .B2(\u_multiplier/K [2]),
    .ZN(\u_multiplier/_0511_ ));
 MUX2_X1 \u_multiplier/_0904_  (.A(\u_multiplier/_0409_ ),
    .B(\u_multiplier/_0403_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_0512_ ));
 NOR2_X1 \u_multiplier/_0905_  (.A1(\u_multiplier/code_x [1]),
    .A2(\u_multiplier/_0512_ ),
    .ZN(\u_multiplier/_0513_ ));
 AOI21_X2 \u_multiplier/_0906_  (.A(\u_multiplier/_0513_ ),
    .B1(\u_multiplier/_0465_ ),
    .B2(\u_multiplier/code_x [1]),
    .ZN(\u_multiplier/_0514_ ));
 MUX2_X1 \u_multiplier/_0907_  (.A(\u_multiplier/_0430_ ),
    .B(\u_multiplier/_0514_ ),
    .S(\u_multiplier/_0708_ ),
    .Z(\u_multiplier/_0515_ ));
 MUX2_X1 \u_multiplier/_0908_  (.A(\u_multiplier/_0411_ ),
    .B(\u_multiplier/_0405_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_0516_ ));
 NOR2_X1 \u_multiplier/_0909_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_0516_ ),
    .ZN(\u_multiplier/_0517_ ));
 AOI21_X2 \u_multiplier/_0910_  (.A(\u_multiplier/_0517_ ),
    .B1(\u_multiplier/_0469_ ),
    .B2(\u_multiplier/code_y [1]),
    .ZN(\u_multiplier/_0518_ ));
 NOR2_X1 \u_multiplier/_0911_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_0518_ ),
    .ZN(\u_multiplier/_0519_ ));
 AOI21_X2 \u_multiplier/_0912_  (.A(\u_multiplier/_0519_ ),
    .B1(\u_multiplier/_0433_ ),
    .B2(\u_multiplier/code_y [2]),
    .ZN(\u_multiplier/_0520_ ));
 NAND2_X1 \u_multiplier/_0913_  (.A1(\u_multiplier/_0515_ ),
    .A2(\u_multiplier/_0520_ ),
    .ZN(\u_multiplier/_0521_ ));
 XOR2_X2 \u_multiplier/_0914_  (.A(\u_multiplier/_0515_ ),
    .B(\u_multiplier/_0520_ ),
    .Z(\u_multiplier/_0522_ ));
 NAND2_X1 \u_multiplier/_0915_  (.A1(\u_multiplier/_0511_ ),
    .A2(\u_multiplier/_0522_ ),
    .ZN(\u_multiplier/_0523_ ));
 XNOR2_X2 \u_multiplier/_0916_  (.A(\u_multiplier/_0511_ ),
    .B(\u_multiplier/_0522_ ),
    .ZN(\u_multiplier/_0524_ ));
 OR2_X1 \u_multiplier/_0917_  (.A1(\u_multiplier/_0504_ ),
    .A2(\u_multiplier/_0524_ ),
    .ZN(\u_multiplier/_0525_ ));
 XNOR2_X2 \u_multiplier/_0918_  (.A(\u_multiplier/_0504_ ),
    .B(\u_multiplier/_0524_ ),
    .ZN(\u_multiplier/_0526_ ));
 AOI21_X1 \u_multiplier/_0919_  (.A(\u_multiplier/_0440_ ),
    .B1(\u_multiplier/_0503_ ),
    .B2(\u_multiplier/_0526_ ),
    .ZN(\u_multiplier/_0527_ ));
 OAI21_X1 \u_multiplier/_0920_  (.A(\u_multiplier/_0527_ ),
    .B1(\u_multiplier/_0526_ ),
    .B2(\u_multiplier/_0503_ ),
    .ZN(\u_multiplier/_0528_ ));
 INV_X1 \u_multiplier/_0921_  (.A(\u_multiplier/_0528_ ),
    .ZN(product[4]));
 OAI21_X2 \u_multiplier/_0922_  (.A(\u_multiplier/_0525_ ),
    .B1(\u_multiplier/_0526_ ),
    .B2(\u_multiplier/_0503_ ),
    .ZN(\u_multiplier/_0529_ ));
 MUX2_X1 \u_multiplier/_0923_  (.A(\u_multiplier/_0414_ ),
    .B(\u_multiplier/_0416_ ),
    .S(\u_multiplier/_0424_ ),
    .Z(\u_multiplier/_0530_ ));
 MUX2_X1 \u_multiplier/_0924_  (.A(\u_multiplier/_0505_ ),
    .B(\u_multiplier/_0530_ ),
    .S(\u_multiplier/_0709_ ),
    .Z(\u_multiplier/_0531_ ));
 MUX2_X1 \u_multiplier/_0925_  (.A(\u_multiplier/_0485_ ),
    .B(\u_multiplier/_0531_ ),
    .S(\u_multiplier/_0710_ ),
    .Z(\u_multiplier/_0532_ ));
 INV_X1 \u_multiplier/_0926_  (.A(\u_multiplier/_0532_ ),
    .ZN(\u_multiplier/_0533_ ));
 AOI21_X1 \u_multiplier/_0927_  (.A(\u_multiplier/dec_out [5]),
    .B1(\u_multiplier/_0445_ ),
    .B2(\u_multiplier/K [2]),
    .ZN(\u_multiplier/_0534_ ));
 OAI21_X2 \u_multiplier/_0928_  (.A(\u_multiplier/_0534_ ),
    .B1(\u_multiplier/_0533_ ),
    .B2(\u_multiplier/K [2]),
    .ZN(\u_multiplier/_0535_ ));
 INV_X1 \u_multiplier/_0929_  (.A(\u_multiplier/_0535_ ),
    .ZN(\u_multiplier/_0536_ ));
 MUX2_X1 \u_multiplier/_0930_  (.A(\u_multiplier/_0416_ ),
    .B(\u_multiplier/_0409_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_0537_ ));
 MUX2_X1 \u_multiplier/_0931_  (.A(\u_multiplier/_0537_ ),
    .B(\u_multiplier/_0488_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_0538_ ));
 NOR2_X1 \u_multiplier/_0932_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_0538_ ),
    .ZN(\u_multiplier/_0539_ ));
 AOI21_X2 \u_multiplier/_0933_  (.A(\u_multiplier/_0539_ ),
    .B1(\u_multiplier/_0448_ ),
    .B2(\u_multiplier/code_x [2]),
    .ZN(\u_multiplier/_0540_ ));
 MUX2_X1 \u_multiplier/_0934_  (.A(\u_multiplier/_0414_ ),
    .B(\u_multiplier/_0411_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_0541_ ));
 NOR2_X1 \u_multiplier/_0935_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_0541_ ),
    .ZN(\u_multiplier/_0542_ ));
 AOI21_X2 \u_multiplier/_0936_  (.A(\u_multiplier/_0542_ ),
    .B1(\u_multiplier/_0492_ ),
    .B2(\u_multiplier/code_y [1]),
    .ZN(\u_multiplier/_0543_ ));
 NOR2_X1 \u_multiplier/_0937_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_0543_ ),
    .ZN(\u_multiplier/_0544_ ));
 AOI21_X2 \u_multiplier/_0938_  (.A(\u_multiplier/_0544_ ),
    .B1(\u_multiplier/_0450_ ),
    .B2(\u_multiplier/code_y [2]),
    .ZN(\u_multiplier/_0545_ ));
 XNOR2_X2 \u_multiplier/_0939_  (.A(\u_multiplier/_0540_ ),
    .B(\u_multiplier/_0545_ ),
    .ZN(\u_multiplier/_0546_ ));
 NOR2_X1 \u_multiplier/_0940_  (.A1(\u_multiplier/_0536_ ),
    .A2(\u_multiplier/_0546_ ),
    .ZN(\u_multiplier/_0547_ ));
 XOR2_X2 \u_multiplier/_0941_  (.A(\u_multiplier/_0535_ ),
    .B(\u_multiplier/_0546_ ),
    .Z(\u_multiplier/_0548_ ));
 AOI21_X2 \u_multiplier/_0942_  (.A(\u_multiplier/_0548_ ),
    .B1(\u_multiplier/_0523_ ),
    .B2(\u_multiplier/_0521_ ),
    .ZN(\u_multiplier/_0549_ ));
 AND3_X1 \u_multiplier/_0943_  (.A1(\u_multiplier/_0521_ ),
    .A2(\u_multiplier/_0523_ ),
    .A3(\u_multiplier/_0548_ ),
    .ZN(\u_multiplier/_0550_ ));
 NOR2_X2 \u_multiplier/_0944_  (.A1(\u_multiplier/_0549_ ),
    .A2(\u_multiplier/_0550_ ),
    .ZN(\u_multiplier/_0551_ ));
 OAI21_X1 \u_multiplier/_0945_  (.A(\u_multiplier/_0439_ ),
    .B1(\u_multiplier/_0529_ ),
    .B2(\u_multiplier/_0551_ ),
    .ZN(\u_multiplier/_0552_ ));
 AOI21_X1 \u_multiplier/_0946_  (.A(\u_multiplier/_0552_ ),
    .B1(\u_multiplier/_0551_ ),
    .B2(\u_multiplier/_0529_ ),
    .ZN(product[5]));
 AOI21_X2 \u_multiplier/_0947_  (.A(\u_multiplier/_0549_ ),
    .B1(\u_multiplier/_0551_ ),
    .B2(\u_multiplier/_0529_ ),
    .ZN(\u_multiplier/_0553_ ));
 AOI21_X2 \u_multiplier/_0948_  (.A(\u_multiplier/_0547_ ),
    .B1(\u_multiplier/_0545_ ),
    .B2(\u_multiplier/_0540_ ),
    .ZN(\u_multiplier/_0554_ ));
 NOR2_X1 \u_multiplier/_0949_  (.A1(\u_multiplier/_0717_ ),
    .A2(\u_multiplier/_0719_ ),
    .ZN(\u_multiplier/_0555_ ));
 MUX2_X1 \u_multiplier/_0950_  (.A(\u_multiplier/_0530_ ),
    .B(\u_multiplier/_0555_ ),
    .S(\u_multiplier/_0709_ ),
    .Z(\u_multiplier/_0556_ ));
 MUX2_X1 \u_multiplier/_0951_  (.A(\u_multiplier/_0506_ ),
    .B(\u_multiplier/_0556_ ),
    .S(\u_multiplier/_0710_ ),
    .Z(\u_multiplier/_0557_ ));
 AND3_X1 \u_multiplier/_0952_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/_0462_ ),
    .A3(\u_multiplier/_0463_ ),
    .ZN(\u_multiplier/_0558_ ));
 AOI211_X2 \u_multiplier/_0953_  (.A(\u_multiplier/dec_out [6]),
    .B(\u_multiplier/_0558_ ),
    .C1(\u_multiplier/_0557_ ),
    .C2(\u_multiplier/_0711_ ),
    .ZN(\u_multiplier/_0559_ ));
 MUX2_X1 \u_multiplier/_0954_  (.A(\u_multiplier/_0718_ ),
    .B(\u_multiplier/_0416_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_0560_ ));
 MUX2_X1 \u_multiplier/_0955_  (.A(\u_multiplier/_0560_ ),
    .B(\u_multiplier/_0512_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_0561_ ));
 NOR2_X1 \u_multiplier/_0956_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_0561_ ),
    .ZN(\u_multiplier/_0562_ ));
 AOI21_X1 \u_multiplier/_0957_  (.A(\u_multiplier/_0562_ ),
    .B1(\u_multiplier/_0467_ ),
    .B2(\u_multiplier/code_x [2]),
    .ZN(\u_multiplier/_0563_ ));
 MUX2_X1 \u_multiplier/_0958_  (.A(\u_multiplier/_0716_ ),
    .B(\u_multiplier/_0414_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_0564_ ));
 MUX2_X1 \u_multiplier/_0959_  (.A(\u_multiplier/_0564_ ),
    .B(\u_multiplier/_0516_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_0565_ ));
 NAND2_X1 \u_multiplier/_0960_  (.A1(\u_multiplier/_0707_ ),
    .A2(\u_multiplier/_0565_ ),
    .ZN(\u_multiplier/_0566_ ));
 OAI21_X1 \u_multiplier/_0961_  (.A(\u_multiplier/_0566_ ),
    .B1(\u_multiplier/_0471_ ),
    .B2(\u_multiplier/_0707_ ),
    .ZN(\u_multiplier/_0567_ ));
 NAND2_X1 \u_multiplier/_0962_  (.A1(\u_multiplier/_0563_ ),
    .A2(\u_multiplier/_0567_ ),
    .ZN(\u_multiplier/_0568_ ));
 XOR2_X1 \u_multiplier/_0963_  (.A(\u_multiplier/_0563_ ),
    .B(\u_multiplier/_0567_ ),
    .Z(\u_multiplier/_0569_ ));
 INV_X1 \u_multiplier/_0964_  (.A(\u_multiplier/_0569_ ),
    .ZN(\u_multiplier/_0570_ ));
 XNOR2_X2 \u_multiplier/_0965_  (.A(\u_multiplier/_0559_ ),
    .B(\u_multiplier/_0570_ ),
    .ZN(\u_multiplier/_0571_ ));
 OR2_X1 \u_multiplier/_0966_  (.A1(\u_multiplier/_0554_ ),
    .A2(\u_multiplier/_0571_ ),
    .ZN(\u_multiplier/_0572_ ));
 XNOR2_X2 \u_multiplier/_0967_  (.A(\u_multiplier/_0554_ ),
    .B(\u_multiplier/_0571_ ),
    .ZN(\u_multiplier/_0573_ ));
 OAI21_X1 \u_multiplier/_0968_  (.A(\u_multiplier/_0439_ ),
    .B1(\u_multiplier/_0553_ ),
    .B2(\u_multiplier/_0573_ ),
    .ZN(\u_multiplier/_0574_ ));
 AOI21_X1 \u_multiplier/_0969_  (.A(\u_multiplier/_0574_ ),
    .B1(\u_multiplier/_0573_ ),
    .B2(\u_multiplier/_0553_ ),
    .ZN(product[6]));
 OAI21_X2 \u_multiplier/_0970_  (.A(\u_multiplier/_0572_ ),
    .B1(\u_multiplier/_0573_ ),
    .B2(\u_multiplier/_0553_ ),
    .ZN(\u_multiplier/_0575_ ));
 OAI21_X1 \u_multiplier/_0971_  (.A(\u_multiplier/_0568_ ),
    .B1(\u_multiplier/_0570_ ),
    .B2(\u_multiplier/_0559_ ),
    .ZN(\u_multiplier/_0576_ ));
 NOR3_X1 \u_multiplier/_0972_  (.A1(\u_multiplier/_0709_ ),
    .A2(\u_multiplier/_0717_ ),
    .A3(\u_multiplier/_0719_ ),
    .ZN(\u_multiplier/_0577_ ));
 MUX2_X1 \u_multiplier/_0973_  (.A(\u_multiplier/_0531_ ),
    .B(\u_multiplier/_0577_ ),
    .S(\u_multiplier/_0710_ ),
    .Z(\u_multiplier/_0578_ ));
 AND2_X1 \u_multiplier/_0974_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/_0486_ ),
    .ZN(\u_multiplier/_0579_ ));
 AOI211_X2 \u_multiplier/_0975_  (.A(\u_multiplier/dec_out [7]),
    .B(\u_multiplier/_0579_ ),
    .C1(\u_multiplier/_0578_ ),
    .C2(\u_multiplier/_0711_ ),
    .ZN(\u_multiplier/_0580_ ));
 INV_X1 \u_multiplier/_0976_  (.A(\u_multiplier/_0580_ ),
    .ZN(\u_multiplier/_0581_ ));
 NAND2_X1 \u_multiplier/_0977_  (.A1(\u_multiplier/code_x [0]),
    .A2(\u_multiplier/_0718_ ),
    .ZN(\u_multiplier/_0582_ ));
 NAND2_X1 \u_multiplier/_0978_  (.A1(\u_multiplier/code_x [1]),
    .A2(\u_multiplier/_0537_ ),
    .ZN(\u_multiplier/_0583_ ));
 OAI21_X2 \u_multiplier/_0979_  (.A(\u_multiplier/_0583_ ),
    .B1(\u_multiplier/_0582_ ),
    .B2(\u_multiplier/code_x [1]),
    .ZN(\u_multiplier/_0584_ ));
 NAND2_X1 \u_multiplier/_0980_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_0490_ ),
    .ZN(\u_multiplier/_0585_ ));
 OAI21_X2 \u_multiplier/_0981_  (.A(\u_multiplier/_0585_ ),
    .B1(\u_multiplier/_0584_ ),
    .B2(\u_multiplier/code_x [2]),
    .ZN(\u_multiplier/_0586_ ));
 NAND2_X1 \u_multiplier/_0982_  (.A1(\u_multiplier/code_y [0]),
    .A2(\u_multiplier/_0716_ ),
    .ZN(\u_multiplier/_0587_ ));
 NAND2_X1 \u_multiplier/_0983_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_0541_ ),
    .ZN(\u_multiplier/_0588_ ));
 OAI21_X2 \u_multiplier/_0984_  (.A(\u_multiplier/_0588_ ),
    .B1(\u_multiplier/_0587_ ),
    .B2(\u_multiplier/code_y [1]),
    .ZN(\u_multiplier/_0589_ ));
 NAND2_X1 \u_multiplier/_0985_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_0493_ ),
    .ZN(\u_multiplier/_0590_ ));
 OAI21_X2 \u_multiplier/_0986_  (.A(\u_multiplier/_0590_ ),
    .B1(\u_multiplier/_0589_ ),
    .B2(\u_multiplier/code_y [2]),
    .ZN(\u_multiplier/_0591_ ));
 XOR2_X2 \u_multiplier/_0987_  (.A(\u_multiplier/_0586_ ),
    .B(\u_multiplier/_0591_ ),
    .Z(\u_multiplier/_0592_ ));
 NAND2_X1 \u_multiplier/_0988_  (.A1(\u_multiplier/_0581_ ),
    .A2(\u_multiplier/_0592_ ),
    .ZN(\u_multiplier/_0593_ ));
 XNOR2_X1 \u_multiplier/_0989_  (.A(\u_multiplier/_0580_ ),
    .B(\u_multiplier/_0592_ ),
    .ZN(\u_multiplier/_0594_ ));
 AND2_X1 \u_multiplier/_0990_  (.A1(\u_multiplier/_0576_ ),
    .A2(\u_multiplier/_0594_ ),
    .ZN(\u_multiplier/_0595_ ));
 XNOR2_X1 \u_multiplier/_0991_  (.A(\u_multiplier/_0576_ ),
    .B(\u_multiplier/_0594_ ),
    .ZN(\u_multiplier/_0596_ ));
 INV_X1 \u_multiplier/_0992_  (.A(\u_multiplier/_0596_ ),
    .ZN(\u_multiplier/_0597_ ));
 OAI21_X1 \u_multiplier/_0993_  (.A(\u_multiplier/_0439_ ),
    .B1(\u_multiplier/_0575_ ),
    .B2(\u_multiplier/_0597_ ),
    .ZN(\u_multiplier/_0598_ ));
 AOI21_X1 \u_multiplier/_0994_  (.A(\u_multiplier/_0598_ ),
    .B1(\u_multiplier/_0597_ ),
    .B2(\u_multiplier/_0575_ ),
    .ZN(product[7]));
 AOI21_X2 \u_multiplier/_0995_  (.A(\u_multiplier/_0595_ ),
    .B1(\u_multiplier/_0597_ ),
    .B2(\u_multiplier/_0575_ ),
    .ZN(\u_multiplier/_0599_ ));
 OAI21_X1 \u_multiplier/_0996_  (.A(\u_multiplier/_0593_ ),
    .B1(\u_multiplier/_0591_ ),
    .B2(\u_multiplier/_0586_ ),
    .ZN(\u_multiplier/_0600_ ));
 NAND2_X1 \u_multiplier/_0997_  (.A1(\u_multiplier/K [1]),
    .A2(\u_multiplier/_0556_ ),
    .ZN(\u_multiplier/_0601_ ));
 NOR2_X1 \u_multiplier/_0998_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/_0601_ ),
    .ZN(\u_multiplier/_0602_ ));
 NOR2_X1 \u_multiplier/_0999_  (.A1(\u_multiplier/dec_out [8]),
    .A2(\u_multiplier/_0602_ ),
    .ZN(\u_multiplier/_0603_ ));
 OAI21_X2 \u_multiplier/_1000_  (.A(\u_multiplier/_0603_ ),
    .B1(\u_multiplier/_0509_ ),
    .B2(\u_multiplier/_0711_ ),
    .ZN(\u_multiplier/_0604_ ));
 AND2_X1 \u_multiplier/_1001_  (.A1(\u_multiplier/code_x [1]),
    .A2(\u_multiplier/_0560_ ),
    .ZN(\u_multiplier/_0605_ ));
 OR2_X1 \u_multiplier/_1002_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_0605_ ),
    .ZN(\u_multiplier/_0606_ ));
 OAI21_X2 \u_multiplier/_1003_  (.A(\u_multiplier/_0606_ ),
    .B1(\u_multiplier/_0514_ ),
    .B2(\u_multiplier/_0708_ ),
    .ZN(\u_multiplier/_0607_ ));
 AND2_X1 \u_multiplier/_1004_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_0564_ ),
    .ZN(\u_multiplier/_0608_ ));
 OR2_X1 \u_multiplier/_1005_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_0608_ ),
    .ZN(\u_multiplier/_0609_ ));
 OAI21_X2 \u_multiplier/_1006_  (.A(\u_multiplier/_0609_ ),
    .B1(\u_multiplier/_0518_ ),
    .B2(\u_multiplier/_0707_ ),
    .ZN(\u_multiplier/_0610_ ));
 NOR2_X1 \u_multiplier/_1007_  (.A1(\u_multiplier/_0607_ ),
    .A2(\u_multiplier/_0610_ ),
    .ZN(\u_multiplier/_0611_ ));
 XOR2_X2 \u_multiplier/_1008_  (.A(\u_multiplier/_0607_ ),
    .B(\u_multiplier/_0610_ ),
    .Z(\u_multiplier/_0612_ ));
 XNOR2_X1 \u_multiplier/_1009_  (.A(\u_multiplier/_0604_ ),
    .B(\u_multiplier/_0612_ ),
    .ZN(\u_multiplier/_0613_ ));
 INV_X1 \u_multiplier/_1010_  (.A(\u_multiplier/_0613_ ),
    .ZN(\u_multiplier/_0614_ ));
 NAND2_X1 \u_multiplier/_1011_  (.A1(\u_multiplier/_0600_ ),
    .A2(\u_multiplier/_0614_ ),
    .ZN(\u_multiplier/_0615_ ));
 XNOR2_X1 \u_multiplier/_1012_  (.A(\u_multiplier/_0600_ ),
    .B(\u_multiplier/_0613_ ),
    .ZN(\u_multiplier/_0616_ ));
 INV_X1 \u_multiplier/_1013_  (.A(\u_multiplier/_0616_ ),
    .ZN(\u_multiplier/_0617_ ));
 OAI21_X1 \u_multiplier/_1014_  (.A(\u_multiplier/_0439_ ),
    .B1(\u_multiplier/_0599_ ),
    .B2(\u_multiplier/_0617_ ),
    .ZN(\u_multiplier/_0618_ ));
 AOI21_X2 \u_multiplier/_1015_  (.A(\u_multiplier/_0618_ ),
    .B1(\u_multiplier/_0617_ ),
    .B2(\u_multiplier/_0599_ ),
    .ZN(product[8]));
 OAI21_X2 \u_multiplier/_1016_  (.A(\u_multiplier/_0615_ ),
    .B1(\u_multiplier/_0617_ ),
    .B2(\u_multiplier/_0599_ ),
    .ZN(\u_multiplier/_0619_ ));
 AOI21_X2 \u_multiplier/_1017_  (.A(\u_multiplier/_0611_ ),
    .B1(\u_multiplier/_0612_ ),
    .B2(\u_multiplier/_0604_ ),
    .ZN(\u_multiplier/_0620_ ));
 NOR2_X1 \u_multiplier/_1018_  (.A1(\u_multiplier/_0711_ ),
    .A2(\u_multiplier/_0533_ ),
    .ZN(\u_multiplier/_0621_ ));
 AND2_X1 \u_multiplier/_1019_  (.A1(\u_multiplier/K [1]),
    .A2(\u_multiplier/_0577_ ),
    .ZN(\u_multiplier/_0622_ ));
 AOI211_X2 \u_multiplier/_1020_  (.A(\u_multiplier/dec_out [9]),
    .B(\u_multiplier/_0621_ ),
    .C1(\u_multiplier/_0622_ ),
    .C2(\u_multiplier/_0711_ ),
    .ZN(\u_multiplier/_0623_ ));
 INV_X1 \u_multiplier/_1021_  (.A(\u_multiplier/_0623_ ),
    .ZN(\u_multiplier/_0624_ ));
 AND3_X1 \u_multiplier/_1022_  (.A1(\u_multiplier/code_x [0]),
    .A2(\u_multiplier/code_x [1]),
    .A3(\u_multiplier/_0718_ ),
    .ZN(\u_multiplier/_0625_ ));
 OR2_X1 \u_multiplier/_1023_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_0625_ ),
    .ZN(\u_multiplier/_0626_ ));
 OAI21_X2 \u_multiplier/_1024_  (.A(\u_multiplier/_0626_ ),
    .B1(\u_multiplier/_0538_ ),
    .B2(\u_multiplier/_0708_ ),
    .ZN(\u_multiplier/_0627_ ));
 AND3_X1 \u_multiplier/_1025_  (.A1(\u_multiplier/code_y [0]),
    .A2(\u_multiplier/code_y [1]),
    .A3(\u_multiplier/_0716_ ),
    .ZN(\u_multiplier/_0628_ ));
 OR2_X1 \u_multiplier/_1026_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_0628_ ),
    .ZN(\u_multiplier/_0629_ ));
 OAI21_X2 \u_multiplier/_1027_  (.A(\u_multiplier/_0629_ ),
    .B1(\u_multiplier/_0543_ ),
    .B2(\u_multiplier/_0707_ ),
    .ZN(\u_multiplier/_0630_ ));
 NOR2_X1 \u_multiplier/_1028_  (.A1(\u_multiplier/_0627_ ),
    .A2(\u_multiplier/_0630_ ),
    .ZN(\u_multiplier/_0631_ ));
 XOR2_X2 \u_multiplier/_1029_  (.A(\u_multiplier/_0627_ ),
    .B(\u_multiplier/_0630_ ),
    .Z(\u_multiplier/_0632_ ));
 XNOR2_X1 \u_multiplier/_1030_  (.A(\u_multiplier/_0623_ ),
    .B(\u_multiplier/_0632_ ),
    .ZN(\u_multiplier/_0633_ ));
 INV_X1 \u_multiplier/_1031_  (.A(\u_multiplier/_0633_ ),
    .ZN(\u_multiplier/_0634_ ));
 NOR2_X1 \u_multiplier/_1032_  (.A1(\u_multiplier/_0620_ ),
    .A2(\u_multiplier/_0634_ ),
    .ZN(\u_multiplier/_0635_ ));
 XOR2_X1 \u_multiplier/_1033_  (.A(\u_multiplier/_0620_ ),
    .B(\u_multiplier/_0633_ ),
    .Z(\u_multiplier/_0636_ ));
 INV_X1 \u_multiplier/_1034_  (.A(\u_multiplier/_0636_ ),
    .ZN(\u_multiplier/_0637_ ));
 OAI21_X1 \u_multiplier/_1035_  (.A(\u_multiplier/_0439_ ),
    .B1(\u_multiplier/_0619_ ),
    .B2(\u_multiplier/_0637_ ),
    .ZN(\u_multiplier/_0638_ ));
 AOI21_X1 \u_multiplier/_1036_  (.A(\u_multiplier/_0638_ ),
    .B1(\u_multiplier/_0637_ ),
    .B2(\u_multiplier/_0619_ ),
    .ZN(product[9]));
 AOI21_X2 \u_multiplier/_1037_  (.A(\u_multiplier/_0635_ ),
    .B1(\u_multiplier/_0637_ ),
    .B2(\u_multiplier/_0619_ ),
    .ZN(\u_multiplier/_0639_ ));
 AOI21_X1 \u_multiplier/_1038_  (.A(\u_multiplier/_0631_ ),
    .B1(\u_multiplier/_0632_ ),
    .B2(\u_multiplier/_0624_ ),
    .ZN(\u_multiplier/_0640_ ));
 AOI21_X2 \u_multiplier/_1039_  (.A(\u_multiplier/dec_out [10]),
    .B1(\u_multiplier/_0557_ ),
    .B2(\u_multiplier/K [2]),
    .ZN(\u_multiplier/_0641_ ));
 NAND2_X1 \u_multiplier/_1040_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_0561_ ),
    .ZN(\u_multiplier/_0642_ ));
 NAND2_X1 \u_multiplier/_1041_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_0565_ ),
    .ZN(\u_multiplier/_0643_ ));
 OR2_X1 \u_multiplier/_1042_  (.A1(\u_multiplier/_0642_ ),
    .A2(\u_multiplier/_0643_ ),
    .ZN(\u_multiplier/_0644_ ));
 XOR2_X1 \u_multiplier/_1043_  (.A(\u_multiplier/_0642_ ),
    .B(\u_multiplier/_0643_ ),
    .Z(\u_multiplier/_0645_ ));
 INV_X1 \u_multiplier/_1044_  (.A(\u_multiplier/_0645_ ),
    .ZN(\u_multiplier/_0646_ ));
 XNOR2_X1 \u_multiplier/_1045_  (.A(\u_multiplier/_0641_ ),
    .B(\u_multiplier/_0646_ ),
    .ZN(\u_multiplier/_0647_ ));
 OR2_X1 \u_multiplier/_1046_  (.A1(\u_multiplier/_0640_ ),
    .A2(\u_multiplier/_0647_ ),
    .ZN(\u_multiplier/_0648_ ));
 XOR2_X1 \u_multiplier/_1047_  (.A(\u_multiplier/_0640_ ),
    .B(\u_multiplier/_0647_ ),
    .Z(\u_multiplier/_0649_ ));
 INV_X1 \u_multiplier/_1048_  (.A(\u_multiplier/_0649_ ),
    .ZN(\u_multiplier/_0650_ ));
 NOR2_X1 \u_multiplier/_1049_  (.A1(\u_multiplier/_0639_ ),
    .A2(\u_multiplier/_0650_ ),
    .ZN(\u_multiplier/_0651_ ));
 AND2_X1 \u_multiplier/_1050_  (.A1(\u_multiplier/_0639_ ),
    .A2(\u_multiplier/_0650_ ),
    .ZN(\u_multiplier/_0652_ ));
 NOR3_X1 \u_multiplier/_1051_  (.A1(\u_multiplier/_0440_ ),
    .A2(\u_multiplier/_0651_ ),
    .A3(\u_multiplier/_0652_ ),
    .ZN(product[10]));
 OAI21_X2 \u_multiplier/_1052_  (.A(\u_multiplier/_0648_ ),
    .B1(\u_multiplier/_0650_ ),
    .B2(\u_multiplier/_0639_ ),
    .ZN(\u_multiplier/_0653_ ));
 OAI21_X2 \u_multiplier/_1053_  (.A(\u_multiplier/_0644_ ),
    .B1(\u_multiplier/_0646_ ),
    .B2(\u_multiplier/_0641_ ),
    .ZN(\u_multiplier/_0654_ ));
 INV_X1 \u_multiplier/_1054_  (.A(\u_multiplier/_0654_ ),
    .ZN(\u_multiplier/_0655_ ));
 AOI21_X2 \u_multiplier/_1055_  (.A(\u_multiplier/dec_out [11]),
    .B1(\u_multiplier/_0578_ ),
    .B2(\u_multiplier/K [2]),
    .ZN(\u_multiplier/_0656_ ));
 NAND2_X1 \u_multiplier/_1056_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_0584_ ),
    .ZN(\u_multiplier/_0657_ ));
 NAND2_X2 \u_multiplier/_1057_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_0589_ ),
    .ZN(\u_multiplier/_0658_ ));
 XNOR2_X2 \u_multiplier/_1058_  (.A(\u_multiplier/_0657_ ),
    .B(\u_multiplier/_0658_ ),
    .ZN(\u_multiplier/_0659_ ));
 OR2_X1 \u_multiplier/_1059_  (.A1(\u_multiplier/_0656_ ),
    .A2(\u_multiplier/_0659_ ),
    .ZN(\u_multiplier/_0660_ ));
 XNOR2_X2 \u_multiplier/_1060_  (.A(\u_multiplier/_0656_ ),
    .B(\u_multiplier/_0659_ ),
    .ZN(\u_multiplier/_0661_ ));
 NOR2_X1 \u_multiplier/_1061_  (.A1(\u_multiplier/_0655_ ),
    .A2(\u_multiplier/_0661_ ),
    .ZN(\u_multiplier/_0662_ ));
 XNOR2_X2 \u_multiplier/_1062_  (.A(\u_multiplier/_0654_ ),
    .B(\u_multiplier/_0661_ ),
    .ZN(\u_multiplier/_0663_ ));
 OAI21_X1 \u_multiplier/_1063_  (.A(\u_multiplier/_0439_ ),
    .B1(\u_multiplier/_0653_ ),
    .B2(\u_multiplier/_0663_ ),
    .ZN(\u_multiplier/_0664_ ));
 AOI21_X1 \u_multiplier/_1064_  (.A(\u_multiplier/_0664_ ),
    .B1(\u_multiplier/_0663_ ),
    .B2(\u_multiplier/_0653_ ),
    .ZN(product[11]));
 AOI21_X2 \u_multiplier/_1065_  (.A(\u_multiplier/_0662_ ),
    .B1(\u_multiplier/_0663_ ),
    .B2(\u_multiplier/_0653_ ),
    .ZN(\u_multiplier/_0665_ ));
 OAI21_X2 \u_multiplier/_1066_  (.A(\u_multiplier/_0660_ ),
    .B1(\u_multiplier/_0658_ ),
    .B2(\u_multiplier/_0657_ ),
    .ZN(\u_multiplier/_0666_ ));
 OAI21_X2 \u_multiplier/_1067_  (.A(\u_multiplier/_0712_ ),
    .B1(\u_multiplier/_0601_ ),
    .B2(\u_multiplier/_0711_ ),
    .ZN(\u_multiplier/_0667_ ));
 AND4_X1 \u_multiplier/_1068_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/code_x [2]),
    .A3(\u_multiplier/_0605_ ),
    .A4(\u_multiplier/_0608_ ),
    .ZN(\u_multiplier/_0668_ ));
 AOI22_X1 \u_multiplier/_1069_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_0605_ ),
    .B1(\u_multiplier/_0608_ ),
    .B2(\u_multiplier/code_y [2]),
    .ZN(\u_multiplier/_0669_ ));
 NOR2_X1 \u_multiplier/_1070_  (.A1(\u_multiplier/_0668_ ),
    .A2(\u_multiplier/_0669_ ),
    .ZN(\u_multiplier/_0670_ ));
 XNOR2_X1 \u_multiplier/_1071_  (.A(\u_multiplier/_0667_ ),
    .B(\u_multiplier/_0670_ ),
    .ZN(\u_multiplier/_0671_ ));
 INV_X1 \u_multiplier/_1072_  (.A(\u_multiplier/_0671_ ),
    .ZN(\u_multiplier/_0672_ ));
 NAND2_X1 \u_multiplier/_1073_  (.A1(\u_multiplier/_0666_ ),
    .A2(\u_multiplier/_0672_ ),
    .ZN(\u_multiplier/_0673_ ));
 XNOR2_X2 \u_multiplier/_1074_  (.A(\u_multiplier/_0666_ ),
    .B(\u_multiplier/_0672_ ),
    .ZN(\u_multiplier/_0674_ ));
 AOI21_X1 \u_multiplier/_1075_  (.A(\u_multiplier/_0440_ ),
    .B1(\u_multiplier/_0665_ ),
    .B2(\u_multiplier/_0674_ ),
    .ZN(\u_multiplier/_0675_ ));
 OAI21_X1 \u_multiplier/_1076_  (.A(\u_multiplier/_0675_ ),
    .B1(\u_multiplier/_0674_ ),
    .B2(\u_multiplier/_0665_ ),
    .ZN(\u_multiplier/_0676_ ));
 INV_X1 \u_multiplier/_1077_  (.A(\u_multiplier/_0676_ ),
    .ZN(product[12]));
 OAI21_X2 \u_multiplier/_1078_  (.A(\u_multiplier/_0673_ ),
    .B1(\u_multiplier/_0674_ ),
    .B2(\u_multiplier/_0665_ ),
    .ZN(\u_multiplier/_0677_ ));
 AOI21_X2 \u_multiplier/_1079_  (.A(\u_multiplier/_0668_ ),
    .B1(\u_multiplier/_0670_ ),
    .B2(\u_multiplier/_0667_ ),
    .ZN(\u_multiplier/_0678_ ));
 INV_X1 \u_multiplier/_1080_  (.A(\u_multiplier/_0678_ ),
    .ZN(\u_multiplier/_0679_ ));
 AOI21_X2 \u_multiplier/_1081_  (.A(\u_multiplier/dec_out [13]),
    .B1(\u_multiplier/_0622_ ),
    .B2(\u_multiplier/K [2]),
    .ZN(\u_multiplier/_0680_ ));
 INV_X1 \u_multiplier/_1082_  (.A(\u_multiplier/_0680_ ),
    .ZN(\u_multiplier/_0681_ ));
 AND4_X1 \u_multiplier/_1083_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/code_x [2]),
    .A3(\u_multiplier/_0625_ ),
    .A4(\u_multiplier/_0628_ ),
    .ZN(\u_multiplier/_0682_ ));
 AOI22_X2 \u_multiplier/_1084_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_0625_ ),
    .B1(\u_multiplier/_0628_ ),
    .B2(\u_multiplier/code_y [2]),
    .ZN(\u_multiplier/_0683_ ));
 NOR2_X2 \u_multiplier/_1085_  (.A1(\u_multiplier/_0682_ ),
    .A2(\u_multiplier/_0683_ ),
    .ZN(\u_multiplier/_0684_ ));
 XNOR2_X2 \u_multiplier/_1086_  (.A(\u_multiplier/_0680_ ),
    .B(\u_multiplier/_0684_ ),
    .ZN(\u_multiplier/_0685_ ));
 NAND2_X1 \u_multiplier/_1087_  (.A1(\u_multiplier/_0679_ ),
    .A2(\u_multiplier/_0685_ ),
    .ZN(\u_multiplier/_0686_ ));
 INV_X1 \u_multiplier/_1088_  (.A(\u_multiplier/_0686_ ),
    .ZN(\u_multiplier/_0687_ ));
 XNOR2_X2 \u_multiplier/_1089_  (.A(\u_multiplier/_0678_ ),
    .B(\u_multiplier/_0685_ ),
    .ZN(\u_multiplier/_0688_ ));
 OAI21_X1 \u_multiplier/_1090_  (.A(\u_multiplier/_0439_ ),
    .B1(\u_multiplier/_0677_ ),
    .B2(\u_multiplier/_0688_ ),
    .ZN(\u_multiplier/_0689_ ));
 AOI21_X1 \u_multiplier/_1091_  (.A(\u_multiplier/_0689_ ),
    .B1(\u_multiplier/_0688_ ),
    .B2(\u_multiplier/_0677_ ),
    .ZN(product[13]));
 AOI21_X2 \u_multiplier/_1092_  (.A(\u_multiplier/_0687_ ),
    .B1(\u_multiplier/_0688_ ),
    .B2(\u_multiplier/_0677_ ),
    .ZN(\u_multiplier/_0690_ ));
 AOI21_X2 \u_multiplier/_1093_  (.A(\u_multiplier/_0682_ ),
    .B1(\u_multiplier/_0684_ ),
    .B2(\u_multiplier/_0681_ ),
    .ZN(\u_multiplier/_0691_ ));
 INV_X1 \u_multiplier/_1094_  (.A(\u_multiplier/_0691_ ),
    .ZN(\u_multiplier/_0692_ ));
 NAND2_X1 \u_multiplier/_1095_  (.A1(\u_multiplier/dec_out [14]),
    .A2(\u_multiplier/_0692_ ),
    .ZN(\u_multiplier/_0693_ ));
 XOR2_X2 \u_multiplier/_1096_  (.A(\u_multiplier/dec_out [14]),
    .B(\u_multiplier/_0691_ ),
    .Z(\u_multiplier/_0694_ ));
 OR2_X1 \u_multiplier/_1097_  (.A1(\u_multiplier/_0690_ ),
    .A2(\u_multiplier/_0694_ ),
    .ZN(\u_multiplier/_0695_ ));
 NAND2_X1 \u_multiplier/_1098_  (.A1(\u_multiplier/_0439_ ),
    .A2(\u_multiplier/_0695_ ),
    .ZN(\u_multiplier/_0696_ ));
 AOI21_X4 \u_multiplier/_1099_  (.A(\u_multiplier/_0696_ ),
    .B1(\u_multiplier/_0694_ ),
    .B2(\u_multiplier/_0690_ ),
    .ZN(product[14]));
 AOI21_X1 \u_multiplier/_1100_  (.A(\u_multiplier/_0713_ ),
    .B1(\u_multiplier/_0693_ ),
    .B2(\u_multiplier/_0695_ ),
    .ZN(\u_multiplier/_0697_ ));
 AND3_X1 \u_multiplier/_1101_  (.A1(\u_multiplier/_0713_ ),
    .A2(\u_multiplier/_0693_ ),
    .A3(\u_multiplier/_0695_ ),
    .ZN(\u_multiplier/_0698_ ));
 NOR3_X1 \u_multiplier/_1102_  (.A1(\u_multiplier/_0440_ ),
    .A2(\u_multiplier/_0697_ ),
    .A3(\u_multiplier/_0698_ ),
    .ZN(product[15]));
 NAND2_X1 \u_multiplier/_1103_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/code_x [2]),
    .ZN(\u_multiplier/_0699_ ));
 NAND2_X1 \u_multiplier/_1104_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/code_x [1]),
    .ZN(\u_multiplier/_0700_ ));
 NAND2_X1 \u_multiplier/_1105_  (.A1(\u_multiplier/code_y [0]),
    .A2(\u_multiplier/code_x [0]),
    .ZN(\u_multiplier/_0701_ ));
 NOR2_X1 \u_multiplier/_1106_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/code_x [1]),
    .ZN(\u_multiplier/_0702_ ));
 XOR2_X2 \u_multiplier/_1107_  (.A(\u_multiplier/code_y [1]),
    .B(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_0703_ ));
 OAI21_X2 \u_multiplier/_1108_  (.A(\u_multiplier/_0700_ ),
    .B1(\u_multiplier/_0701_ ),
    .B2(\u_multiplier/_0702_ ),
    .ZN(\u_multiplier/_0704_ ));
 INV_X1 \u_multiplier/_1109_  (.A(\u_multiplier/_0704_ ),
    .ZN(\u_multiplier/_0705_ ));
 XNOR2_X2 \u_multiplier/_1110_  (.A(\u_multiplier/code_y [2]),
    .B(\u_multiplier/code_x [2]),
    .ZN(\u_multiplier/_0706_ ));
 OAI21_X4 \u_multiplier/_1111_  (.A(\u_multiplier/_0699_ ),
    .B1(\u_multiplier/_0705_ ),
    .B2(\u_multiplier/_0706_ ),
    .ZN(\u_multiplier/_0355_ ));
 XNOR2_X2 \u_multiplier/_1112_  (.A(\u_multiplier/_0701_ ),
    .B(\u_multiplier/_0703_ ),
    .ZN(\u_multiplier/_0353_ ));
 XNOR2_X2 \u_multiplier/_1113_  (.A(\u_multiplier/_0704_ ),
    .B(\u_multiplier/_0706_ ),
    .ZN(\u_multiplier/_0354_ ));
 XOR2_X2 \u_multiplier/_1114_  (.A(\u_multiplier/code_y [0]),
    .B(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_0352_ ));
 INV_X2 \u_multiplier/dec/_40_  (.A(\u_multiplier/_0355_ ),
    .ZN(\u_multiplier/dec/_34_ ));
 INV_X1 \u_multiplier/dec/_41_  (.A(\u_multiplier/_0352_ ),
    .ZN(\u_multiplier/dec/_35_ ));
 INV_X2 \u_multiplier/dec/_42_  (.A(\u_multiplier/_0353_ ),
    .ZN(\u_multiplier/dec/_36_ ));
 INV_X2 \u_multiplier/dec/_43_  (.A(\u_multiplier/_0354_ ),
    .ZN(\u_multiplier/dec/_37_ ));
 NOR4_X1 \u_multiplier/dec/_44_  (.A1(\u_multiplier/_0355_ ),
    .A2(\u_multiplier/_0352_ ),
    .A3(\u_multiplier/_0353_ ),
    .A4(\u_multiplier/_0354_ ),
    .ZN(\u_multiplier/dec_out [0]));
 NOR4_X2 \u_multiplier/dec/_45_  (.A1(\u_multiplier/_0355_ ),
    .A2(\u_multiplier/dec/_35_ ),
    .A3(\u_multiplier/_0353_ ),
    .A4(\u_multiplier/_0354_ ),
    .ZN(\u_multiplier/dec_out [1]));
 NOR4_X2 \u_multiplier/dec/_46_  (.A1(\u_multiplier/_0355_ ),
    .A2(\u_multiplier/_0352_ ),
    .A3(\u_multiplier/dec/_36_ ),
    .A4(\u_multiplier/_0354_ ),
    .ZN(\u_multiplier/dec_out [2]));
 NAND2_X1 \u_multiplier/dec/_47_  (.A1(\u_multiplier/_0352_ ),
    .A2(\u_multiplier/_0353_ ),
    .ZN(\u_multiplier/dec/_38_ ));
 NOR3_X1 \u_multiplier/dec/_48_  (.A1(\u_multiplier/_0355_ ),
    .A2(\u_multiplier/_0354_ ),
    .A3(\u_multiplier/dec/_38_ ),
    .ZN(\u_multiplier/dec_out [3]));
 NOR4_X1 \u_multiplier/dec/_49_  (.A1(\u_multiplier/_0355_ ),
    .A2(\u_multiplier/_0352_ ),
    .A3(\u_multiplier/_0353_ ),
    .A4(\u_multiplier/dec/_37_ ),
    .ZN(\u_multiplier/dec_out [4]));
 NOR4_X1 \u_multiplier/dec/_50_  (.A1(\u_multiplier/_0355_ ),
    .A2(\u_multiplier/dec/_35_ ),
    .A3(\u_multiplier/_0353_ ),
    .A4(\u_multiplier/dec/_37_ ),
    .ZN(\u_multiplier/dec_out [5]));
 NOR4_X1 \u_multiplier/dec/_51_  (.A1(\u_multiplier/_0355_ ),
    .A2(\u_multiplier/_0352_ ),
    .A3(\u_multiplier/dec/_36_ ),
    .A4(\u_multiplier/dec/_37_ ),
    .ZN(\u_multiplier/dec_out [6]));
 NAND3_X1 \u_multiplier/dec/_52_  (.A1(\u_multiplier/_0352_ ),
    .A2(\u_multiplier/_0353_ ),
    .A3(\u_multiplier/_0354_ ),
    .ZN(\u_multiplier/dec/_39_ ));
 NOR2_X1 \u_multiplier/dec/_53_  (.A1(\u_multiplier/_0355_ ),
    .A2(\u_multiplier/dec/_39_ ),
    .ZN(\u_multiplier/dec_out [7]));
 NOR4_X1 \u_multiplier/dec/_54_  (.A1(\u_multiplier/dec/_34_ ),
    .A2(\u_multiplier/_0352_ ),
    .A3(\u_multiplier/_0353_ ),
    .A4(\u_multiplier/_0354_ ),
    .ZN(\u_multiplier/dec_out [8]));
 NOR4_X1 \u_multiplier/dec/_55_  (.A1(\u_multiplier/dec/_34_ ),
    .A2(\u_multiplier/dec/_35_ ),
    .A3(\u_multiplier/_0353_ ),
    .A4(\u_multiplier/_0354_ ),
    .ZN(\u_multiplier/dec_out [9]));
 NOR4_X2 \u_multiplier/dec/_56_  (.A1(\u_multiplier/dec/_34_ ),
    .A2(\u_multiplier/_0352_ ),
    .A3(\u_multiplier/dec/_36_ ),
    .A4(\u_multiplier/_0354_ ),
    .ZN(\u_multiplier/dec_out [10]));
 NOR3_X1 \u_multiplier/dec/_57_  (.A1(\u_multiplier/dec/_34_ ),
    .A2(\u_multiplier/_0354_ ),
    .A3(\u_multiplier/dec/_38_ ),
    .ZN(\u_multiplier/dec_out [11]));
 NOR4_X1 \u_multiplier/dec/_58_  (.A1(\u_multiplier/dec/_34_ ),
    .A2(\u_multiplier/_0352_ ),
    .A3(\u_multiplier/_0353_ ),
    .A4(\u_multiplier/dec/_37_ ),
    .ZN(\u_multiplier/dec_out [12]));
 NOR4_X1 \u_multiplier/dec/_59_  (.A1(\u_multiplier/dec/_34_ ),
    .A2(\u_multiplier/dec/_35_ ),
    .A3(\u_multiplier/_0353_ ),
    .A4(\u_multiplier/dec/_37_ ),
    .ZN(\u_multiplier/dec_out [13]));
 NOR4_X4 \u_multiplier/dec/_60_  (.A1(\u_multiplier/dec/_34_ ),
    .A2(\u_multiplier/_0352_ ),
    .A3(\u_multiplier/dec/_36_ ),
    .A4(\u_multiplier/dec/_37_ ),
    .ZN(\u_multiplier/dec_out [14]));
 NOR2_X1 \u_multiplier/dec/_61_  (.A1(\u_multiplier/dec/_34_ ),
    .A2(\u_multiplier/dec/_39_ ),
    .ZN(\u_multiplier/dec_out [15]));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_2_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_2_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_2_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_2_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_2_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_2_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_2_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_2_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_2_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_2_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_2_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_2_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_2_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_2_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_2_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_2_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_2_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_2_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_2_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_2_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_2_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_2_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_2_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_2_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_2_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_2_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_2_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_2_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_2_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_2_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_2_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_2_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_2_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_2_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_2_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_2_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_2_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_2_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_2_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_2_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_2_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_2_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_2_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_2_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_2_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_2_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_2_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_2_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_2_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_2_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_2_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_2_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_2_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_2_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_2_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_2_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_2_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_2_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_2_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_2_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_2_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_2_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_2_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_2_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_2_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_2_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_2_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_2_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_2_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_2_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_2_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_2_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_2_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_2_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_1_Left_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_1_Left_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_1_Left_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_1_Left_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_1_Left_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_1_Left_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_1_Left_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_1_Left_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_1_Left_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_1_Left_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_1_Left_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_1_Left_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_1_Left_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_1_Left_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_1_Left_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_1_Left_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_1_Left_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_1_Left_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_1_Left_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_1_Left_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_1_Left_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_1_Left_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_1_Left_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_1_Left_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_1_Left_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_1_Left_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_1_Left_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_1_Left_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_1_Left_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_1_Left_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_1_Left_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_1_Left_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_1_Left_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_1_Left_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_1_Left_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_1_Left_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_1_Left_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_1_Left_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_1_Left_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_1_Left_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_1_Left_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_1_Left_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_1_Left_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_1_Left_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_1_Left_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_1_Left_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_1_Left_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_1_Left_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_1_Left_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_1_Left_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_1_Left_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_1_Left_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_1_Left_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_1_Left_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_1_Left_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_1_Left_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_1_Left_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_1_Left_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_1_Left_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_1_Left_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_1_Left_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_1_Left_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_1_Left_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_1_Left_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_1_Left_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_1_Left_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_1_Left_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_1_Left_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_1_Left_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_1_Left_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_1_Left_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_1_Left_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_1_Left_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Left_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Left_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Left_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Left_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Left_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Left_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Left_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Left_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Left_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Left_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_1_Left_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_2_Left_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_2_Left_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_2_Left_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_2_Left_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_2_Left_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_2_Left_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_2_Left_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_2_Left_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_2_Left_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_2_Left_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_2_Left_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_2_Left_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_2_Left_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_2_Left_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_2_Left_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_2_Left_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_2_Left_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_2_Left_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_2_Left_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_2_Left_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_2_Left_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_2_Left_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_2_Left_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_2_Left_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_2_Left_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_2_Left_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_2_Left_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_2_Left_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_2_Left_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_2_Left_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_2_Left_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_2_Left_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_2_Left_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_2_Left_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_2_Left_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_2_Left_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_2_Left_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_2_Left_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_2_Left_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_2_Left_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_2_Left_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_2_Left_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_2_Left_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_2_Left_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_2_Left_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_2_Left_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_2_Left_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_2_Left_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_2_Left_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_2_Left_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_2_Left_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_2_Left_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_2_Left_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_2_Left_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_2_Left_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_2_Left_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_2_Left_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_2_Left_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_2_Left_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_2_Left_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_2_Left_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_2_Left_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_2_Left_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_2_Left_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_2_Left_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_2_Left_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_2_Left_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_2_Left_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_2_Left_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_2_Left_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_2_Left_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_2_Left_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_2_Left_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_2_Left_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_1_Right_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_1_Right_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_1_Right_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_1_Right_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_1_Right_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_1_Right_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_1_Right_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_1_Right_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_1_Right_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_1_Right_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_1_Right_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_1_Right_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_1_Right_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_1_Right_265 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_1_Right_266 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_1_Right_267 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_1_Right_268 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_1_Right_269 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_1_Right_270 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_1_Right_271 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_1_Right_272 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_1_Right_273 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_1_Right_274 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_1_Right_275 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_1_Right_276 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_1_Right_277 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_1_Right_278 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_1_Right_279 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_1_Right_280 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_1_Right_281 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_1_Right_282 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_1_Right_283 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_1_Right_284 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_1_Right_285 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_1_Right_286 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_1_Right_287 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_1_Right_288 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_1_Right_289 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_1_Right_290 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_1_Right_291 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_1_Right_292 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_1_Right_293 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_1_Right_294 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_1_Right_295 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_1_Right_296 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_1_Right_297 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_1_Right_298 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_1_Right_299 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_1_Right_300 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_1_Right_301 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_1_Right_302 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_1_Right_303 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_1_Right_304 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_1_Right_305 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_1_Right_306 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_1_Right_307 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_1_Right_308 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_1_Right_309 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_1_Right_310 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_1_Right_311 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_1_Right_312 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_1_Right_313 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_1_Right_314 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_1_Right_315 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_1_Right_316 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_1_Right_317 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_1_Right_318 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_1_Right_319 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_1_Right_320 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_1_Right_321 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_1_Right_322 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_1_Right_323 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_1_Right_324 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_1_Right_325 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_326 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_327 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_328 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_79_329 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_330 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_331 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_332 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_333 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_334 ();
 LOGIC1_X1 \u_multiplier/NOD/nod_cels[5].Nod_bits/_07__30  (.Z(net30));
 CLKBUF_X1 hold31 (.A(net56),
    .Z(net31));
 BUF_X2 input1 (.A(data_in[0]),
    .Z(net1));
 BUF_X1 input2 (.A(data_in[1]),
    .Z(net2));
 BUF_X1 input3 (.A(data_in[2]),
    .Z(net3));
 CLKBUF_X2 input4 (.A(data_in[3]),
    .Z(net4));
 CLKBUF_X2 input5 (.A(data_in[4]),
    .Z(net5));
 BUF_X1 input6 (.A(data_in[5]),
    .Z(net6));
 BUF_X2 input7 (.A(data_in[6]),
    .Z(net7));
 BUF_X1 input8 (.A(data_in[7]),
    .Z(net8));
 BUF_X2 input9 (.A(init_enable),
    .Z(net9));
 BUF_X2 input10 (.A(pe_ce),
    .Z(net10));
 BUF_X8 input11 (.A(rst_n),
    .Z(net11));
 BUF_X1 output12 (.A(net12),
    .Z(curr_state[1]));
 BUF_X1 output13 (.A(net13),
    .Z(data_out[0]));
 BUF_X1 output14 (.A(net14),
    .Z(data_out[10]));
 BUF_X1 output15 (.A(net15),
    .Z(data_out[11]));
 BUF_X1 output16 (.A(net16),
    .Z(data_out[12]));
 BUF_X1 output17 (.A(net17),
    .Z(data_out[13]));
 BUF_X1 output18 (.A(net18),
    .Z(data_out[14]));
 BUF_X1 output19 (.A(net19),
    .Z(data_out[15]));
 BUF_X1 output20 (.A(net20),
    .Z(data_out[1]));
 BUF_X1 output21 (.A(net21),
    .Z(data_out[2]));
 BUF_X1 output22 (.A(net22),
    .Z(data_out[3]));
 BUF_X1 output23 (.A(net23),
    .Z(data_out[4]));
 BUF_X1 output24 (.A(net24),
    .Z(data_out[5]));
 BUF_X1 output25 (.A(net25),
    .Z(data_out[6]));
 BUF_X1 output26 (.A(net26),
    .Z(data_out[7]));
 BUF_X1 output27 (.A(net27),
    .Z(data_out[8]));
 BUF_X1 output28 (.A(net28),
    .Z(data_out[9]));
 BUF_X1 output29 (.A(net29),
    .Z(valid_reg_out));
 CLKBUF_X1 hold32 (.A(net60),
    .Z(net32));
 CLKBUF_X1 hold33 (.A(net67),
    .Z(net33));
 CLKBUF_X1 hold34 (.A(net53),
    .Z(net34));
 CLKBUF_X1 hold35 (.A(net65),
    .Z(net35));
 CLKBUF_X1 hold36 (.A(net69),
    .Z(net36));
 CLKBUF_X1 hold37 (.A(net71),
    .Z(net37));
 CLKBUF_X1 hold38 (.A(net78),
    .Z(net38));
 CLKBUF_X1 hold39 (.A(net76),
    .Z(net39));
 CLKBUF_X1 hold40 (.A(net63),
    .Z(net40));
 CLKBUF_X1 hold41 (.A(net74),
    .Z(net41));
 CLKBUF_X1 hold42 (.A(net81),
    .Z(net42));
 CLKBUF_X1 hold43 (.A(net83),
    .Z(net43));
 CLKBUF_X1 hold44 (.A(net84),
    .Z(net44));
 CLKBUF_X1 hold45 (.A(net86),
    .Z(net45));
 CLKBUF_X1 hold46 (.A(net87),
    .Z(net46));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 CLKBUF_X3 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 CLKBUF_X3 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 CLKBUF_X3 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 INV_X2 clkload0 (.A(clknet_2_0__leaf_clk));
 CLKBUF_X1 clkload1 (.A(clknet_2_2__leaf_clk));
 INV_X1 clkload2 (.A(clknet_2_3__leaf_clk));
 CLKBUF_X1 hold1 (.A(_265_),
    .Z(net47));
 CLKBUF_X1 hold2 (.A(_194_),
    .Z(net48));
 CLKBUF_X1 hold3 (.A(_266_),
    .Z(net49));
 CLKBUF_X1 hold4 (.A(_197_),
    .Z(net50));
 CLKBUF_X1 hold5 (.A(net89),
    .Z(net51));
 CLKBUF_X1 hold6 (.A(net88),
    .Z(net52));
 CLKBUF_X1 hold7 (.A(_267_),
    .Z(net53));
 CLKBUF_X1 hold8 (.A(_201_),
    .Z(net54));
 CLKBUF_X1 hold9 (.A(_093_),
    .Z(net55));
 CLKBUF_X1 hold10 (.A(_244_),
    .Z(net56));
 CLKBUF_X1 hold11 (.A(net31),
    .Z(net57));
 CLKBUF_X1 hold12 (.A(_133_),
    .Z(net58));
 CLKBUF_X1 hold13 (.A(net90),
    .Z(net59));
 CLKBUF_X1 hold14 (.A(_268_),
    .Z(net60));
 CLKBUF_X1 hold15 (.A(net32),
    .Z(net61));
 CLKBUF_X1 hold16 (.A(_118_),
    .Z(net62));
 CLKBUF_X1 hold17 (.A(_264_),
    .Z(net63));
 CLKBUF_X1 hold18 (.A(_188_),
    .Z(net64));
 CLKBUF_X1 hold19 (.A(addr_ptr[1]),
    .Z(net65));
 CLKBUF_X1 hold20 (.A(net35),
    .Z(net66));
 CLKBUF_X1 hold21 (.A(addr_ptr[3]),
    .Z(net67));
 CLKBUF_X1 hold22 (.A(net33),
    .Z(net68));
 CLKBUF_X1 hold23 (.A(addr_ptr[2]),
    .Z(net69));
 CLKBUF_X1 hold24 (.A(net36),
    .Z(net70));
 CLKBUF_X1 hold25 (.A(_270_),
    .Z(net71));
 CLKBUF_X1 hold26 (.A(net37),
    .Z(net72));
 CLKBUF_X1 hold27 (.A(_120_),
    .Z(net73));
 CLKBUF_X1 hold28 (.A(addr_ptr[0]),
    .Z(net74));
 CLKBUF_X1 hold29 (.A(net41),
    .Z(net75));
 CLKBUF_X1 hold30 (.A(_271_),
    .Z(net76));
 CLKBUF_X1 hold47 (.A(_121_),
    .Z(net77));
 CLKBUF_X1 hold48 (.A(_269_),
    .Z(net78));
 CLKBUF_X1 hold49 (.A(net38),
    .Z(net79));
 CLKBUF_X1 hold50 (.A(_119_),
    .Z(net80));
 CLKBUF_X1 hold51 (.A(\u_multiplier/LODx/z [7]),
    .Z(net81));
 CLKBUF_X1 hold52 (.A(curr_state[2]),
    .Z(net82));
 CLKBUF_X1 hold53 (.A(data_in_reg[5]),
    .Z(net83));
 CLKBUF_X1 hold54 (.A(data_in_reg[4]),
    .Z(net84));
 CLKBUF_X1 hold55 (.A(curr_state[0]),
    .Z(net85));
 CLKBUF_X1 hold56 (.A(data_in_reg[0]),
    .Z(net86));
 CLKBUF_X1 hold57 (.A(data_in_reg[1]),
    .Z(net87));
 CLKBUF_X1 hold58 (.A(\u_multiplier/LODx/z [3]),
    .Z(net88));
 CLKBUF_X1 hold59 (.A(data_in_reg[2]),
    .Z(net89));
 CLKBUF_X1 hold60 (.A(data_in_reg[6]),
    .Z(net90));
 FILLCELL_X4 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_8 ();
 FILLCELL_X16 FILLER_0_40 ();
 FILLCELL_X8 FILLER_0_56 ();
 FILLCELL_X4 FILLER_0_64 ();
 FILLCELL_X32 FILLER_0_71 ();
 FILLCELL_X32 FILLER_0_103 ();
 FILLCELL_X16 FILLER_0_135 ();
 FILLCELL_X8 FILLER_0_151 ();
 FILLCELL_X2 FILLER_0_159 ();
 FILLCELL_X1 FILLER_0_161 ();
 FILLCELL_X32 FILLER_0_165 ();
 FILLCELL_X32 FILLER_0_197 ();
 FILLCELL_X16 FILLER_0_229 ();
 FILLCELL_X8 FILLER_0_245 ();
 FILLCELL_X2 FILLER_0_253 ();
 FILLCELL_X1 FILLER_0_255 ();
 FILLCELL_X16 FILLER_0_259 ();
 FILLCELL_X8 FILLER_0_275 ();
 FILLCELL_X4 FILLER_0_283 ();
 FILLCELL_X2 FILLER_0_287 ();
 FILLCELL_X1 FILLER_0_289 ();
 FILLCELL_X32 FILLER_0_294 ();
 FILLCELL_X16 FILLER_0_326 ();
 FILLCELL_X8 FILLER_0_342 ();
 FILLCELL_X1 FILLER_0_350 ();
 FILLCELL_X32 FILLER_0_355 ();
 FILLCELL_X32 FILLER_0_387 ();
 FILLCELL_X16 FILLER_0_419 ();
 FILLCELL_X1 FILLER_0_435 ();
 FILLCELL_X4 FILLER_0_440 ();
 FILLCELL_X4 FILLER_0_448 ();
 FILLCELL_X32 FILLER_0_455 ();
 FILLCELL_X32 FILLER_0_487 ();
 FILLCELL_X16 FILLER_0_519 ();
 FILLCELL_X4 FILLER_0_535 ();
 FILLCELL_X32 FILLER_0_542 ();
 FILLCELL_X32 FILLER_0_574 ();
 FILLCELL_X16 FILLER_0_606 ();
 FILLCELL_X8 FILLER_0_622 ();
 FILLCELL_X1 FILLER_0_630 ();
 FILLCELL_X4 FILLER_0_632 ();
 FILLCELL_X16 FILLER_0_639 ();
 FILLCELL_X2 FILLER_0_655 ();
 FILLCELL_X1 FILLER_0_657 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X8 FILLER_1_257 ();
 FILLCELL_X1 FILLER_1_265 ();
 FILLCELL_X4 FILLER_1_270 ();
 FILLCELL_X4 FILLER_1_293 ();
 FILLCELL_X16 FILLER_1_316 ();
 FILLCELL_X1 FILLER_1_332 ();
 FILLCELL_X4 FILLER_1_337 ();
 FILLCELL_X32 FILLER_1_360 ();
 FILLCELL_X16 FILLER_1_392 ();
 FILLCELL_X2 FILLER_1_408 ();
 FILLCELL_X8 FILLER_1_414 ();
 FILLCELL_X4 FILLER_1_422 ();
 FILLCELL_X2 FILLER_1_426 ();
 FILLCELL_X8 FILLER_1_432 ();
 FILLCELL_X2 FILLER_1_440 ();
 FILLCELL_X32 FILLER_1_461 ();
 FILLCELL_X32 FILLER_1_493 ();
 FILLCELL_X32 FILLER_1_525 ();
 FILLCELL_X32 FILLER_1_557 ();
 FILLCELL_X32 FILLER_1_589 ();
 FILLCELL_X32 FILLER_1_621 ();
 FILLCELL_X4 FILLER_1_653 ();
 FILLCELL_X1 FILLER_1_657 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X16 FILLER_2_289 ();
 FILLCELL_X8 FILLER_2_305 ();
 FILLCELL_X4 FILLER_2_317 ();
 FILLCELL_X4 FILLER_2_340 ();
 FILLCELL_X2 FILLER_2_344 ();
 FILLCELL_X1 FILLER_2_346 ();
 FILLCELL_X4 FILLER_2_366 ();
 FILLCELL_X4 FILLER_2_373 ();
 FILLCELL_X16 FILLER_2_380 ();
 FILLCELL_X8 FILLER_2_396 ();
 FILLCELL_X4 FILLER_2_404 ();
 FILLCELL_X4 FILLER_2_427 ();
 FILLCELL_X2 FILLER_2_431 ();
 FILLCELL_X1 FILLER_2_433 ();
 FILLCELL_X4 FILLER_2_453 ();
 FILLCELL_X1 FILLER_2_457 ();
 FILLCELL_X4 FILLER_2_462 ();
 FILLCELL_X32 FILLER_2_469 ();
 FILLCELL_X32 FILLER_2_501 ();
 FILLCELL_X32 FILLER_2_533 ();
 FILLCELL_X16 FILLER_2_565 ();
 FILLCELL_X1 FILLER_2_581 ();
 FILLCELL_X32 FILLER_2_584 ();
 FILLCELL_X8 FILLER_2_616 ();
 FILLCELL_X4 FILLER_2_624 ();
 FILLCELL_X2 FILLER_2_628 ();
 FILLCELL_X1 FILLER_2_630 ();
 FILLCELL_X16 FILLER_2_632 ();
 FILLCELL_X2 FILLER_2_648 ();
 FILLCELL_X1 FILLER_2_650 ();
 FILLCELL_X4 FILLER_2_654 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X16 FILLER_3_257 ();
 FILLCELL_X4 FILLER_3_273 ();
 FILLCELL_X4 FILLER_3_280 ();
 FILLCELL_X8 FILLER_3_288 ();
 FILLCELL_X4 FILLER_3_296 ();
 FILLCELL_X1 FILLER_3_300 ();
 FILLCELL_X4 FILLER_3_320 ();
 FILLCELL_X4 FILLER_3_343 ();
 FILLCELL_X8 FILLER_3_351 ();
 FILLCELL_X4 FILLER_3_362 ();
 FILLCELL_X16 FILLER_3_385 ();
 FILLCELL_X8 FILLER_3_401 ();
 FILLCELL_X8 FILLER_3_412 ();
 FILLCELL_X4 FILLER_3_420 ();
 FILLCELL_X2 FILLER_3_424 ();
 FILLCELL_X8 FILLER_3_445 ();
 FILLCELL_X2 FILLER_3_453 ();
 FILLCELL_X1 FILLER_3_455 ();
 FILLCELL_X32 FILLER_3_475 ();
 FILLCELL_X16 FILLER_3_507 ();
 FILLCELL_X8 FILLER_3_523 ();
 FILLCELL_X8 FILLER_3_533 ();
 FILLCELL_X4 FILLER_3_541 ();
 FILLCELL_X2 FILLER_3_545 ();
 FILLCELL_X16 FILLER_3_549 ();
 FILLCELL_X8 FILLER_3_567 ();
 FILLCELL_X2 FILLER_3_575 ();
 FILLCELL_X1 FILLER_3_577 ();
 FILLCELL_X4 FILLER_3_580 ();
 FILLCELL_X1 FILLER_3_584 ();
 FILLCELL_X32 FILLER_3_588 ();
 FILLCELL_X32 FILLER_3_620 ();
 FILLCELL_X4 FILLER_3_652 ();
 FILLCELL_X2 FILLER_3_656 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X8 FILLER_4_257 ();
 FILLCELL_X4 FILLER_4_265 ();
 FILLCELL_X2 FILLER_4_269 ();
 FILLCELL_X4 FILLER_4_274 ();
 FILLCELL_X4 FILLER_4_297 ();
 FILLCELL_X8 FILLER_4_305 ();
 FILLCELL_X4 FILLER_4_313 ();
 FILLCELL_X2 FILLER_4_317 ();
 FILLCELL_X8 FILLER_4_323 ();
 FILLCELL_X2 FILLER_4_331 ();
 FILLCELL_X1 FILLER_4_333 ();
 FILLCELL_X4 FILLER_4_337 ();
 FILLCELL_X4 FILLER_4_344 ();
 FILLCELL_X4 FILLER_4_352 ();
 FILLCELL_X4 FILLER_4_360 ();
 FILLCELL_X1 FILLER_4_364 ();
 FILLCELL_X4 FILLER_4_368 ();
 FILLCELL_X4 FILLER_4_391 ();
 FILLCELL_X2 FILLER_4_395 ();
 FILLCELL_X16 FILLER_4_400 ();
 FILLCELL_X4 FILLER_4_416 ();
 FILLCELL_X2 FILLER_4_420 ();
 FILLCELL_X4 FILLER_4_425 ();
 FILLCELL_X4 FILLER_4_432 ();
 FILLCELL_X1 FILLER_4_436 ();
 FILLCELL_X8 FILLER_4_440 ();
 FILLCELL_X8 FILLER_4_451 ();
 FILLCELL_X32 FILLER_4_462 ();
 FILLCELL_X16 FILLER_4_494 ();
 FILLCELL_X8 FILLER_4_510 ();
 FILLCELL_X4 FILLER_4_518 ();
 FILLCELL_X1 FILLER_4_522 ();
 FILLCELL_X4 FILLER_4_525 ();
 FILLCELL_X4 FILLER_4_533 ();
 FILLCELL_X8 FILLER_4_543 ();
 FILLCELL_X1 FILLER_4_551 ();
 FILLCELL_X4 FILLER_4_555 ();
 FILLCELL_X2 FILLER_4_559 ();
 FILLCELL_X1 FILLER_4_561 ();
 FILLCELL_X4 FILLER_4_566 ();
 FILLCELL_X4 FILLER_4_575 ();
 FILLCELL_X4 FILLER_4_584 ();
 FILLCELL_X32 FILLER_4_592 ();
 FILLCELL_X4 FILLER_4_624 ();
 FILLCELL_X2 FILLER_4_628 ();
 FILLCELL_X1 FILLER_4_630 ();
 FILLCELL_X16 FILLER_4_632 ();
 FILLCELL_X8 FILLER_4_648 ();
 FILLCELL_X2 FILLER_4_656 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X16 FILLER_5_97 ();
 FILLCELL_X4 FILLER_5_113 ();
 FILLCELL_X1 FILLER_5_117 ();
 FILLCELL_X4 FILLER_5_516 ();
 FILLCELL_X4 FILLER_5_523 ();
 FILLCELL_X4 FILLER_5_534 ();
 FILLCELL_X4 FILLER_5_543 ();
 FILLCELL_X4 FILLER_5_552 ();
 FILLCELL_X16 FILLER_5_560 ();
 FILLCELL_X8 FILLER_5_581 ();
 FILLCELL_X2 FILLER_5_589 ();
 FILLCELL_X1 FILLER_5_591 ();
 FILLCELL_X32 FILLER_5_601 ();
 FILLCELL_X16 FILLER_5_633 ();
 FILLCELL_X8 FILLER_5_649 ();
 FILLCELL_X1 FILLER_5_657 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X16 FILLER_6_97 ();
 FILLCELL_X4 FILLER_6_113 ();
 FILLCELL_X1 FILLER_6_117 ();
 FILLCELL_X8 FILLER_6_516 ();
 FILLCELL_X1 FILLER_6_524 ();
 FILLCELL_X4 FILLER_6_527 ();
 FILLCELL_X4 FILLER_6_536 ();
 FILLCELL_X4 FILLER_6_545 ();
 FILLCELL_X8 FILLER_6_554 ();
 FILLCELL_X2 FILLER_6_562 ();
 FILLCELL_X1 FILLER_6_564 ();
 FILLCELL_X4 FILLER_6_570 ();
 FILLCELL_X4 FILLER_6_584 ();
 FILLCELL_X2 FILLER_6_588 ();
 FILLCELL_X32 FILLER_6_600 ();
 FILLCELL_X16 FILLER_6_632 ();
 FILLCELL_X8 FILLER_6_648 ();
 FILLCELL_X2 FILLER_6_656 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X16 FILLER_7_97 ();
 FILLCELL_X4 FILLER_7_113 ();
 FILLCELL_X1 FILLER_7_117 ();
 FILLCELL_X4 FILLER_7_516 ();
 FILLCELL_X4 FILLER_7_525 ();
 FILLCELL_X8 FILLER_7_531 ();
 FILLCELL_X4 FILLER_7_539 ();
 FILLCELL_X2 FILLER_7_543 ();
 FILLCELL_X8 FILLER_7_554 ();
 FILLCELL_X4 FILLER_7_575 ();
 FILLCELL_X2 FILLER_7_579 ();
 FILLCELL_X4 FILLER_7_591 ();
 FILLCELL_X4 FILLER_7_604 ();
 FILLCELL_X32 FILLER_7_617 ();
 FILLCELL_X8 FILLER_7_649 ();
 FILLCELL_X1 FILLER_7_657 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X16 FILLER_8_97 ();
 FILLCELL_X4 FILLER_8_113 ();
 FILLCELL_X1 FILLER_8_117 ();
 FILLCELL_X4 FILLER_8_516 ();
 FILLCELL_X4 FILLER_8_524 ();
 FILLCELL_X4 FILLER_8_532 ();
 FILLCELL_X8 FILLER_8_538 ();
 FILLCELL_X2 FILLER_8_546 ();
 FILLCELL_X1 FILLER_8_548 ();
 FILLCELL_X4 FILLER_8_562 ();
 FILLCELL_X4 FILLER_8_579 ();
 FILLCELL_X4 FILLER_8_593 ();
 FILLCELL_X8 FILLER_8_606 ();
 FILLCELL_X4 FILLER_8_614 ();
 FILLCELL_X1 FILLER_8_618 ();
 FILLCELL_X4 FILLER_8_621 ();
 FILLCELL_X4 FILLER_8_627 ();
 FILLCELL_X8 FILLER_8_633 ();
 FILLCELL_X4 FILLER_8_641 ();
 FILLCELL_X8 FILLER_8_647 ();
 FILLCELL_X2 FILLER_8_655 ();
 FILLCELL_X1 FILLER_8_657 ();
 FILLCELL_X4 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_8 ();
 FILLCELL_X32 FILLER_9_40 ();
 FILLCELL_X32 FILLER_9_72 ();
 FILLCELL_X8 FILLER_9_104 ();
 FILLCELL_X4 FILLER_9_112 ();
 FILLCELL_X2 FILLER_9_116 ();
 FILLCELL_X4 FILLER_9_516 ();
 FILLCELL_X1 FILLER_9_520 ();
 FILLCELL_X4 FILLER_9_527 ();
 FILLCELL_X1 FILLER_9_531 ();
 FILLCELL_X8 FILLER_9_541 ();
 FILLCELL_X2 FILLER_9_549 ();
 FILLCELL_X1 FILLER_9_551 ();
 FILLCELL_X4 FILLER_9_562 ();
 FILLCELL_X32 FILLER_9_575 ();
 FILLCELL_X4 FILLER_9_607 ();
 FILLCELL_X2 FILLER_9_611 ();
 FILLCELL_X4 FILLER_9_617 ();
 FILLCELL_X4 FILLER_9_626 ();
 FILLCELL_X4 FILLER_9_634 ();
 FILLCELL_X4 FILLER_9_642 ();
 FILLCELL_X8 FILLER_9_649 ();
 FILLCELL_X1 FILLER_9_657 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X16 FILLER_10_97 ();
 FILLCELL_X4 FILLER_10_113 ();
 FILLCELL_X1 FILLER_10_117 ();
 FILLCELL_X4 FILLER_10_516 ();
 FILLCELL_X2 FILLER_10_520 ();
 FILLCELL_X4 FILLER_10_525 ();
 FILLCELL_X16 FILLER_10_539 ();
 FILLCELL_X2 FILLER_10_555 ();
 FILLCELL_X8 FILLER_10_566 ();
 FILLCELL_X4 FILLER_10_574 ();
 FILLCELL_X1 FILLER_10_578 ();
 FILLCELL_X4 FILLER_10_584 ();
 FILLCELL_X4 FILLER_10_595 ();
 FILLCELL_X4 FILLER_10_608 ();
 FILLCELL_X2 FILLER_10_612 ();
 FILLCELL_X1 FILLER_10_614 ();
 FILLCELL_X4 FILLER_10_619 ();
 FILLCELL_X4 FILLER_10_632 ();
 FILLCELL_X4 FILLER_10_653 ();
 FILLCELL_X1 FILLER_10_657 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X16 FILLER_11_97 ();
 FILLCELL_X4 FILLER_11_113 ();
 FILLCELL_X1 FILLER_11_117 ();
 FILLCELL_X8 FILLER_11_516 ();
 FILLCELL_X4 FILLER_11_529 ();
 FILLCELL_X4 FILLER_11_538 ();
 FILLCELL_X2 FILLER_11_542 ();
 FILLCELL_X4 FILLER_11_553 ();
 FILLCELL_X8 FILLER_11_567 ();
 FILLCELL_X4 FILLER_11_575 ();
 FILLCELL_X1 FILLER_11_579 ();
 FILLCELL_X8 FILLER_11_585 ();
 FILLCELL_X2 FILLER_11_593 ();
 FILLCELL_X1 FILLER_11_595 ();
 FILLCELL_X4 FILLER_11_601 ();
 FILLCELL_X4 FILLER_11_614 ();
 FILLCELL_X8 FILLER_11_620 ();
 FILLCELL_X4 FILLER_11_632 ();
 FILLCELL_X4 FILLER_11_640 ();
 FILLCELL_X4 FILLER_11_647 ();
 FILLCELL_X4 FILLER_11_653 ();
 FILLCELL_X1 FILLER_11_657 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X16 FILLER_12_97 ();
 FILLCELL_X4 FILLER_12_113 ();
 FILLCELL_X1 FILLER_12_117 ();
 FILLCELL_X4 FILLER_12_516 ();
 FILLCELL_X4 FILLER_12_522 ();
 FILLCELL_X8 FILLER_12_531 ();
 FILLCELL_X1 FILLER_12_539 ();
 FILLCELL_X8 FILLER_12_550 ();
 FILLCELL_X2 FILLER_12_558 ();
 FILLCELL_X1 FILLER_12_560 ();
 FILLCELL_X4 FILLER_12_563 ();
 FILLCELL_X4 FILLER_12_570 ();
 FILLCELL_X4 FILLER_12_578 ();
 FILLCELL_X4 FILLER_12_587 ();
 FILLCELL_X8 FILLER_12_596 ();
 FILLCELL_X1 FILLER_12_604 ();
 FILLCELL_X8 FILLER_12_614 ();
 FILLCELL_X1 FILLER_12_622 ();
 FILLCELL_X4 FILLER_12_625 ();
 FILLCELL_X4 FILLER_12_633 ();
 FILLCELL_X4 FILLER_12_644 ();
 FILLCELL_X2 FILLER_12_648 ();
 FILLCELL_X1 FILLER_12_650 ();
 FILLCELL_X4 FILLER_12_654 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X16 FILLER_13_97 ();
 FILLCELL_X4 FILLER_13_113 ();
 FILLCELL_X1 FILLER_13_117 ();
 FILLCELL_X8 FILLER_13_516 ();
 FILLCELL_X4 FILLER_13_524 ();
 FILLCELL_X4 FILLER_13_531 ();
 FILLCELL_X4 FILLER_13_537 ();
 FILLCELL_X4 FILLER_13_551 ();
 FILLCELL_X8 FILLER_13_564 ();
 FILLCELL_X1 FILLER_13_572 ();
 FILLCELL_X4 FILLER_13_582 ();
 FILLCELL_X4 FILLER_13_600 ();
 FILLCELL_X2 FILLER_13_604 ();
 FILLCELL_X1 FILLER_13_606 ();
 FILLCELL_X4 FILLER_13_616 ();
 FILLCELL_X2 FILLER_13_620 ();
 FILLCELL_X4 FILLER_13_624 ();
 FILLCELL_X4 FILLER_13_632 ();
 FILLCELL_X1 FILLER_13_636 ();
 FILLCELL_X4 FILLER_13_641 ();
 FILLCELL_X4 FILLER_13_648 ();
 FILLCELL_X4 FILLER_13_654 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X16 FILLER_14_97 ();
 FILLCELL_X4 FILLER_14_113 ();
 FILLCELL_X1 FILLER_14_117 ();
 FILLCELL_X4 FILLER_14_516 ();
 FILLCELL_X16 FILLER_14_522 ();
 FILLCELL_X1 FILLER_14_538 ();
 FILLCELL_X16 FILLER_14_548 ();
 FILLCELL_X2 FILLER_14_564 ();
 FILLCELL_X1 FILLER_14_566 ();
 FILLCELL_X4 FILLER_14_570 ();
 FILLCELL_X4 FILLER_14_585 ();
 FILLCELL_X16 FILLER_14_600 ();
 FILLCELL_X8 FILLER_14_616 ();
 FILLCELL_X4 FILLER_14_624 ();
 FILLCELL_X4 FILLER_14_632 ();
 FILLCELL_X8 FILLER_14_649 ();
 FILLCELL_X1 FILLER_14_657 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X16 FILLER_15_97 ();
 FILLCELL_X4 FILLER_15_113 ();
 FILLCELL_X1 FILLER_15_117 ();
 FILLCELL_X8 FILLER_15_516 ();
 FILLCELL_X4 FILLER_15_529 ();
 FILLCELL_X8 FILLER_15_538 ();
 FILLCELL_X1 FILLER_15_546 ();
 FILLCELL_X32 FILLER_15_557 ();
 FILLCELL_X1 FILLER_15_589 ();
 FILLCELL_X16 FILLER_15_595 ();
 FILLCELL_X8 FILLER_15_611 ();
 FILLCELL_X1 FILLER_15_619 ();
 FILLCELL_X4 FILLER_15_622 ();
 FILLCELL_X4 FILLER_15_633 ();
 FILLCELL_X8 FILLER_15_650 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X16 FILLER_16_97 ();
 FILLCELL_X4 FILLER_16_113 ();
 FILLCELL_X1 FILLER_16_117 ();
 FILLCELL_X4 FILLER_16_516 ();
 FILLCELL_X4 FILLER_16_527 ();
 FILLCELL_X4 FILLER_16_540 ();
 FILLCELL_X8 FILLER_16_557 ();
 FILLCELL_X4 FILLER_16_565 ();
 FILLCELL_X4 FILLER_16_572 ();
 FILLCELL_X2 FILLER_16_576 ();
 FILLCELL_X4 FILLER_16_595 ();
 FILLCELL_X8 FILLER_16_612 ();
 FILLCELL_X4 FILLER_16_620 ();
 FILLCELL_X1 FILLER_16_624 ();
 FILLCELL_X4 FILLER_16_629 ();
 FILLCELL_X4 FILLER_16_646 ();
 FILLCELL_X4 FILLER_16_654 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X16 FILLER_17_97 ();
 FILLCELL_X4 FILLER_17_113 ();
 FILLCELL_X1 FILLER_17_117 ();
 FILLCELL_X4 FILLER_17_516 ();
 FILLCELL_X4 FILLER_17_524 ();
 FILLCELL_X2 FILLER_17_528 ();
 FILLCELL_X1 FILLER_17_530 ();
 FILLCELL_X4 FILLER_17_536 ();
 FILLCELL_X2 FILLER_17_540 ();
 FILLCELL_X4 FILLER_17_555 ();
 FILLCELL_X8 FILLER_17_568 ();
 FILLCELL_X2 FILLER_17_576 ();
 FILLCELL_X4 FILLER_17_595 ();
 FILLCELL_X4 FILLER_17_608 ();
 FILLCELL_X1 FILLER_17_612 ();
 FILLCELL_X4 FILLER_17_622 ();
 FILLCELL_X2 FILLER_17_626 ();
 FILLCELL_X1 FILLER_17_628 ();
 FILLCELL_X4 FILLER_17_634 ();
 FILLCELL_X4 FILLER_17_645 ();
 FILLCELL_X4 FILLER_17_652 ();
 FILLCELL_X2 FILLER_17_656 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X16 FILLER_18_97 ();
 FILLCELL_X4 FILLER_18_113 ();
 FILLCELL_X1 FILLER_18_117 ();
 FILLCELL_X4 FILLER_18_516 ();
 FILLCELL_X1 FILLER_18_520 ();
 FILLCELL_X4 FILLER_18_525 ();
 FILLCELL_X4 FILLER_18_533 ();
 FILLCELL_X4 FILLER_18_550 ();
 FILLCELL_X4 FILLER_18_556 ();
 FILLCELL_X1 FILLER_18_560 ();
 FILLCELL_X4 FILLER_18_568 ();
 FILLCELL_X4 FILLER_18_591 ();
 FILLCELL_X1 FILLER_18_595 ();
 FILLCELL_X4 FILLER_18_605 ();
 FILLCELL_X2 FILLER_18_609 ();
 FILLCELL_X4 FILLER_18_618 ();
 FILLCELL_X4 FILLER_18_629 ();
 FILLCELL_X8 FILLER_18_635 ();
 FILLCELL_X4 FILLER_18_643 ();
 FILLCELL_X8 FILLER_18_649 ();
 FILLCELL_X1 FILLER_18_657 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X16 FILLER_19_97 ();
 FILLCELL_X4 FILLER_19_113 ();
 FILLCELL_X1 FILLER_19_117 ();
 FILLCELL_X4 FILLER_19_516 ();
 FILLCELL_X4 FILLER_19_523 ();
 FILLCELL_X2 FILLER_19_527 ();
 FILLCELL_X1 FILLER_19_529 ();
 FILLCELL_X4 FILLER_19_535 ();
 FILLCELL_X2 FILLER_19_539 ();
 FILLCELL_X1 FILLER_19_541 ();
 FILLCELL_X16 FILLER_19_552 ();
 FILLCELL_X4 FILLER_19_568 ();
 FILLCELL_X16 FILLER_19_579 ();
 FILLCELL_X8 FILLER_19_595 ();
 FILLCELL_X2 FILLER_19_603 ();
 FILLCELL_X4 FILLER_19_614 ();
 FILLCELL_X4 FILLER_19_627 ();
 FILLCELL_X1 FILLER_19_631 ();
 FILLCELL_X4 FILLER_19_636 ();
 FILLCELL_X8 FILLER_19_643 ();
 FILLCELL_X4 FILLER_19_651 ();
 FILLCELL_X2 FILLER_19_655 ();
 FILLCELL_X1 FILLER_19_657 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X16 FILLER_20_97 ();
 FILLCELL_X4 FILLER_20_113 ();
 FILLCELL_X1 FILLER_20_117 ();
 FILLCELL_X4 FILLER_20_516 ();
 FILLCELL_X4 FILLER_20_525 ();
 FILLCELL_X4 FILLER_20_532 ();
 FILLCELL_X1 FILLER_20_536 ();
 FILLCELL_X16 FILLER_20_546 ();
 FILLCELL_X8 FILLER_20_562 ();
 FILLCELL_X4 FILLER_20_570 ();
 FILLCELL_X2 FILLER_20_574 ();
 FILLCELL_X4 FILLER_20_583 ();
 FILLCELL_X8 FILLER_20_594 ();
 FILLCELL_X2 FILLER_20_602 ();
 FILLCELL_X4 FILLER_20_611 ();
 FILLCELL_X8 FILLER_20_624 ();
 FILLCELL_X1 FILLER_20_632 ();
 FILLCELL_X4 FILLER_20_640 ();
 FILLCELL_X4 FILLER_20_651 ();
 FILLCELL_X2 FILLER_20_655 ();
 FILLCELL_X1 FILLER_20_657 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X16 FILLER_21_97 ();
 FILLCELL_X4 FILLER_21_113 ();
 FILLCELL_X1 FILLER_21_117 ();
 FILLCELL_X16 FILLER_21_516 ();
 FILLCELL_X8 FILLER_21_534 ();
 FILLCELL_X2 FILLER_21_542 ();
 FILLCELL_X4 FILLER_21_551 ();
 FILLCELL_X8 FILLER_21_562 ();
 FILLCELL_X4 FILLER_21_577 ();
 FILLCELL_X4 FILLER_21_588 ();
 FILLCELL_X8 FILLER_21_599 ();
 FILLCELL_X4 FILLER_21_607 ();
 FILLCELL_X1 FILLER_21_611 ();
 FILLCELL_X4 FILLER_21_619 ();
 FILLCELL_X2 FILLER_21_623 ();
 FILLCELL_X1 FILLER_21_625 ();
 FILLCELL_X4 FILLER_21_633 ();
 FILLCELL_X4 FILLER_21_644 ();
 FILLCELL_X4 FILLER_21_651 ();
 FILLCELL_X2 FILLER_21_655 ();
 FILLCELL_X1 FILLER_21_657 ();
 FILLCELL_X4 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_9 ();
 FILLCELL_X32 FILLER_22_41 ();
 FILLCELL_X32 FILLER_22_73 ();
 FILLCELL_X8 FILLER_22_105 ();
 FILLCELL_X4 FILLER_22_113 ();
 FILLCELL_X1 FILLER_22_117 ();
 FILLCELL_X16 FILLER_22_516 ();
 FILLCELL_X8 FILLER_22_532 ();
 FILLCELL_X2 FILLER_22_540 ();
 FILLCELL_X4 FILLER_22_549 ();
 FILLCELL_X8 FILLER_22_560 ();
 FILLCELL_X2 FILLER_22_568 ();
 FILLCELL_X4 FILLER_22_573 ();
 FILLCELL_X4 FILLER_22_580 ();
 FILLCELL_X1 FILLER_22_584 ();
 FILLCELL_X4 FILLER_22_592 ();
 FILLCELL_X4 FILLER_22_599 ();
 FILLCELL_X16 FILLER_22_606 ();
 FILLCELL_X4 FILLER_22_622 ();
 FILLCELL_X1 FILLER_22_626 ();
 FILLCELL_X4 FILLER_22_630 ();
 FILLCELL_X4 FILLER_22_637 ();
 FILLCELL_X8 FILLER_22_648 ();
 FILLCELL_X2 FILLER_22_656 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X16 FILLER_23_97 ();
 FILLCELL_X4 FILLER_23_113 ();
 FILLCELL_X1 FILLER_23_117 ();
 FILLCELL_X16 FILLER_23_516 ();
 FILLCELL_X4 FILLER_23_532 ();
 FILLCELL_X2 FILLER_23_536 ();
 FILLCELL_X4 FILLER_23_545 ();
 FILLCELL_X1 FILLER_23_549 ();
 FILLCELL_X4 FILLER_23_557 ();
 FILLCELL_X2 FILLER_23_561 ();
 FILLCELL_X1 FILLER_23_563 ();
 FILLCELL_X4 FILLER_23_571 ();
 FILLCELL_X4 FILLER_23_582 ();
 FILLCELL_X4 FILLER_23_593 ();
 FILLCELL_X8 FILLER_23_606 ();
 FILLCELL_X4 FILLER_23_614 ();
 FILLCELL_X2 FILLER_23_618 ();
 FILLCELL_X1 FILLER_23_620 ();
 FILLCELL_X4 FILLER_23_626 ();
 FILLCELL_X4 FILLER_23_634 ();
 FILLCELL_X4 FILLER_23_640 ();
 FILLCELL_X4 FILLER_23_651 ();
 FILLCELL_X2 FILLER_23_655 ();
 FILLCELL_X1 FILLER_23_657 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X8 FILLER_24_97 ();
 FILLCELL_X4 FILLER_24_105 ();
 FILLCELL_X2 FILLER_24_109 ();
 FILLCELL_X4 FILLER_24_114 ();
 FILLCELL_X4 FILLER_24_516 ();
 FILLCELL_X32 FILLER_24_539 ();
 FILLCELL_X4 FILLER_24_571 ();
 FILLCELL_X2 FILLER_24_575 ();
 FILLCELL_X4 FILLER_24_584 ();
 FILLCELL_X4 FILLER_24_592 ();
 FILLCELL_X16 FILLER_24_599 ();
 FILLCELL_X2 FILLER_24_615 ();
 FILLCELL_X1 FILLER_24_617 ();
 FILLCELL_X4 FILLER_24_622 ();
 FILLCELL_X4 FILLER_24_633 ();
 FILLCELL_X4 FILLER_24_644 ();
 FILLCELL_X4 FILLER_24_651 ();
 FILLCELL_X2 FILLER_24_655 ();
 FILLCELL_X1 FILLER_24_657 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X8 FILLER_25_97 ();
 FILLCELL_X4 FILLER_25_105 ();
 FILLCELL_X4 FILLER_25_114 ();
 FILLCELL_X16 FILLER_25_516 ();
 FILLCELL_X2 FILLER_25_532 ();
 FILLCELL_X1 FILLER_25_534 ();
 FILLCELL_X4 FILLER_25_538 ();
 FILLCELL_X4 FILLER_25_549 ();
 FILLCELL_X4 FILLER_25_560 ();
 FILLCELL_X8 FILLER_25_568 ();
 FILLCELL_X1 FILLER_25_576 ();
 FILLCELL_X4 FILLER_25_580 ();
 FILLCELL_X4 FILLER_25_591 ();
 FILLCELL_X16 FILLER_25_598 ();
 FILLCELL_X1 FILLER_25_614 ();
 FILLCELL_X4 FILLER_25_619 ();
 FILLCELL_X4 FILLER_25_632 ();
 FILLCELL_X4 FILLER_25_640 ();
 FILLCELL_X4 FILLER_25_648 ();
 FILLCELL_X4 FILLER_25_654 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X16 FILLER_26_97 ();
 FILLCELL_X4 FILLER_26_113 ();
 FILLCELL_X1 FILLER_26_117 ();
 FILLCELL_X4 FILLER_26_516 ();
 FILLCELL_X8 FILLER_26_524 ();
 FILLCELL_X4 FILLER_26_532 ();
 FILLCELL_X1 FILLER_26_536 ();
 FILLCELL_X4 FILLER_26_541 ();
 FILLCELL_X1 FILLER_26_545 ();
 FILLCELL_X4 FILLER_26_549 ();
 FILLCELL_X4 FILLER_26_556 ();
 FILLCELL_X4 FILLER_26_563 ();
 FILLCELL_X4 FILLER_26_570 ();
 FILLCELL_X2 FILLER_26_574 ();
 FILLCELL_X1 FILLER_26_576 ();
 FILLCELL_X4 FILLER_26_582 ();
 FILLCELL_X16 FILLER_26_591 ();
 FILLCELL_X8 FILLER_26_607 ();
 FILLCELL_X2 FILLER_26_615 ();
 FILLCELL_X1 FILLER_26_617 ();
 FILLCELL_X4 FILLER_26_627 ();
 FILLCELL_X4 FILLER_26_635 ();
 FILLCELL_X1 FILLER_26_639 ();
 FILLCELL_X8 FILLER_26_643 ();
 FILLCELL_X4 FILLER_26_654 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X16 FILLER_27_97 ();
 FILLCELL_X4 FILLER_27_113 ();
 FILLCELL_X1 FILLER_27_117 ();
 FILLCELL_X16 FILLER_27_516 ();
 FILLCELL_X4 FILLER_27_532 ();
 FILLCELL_X2 FILLER_27_536 ();
 FILLCELL_X4 FILLER_27_541 ();
 FILLCELL_X4 FILLER_27_552 ();
 FILLCELL_X4 FILLER_27_563 ();
 FILLCELL_X4 FILLER_27_574 ();
 FILLCELL_X4 FILLER_27_582 ();
 FILLCELL_X1 FILLER_27_586 ();
 FILLCELL_X4 FILLER_27_596 ();
 FILLCELL_X4 FILLER_27_603 ();
 FILLCELL_X4 FILLER_27_610 ();
 FILLCELL_X4 FILLER_27_619 ();
 FILLCELL_X8 FILLER_27_628 ();
 FILLCELL_X1 FILLER_27_636 ();
 FILLCELL_X4 FILLER_27_642 ();
 FILLCELL_X4 FILLER_27_651 ();
 FILLCELL_X2 FILLER_27_655 ();
 FILLCELL_X1 FILLER_27_657 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X16 FILLER_28_97 ();
 FILLCELL_X4 FILLER_28_113 ();
 FILLCELL_X1 FILLER_28_117 ();
 FILLCELL_X16 FILLER_28_516 ();
 FILLCELL_X4 FILLER_28_532 ();
 FILLCELL_X2 FILLER_28_536 ();
 FILLCELL_X1 FILLER_28_538 ();
 FILLCELL_X4 FILLER_28_545 ();
 FILLCELL_X4 FILLER_28_554 ();
 FILLCELL_X4 FILLER_28_565 ();
 FILLCELL_X2 FILLER_28_569 ();
 FILLCELL_X4 FILLER_28_576 ();
 FILLCELL_X2 FILLER_28_580 ();
 FILLCELL_X4 FILLER_28_591 ();
 FILLCELL_X4 FILLER_28_605 ();
 FILLCELL_X8 FILLER_28_616 ();
 FILLCELL_X2 FILLER_28_624 ();
 FILLCELL_X4 FILLER_28_630 ();
 FILLCELL_X8 FILLER_28_638 ();
 FILLCELL_X4 FILLER_28_651 ();
 FILLCELL_X2 FILLER_28_655 ();
 FILLCELL_X1 FILLER_28_657 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X16 FILLER_29_97 ();
 FILLCELL_X4 FILLER_29_113 ();
 FILLCELL_X1 FILLER_29_117 ();
 FILLCELL_X16 FILLER_29_516 ();
 FILLCELL_X4 FILLER_29_532 ();
 FILLCELL_X2 FILLER_29_536 ();
 FILLCELL_X4 FILLER_29_545 ();
 FILLCELL_X4 FILLER_29_556 ();
 FILLCELL_X4 FILLER_29_563 ();
 FILLCELL_X2 FILLER_29_567 ();
 FILLCELL_X1 FILLER_29_569 ();
 FILLCELL_X8 FILLER_29_574 ();
 FILLCELL_X4 FILLER_29_582 ();
 FILLCELL_X2 FILLER_29_586 ();
 FILLCELL_X1 FILLER_29_588 ();
 FILLCELL_X4 FILLER_29_591 ();
 FILLCELL_X4 FILLER_29_605 ();
 FILLCELL_X2 FILLER_29_609 ();
 FILLCELL_X4 FILLER_29_618 ();
 FILLCELL_X4 FILLER_29_635 ();
 FILLCELL_X4 FILLER_29_646 ();
 FILLCELL_X4 FILLER_29_653 ();
 FILLCELL_X1 FILLER_29_657 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X16 FILLER_30_97 ();
 FILLCELL_X4 FILLER_30_113 ();
 FILLCELL_X1 FILLER_30_117 ();
 FILLCELL_X16 FILLER_30_516 ();
 FILLCELL_X1 FILLER_30_532 ();
 FILLCELL_X4 FILLER_30_542 ();
 FILLCELL_X4 FILLER_30_553 ();
 FILLCELL_X4 FILLER_30_560 ();
 FILLCELL_X16 FILLER_30_567 ();
 FILLCELL_X4 FILLER_30_593 ();
 FILLCELL_X8 FILLER_30_610 ();
 FILLCELL_X4 FILLER_30_625 ();
 FILLCELL_X1 FILLER_30_629 ();
 FILLCELL_X4 FILLER_30_639 ();
 FILLCELL_X4 FILLER_30_652 ();
 FILLCELL_X2 FILLER_30_656 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X16 FILLER_31_97 ();
 FILLCELL_X4 FILLER_31_113 ();
 FILLCELL_X1 FILLER_31_117 ();
 FILLCELL_X4 FILLER_31_516 ();
 FILLCELL_X8 FILLER_31_525 ();
 FILLCELL_X4 FILLER_31_543 ();
 FILLCELL_X4 FILLER_31_554 ();
 FILLCELL_X8 FILLER_31_561 ();
 FILLCELL_X4 FILLER_31_569 ();
 FILLCELL_X2 FILLER_31_573 ();
 FILLCELL_X4 FILLER_31_579 ();
 FILLCELL_X4 FILLER_31_586 ();
 FILLCELL_X4 FILLER_31_593 ();
 FILLCELL_X16 FILLER_31_600 ();
 FILLCELL_X8 FILLER_31_616 ();
 FILLCELL_X1 FILLER_31_624 ();
 FILLCELL_X4 FILLER_31_628 ();
 FILLCELL_X4 FILLER_31_637 ();
 FILLCELL_X4 FILLER_31_646 ();
 FILLCELL_X4 FILLER_31_652 ();
 FILLCELL_X2 FILLER_31_656 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X16 FILLER_32_97 ();
 FILLCELL_X4 FILLER_32_113 ();
 FILLCELL_X1 FILLER_32_117 ();
 FILLCELL_X8 FILLER_32_516 ();
 FILLCELL_X2 FILLER_32_524 ();
 FILLCELL_X4 FILLER_32_531 ();
 FILLCELL_X2 FILLER_32_535 ();
 FILLCELL_X4 FILLER_32_546 ();
 FILLCELL_X4 FILLER_32_553 ();
 FILLCELL_X4 FILLER_32_560 ();
 FILLCELL_X2 FILLER_32_564 ();
 FILLCELL_X4 FILLER_32_573 ();
 FILLCELL_X4 FILLER_32_584 ();
 FILLCELL_X4 FILLER_32_592 ();
 FILLCELL_X16 FILLER_32_600 ();
 FILLCELL_X2 FILLER_32_616 ();
 FILLCELL_X1 FILLER_32_618 ();
 FILLCELL_X4 FILLER_32_622 ();
 FILLCELL_X4 FILLER_32_629 ();
 FILLCELL_X4 FILLER_32_636 ();
 FILLCELL_X4 FILLER_32_647 ();
 FILLCELL_X4 FILLER_32_654 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X16 FILLER_33_97 ();
 FILLCELL_X4 FILLER_33_113 ();
 FILLCELL_X1 FILLER_33_117 ();
 FILLCELL_X16 FILLER_33_516 ();
 FILLCELL_X4 FILLER_33_532 ();
 FILLCELL_X8 FILLER_33_545 ();
 FILLCELL_X4 FILLER_33_562 ();
 FILLCELL_X1 FILLER_33_566 ();
 FILLCELL_X4 FILLER_33_570 ();
 FILLCELL_X4 FILLER_33_581 ();
 FILLCELL_X8 FILLER_33_591 ();
 FILLCELL_X2 FILLER_33_599 ();
 FILLCELL_X1 FILLER_33_601 ();
 FILLCELL_X4 FILLER_33_607 ();
 FILLCELL_X4 FILLER_33_616 ();
 FILLCELL_X8 FILLER_33_624 ();
 FILLCELL_X2 FILLER_33_632 ();
 FILLCELL_X4 FILLER_33_641 ();
 FILLCELL_X8 FILLER_33_650 ();
 FILLCELL_X4 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_9 ();
 FILLCELL_X32 FILLER_34_41 ();
 FILLCELL_X32 FILLER_34_73 ();
 FILLCELL_X8 FILLER_34_105 ();
 FILLCELL_X4 FILLER_34_113 ();
 FILLCELL_X1 FILLER_34_117 ();
 FILLCELL_X4 FILLER_34_516 ();
 FILLCELL_X2 FILLER_34_520 ();
 FILLCELL_X4 FILLER_34_526 ();
 FILLCELL_X8 FILLER_34_534 ();
 FILLCELL_X1 FILLER_34_542 ();
 FILLCELL_X4 FILLER_34_553 ();
 FILLCELL_X4 FILLER_34_559 ();
 FILLCELL_X2 FILLER_34_563 ();
 FILLCELL_X8 FILLER_34_567 ();
 FILLCELL_X4 FILLER_34_582 ();
 FILLCELL_X8 FILLER_34_590 ();
 FILLCELL_X4 FILLER_34_598 ();
 FILLCELL_X2 FILLER_34_602 ();
 FILLCELL_X1 FILLER_34_604 ();
 FILLCELL_X4 FILLER_34_610 ();
 FILLCELL_X2 FILLER_34_614 ();
 FILLCELL_X4 FILLER_34_625 ();
 FILLCELL_X4 FILLER_34_634 ();
 FILLCELL_X4 FILLER_34_642 ();
 FILLCELL_X2 FILLER_34_646 ();
 FILLCELL_X1 FILLER_34_648 ();
 FILLCELL_X4 FILLER_34_654 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X16 FILLER_35_97 ();
 FILLCELL_X4 FILLER_35_113 ();
 FILLCELL_X1 FILLER_35_117 ();
 FILLCELL_X4 FILLER_35_516 ();
 FILLCELL_X4 FILLER_35_525 ();
 FILLCELL_X2 FILLER_35_529 ();
 FILLCELL_X1 FILLER_35_531 ();
 FILLCELL_X4 FILLER_35_537 ();
 FILLCELL_X4 FILLER_35_548 ();
 FILLCELL_X16 FILLER_35_557 ();
 FILLCELL_X4 FILLER_35_573 ();
 FILLCELL_X2 FILLER_35_577 ();
 FILLCELL_X16 FILLER_35_582 ();
 FILLCELL_X8 FILLER_35_598 ();
 FILLCELL_X1 FILLER_35_606 ();
 FILLCELL_X8 FILLER_35_616 ();
 FILLCELL_X1 FILLER_35_624 ();
 FILLCELL_X4 FILLER_35_634 ();
 FILLCELL_X4 FILLER_35_642 ();
 FILLCELL_X8 FILLER_35_650 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X16 FILLER_36_97 ();
 FILLCELL_X4 FILLER_36_113 ();
 FILLCELL_X1 FILLER_36_117 ();
 FILLCELL_X4 FILLER_36_516 ();
 FILLCELL_X16 FILLER_36_522 ();
 FILLCELL_X2 FILLER_36_538 ();
 FILLCELL_X4 FILLER_36_544 ();
 FILLCELL_X4 FILLER_36_552 ();
 FILLCELL_X4 FILLER_36_559 ();
 FILLCELL_X4 FILLER_36_570 ();
 FILLCELL_X4 FILLER_36_579 ();
 FILLCELL_X4 FILLER_36_587 ();
 FILLCELL_X8 FILLER_36_597 ();
 FILLCELL_X4 FILLER_36_605 ();
 FILLCELL_X2 FILLER_36_609 ();
 FILLCELL_X1 FILLER_36_611 ();
 FILLCELL_X4 FILLER_36_619 ();
 FILLCELL_X4 FILLER_36_632 ();
 FILLCELL_X4 FILLER_36_654 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X16 FILLER_37_97 ();
 FILLCELL_X4 FILLER_37_113 ();
 FILLCELL_X1 FILLER_37_117 ();
 FILLCELL_X8 FILLER_37_516 ();
 FILLCELL_X2 FILLER_37_524 ();
 FILLCELL_X4 FILLER_37_530 ();
 FILLCELL_X4 FILLER_37_540 ();
 FILLCELL_X8 FILLER_37_548 ();
 FILLCELL_X2 FILLER_37_556 ();
 FILLCELL_X4 FILLER_37_567 ();
 FILLCELL_X4 FILLER_37_574 ();
 FILLCELL_X1 FILLER_37_578 ();
 FILLCELL_X4 FILLER_37_586 ();
 FILLCELL_X4 FILLER_37_599 ();
 FILLCELL_X8 FILLER_37_607 ();
 FILLCELL_X4 FILLER_37_615 ();
 FILLCELL_X1 FILLER_37_619 ();
 FILLCELL_X4 FILLER_37_627 ();
 FILLCELL_X4 FILLER_37_638 ();
 FILLCELL_X4 FILLER_37_645 ();
 FILLCELL_X1 FILLER_37_649 ();
 FILLCELL_X4 FILLER_37_653 ();
 FILLCELL_X1 FILLER_37_657 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X16 FILLER_38_97 ();
 FILLCELL_X4 FILLER_38_113 ();
 FILLCELL_X1 FILLER_38_117 ();
 FILLCELL_X8 FILLER_38_516 ();
 FILLCELL_X2 FILLER_38_524 ();
 FILLCELL_X1 FILLER_38_526 ();
 FILLCELL_X4 FILLER_38_534 ();
 FILLCELL_X4 FILLER_38_545 ();
 FILLCELL_X4 FILLER_38_554 ();
 FILLCELL_X4 FILLER_38_561 ();
 FILLCELL_X4 FILLER_38_568 ();
 FILLCELL_X1 FILLER_38_572 ();
 FILLCELL_X4 FILLER_38_576 ();
 FILLCELL_X4 FILLER_38_587 ();
 FILLCELL_X1 FILLER_38_591 ();
 FILLCELL_X4 FILLER_38_598 ();
 FILLCELL_X4 FILLER_38_607 ();
 FILLCELL_X4 FILLER_38_616 ();
 FILLCELL_X1 FILLER_38_620 ();
 FILLCELL_X4 FILLER_38_623 ();
 FILLCELL_X4 FILLER_38_630 ();
 FILLCELL_X4 FILLER_38_637 ();
 FILLCELL_X4 FILLER_38_644 ();
 FILLCELL_X4 FILLER_38_652 ();
 FILLCELL_X2 FILLER_38_656 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X8 FILLER_39_97 ();
 FILLCELL_X4 FILLER_39_105 ();
 FILLCELL_X4 FILLER_39_114 ();
 FILLCELL_X32 FILLER_39_516 ();
 FILLCELL_X16 FILLER_39_548 ();
 FILLCELL_X4 FILLER_39_564 ();
 FILLCELL_X2 FILLER_39_568 ();
 FILLCELL_X4 FILLER_39_572 ();
 FILLCELL_X4 FILLER_39_580 ();
 FILLCELL_X2 FILLER_39_584 ();
 FILLCELL_X16 FILLER_39_589 ();
 FILLCELL_X2 FILLER_39_605 ();
 FILLCELL_X8 FILLER_39_610 ();
 FILLCELL_X4 FILLER_39_625 ();
 FILLCELL_X4 FILLER_39_639 ();
 FILLCELL_X2 FILLER_39_643 ();
 FILLCELL_X8 FILLER_39_649 ();
 FILLCELL_X1 FILLER_39_657 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X16 FILLER_40_97 ();
 FILLCELL_X4 FILLER_40_113 ();
 FILLCELL_X1 FILLER_40_117 ();
 FILLCELL_X16 FILLER_40_516 ();
 FILLCELL_X4 FILLER_40_532 ();
 FILLCELL_X1 FILLER_40_536 ();
 FILLCELL_X4 FILLER_40_541 ();
 FILLCELL_X1 FILLER_40_545 ();
 FILLCELL_X4 FILLER_40_551 ();
 FILLCELL_X4 FILLER_40_558 ();
 FILLCELL_X2 FILLER_40_562 ();
 FILLCELL_X4 FILLER_40_568 ();
 FILLCELL_X8 FILLER_40_575 ();
 FILLCELL_X16 FILLER_40_592 ();
 FILLCELL_X8 FILLER_40_608 ();
 FILLCELL_X1 FILLER_40_616 ();
 FILLCELL_X4 FILLER_40_624 ();
 FILLCELL_X4 FILLER_40_634 ();
 FILLCELL_X1 FILLER_40_638 ();
 FILLCELL_X4 FILLER_40_648 ();
 FILLCELL_X4 FILLER_40_654 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X8 FILLER_41_97 ();
 FILLCELL_X4 FILLER_41_105 ();
 FILLCELL_X1 FILLER_41_109 ();
 FILLCELL_X4 FILLER_41_114 ();
 FILLCELL_X16 FILLER_41_516 ();
 FILLCELL_X2 FILLER_41_532 ();
 FILLCELL_X4 FILLER_41_543 ();
 FILLCELL_X4 FILLER_41_556 ();
 FILLCELL_X8 FILLER_41_565 ();
 FILLCELL_X1 FILLER_41_573 ();
 FILLCELL_X4 FILLER_41_577 ();
 FILLCELL_X4 FILLER_41_584 ();
 FILLCELL_X1 FILLER_41_588 ();
 FILLCELL_X4 FILLER_41_598 ();
 FILLCELL_X8 FILLER_41_609 ();
 FILLCELL_X4 FILLER_41_617 ();
 FILLCELL_X2 FILLER_41_621 ();
 FILLCELL_X4 FILLER_41_625 ();
 FILLCELL_X4 FILLER_41_639 ();
 FILLCELL_X4 FILLER_41_648 ();
 FILLCELL_X4 FILLER_41_654 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X16 FILLER_42_65 ();
 FILLCELL_X8 FILLER_42_81 ();
 FILLCELL_X2 FILLER_42_89 ();
 FILLCELL_X1 FILLER_42_91 ();
 FILLCELL_X8 FILLER_42_109 ();
 FILLCELL_X1 FILLER_42_117 ();
 FILLCELL_X8 FILLER_42_516 ();
 FILLCELL_X1 FILLER_42_524 ();
 FILLCELL_X4 FILLER_42_528 ();
 FILLCELL_X4 FILLER_42_539 ();
 FILLCELL_X4 FILLER_42_553 ();
 FILLCELL_X4 FILLER_42_561 ();
 FILLCELL_X4 FILLER_42_569 ();
 FILLCELL_X4 FILLER_42_576 ();
 FILLCELL_X4 FILLER_42_583 ();
 FILLCELL_X4 FILLER_42_593 ();
 FILLCELL_X4 FILLER_42_600 ();
 FILLCELL_X4 FILLER_42_607 ();
 FILLCELL_X8 FILLER_42_613 ();
 FILLCELL_X1 FILLER_42_621 ();
 FILLCELL_X4 FILLER_42_626 ();
 FILLCELL_X4 FILLER_42_643 ();
 FILLCELL_X4 FILLER_42_651 ();
 FILLCELL_X2 FILLER_42_655 ();
 FILLCELL_X1 FILLER_42_657 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X16 FILLER_43_65 ();
 FILLCELL_X4 FILLER_43_81 ();
 FILLCELL_X1 FILLER_43_85 ();
 FILLCELL_X8 FILLER_43_103 ();
 FILLCELL_X4 FILLER_43_111 ();
 FILLCELL_X2 FILLER_43_115 ();
 FILLCELL_X1 FILLER_43_117 ();
 FILLCELL_X8 FILLER_43_516 ();
 FILLCELL_X2 FILLER_43_524 ();
 FILLCELL_X4 FILLER_43_530 ();
 FILLCELL_X4 FILLER_43_541 ();
 FILLCELL_X4 FILLER_43_552 ();
 FILLCELL_X8 FILLER_43_560 ();
 FILLCELL_X4 FILLER_43_575 ();
 FILLCELL_X4 FILLER_43_586 ();
 FILLCELL_X1 FILLER_43_590 ();
 FILLCELL_X4 FILLER_43_596 ();
 FILLCELL_X4 FILLER_43_606 ();
 FILLCELL_X4 FILLER_43_614 ();
 FILLCELL_X1 FILLER_43_618 ();
 FILLCELL_X4 FILLER_43_621 ();
 FILLCELL_X8 FILLER_43_628 ();
 FILLCELL_X1 FILLER_43_636 ();
 FILLCELL_X4 FILLER_43_644 ();
 FILLCELL_X4 FILLER_43_652 ();
 FILLCELL_X2 FILLER_43_656 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X32 FILLER_44_33 ();
 FILLCELL_X16 FILLER_44_65 ();
 FILLCELL_X4 FILLER_44_81 ();
 FILLCELL_X2 FILLER_44_85 ();
 FILLCELL_X1 FILLER_44_87 ();
 FILLCELL_X4 FILLER_44_105 ();
 FILLCELL_X4 FILLER_44_113 ();
 FILLCELL_X1 FILLER_44_117 ();
 FILLCELL_X4 FILLER_44_516 ();
 FILLCELL_X8 FILLER_44_522 ();
 FILLCELL_X4 FILLER_44_534 ();
 FILLCELL_X1 FILLER_44_538 ();
 FILLCELL_X4 FILLER_44_546 ();
 FILLCELL_X16 FILLER_44_554 ();
 FILLCELL_X4 FILLER_44_576 ();
 FILLCELL_X8 FILLER_44_583 ();
 FILLCELL_X2 FILLER_44_591 ();
 FILLCELL_X1 FILLER_44_593 ();
 FILLCELL_X16 FILLER_44_600 ();
 FILLCELL_X2 FILLER_44_616 ();
 FILLCELL_X1 FILLER_44_618 ();
 FILLCELL_X4 FILLER_44_623 ();
 FILLCELL_X4 FILLER_44_629 ();
 FILLCELL_X2 FILLER_44_633 ();
 FILLCELL_X1 FILLER_44_635 ();
 FILLCELL_X4 FILLER_44_640 ();
 FILLCELL_X8 FILLER_44_648 ();
 FILLCELL_X2 FILLER_44_656 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X32 FILLER_45_33 ();
 FILLCELL_X32 FILLER_45_65 ();
 FILLCELL_X4 FILLER_45_97 ();
 FILLCELL_X1 FILLER_45_101 ();
 FILLCELL_X8 FILLER_45_106 ();
 FILLCELL_X4 FILLER_45_114 ();
 FILLCELL_X8 FILLER_45_516 ();
 FILLCELL_X4 FILLER_45_524 ();
 FILLCELL_X2 FILLER_45_528 ();
 FILLCELL_X4 FILLER_45_534 ();
 FILLCELL_X16 FILLER_45_548 ();
 FILLCELL_X4 FILLER_45_564 ();
 FILLCELL_X1 FILLER_45_568 ();
 FILLCELL_X4 FILLER_45_571 ();
 FILLCELL_X8 FILLER_45_584 ();
 FILLCELL_X4 FILLER_45_592 ();
 FILLCELL_X2 FILLER_45_596 ();
 FILLCELL_X1 FILLER_45_598 ();
 FILLCELL_X4 FILLER_45_603 ();
 FILLCELL_X1 FILLER_45_607 ();
 FILLCELL_X4 FILLER_45_618 ();
 FILLCELL_X4 FILLER_45_629 ();
 FILLCELL_X2 FILLER_45_633 ();
 FILLCELL_X1 FILLER_45_635 ();
 FILLCELL_X4 FILLER_45_653 ();
 FILLCELL_X1 FILLER_45_657 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X16 FILLER_46_33 ();
 FILLCELL_X4 FILLER_46_49 ();
 FILLCELL_X2 FILLER_46_53 ();
 FILLCELL_X4 FILLER_46_58 ();
 FILLCELL_X4 FILLER_46_65 ();
 FILLCELL_X32 FILLER_46_73 ();
 FILLCELL_X1 FILLER_46_105 ();
 FILLCELL_X8 FILLER_46_110 ();
 FILLCELL_X16 FILLER_46_516 ();
 FILLCELL_X4 FILLER_46_532 ();
 FILLCELL_X1 FILLER_46_536 ();
 FILLCELL_X16 FILLER_46_541 ();
 FILLCELL_X8 FILLER_46_557 ();
 FILLCELL_X4 FILLER_46_565 ();
 FILLCELL_X2 FILLER_46_569 ();
 FILLCELL_X4 FILLER_46_575 ();
 FILLCELL_X4 FILLER_46_583 ();
 FILLCELL_X4 FILLER_46_590 ();
 FILLCELL_X8 FILLER_46_596 ();
 FILLCELL_X1 FILLER_46_604 ();
 FILLCELL_X4 FILLER_46_607 ();
 FILLCELL_X4 FILLER_46_618 ();
 FILLCELL_X4 FILLER_46_632 ();
 FILLCELL_X16 FILLER_46_639 ();
 FILLCELL_X2 FILLER_46_655 ();
 FILLCELL_X1 FILLER_46_657 ();
 FILLCELL_X4 FILLER_47_1 ();
 FILLCELL_X32 FILLER_47_9 ();
 FILLCELL_X8 FILLER_47_41 ();
 FILLCELL_X4 FILLER_47_52 ();
 FILLCELL_X8 FILLER_47_62 ();
 FILLCELL_X2 FILLER_47_70 ();
 FILLCELL_X4 FILLER_47_89 ();
 FILLCELL_X8 FILLER_47_110 ();
 FILLCELL_X8 FILLER_47_516 ();
 FILLCELL_X2 FILLER_47_524 ();
 FILLCELL_X1 FILLER_47_526 ();
 FILLCELL_X4 FILLER_47_529 ();
 FILLCELL_X4 FILLER_47_537 ();
 FILLCELL_X4 FILLER_47_545 ();
 FILLCELL_X8 FILLER_47_553 ();
 FILLCELL_X1 FILLER_47_561 ();
 FILLCELL_X4 FILLER_47_572 ();
 FILLCELL_X1 FILLER_47_576 ();
 FILLCELL_X4 FILLER_47_583 ();
 FILLCELL_X4 FILLER_47_593 ();
 FILLCELL_X8 FILLER_47_599 ();
 FILLCELL_X2 FILLER_47_607 ();
 FILLCELL_X8 FILLER_47_615 ();
 FILLCELL_X4 FILLER_47_623 ();
 FILLCELL_X2 FILLER_47_627 ();
 FILLCELL_X4 FILLER_47_639 ();
 FILLCELL_X8 FILLER_47_650 ();
 FILLCELL_X32 FILLER_48_1 ();
 FILLCELL_X8 FILLER_48_33 ();
 FILLCELL_X4 FILLER_48_41 ();
 FILLCELL_X2 FILLER_48_45 ();
 FILLCELL_X1 FILLER_48_47 ();
 FILLCELL_X4 FILLER_48_67 ();
 FILLCELL_X2 FILLER_48_71 ();
 FILLCELL_X4 FILLER_48_77 ();
 FILLCELL_X2 FILLER_48_81 ();
 FILLCELL_X1 FILLER_48_83 ();
 FILLCELL_X4 FILLER_48_103 ();
 FILLCELL_X4 FILLER_48_111 ();
 FILLCELL_X2 FILLER_48_115 ();
 FILLCELL_X1 FILLER_48_117 ();
 FILLCELL_X8 FILLER_48_516 ();
 FILLCELL_X4 FILLER_48_524 ();
 FILLCELL_X2 FILLER_48_528 ();
 FILLCELL_X4 FILLER_48_547 ();
 FILLCELL_X4 FILLER_48_561 ();
 FILLCELL_X4 FILLER_48_572 ();
 FILLCELL_X4 FILLER_48_580 ();
 FILLCELL_X4 FILLER_48_587 ();
 FILLCELL_X4 FILLER_48_593 ();
 FILLCELL_X2 FILLER_48_597 ();
 FILLCELL_X1 FILLER_48_599 ();
 FILLCELL_X16 FILLER_48_603 ();
 FILLCELL_X4 FILLER_48_619 ();
 FILLCELL_X8 FILLER_48_626 ();
 FILLCELL_X4 FILLER_48_638 ();
 FILLCELL_X8 FILLER_48_644 ();
 FILLCELL_X4 FILLER_48_652 ();
 FILLCELL_X2 FILLER_48_656 ();
 FILLCELL_X16 FILLER_49_1 ();
 FILLCELL_X8 FILLER_49_17 ();
 FILLCELL_X4 FILLER_49_25 ();
 FILLCELL_X2 FILLER_49_29 ();
 FILLCELL_X1 FILLER_49_31 ();
 FILLCELL_X4 FILLER_49_34 ();
 FILLCELL_X4 FILLER_49_41 ();
 FILLCELL_X4 FILLER_49_64 ();
 FILLCELL_X8 FILLER_49_73 ();
 FILLCELL_X1 FILLER_49_81 ();
 FILLCELL_X4 FILLER_49_86 ();
 FILLCELL_X4 FILLER_49_95 ();
 FILLCELL_X4 FILLER_49_104 ();
 FILLCELL_X2 FILLER_49_108 ();
 FILLCELL_X1 FILLER_49_110 ();
 FILLCELL_X4 FILLER_49_114 ();
 FILLCELL_X8 FILLER_49_516 ();
 FILLCELL_X4 FILLER_49_524 ();
 FILLCELL_X8 FILLER_49_545 ();
 FILLCELL_X2 FILLER_49_553 ();
 FILLCELL_X1 FILLER_49_555 ();
 FILLCELL_X4 FILLER_49_560 ();
 FILLCELL_X4 FILLER_49_570 ();
 FILLCELL_X4 FILLER_49_581 ();
 FILLCELL_X1 FILLER_49_585 ();
 FILLCELL_X4 FILLER_49_588 ();
 FILLCELL_X4 FILLER_49_598 ();
 FILLCELL_X2 FILLER_49_602 ();
 FILLCELL_X1 FILLER_49_604 ();
 FILLCELL_X4 FILLER_49_611 ();
 FILLCELL_X8 FILLER_49_619 ();
 FILLCELL_X1 FILLER_49_627 ();
 FILLCELL_X4 FILLER_49_638 ();
 FILLCELL_X8 FILLER_49_649 ();
 FILLCELL_X1 FILLER_49_657 ();
 FILLCELL_X32 FILLER_50_1 ();
 FILLCELL_X4 FILLER_50_33 ();
 FILLCELL_X2 FILLER_50_37 ();
 FILLCELL_X1 FILLER_50_39 ();
 FILLCELL_X4 FILLER_50_43 ();
 FILLCELL_X4 FILLER_50_50 ();
 FILLCELL_X4 FILLER_50_60 ();
 FILLCELL_X4 FILLER_50_68 ();
 FILLCELL_X4 FILLER_50_75 ();
 FILLCELL_X2 FILLER_50_79 ();
 FILLCELL_X4 FILLER_50_84 ();
 FILLCELL_X4 FILLER_50_91 ();
 FILLCELL_X4 FILLER_50_99 ();
 FILLCELL_X4 FILLER_50_106 ();
 FILLCELL_X4 FILLER_50_113 ();
 FILLCELL_X1 FILLER_50_117 ();
 FILLCELL_X16 FILLER_50_516 ();
 FILLCELL_X4 FILLER_50_532 ();
 FILLCELL_X4 FILLER_50_540 ();
 FILLCELL_X8 FILLER_50_551 ();
 FILLCELL_X4 FILLER_50_559 ();
 FILLCELL_X2 FILLER_50_563 ();
 FILLCELL_X4 FILLER_50_572 ();
 FILLCELL_X4 FILLER_50_578 ();
 FILLCELL_X2 FILLER_50_582 ();
 FILLCELL_X1 FILLER_50_584 ();
 FILLCELL_X4 FILLER_50_587 ();
 FILLCELL_X8 FILLER_50_593 ();
 FILLCELL_X1 FILLER_50_601 ();
 FILLCELL_X4 FILLER_50_605 ();
 FILLCELL_X1 FILLER_50_609 ();
 FILLCELL_X4 FILLER_50_617 ();
 FILLCELL_X2 FILLER_50_621 ();
 FILLCELL_X4 FILLER_50_627 ();
 FILLCELL_X2 FILLER_50_631 ();
 FILLCELL_X1 FILLER_50_633 ();
 FILLCELL_X4 FILLER_50_638 ();
 FILLCELL_X4 FILLER_50_646 ();
 FILLCELL_X4 FILLER_50_652 ();
 FILLCELL_X2 FILLER_50_656 ();
 FILLCELL_X32 FILLER_51_1 ();
 FILLCELL_X8 FILLER_51_33 ();
 FILLCELL_X2 FILLER_51_41 ();
 FILLCELL_X1 FILLER_51_43 ();
 FILLCELL_X4 FILLER_51_47 ();
 FILLCELL_X4 FILLER_51_54 ();
 FILLCELL_X4 FILLER_51_62 ();
 FILLCELL_X16 FILLER_51_69 ();
 FILLCELL_X1 FILLER_51_85 ();
 FILLCELL_X4 FILLER_51_89 ();
 FILLCELL_X8 FILLER_51_97 ();
 FILLCELL_X4 FILLER_51_114 ();
 FILLCELL_X16 FILLER_51_516 ();
 FILLCELL_X4 FILLER_51_532 ();
 FILLCELL_X2 FILLER_51_536 ();
 FILLCELL_X16 FILLER_51_542 ();
 FILLCELL_X2 FILLER_51_558 ();
 FILLCELL_X1 FILLER_51_560 ();
 FILLCELL_X16 FILLER_51_565 ();
 FILLCELL_X4 FILLER_51_585 ();
 FILLCELL_X4 FILLER_51_596 ();
 FILLCELL_X2 FILLER_51_600 ();
 FILLCELL_X4 FILLER_51_606 ();
 FILLCELL_X8 FILLER_51_614 ();
 FILLCELL_X1 FILLER_51_622 ();
 FILLCELL_X8 FILLER_51_627 ();
 FILLCELL_X1 FILLER_51_635 ();
 FILLCELL_X4 FILLER_51_653 ();
 FILLCELL_X1 FILLER_51_657 ();
 FILLCELL_X32 FILLER_52_1 ();
 FILLCELL_X8 FILLER_52_33 ();
 FILLCELL_X4 FILLER_52_41 ();
 FILLCELL_X1 FILLER_52_45 ();
 FILLCELL_X4 FILLER_52_49 ();
 FILLCELL_X4 FILLER_52_57 ();
 FILLCELL_X4 FILLER_52_79 ();
 FILLCELL_X1 FILLER_52_83 ();
 FILLCELL_X4 FILLER_52_103 ();
 FILLCELL_X8 FILLER_52_110 ();
 FILLCELL_X8 FILLER_52_516 ();
 FILLCELL_X4 FILLER_52_524 ();
 FILLCELL_X2 FILLER_52_528 ();
 FILLCELL_X1 FILLER_52_530 ();
 FILLCELL_X8 FILLER_52_548 ();
 FILLCELL_X2 FILLER_52_556 ();
 FILLCELL_X1 FILLER_52_558 ();
 FILLCELL_X16 FILLER_52_563 ();
 FILLCELL_X2 FILLER_52_579 ();
 FILLCELL_X32 FILLER_52_585 ();
 FILLCELL_X2 FILLER_52_617 ();
 FILLCELL_X1 FILLER_52_619 ();
 FILLCELL_X4 FILLER_52_624 ();
 FILLCELL_X4 FILLER_52_632 ();
 FILLCELL_X4 FILLER_52_653 ();
 FILLCELL_X1 FILLER_52_657 ();
 FILLCELL_X32 FILLER_53_1 ();
 FILLCELL_X16 FILLER_53_33 ();
 FILLCELL_X4 FILLER_53_53 ();
 FILLCELL_X4 FILLER_53_63 ();
 FILLCELL_X4 FILLER_53_72 ();
 FILLCELL_X16 FILLER_53_80 ();
 FILLCELL_X1 FILLER_53_96 ();
 FILLCELL_X4 FILLER_53_101 ();
 FILLCELL_X2 FILLER_53_105 ();
 FILLCELL_X8 FILLER_53_110 ();
 FILLCELL_X16 FILLER_53_516 ();
 FILLCELL_X2 FILLER_53_532 ();
 FILLCELL_X1 FILLER_53_534 ();
 FILLCELL_X16 FILLER_53_539 ();
 FILLCELL_X2 FILLER_53_555 ();
 FILLCELL_X8 FILLER_53_561 ();
 FILLCELL_X4 FILLER_53_569 ();
 FILLCELL_X8 FILLER_53_592 ();
 FILLCELL_X2 FILLER_53_600 ();
 FILLCELL_X1 FILLER_53_602 ();
 FILLCELL_X32 FILLER_53_607 ();
 FILLCELL_X16 FILLER_53_639 ();
 FILLCELL_X2 FILLER_53_655 ();
 FILLCELL_X1 FILLER_53_657 ();
 FILLCELL_X32 FILLER_54_1 ();
 FILLCELL_X4 FILLER_54_33 ();
 FILLCELL_X2 FILLER_54_37 ();
 FILLCELL_X1 FILLER_54_39 ();
 FILLCELL_X4 FILLER_54_43 ();
 FILLCELL_X4 FILLER_54_66 ();
 FILLCELL_X4 FILLER_54_81 ();
 FILLCELL_X1 FILLER_54_85 ();
 FILLCELL_X4 FILLER_54_89 ();
 FILLCELL_X4 FILLER_54_97 ();
 FILLCELL_X4 FILLER_54_106 ();
 FILLCELL_X4 FILLER_54_114 ();
 FILLCELL_X8 FILLER_54_516 ();
 FILLCELL_X4 FILLER_54_524 ();
 FILLCELL_X2 FILLER_54_528 ();
 FILLCELL_X1 FILLER_54_530 ();
 FILLCELL_X4 FILLER_54_548 ();
 FILLCELL_X2 FILLER_54_552 ();
 FILLCELL_X1 FILLER_54_554 ();
 FILLCELL_X4 FILLER_54_572 ();
 FILLCELL_X2 FILLER_54_576 ();
 FILLCELL_X32 FILLER_54_582 ();
 FILLCELL_X4 FILLER_54_614 ();
 FILLCELL_X2 FILLER_54_618 ();
 FILLCELL_X16 FILLER_54_637 ();
 FILLCELL_X4 FILLER_54_653 ();
 FILLCELL_X1 FILLER_54_657 ();
 FILLCELL_X32 FILLER_55_1 ();
 FILLCELL_X4 FILLER_55_33 ();
 FILLCELL_X2 FILLER_55_37 ();
 FILLCELL_X1 FILLER_55_39 ();
 FILLCELL_X4 FILLER_55_43 ();
 FILLCELL_X4 FILLER_55_66 ();
 FILLCELL_X4 FILLER_55_73 ();
 FILLCELL_X4 FILLER_55_81 ();
 FILLCELL_X4 FILLER_55_87 ();
 FILLCELL_X4 FILLER_55_98 ();
 FILLCELL_X4 FILLER_55_108 ();
 FILLCELL_X4 FILLER_55_114 ();
 FILLCELL_X32 FILLER_55_516 ();
 FILLCELL_X32 FILLER_55_548 ();
 FILLCELL_X16 FILLER_55_580 ();
 FILLCELL_X4 FILLER_55_596 ();
 FILLCELL_X2 FILLER_55_600 ();
 FILLCELL_X32 FILLER_55_619 ();
 FILLCELL_X4 FILLER_55_651 ();
 FILLCELL_X2 FILLER_55_655 ();
 FILLCELL_X1 FILLER_55_657 ();
 FILLCELL_X32 FILLER_56_1 ();
 FILLCELL_X8 FILLER_56_33 ();
 FILLCELL_X2 FILLER_56_41 ();
 FILLCELL_X4 FILLER_56_46 ();
 FILLCELL_X4 FILLER_56_53 ();
 FILLCELL_X4 FILLER_56_62 ();
 FILLCELL_X1 FILLER_56_66 ();
 FILLCELL_X4 FILLER_56_70 ();
 FILLCELL_X4 FILLER_56_80 ();
 FILLCELL_X8 FILLER_56_88 ();
 FILLCELL_X4 FILLER_56_113 ();
 FILLCELL_X1 FILLER_56_117 ();
 FILLCELL_X32 FILLER_56_516 ();
 FILLCELL_X32 FILLER_56_548 ();
 FILLCELL_X32 FILLER_56_580 ();
 FILLCELL_X32 FILLER_56_612 ();
 FILLCELL_X8 FILLER_56_644 ();
 FILLCELL_X4 FILLER_56_652 ();
 FILLCELL_X2 FILLER_56_656 ();
 FILLCELL_X32 FILLER_57_1 ();
 FILLCELL_X16 FILLER_57_33 ();
 FILLCELL_X1 FILLER_57_49 ();
 FILLCELL_X4 FILLER_57_53 ();
 FILLCELL_X4 FILLER_57_60 ();
 FILLCELL_X8 FILLER_57_83 ();
 FILLCELL_X1 FILLER_57_91 ();
 FILLCELL_X4 FILLER_57_96 ();
 FILLCELL_X4 FILLER_57_104 ();
 FILLCELL_X2 FILLER_57_108 ();
 FILLCELL_X1 FILLER_57_110 ();
 FILLCELL_X4 FILLER_57_114 ();
 FILLCELL_X32 FILLER_57_516 ();
 FILLCELL_X32 FILLER_57_548 ();
 FILLCELL_X32 FILLER_57_580 ();
 FILLCELL_X32 FILLER_57_612 ();
 FILLCELL_X8 FILLER_57_644 ();
 FILLCELL_X4 FILLER_57_652 ();
 FILLCELL_X2 FILLER_57_656 ();
 FILLCELL_X32 FILLER_58_1 ();
 FILLCELL_X16 FILLER_58_33 ();
 FILLCELL_X8 FILLER_58_49 ();
 FILLCELL_X1 FILLER_58_57 ();
 FILLCELL_X4 FILLER_58_61 ();
 FILLCELL_X4 FILLER_58_68 ();
 FILLCELL_X2 FILLER_58_72 ();
 FILLCELL_X1 FILLER_58_74 ();
 FILLCELL_X4 FILLER_58_78 ();
 FILLCELL_X4 FILLER_58_86 ();
 FILLCELL_X4 FILLER_58_94 ();
 FILLCELL_X8 FILLER_58_102 ();
 FILLCELL_X4 FILLER_58_114 ();
 FILLCELL_X32 FILLER_58_516 ();
 FILLCELL_X32 FILLER_58_548 ();
 FILLCELL_X32 FILLER_58_580 ();
 FILLCELL_X32 FILLER_58_612 ();
 FILLCELL_X8 FILLER_58_644 ();
 FILLCELL_X4 FILLER_58_652 ();
 FILLCELL_X2 FILLER_58_656 ();
 FILLCELL_X32 FILLER_59_1 ();
 FILLCELL_X32 FILLER_59_33 ();
 FILLCELL_X1 FILLER_59_65 ();
 FILLCELL_X4 FILLER_59_69 ();
 FILLCELL_X2 FILLER_59_73 ();
 FILLCELL_X4 FILLER_59_79 ();
 FILLCELL_X4 FILLER_59_100 ();
 FILLCELL_X8 FILLER_59_109 ();
 FILLCELL_X1 FILLER_59_117 ();
 FILLCELL_X32 FILLER_59_516 ();
 FILLCELL_X32 FILLER_59_548 ();
 FILLCELL_X32 FILLER_59_580 ();
 FILLCELL_X32 FILLER_59_612 ();
 FILLCELL_X8 FILLER_59_644 ();
 FILLCELL_X4 FILLER_59_652 ();
 FILLCELL_X2 FILLER_59_656 ();
 FILLCELL_X4 FILLER_60_1 ();
 FILLCELL_X32 FILLER_60_8 ();
 FILLCELL_X32 FILLER_60_40 ();
 FILLCELL_X4 FILLER_60_75 ();
 FILLCELL_X4 FILLER_60_82 ();
 FILLCELL_X4 FILLER_60_103 ();
 FILLCELL_X4 FILLER_60_113 ();
 FILLCELL_X1 FILLER_60_117 ();
 FILLCELL_X32 FILLER_60_516 ();
 FILLCELL_X32 FILLER_60_548 ();
 FILLCELL_X32 FILLER_60_580 ();
 FILLCELL_X32 FILLER_60_612 ();
 FILLCELL_X8 FILLER_60_644 ();
 FILLCELL_X4 FILLER_60_652 ();
 FILLCELL_X2 FILLER_60_656 ();
 FILLCELL_X32 FILLER_61_1 ();
 FILLCELL_X32 FILLER_61_33 ();
 FILLCELL_X8 FILLER_61_65 ();
 FILLCELL_X4 FILLER_61_73 ();
 FILLCELL_X2 FILLER_61_77 ();
 FILLCELL_X1 FILLER_61_79 ();
 FILLCELL_X8 FILLER_61_83 ();
 FILLCELL_X4 FILLER_61_94 ();
 FILLCELL_X4 FILLER_61_104 ();
 FILLCELL_X4 FILLER_61_111 ();
 FILLCELL_X2 FILLER_61_115 ();
 FILLCELL_X1 FILLER_61_117 ();
 FILLCELL_X32 FILLER_61_516 ();
 FILLCELL_X32 FILLER_61_548 ();
 FILLCELL_X32 FILLER_61_580 ();
 FILLCELL_X32 FILLER_61_612 ();
 FILLCELL_X8 FILLER_61_644 ();
 FILLCELL_X4 FILLER_61_652 ();
 FILLCELL_X2 FILLER_61_656 ();
 FILLCELL_X32 FILLER_62_1 ();
 FILLCELL_X32 FILLER_62_33 ();
 FILLCELL_X16 FILLER_62_65 ();
 FILLCELL_X8 FILLER_62_81 ();
 FILLCELL_X4 FILLER_62_89 ();
 FILLCELL_X2 FILLER_62_93 ();
 FILLCELL_X1 FILLER_62_95 ();
 FILLCELL_X4 FILLER_62_99 ();
 FILLCELL_X1 FILLER_62_103 ();
 FILLCELL_X4 FILLER_62_107 ();
 FILLCELL_X4 FILLER_62_114 ();
 FILLCELL_X32 FILLER_62_516 ();
 FILLCELL_X32 FILLER_62_548 ();
 FILLCELL_X32 FILLER_62_580 ();
 FILLCELL_X32 FILLER_62_612 ();
 FILLCELL_X8 FILLER_62_644 ();
 FILLCELL_X4 FILLER_62_652 ();
 FILLCELL_X2 FILLER_62_656 ();
 FILLCELL_X32 FILLER_63_1 ();
 FILLCELL_X32 FILLER_63_33 ();
 FILLCELL_X32 FILLER_63_65 ();
 FILLCELL_X4 FILLER_63_100 ();
 FILLCELL_X4 FILLER_63_107 ();
 FILLCELL_X4 FILLER_63_114 ();
 FILLCELL_X32 FILLER_63_516 ();
 FILLCELL_X32 FILLER_63_548 ();
 FILLCELL_X32 FILLER_63_580 ();
 FILLCELL_X32 FILLER_63_612 ();
 FILLCELL_X8 FILLER_63_644 ();
 FILLCELL_X4 FILLER_63_652 ();
 FILLCELL_X2 FILLER_63_656 ();
 FILLCELL_X32 FILLER_64_1 ();
 FILLCELL_X32 FILLER_64_33 ();
 FILLCELL_X32 FILLER_64_65 ();
 FILLCELL_X8 FILLER_64_97 ();
 FILLCELL_X1 FILLER_64_105 ();
 FILLCELL_X8 FILLER_64_109 ();
 FILLCELL_X1 FILLER_64_117 ();
 FILLCELL_X32 FILLER_64_516 ();
 FILLCELL_X32 FILLER_64_548 ();
 FILLCELL_X32 FILLER_64_580 ();
 FILLCELL_X32 FILLER_64_612 ();
 FILLCELL_X8 FILLER_64_644 ();
 FILLCELL_X4 FILLER_64_652 ();
 FILLCELL_X2 FILLER_64_656 ();
 FILLCELL_X32 FILLER_65_1 ();
 FILLCELL_X32 FILLER_65_33 ();
 FILLCELL_X32 FILLER_65_65 ();
 FILLCELL_X4 FILLER_65_97 ();
 FILLCELL_X2 FILLER_65_101 ();
 FILLCELL_X1 FILLER_65_103 ();
 FILLCELL_X4 FILLER_65_107 ();
 FILLCELL_X4 FILLER_65_114 ();
 FILLCELL_X32 FILLER_65_516 ();
 FILLCELL_X32 FILLER_65_548 ();
 FILLCELL_X32 FILLER_65_580 ();
 FILLCELL_X32 FILLER_65_612 ();
 FILLCELL_X8 FILLER_65_644 ();
 FILLCELL_X4 FILLER_65_652 ();
 FILLCELL_X2 FILLER_65_656 ();
 FILLCELL_X32 FILLER_66_1 ();
 FILLCELL_X32 FILLER_66_33 ();
 FILLCELL_X32 FILLER_66_65 ();
 FILLCELL_X16 FILLER_66_97 ();
 FILLCELL_X4 FILLER_66_113 ();
 FILLCELL_X1 FILLER_66_117 ();
 FILLCELL_X32 FILLER_66_516 ();
 FILLCELL_X32 FILLER_66_548 ();
 FILLCELL_X32 FILLER_66_580 ();
 FILLCELL_X32 FILLER_66_612 ();
 FILLCELL_X4 FILLER_66_644 ();
 FILLCELL_X2 FILLER_66_648 ();
 FILLCELL_X1 FILLER_66_650 ();
 FILLCELL_X4 FILLER_66_654 ();
 FILLCELL_X32 FILLER_67_1 ();
 FILLCELL_X32 FILLER_67_33 ();
 FILLCELL_X32 FILLER_67_65 ();
 FILLCELL_X8 FILLER_67_97 ();
 FILLCELL_X4 FILLER_67_105 ();
 FILLCELL_X2 FILLER_67_109 ();
 FILLCELL_X4 FILLER_67_114 ();
 FILLCELL_X32 FILLER_67_516 ();
 FILLCELL_X32 FILLER_67_548 ();
 FILLCELL_X32 FILLER_67_580 ();
 FILLCELL_X32 FILLER_67_612 ();
 FILLCELL_X8 FILLER_67_644 ();
 FILLCELL_X4 FILLER_67_652 ();
 FILLCELL_X2 FILLER_67_656 ();
 FILLCELL_X32 FILLER_68_1 ();
 FILLCELL_X32 FILLER_68_33 ();
 FILLCELL_X32 FILLER_68_65 ();
 FILLCELL_X16 FILLER_68_97 ();
 FILLCELL_X4 FILLER_68_113 ();
 FILLCELL_X1 FILLER_68_117 ();
 FILLCELL_X32 FILLER_68_516 ();
 FILLCELL_X32 FILLER_68_548 ();
 FILLCELL_X32 FILLER_68_580 ();
 FILLCELL_X32 FILLER_68_612 ();
 FILLCELL_X8 FILLER_68_644 ();
 FILLCELL_X4 FILLER_68_652 ();
 FILLCELL_X2 FILLER_68_656 ();
 FILLCELL_X32 FILLER_69_1 ();
 FILLCELL_X32 FILLER_69_33 ();
 FILLCELL_X32 FILLER_69_65 ();
 FILLCELL_X8 FILLER_69_97 ();
 FILLCELL_X4 FILLER_69_105 ();
 FILLCELL_X2 FILLER_69_109 ();
 FILLCELL_X4 FILLER_69_114 ();
 FILLCELL_X32 FILLER_69_516 ();
 FILLCELL_X32 FILLER_69_548 ();
 FILLCELL_X32 FILLER_69_580 ();
 FILLCELL_X32 FILLER_69_612 ();
 FILLCELL_X8 FILLER_69_644 ();
 FILLCELL_X4 FILLER_69_652 ();
 FILLCELL_X2 FILLER_69_656 ();
 FILLCELL_X32 FILLER_70_1 ();
 FILLCELL_X32 FILLER_70_33 ();
 FILLCELL_X32 FILLER_70_65 ();
 FILLCELL_X16 FILLER_70_97 ();
 FILLCELL_X4 FILLER_70_113 ();
 FILLCELL_X1 FILLER_70_117 ();
 FILLCELL_X32 FILLER_70_516 ();
 FILLCELL_X32 FILLER_70_548 ();
 FILLCELL_X32 FILLER_70_580 ();
 FILLCELL_X32 FILLER_70_612 ();
 FILLCELL_X8 FILLER_70_644 ();
 FILLCELL_X4 FILLER_70_652 ();
 FILLCELL_X2 FILLER_70_656 ();
 FILLCELL_X32 FILLER_71_1 ();
 FILLCELL_X32 FILLER_71_33 ();
 FILLCELL_X32 FILLER_71_65 ();
 FILLCELL_X16 FILLER_71_97 ();
 FILLCELL_X4 FILLER_71_113 ();
 FILLCELL_X1 FILLER_71_117 ();
 FILLCELL_X32 FILLER_71_516 ();
 FILLCELL_X32 FILLER_71_548 ();
 FILLCELL_X32 FILLER_71_580 ();
 FILLCELL_X32 FILLER_71_612 ();
 FILLCELL_X8 FILLER_71_644 ();
 FILLCELL_X4 FILLER_71_652 ();
 FILLCELL_X2 FILLER_71_656 ();
 FILLCELL_X32 FILLER_72_1 ();
 FILLCELL_X32 FILLER_72_33 ();
 FILLCELL_X32 FILLER_72_65 ();
 FILLCELL_X8 FILLER_72_97 ();
 FILLCELL_X4 FILLER_72_105 ();
 FILLCELL_X2 FILLER_72_109 ();
 FILLCELL_X4 FILLER_72_114 ();
 FILLCELL_X32 FILLER_72_516 ();
 FILLCELL_X32 FILLER_72_548 ();
 FILLCELL_X32 FILLER_72_580 ();
 FILLCELL_X32 FILLER_72_612 ();
 FILLCELL_X8 FILLER_72_644 ();
 FILLCELL_X4 FILLER_72_652 ();
 FILLCELL_X2 FILLER_72_656 ();
 FILLCELL_X4 FILLER_73_1 ();
 FILLCELL_X32 FILLER_73_9 ();
 FILLCELL_X32 FILLER_73_41 ();
 FILLCELL_X32 FILLER_73_73 ();
 FILLCELL_X4 FILLER_73_105 ();
 FILLCELL_X2 FILLER_73_109 ();
 FILLCELL_X4 FILLER_73_114 ();
 FILLCELL_X32 FILLER_73_516 ();
 FILLCELL_X32 FILLER_73_548 ();
 FILLCELL_X32 FILLER_73_580 ();
 FILLCELL_X32 FILLER_73_612 ();
 FILLCELL_X8 FILLER_73_644 ();
 FILLCELL_X4 FILLER_73_652 ();
 FILLCELL_X2 FILLER_73_656 ();
 FILLCELL_X32 FILLER_74_1 ();
 FILLCELL_X32 FILLER_74_33 ();
 FILLCELL_X32 FILLER_74_65 ();
 FILLCELL_X16 FILLER_74_97 ();
 FILLCELL_X4 FILLER_74_113 ();
 FILLCELL_X1 FILLER_74_117 ();
 FILLCELL_X32 FILLER_74_516 ();
 FILLCELL_X32 FILLER_74_548 ();
 FILLCELL_X32 FILLER_74_580 ();
 FILLCELL_X32 FILLER_74_612 ();
 FILLCELL_X8 FILLER_74_644 ();
 FILLCELL_X4 FILLER_74_652 ();
 FILLCELL_X2 FILLER_74_656 ();
 FILLCELL_X32 FILLER_75_1 ();
 FILLCELL_X32 FILLER_75_33 ();
 FILLCELL_X32 FILLER_75_65 ();
 FILLCELL_X16 FILLER_75_97 ();
 FILLCELL_X4 FILLER_75_113 ();
 FILLCELL_X1 FILLER_75_117 ();
 FILLCELL_X32 FILLER_75_516 ();
 FILLCELL_X32 FILLER_75_548 ();
 FILLCELL_X32 FILLER_75_580 ();
 FILLCELL_X32 FILLER_75_612 ();
 FILLCELL_X8 FILLER_75_644 ();
 FILLCELL_X4 FILLER_75_652 ();
 FILLCELL_X2 FILLER_75_656 ();
 FILLCELL_X32 FILLER_76_1 ();
 FILLCELL_X32 FILLER_76_33 ();
 FILLCELL_X32 FILLER_76_65 ();
 FILLCELL_X16 FILLER_76_97 ();
 FILLCELL_X4 FILLER_76_113 ();
 FILLCELL_X1 FILLER_76_117 ();
 FILLCELL_X32 FILLER_76_516 ();
 FILLCELL_X32 FILLER_76_548 ();
 FILLCELL_X32 FILLER_76_580 ();
 FILLCELL_X32 FILLER_76_612 ();
 FILLCELL_X8 FILLER_76_644 ();
 FILLCELL_X4 FILLER_76_652 ();
 FILLCELL_X2 FILLER_76_656 ();
 FILLCELL_X32 FILLER_77_1 ();
 FILLCELL_X32 FILLER_77_33 ();
 FILLCELL_X32 FILLER_77_65 ();
 FILLCELL_X16 FILLER_77_97 ();
 FILLCELL_X4 FILLER_77_113 ();
 FILLCELL_X1 FILLER_77_117 ();
 FILLCELL_X32 FILLER_77_516 ();
 FILLCELL_X32 FILLER_77_548 ();
 FILLCELL_X32 FILLER_77_580 ();
 FILLCELL_X32 FILLER_77_612 ();
 FILLCELL_X8 FILLER_77_644 ();
 FILLCELL_X4 FILLER_77_652 ();
 FILLCELL_X2 FILLER_77_656 ();
 FILLCELL_X32 FILLER_78_1 ();
 FILLCELL_X32 FILLER_78_33 ();
 FILLCELL_X32 FILLER_78_65 ();
 FILLCELL_X16 FILLER_78_97 ();
 FILLCELL_X4 FILLER_78_113 ();
 FILLCELL_X1 FILLER_78_117 ();
 FILLCELL_X32 FILLER_78_516 ();
 FILLCELL_X32 FILLER_78_548 ();
 FILLCELL_X32 FILLER_78_580 ();
 FILLCELL_X32 FILLER_78_612 ();
 FILLCELL_X8 FILLER_78_644 ();
 FILLCELL_X4 FILLER_78_652 ();
 FILLCELL_X2 FILLER_78_656 ();
 FILLCELL_X32 FILLER_79_1 ();
 FILLCELL_X32 FILLER_79_33 ();
 FILLCELL_X32 FILLER_79_65 ();
 FILLCELL_X32 FILLER_79_97 ();
 FILLCELL_X32 FILLER_79_129 ();
 FILLCELL_X32 FILLER_79_161 ();
 FILLCELL_X32 FILLER_79_193 ();
 FILLCELL_X32 FILLER_79_225 ();
 FILLCELL_X32 FILLER_79_257 ();
 FILLCELL_X32 FILLER_79_289 ();
 FILLCELL_X32 FILLER_79_321 ();
 FILLCELL_X32 FILLER_79_353 ();
 FILLCELL_X32 FILLER_79_385 ();
 FILLCELL_X32 FILLER_79_417 ();
 FILLCELL_X32 FILLER_79_449 ();
 FILLCELL_X32 FILLER_79_481 ();
 FILLCELL_X32 FILLER_79_513 ();
 FILLCELL_X32 FILLER_79_545 ();
 FILLCELL_X32 FILLER_79_577 ();
 FILLCELL_X16 FILLER_79_609 ();
 FILLCELL_X4 FILLER_79_625 ();
 FILLCELL_X2 FILLER_79_629 ();
 FILLCELL_X16 FILLER_79_632 ();
 FILLCELL_X2 FILLER_79_648 ();
 FILLCELL_X1 FILLER_79_650 ();
 FILLCELL_X4 FILLER_79_654 ();
 FILLCELL_X32 FILLER_80_1 ();
 FILLCELL_X32 FILLER_80_33 ();
 FILLCELL_X32 FILLER_80_65 ();
 FILLCELL_X32 FILLER_80_97 ();
 FILLCELL_X32 FILLER_80_129 ();
 FILLCELL_X32 FILLER_80_161 ();
 FILLCELL_X32 FILLER_80_193 ();
 FILLCELL_X32 FILLER_80_225 ();
 FILLCELL_X32 FILLER_80_257 ();
 FILLCELL_X32 FILLER_80_289 ();
 FILLCELL_X32 FILLER_80_321 ();
 FILLCELL_X32 FILLER_80_353 ();
 FILLCELL_X32 FILLER_80_385 ();
 FILLCELL_X32 FILLER_80_417 ();
 FILLCELL_X32 FILLER_80_449 ();
 FILLCELL_X32 FILLER_80_481 ();
 FILLCELL_X32 FILLER_80_513 ();
 FILLCELL_X32 FILLER_80_545 ();
 FILLCELL_X32 FILLER_80_577 ();
 FILLCELL_X16 FILLER_80_609 ();
 FILLCELL_X4 FILLER_80_625 ();
 FILLCELL_X2 FILLER_80_629 ();
 FILLCELL_X16 FILLER_80_632 ();
 FILLCELL_X8 FILLER_80_648 ();
 FILLCELL_X2 FILLER_80_656 ();
 FILLCELL_X32 FILLER_81_1 ();
 FILLCELL_X32 FILLER_81_33 ();
 FILLCELL_X32 FILLER_81_65 ();
 FILLCELL_X32 FILLER_81_97 ();
 FILLCELL_X32 FILLER_81_129 ();
 FILLCELL_X32 FILLER_81_161 ();
 FILLCELL_X32 FILLER_81_193 ();
 FILLCELL_X32 FILLER_81_225 ();
 FILLCELL_X32 FILLER_81_257 ();
 FILLCELL_X32 FILLER_81_289 ();
 FILLCELL_X32 FILLER_81_321 ();
 FILLCELL_X32 FILLER_81_353 ();
 FILLCELL_X32 FILLER_81_385 ();
 FILLCELL_X32 FILLER_81_417 ();
 FILLCELL_X32 FILLER_81_449 ();
 FILLCELL_X32 FILLER_81_481 ();
 FILLCELL_X32 FILLER_81_513 ();
 FILLCELL_X32 FILLER_81_545 ();
 FILLCELL_X32 FILLER_81_577 ();
 FILLCELL_X32 FILLER_81_609 ();
 FILLCELL_X16 FILLER_81_641 ();
 FILLCELL_X1 FILLER_81_657 ();
 FILLCELL_X32 FILLER_82_1 ();
 FILLCELL_X32 FILLER_82_33 ();
 FILLCELL_X32 FILLER_82_65 ();
 FILLCELL_X32 FILLER_82_97 ();
 FILLCELL_X32 FILLER_82_129 ();
 FILLCELL_X32 FILLER_82_161 ();
 FILLCELL_X32 FILLER_82_193 ();
 FILLCELL_X32 FILLER_82_225 ();
 FILLCELL_X32 FILLER_82_257 ();
 FILLCELL_X32 FILLER_82_289 ();
 FILLCELL_X32 FILLER_82_321 ();
 FILLCELL_X32 FILLER_82_353 ();
 FILLCELL_X32 FILLER_82_385 ();
 FILLCELL_X32 FILLER_82_417 ();
 FILLCELL_X32 FILLER_82_449 ();
 FILLCELL_X32 FILLER_82_481 ();
 FILLCELL_X32 FILLER_82_513 ();
 FILLCELL_X32 FILLER_82_545 ();
 FILLCELL_X32 FILLER_82_577 ();
 FILLCELL_X16 FILLER_82_609 ();
 FILLCELL_X4 FILLER_82_625 ();
 FILLCELL_X2 FILLER_82_629 ();
 FILLCELL_X16 FILLER_82_632 ();
 FILLCELL_X8 FILLER_82_648 ();
 FILLCELL_X2 FILLER_82_656 ();
 FILLCELL_X32 FILLER_83_1 ();
 FILLCELL_X32 FILLER_83_33 ();
 FILLCELL_X32 FILLER_83_65 ();
 FILLCELL_X32 FILLER_83_97 ();
 FILLCELL_X32 FILLER_83_129 ();
 FILLCELL_X32 FILLER_83_161 ();
 FILLCELL_X32 FILLER_83_193 ();
 FILLCELL_X32 FILLER_83_225 ();
 FILLCELL_X32 FILLER_83_257 ();
 FILLCELL_X32 FILLER_83_289 ();
 FILLCELL_X32 FILLER_83_321 ();
 FILLCELL_X32 FILLER_83_353 ();
 FILLCELL_X32 FILLER_83_385 ();
 FILLCELL_X32 FILLER_83_417 ();
 FILLCELL_X32 FILLER_83_449 ();
 FILLCELL_X32 FILLER_83_481 ();
 FILLCELL_X32 FILLER_83_513 ();
 FILLCELL_X32 FILLER_83_545 ();
 FILLCELL_X32 FILLER_83_577 ();
 FILLCELL_X32 FILLER_83_609 ();
 FILLCELL_X16 FILLER_83_641 ();
 FILLCELL_X1 FILLER_83_657 ();
 FILLCELL_X32 FILLER_84_1 ();
 FILLCELL_X32 FILLER_84_33 ();
 FILLCELL_X32 FILLER_84_65 ();
 FILLCELL_X32 FILLER_84_97 ();
 FILLCELL_X32 FILLER_84_129 ();
 FILLCELL_X32 FILLER_84_161 ();
 FILLCELL_X32 FILLER_84_193 ();
 FILLCELL_X32 FILLER_84_225 ();
 FILLCELL_X32 FILLER_84_257 ();
 FILLCELL_X32 FILLER_84_289 ();
 FILLCELL_X32 FILLER_84_321 ();
 FILLCELL_X32 FILLER_84_353 ();
 FILLCELL_X32 FILLER_84_385 ();
 FILLCELL_X32 FILLER_84_417 ();
 FILLCELL_X32 FILLER_84_449 ();
 FILLCELL_X32 FILLER_84_481 ();
 FILLCELL_X32 FILLER_84_513 ();
 FILLCELL_X32 FILLER_84_545 ();
 FILLCELL_X32 FILLER_84_577 ();
 FILLCELL_X16 FILLER_84_609 ();
 FILLCELL_X4 FILLER_84_625 ();
 FILLCELL_X2 FILLER_84_629 ();
 FILLCELL_X16 FILLER_84_632 ();
 FILLCELL_X8 FILLER_84_648 ();
 FILLCELL_X2 FILLER_84_656 ();
 FILLCELL_X32 FILLER_85_1 ();
 FILLCELL_X32 FILLER_85_33 ();
 FILLCELL_X32 FILLER_85_65 ();
 FILLCELL_X32 FILLER_85_97 ();
 FILLCELL_X32 FILLER_85_129 ();
 FILLCELL_X32 FILLER_85_161 ();
 FILLCELL_X32 FILLER_85_193 ();
 FILLCELL_X32 FILLER_85_225 ();
 FILLCELL_X32 FILLER_85_257 ();
 FILLCELL_X32 FILLER_85_289 ();
 FILLCELL_X32 FILLER_85_321 ();
 FILLCELL_X32 FILLER_85_353 ();
 FILLCELL_X32 FILLER_85_385 ();
 FILLCELL_X32 FILLER_85_417 ();
 FILLCELL_X32 FILLER_85_449 ();
 FILLCELL_X32 FILLER_85_481 ();
 FILLCELL_X32 FILLER_85_513 ();
 FILLCELL_X32 FILLER_85_545 ();
 FILLCELL_X32 FILLER_85_577 ();
 FILLCELL_X32 FILLER_85_609 ();
 FILLCELL_X16 FILLER_85_641 ();
 FILLCELL_X1 FILLER_85_657 ();
 FILLCELL_X4 FILLER_86_1 ();
 FILLCELL_X32 FILLER_86_18 ();
 FILLCELL_X32 FILLER_86_50 ();
 FILLCELL_X32 FILLER_86_82 ();
 FILLCELL_X32 FILLER_86_114 ();
 FILLCELL_X32 FILLER_86_146 ();
 FILLCELL_X32 FILLER_86_178 ();
 FILLCELL_X32 FILLER_86_210 ();
 FILLCELL_X32 FILLER_86_242 ();
 FILLCELL_X32 FILLER_86_274 ();
 FILLCELL_X32 FILLER_86_306 ();
 FILLCELL_X32 FILLER_86_338 ();
 FILLCELL_X32 FILLER_86_370 ();
 FILLCELL_X32 FILLER_86_402 ();
 FILLCELL_X32 FILLER_86_434 ();
 FILLCELL_X32 FILLER_86_466 ();
 FILLCELL_X32 FILLER_86_498 ();
 FILLCELL_X32 FILLER_86_530 ();
 FILLCELL_X32 FILLER_86_562 ();
 FILLCELL_X32 FILLER_86_594 ();
 FILLCELL_X4 FILLER_86_626 ();
 FILLCELL_X1 FILLER_86_630 ();
 FILLCELL_X16 FILLER_86_632 ();
 FILLCELL_X8 FILLER_86_648 ();
 FILLCELL_X2 FILLER_86_656 ();
 FILLCELL_X32 FILLER_87_1 ();
 FILLCELL_X32 FILLER_87_33 ();
 FILLCELL_X32 FILLER_87_65 ();
 FILLCELL_X32 FILLER_87_97 ();
 FILLCELL_X32 FILLER_87_129 ();
 FILLCELL_X32 FILLER_87_161 ();
 FILLCELL_X32 FILLER_87_193 ();
 FILLCELL_X32 FILLER_87_225 ();
 FILLCELL_X32 FILLER_87_257 ();
 FILLCELL_X32 FILLER_87_289 ();
 FILLCELL_X32 FILLER_87_321 ();
 FILLCELL_X32 FILLER_87_353 ();
 FILLCELL_X32 FILLER_87_385 ();
 FILLCELL_X32 FILLER_87_417 ();
 FILLCELL_X32 FILLER_87_449 ();
 FILLCELL_X32 FILLER_87_481 ();
 FILLCELL_X32 FILLER_87_513 ();
 FILLCELL_X32 FILLER_87_545 ();
 FILLCELL_X32 FILLER_87_577 ();
 FILLCELL_X32 FILLER_87_609 ();
 FILLCELL_X16 FILLER_87_641 ();
 FILLCELL_X1 FILLER_87_657 ();
 FILLCELL_X16 FILLER_88_1 ();
 FILLCELL_X4 FILLER_88_17 ();
 FILLCELL_X32 FILLER_88_24 ();
 FILLCELL_X32 FILLER_88_56 ();
 FILLCELL_X16 FILLER_88_88 ();
 FILLCELL_X8 FILLER_88_104 ();
 FILLCELL_X2 FILLER_88_112 ();
 FILLCELL_X1 FILLER_88_114 ();
 FILLCELL_X32 FILLER_88_118 ();
 FILLCELL_X32 FILLER_88_150 ();
 FILLCELL_X16 FILLER_88_182 ();
 FILLCELL_X8 FILLER_88_198 ();
 FILLCELL_X2 FILLER_88_206 ();
 FILLCELL_X1 FILLER_88_208 ();
 FILLCELL_X32 FILLER_88_213 ();
 FILLCELL_X32 FILLER_88_245 ();
 FILLCELL_X16 FILLER_88_277 ();
 FILLCELL_X8 FILLER_88_293 ();
 FILLCELL_X2 FILLER_88_301 ();
 FILLCELL_X1 FILLER_88_303 ();
 FILLCELL_X32 FILLER_88_307 ();
 FILLCELL_X32 FILLER_88_339 ();
 FILLCELL_X16 FILLER_88_371 ();
 FILLCELL_X8 FILLER_88_387 ();
 FILLCELL_X2 FILLER_88_395 ();
 FILLCELL_X1 FILLER_88_397 ();
 FILLCELL_X32 FILLER_88_401 ();
 FILLCELL_X32 FILLER_88_433 ();
 FILLCELL_X16 FILLER_88_465 ();
 FILLCELL_X8 FILLER_88_481 ();
 FILLCELL_X2 FILLER_88_489 ();
 FILLCELL_X1 FILLER_88_491 ();
 FILLCELL_X32 FILLER_88_495 ();
 FILLCELL_X32 FILLER_88_527 ();
 FILLCELL_X16 FILLER_88_559 ();
 FILLCELL_X8 FILLER_88_575 ();
 FILLCELL_X4 FILLER_88_583 ();
 FILLCELL_X32 FILLER_88_590 ();
 FILLCELL_X8 FILLER_88_622 ();
 FILLCELL_X1 FILLER_88_630 ();
 FILLCELL_X16 FILLER_88_632 ();
 FILLCELL_X2 FILLER_88_648 ();
 FILLCELL_X1 FILLER_88_650 ();
 FILLCELL_X4 FILLER_88_654 ();
 assign init_done = curr_state[1];
 assign valid_out = valid_reg_out;
endmodule
