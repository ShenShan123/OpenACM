module sram_multiplier_system (clk,
    init_done,
    init_enable,
    pe_ce,
    rst_n,
    valid_out,
    data_in,
    data_out);
 input clk;
 output init_done;
 input init_enable;
 input pe_ce;
 input rst_n;
 output valid_out;
 input [31:0] data_in;
 output [63:0] data_out;

 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire \u_multiplier/_1830_ ;
 wire \u_multiplier/_1831_ ;
 wire \u_multiplier/_1832_ ;
 wire \u_multiplier/_1833_ ;
 wire \u_multiplier/_1834_ ;
 wire \u_multiplier/_1835_ ;
 wire \u_multiplier/_1836_ ;
 wire \u_multiplier/_1837_ ;
 wire \u_multiplier/_1838_ ;
 wire \u_multiplier/_1839_ ;
 wire \u_multiplier/_1840_ ;
 wire \u_multiplier/_1841_ ;
 wire \u_multiplier/_1842_ ;
 wire \u_multiplier/_1843_ ;
 wire \u_multiplier/_1844_ ;
 wire \u_multiplier/_1845_ ;
 wire \u_multiplier/_1846_ ;
 wire \u_multiplier/_1847_ ;
 wire \u_multiplier/_1848_ ;
 wire \u_multiplier/_1849_ ;
 wire \u_multiplier/_1850_ ;
 wire \u_multiplier/_1851_ ;
 wire \u_multiplier/_1852_ ;
 wire \u_multiplier/_1853_ ;
 wire \u_multiplier/_1854_ ;
 wire \u_multiplier/_1855_ ;
 wire \u_multiplier/_1856_ ;
 wire \u_multiplier/_1857_ ;
 wire \u_multiplier/_1858_ ;
 wire \u_multiplier/_1859_ ;
 wire \u_multiplier/_1860_ ;
 wire \u_multiplier/_1861_ ;
 wire \u_multiplier/_1862_ ;
 wire \u_multiplier/_1863_ ;
 wire \u_multiplier/_1864_ ;
 wire \u_multiplier/_1865_ ;
 wire \u_multiplier/_1866_ ;
 wire \u_multiplier/_2003_ ;
 wire \u_multiplier/_2004_ ;
 wire \u_multiplier/_2005_ ;
 wire \u_multiplier/_2006_ ;
 wire \u_multiplier/_2007_ ;
 wire \u_multiplier/_2008_ ;
 wire \u_multiplier/_2009_ ;
 wire \u_multiplier/_2010_ ;
 wire \u_multiplier/_2011_ ;
 wire \u_multiplier/_2012_ ;
 wire \u_multiplier/_2013_ ;
 wire \u_multiplier/_2014_ ;
 wire \u_multiplier/_2015_ ;
 wire \u_multiplier/_2016_ ;
 wire \u_multiplier/_2017_ ;
 wire \u_multiplier/_2018_ ;
 wire \u_multiplier/_2019_ ;
 wire \u_multiplier/_2020_ ;
 wire \u_multiplier/_2021_ ;
 wire \u_multiplier/_2022_ ;
 wire \u_multiplier/_2023_ ;
 wire \u_multiplier/_2024_ ;
 wire \u_multiplier/_2025_ ;
 wire \u_multiplier/_2026_ ;
 wire \u_multiplier/_2027_ ;
 wire \u_multiplier/_2028_ ;
 wire \u_multiplier/_2029_ ;
 wire \u_multiplier/_2030_ ;
 wire \u_multiplier/_2031_ ;
 wire \u_multiplier/_2032_ ;
 wire \u_multiplier/_2033_ ;
 wire \u_multiplier/_2034_ ;
 wire \u_multiplier/_2035_ ;
 wire \u_multiplier/_2036_ ;
 wire \u_multiplier/_2037_ ;
 wire \u_multiplier/_2038_ ;
 wire \u_multiplier/_2039_ ;
 wire \u_multiplier/_2040_ ;
 wire \u_multiplier/_2041_ ;
 wire \u_multiplier/_2042_ ;
 wire \u_multiplier/_2043_ ;
 wire \u_multiplier/_2044_ ;
 wire \u_multiplier/_2045_ ;
 wire \u_multiplier/_2046_ ;
 wire \u_multiplier/_2047_ ;
 wire \u_multiplier/_2048_ ;
 wire \u_multiplier/_2049_ ;
 wire \u_multiplier/_2050_ ;
 wire \u_multiplier/_2051_ ;
 wire \u_multiplier/_2052_ ;
 wire \u_multiplier/_2053_ ;
 wire \u_multiplier/_2054_ ;
 wire \u_multiplier/_2055_ ;
 wire \u_multiplier/_2056_ ;
 wire \u_multiplier/_2057_ ;
 wire \u_multiplier/_2058_ ;
 wire \u_multiplier/_2059_ ;
 wire \u_multiplier/_2060_ ;
 wire \u_multiplier/_2061_ ;
 wire \u_multiplier/_2062_ ;
 wire \u_multiplier/_2063_ ;
 wire \u_multiplier/_2064_ ;
 wire \u_multiplier/_2065_ ;
 wire \u_multiplier/_2066_ ;
 wire \u_multiplier/_2067_ ;
 wire \u_multiplier/_2068_ ;
 wire \u_multiplier/_2069_ ;
 wire \u_multiplier/_2070_ ;
 wire \u_multiplier/_2071_ ;
 wire \u_multiplier/_2072_ ;
 wire \u_multiplier/_2073_ ;
 wire \u_multiplier/_2074_ ;
 wire \u_multiplier/_2075_ ;
 wire \u_multiplier/_2076_ ;
 wire \u_multiplier/_2077_ ;
 wire \u_multiplier/_2078_ ;
 wire \u_multiplier/_2079_ ;
 wire \u_multiplier/_2080_ ;
 wire \u_multiplier/_2081_ ;
 wire \u_multiplier/_2082_ ;
 wire \u_multiplier/_2083_ ;
 wire \u_multiplier/_2084_ ;
 wire \u_multiplier/_2085_ ;
 wire \u_multiplier/_2086_ ;
 wire \u_multiplier/_2087_ ;
 wire \u_multiplier/_2088_ ;
 wire \u_multiplier/_2089_ ;
 wire \u_multiplier/_2090_ ;
 wire \u_multiplier/_2091_ ;
 wire \u_multiplier/_2092_ ;
 wire \u_multiplier/_2093_ ;
 wire \u_multiplier/_2094_ ;
 wire \u_multiplier/_2095_ ;
 wire \u_multiplier/_2096_ ;
 wire \u_multiplier/_2097_ ;
 wire \u_multiplier/_2098_ ;
 wire \u_multiplier/_2099_ ;
 wire \u_multiplier/_2100_ ;
 wire \u_multiplier/_2101_ ;
 wire \u_multiplier/_2102_ ;
 wire \u_multiplier/_2103_ ;
 wire \u_multiplier/_2104_ ;
 wire \u_multiplier/_2105_ ;
 wire \u_multiplier/_2106_ ;
 wire \u_multiplier/_2107_ ;
 wire \u_multiplier/_2108_ ;
 wire \u_multiplier/_2109_ ;
 wire \u_multiplier/_2110_ ;
 wire \u_multiplier/_2111_ ;
 wire \u_multiplier/_2112_ ;
 wire \u_multiplier/_2113_ ;
 wire \u_multiplier/_2114_ ;
 wire \u_multiplier/_2115_ ;
 wire \u_multiplier/_2116_ ;
 wire \u_multiplier/_2117_ ;
 wire \u_multiplier/_2118_ ;
 wire \u_multiplier/_2119_ ;
 wire \u_multiplier/_2120_ ;
 wire \u_multiplier/_2121_ ;
 wire \u_multiplier/_2122_ ;
 wire \u_multiplier/_2123_ ;
 wire \u_multiplier/_2124_ ;
 wire \u_multiplier/_2125_ ;
 wire \u_multiplier/_2126_ ;
 wire \u_multiplier/_2127_ ;
 wire \u_multiplier/_2128_ ;
 wire \u_multiplier/_2129_ ;
 wire \u_multiplier/_2130_ ;
 wire \u_multiplier/_2131_ ;
 wire \u_multiplier/_2132_ ;
 wire \u_multiplier/_2133_ ;
 wire \u_multiplier/_2134_ ;
 wire \u_multiplier/_2135_ ;
 wire \u_multiplier/_2136_ ;
 wire \u_multiplier/_2137_ ;
 wire \u_multiplier/_2138_ ;
 wire \u_multiplier/_2139_ ;
 wire \u_multiplier/_2140_ ;
 wire \u_multiplier/_2141_ ;
 wire \u_multiplier/_2142_ ;
 wire \u_multiplier/_2143_ ;
 wire \u_multiplier/_2144_ ;
 wire \u_multiplier/_2145_ ;
 wire \u_multiplier/_2146_ ;
 wire \u_multiplier/_2147_ ;
 wire \u_multiplier/_2148_ ;
 wire \u_multiplier/_2149_ ;
 wire \u_multiplier/_2150_ ;
 wire \u_multiplier/_2151_ ;
 wire \u_multiplier/_2152_ ;
 wire \u_multiplier/_2153_ ;
 wire \u_multiplier/_2154_ ;
 wire \u_multiplier/_2155_ ;
 wire \u_multiplier/_2156_ ;
 wire \u_multiplier/_2157_ ;
 wire \u_multiplier/_2158_ ;
 wire \u_multiplier/_2159_ ;
 wire \u_multiplier/_2160_ ;
 wire \u_multiplier/_2161_ ;
 wire \u_multiplier/_2162_ ;
 wire \u_multiplier/_2163_ ;
 wire \u_multiplier/_2164_ ;
 wire \u_multiplier/_2165_ ;
 wire \u_multiplier/_2166_ ;
 wire \u_multiplier/_2167_ ;
 wire \u_multiplier/_2168_ ;
 wire \u_multiplier/_2169_ ;
 wire \u_multiplier/_2170_ ;
 wire \u_multiplier/_2171_ ;
 wire \u_multiplier/_2172_ ;
 wire \u_multiplier/_2173_ ;
 wire \u_multiplier/_2174_ ;
 wire \u_multiplier/_2175_ ;
 wire \u_multiplier/_2176_ ;
 wire \u_multiplier/_2177_ ;
 wire \u_multiplier/_2178_ ;
 wire \u_multiplier/_2179_ ;
 wire \u_multiplier/_2180_ ;
 wire \u_multiplier/_2181_ ;
 wire \u_multiplier/_2182_ ;
 wire \u_multiplier/_2183_ ;
 wire \u_multiplier/_2184_ ;
 wire \u_multiplier/_2185_ ;
 wire \u_multiplier/_2186_ ;
 wire \u_multiplier/_2187_ ;
 wire \u_multiplier/_2188_ ;
 wire \u_multiplier/_2189_ ;
 wire \u_multiplier/_2190_ ;
 wire \u_multiplier/_2191_ ;
 wire \u_multiplier/_2192_ ;
 wire \u_multiplier/_2193_ ;
 wire \u_multiplier/_2194_ ;
 wire \u_multiplier/_2195_ ;
 wire \u_multiplier/_2196_ ;
 wire \u_multiplier/_2197_ ;
 wire \u_multiplier/_2198_ ;
 wire \u_multiplier/_2199_ ;
 wire \u_multiplier/_2200_ ;
 wire \u_multiplier/_2201_ ;
 wire \u_multiplier/_2202_ ;
 wire \u_multiplier/_2203_ ;
 wire \u_multiplier/_2204_ ;
 wire \u_multiplier/_2205_ ;
 wire \u_multiplier/_2206_ ;
 wire \u_multiplier/_2207_ ;
 wire \u_multiplier/_2208_ ;
 wire \u_multiplier/_2209_ ;
 wire \u_multiplier/_2210_ ;
 wire \u_multiplier/_2211_ ;
 wire \u_multiplier/_2212_ ;
 wire \u_multiplier/_2213_ ;
 wire \u_multiplier/_2214_ ;
 wire \u_multiplier/_2215_ ;
 wire \u_multiplier/_2216_ ;
 wire \u_multiplier/_2217_ ;
 wire \u_multiplier/_2218_ ;
 wire \u_multiplier/_2219_ ;
 wire \u_multiplier/_2220_ ;
 wire \u_multiplier/_2221_ ;
 wire \u_multiplier/_2222_ ;
 wire \u_multiplier/_2223_ ;
 wire \u_multiplier/_2224_ ;
 wire \u_multiplier/_2225_ ;
 wire \u_multiplier/_2226_ ;
 wire \u_multiplier/_2227_ ;
 wire \u_multiplier/_2228_ ;
 wire \u_multiplier/_2229_ ;
 wire \u_multiplier/_2230_ ;
 wire \u_multiplier/_2231_ ;
 wire \u_multiplier/_2232_ ;
 wire \u_multiplier/_2233_ ;
 wire \u_multiplier/_2234_ ;
 wire \u_multiplier/_2235_ ;
 wire \u_multiplier/_2236_ ;
 wire \u_multiplier/_2237_ ;
 wire \u_multiplier/_2238_ ;
 wire \u_multiplier/_2239_ ;
 wire \u_multiplier/_2240_ ;
 wire \u_multiplier/_2241_ ;
 wire \u_multiplier/_2242_ ;
 wire \u_multiplier/_2243_ ;
 wire \u_multiplier/_2244_ ;
 wire \u_multiplier/_2245_ ;
 wire \u_multiplier/_2246_ ;
 wire \u_multiplier/_2247_ ;
 wire \u_multiplier/_2248_ ;
 wire \u_multiplier/_2249_ ;
 wire \u_multiplier/_2250_ ;
 wire \u_multiplier/_2251_ ;
 wire \u_multiplier/_2252_ ;
 wire \u_multiplier/_2253_ ;
 wire \u_multiplier/_2254_ ;
 wire \u_multiplier/_2255_ ;
 wire \u_multiplier/_2256_ ;
 wire \u_multiplier/_2257_ ;
 wire \u_multiplier/_2258_ ;
 wire \u_multiplier/_2259_ ;
 wire \u_multiplier/_2260_ ;
 wire \u_multiplier/_2261_ ;
 wire \u_multiplier/_2262_ ;
 wire \u_multiplier/_2263_ ;
 wire \u_multiplier/_2264_ ;
 wire \u_multiplier/_2265_ ;
 wire \u_multiplier/_2266_ ;
 wire \u_multiplier/_2267_ ;
 wire \u_multiplier/_2268_ ;
 wire \u_multiplier/_2269_ ;
 wire \u_multiplier/_2270_ ;
 wire \u_multiplier/_2271_ ;
 wire \u_multiplier/_2272_ ;
 wire \u_multiplier/_2273_ ;
 wire \u_multiplier/_2274_ ;
 wire \u_multiplier/_2275_ ;
 wire \u_multiplier/_2276_ ;
 wire \u_multiplier/_2277_ ;
 wire \u_multiplier/_2278_ ;
 wire \u_multiplier/_2279_ ;
 wire \u_multiplier/_2280_ ;
 wire \u_multiplier/_2281_ ;
 wire \u_multiplier/_2282_ ;
 wire \u_multiplier/_2283_ ;
 wire \u_multiplier/_2284_ ;
 wire \u_multiplier/_2285_ ;
 wire \u_multiplier/_2286_ ;
 wire \u_multiplier/_2287_ ;
 wire \u_multiplier/_2288_ ;
 wire \u_multiplier/_2289_ ;
 wire \u_multiplier/_2290_ ;
 wire \u_multiplier/_2291_ ;
 wire \u_multiplier/_2292_ ;
 wire \u_multiplier/_2293_ ;
 wire \u_multiplier/_2294_ ;
 wire \u_multiplier/_2295_ ;
 wire \u_multiplier/_2296_ ;
 wire \u_multiplier/_2297_ ;
 wire \u_multiplier/_2298_ ;
 wire \u_multiplier/_2299_ ;
 wire \u_multiplier/_2300_ ;
 wire \u_multiplier/_2301_ ;
 wire \u_multiplier/_2302_ ;
 wire \u_multiplier/_2303_ ;
 wire \u_multiplier/_2304_ ;
 wire \u_multiplier/_2305_ ;
 wire \u_multiplier/_2306_ ;
 wire \u_multiplier/_2307_ ;
 wire \u_multiplier/_2308_ ;
 wire \u_multiplier/_2309_ ;
 wire \u_multiplier/_2310_ ;
 wire \u_multiplier/_2311_ ;
 wire \u_multiplier/_2312_ ;
 wire \u_multiplier/_2313_ ;
 wire \u_multiplier/_2314_ ;
 wire \u_multiplier/_2315_ ;
 wire \u_multiplier/_2316_ ;
 wire \u_multiplier/_2317_ ;
 wire \u_multiplier/_2318_ ;
 wire \u_multiplier/_2319_ ;
 wire \u_multiplier/_2320_ ;
 wire \u_multiplier/_2321_ ;
 wire \u_multiplier/_2322_ ;
 wire \u_multiplier/_2323_ ;
 wire \u_multiplier/_2324_ ;
 wire \u_multiplier/_2325_ ;
 wire \u_multiplier/_2326_ ;
 wire \u_multiplier/_2327_ ;
 wire \u_multiplier/_2328_ ;
 wire \u_multiplier/_2329_ ;
 wire \u_multiplier/_2330_ ;
 wire \u_multiplier/_2331_ ;
 wire \u_multiplier/_2332_ ;
 wire \u_multiplier/_2333_ ;
 wire \u_multiplier/_2334_ ;
 wire \u_multiplier/_2335_ ;
 wire \u_multiplier/_2336_ ;
 wire \u_multiplier/_2337_ ;
 wire \u_multiplier/_2338_ ;
 wire \u_multiplier/_2339_ ;
 wire \u_multiplier/_2340_ ;
 wire \u_multiplier/_2341_ ;
 wire \u_multiplier/_2342_ ;
 wire \u_multiplier/_2343_ ;
 wire \u_multiplier/_2344_ ;
 wire \u_multiplier/_2345_ ;
 wire \u_multiplier/_2346_ ;
 wire \u_multiplier/_2347_ ;
 wire \u_multiplier/_2348_ ;
 wire \u_multiplier/_2349_ ;
 wire \u_multiplier/_2350_ ;
 wire \u_multiplier/_2351_ ;
 wire \u_multiplier/_2352_ ;
 wire \u_multiplier/_2353_ ;
 wire \u_multiplier/_2354_ ;
 wire \u_multiplier/_2355_ ;
 wire \u_multiplier/_2356_ ;
 wire \u_multiplier/_2357_ ;
 wire \u_multiplier/_2358_ ;
 wire \u_multiplier/_2359_ ;
 wire \u_multiplier/_2360_ ;
 wire \u_multiplier/_2361_ ;
 wire \u_multiplier/_2362_ ;
 wire \u_multiplier/_2363_ ;
 wire \u_multiplier/_2364_ ;
 wire \u_multiplier/_2365_ ;
 wire \u_multiplier/_2366_ ;
 wire \u_multiplier/_2367_ ;
 wire \u_multiplier/_2368_ ;
 wire \u_multiplier/_2369_ ;
 wire \u_multiplier/_2370_ ;
 wire \u_multiplier/_2371_ ;
 wire \u_multiplier/_2372_ ;
 wire \u_multiplier/_2373_ ;
 wire \u_multiplier/_2374_ ;
 wire \u_multiplier/_2375_ ;
 wire \u_multiplier/_2376_ ;
 wire \u_multiplier/_2377_ ;
 wire \u_multiplier/_2378_ ;
 wire \u_multiplier/_2379_ ;
 wire \u_multiplier/_2380_ ;
 wire \u_multiplier/_2381_ ;
 wire \u_multiplier/_2382_ ;
 wire \u_multiplier/_2383_ ;
 wire \u_multiplier/_2384_ ;
 wire \u_multiplier/_2385_ ;
 wire \u_multiplier/_2386_ ;
 wire \u_multiplier/_2387_ ;
 wire \u_multiplier/_2388_ ;
 wire \u_multiplier/_2389_ ;
 wire \u_multiplier/_2390_ ;
 wire \u_multiplier/_2391_ ;
 wire \u_multiplier/_2392_ ;
 wire \u_multiplier/_2393_ ;
 wire \u_multiplier/_2394_ ;
 wire \u_multiplier/_2395_ ;
 wire \u_multiplier/_2396_ ;
 wire \u_multiplier/_2397_ ;
 wire \u_multiplier/_2398_ ;
 wire \u_multiplier/_2399_ ;
 wire \u_multiplier/_2400_ ;
 wire \u_multiplier/_2401_ ;
 wire \u_multiplier/_2402_ ;
 wire \u_multiplier/_2403_ ;
 wire \u_multiplier/_2404_ ;
 wire \u_multiplier/_2405_ ;
 wire \u_multiplier/_2406_ ;
 wire \u_multiplier/_2407_ ;
 wire \u_multiplier/_2408_ ;
 wire \u_multiplier/_2409_ ;
 wire \u_multiplier/_2410_ ;
 wire \u_multiplier/_2411_ ;
 wire \u_multiplier/_2412_ ;
 wire \u_multiplier/_2413_ ;
 wire \u_multiplier/_2414_ ;
 wire \u_multiplier/_2415_ ;
 wire \u_multiplier/_2416_ ;
 wire \u_multiplier/_2417_ ;
 wire \u_multiplier/_2418_ ;
 wire \u_multiplier/_2419_ ;
 wire \u_multiplier/_2420_ ;
 wire \u_multiplier/_2421_ ;
 wire \u_multiplier/_2422_ ;
 wire \u_multiplier/_2423_ ;
 wire \u_multiplier/_2424_ ;
 wire \u_multiplier/_2425_ ;
 wire \u_multiplier/_2426_ ;
 wire \u_multiplier/_2427_ ;
 wire \u_multiplier/_2428_ ;
 wire \u_multiplier/_2429_ ;
 wire \u_multiplier/_2430_ ;
 wire \u_multiplier/_2431_ ;
 wire \u_multiplier/_2432_ ;
 wire \u_multiplier/_2433_ ;
 wire \u_multiplier/_2434_ ;
 wire \u_multiplier/_2435_ ;
 wire \u_multiplier/_2436_ ;
 wire \u_multiplier/_2437_ ;
 wire \u_multiplier/_2438_ ;
 wire \u_multiplier/_2439_ ;
 wire \u_multiplier/_2440_ ;
 wire \u_multiplier/_2441_ ;
 wire \u_multiplier/_2442_ ;
 wire \u_multiplier/_2443_ ;
 wire \u_multiplier/_2444_ ;
 wire \u_multiplier/_2445_ ;
 wire \u_multiplier/_2446_ ;
 wire \u_multiplier/_2447_ ;
 wire \u_multiplier/_2448_ ;
 wire \u_multiplier/_2449_ ;
 wire \u_multiplier/_2450_ ;
 wire \u_multiplier/_2451_ ;
 wire \u_multiplier/_2452_ ;
 wire \u_multiplier/_2453_ ;
 wire \u_multiplier/_2454_ ;
 wire \u_multiplier/_2455_ ;
 wire \u_multiplier/_2456_ ;
 wire \u_multiplier/_2457_ ;
 wire \u_multiplier/_2458_ ;
 wire \u_multiplier/_2459_ ;
 wire \u_multiplier/_2460_ ;
 wire \u_multiplier/_2461_ ;
 wire \u_multiplier/_2462_ ;
 wire \u_multiplier/_2463_ ;
 wire \u_multiplier/_2464_ ;
 wire \u_multiplier/_2465_ ;
 wire \u_multiplier/_2466_ ;
 wire \u_multiplier/_2467_ ;
 wire \u_multiplier/_2468_ ;
 wire \u_multiplier/_2469_ ;
 wire \u_multiplier/_2470_ ;
 wire \u_multiplier/_2471_ ;
 wire \u_multiplier/_2472_ ;
 wire \u_multiplier/_2473_ ;
 wire \u_multiplier/_2474_ ;
 wire \u_multiplier/_2475_ ;
 wire \u_multiplier/_2476_ ;
 wire \u_multiplier/_2477_ ;
 wire \u_multiplier/_2478_ ;
 wire \u_multiplier/_2479_ ;
 wire \u_multiplier/_2480_ ;
 wire \u_multiplier/_2481_ ;
 wire \u_multiplier/_2482_ ;
 wire \u_multiplier/_2483_ ;
 wire \u_multiplier/_2484_ ;
 wire \u_multiplier/_2485_ ;
 wire \u_multiplier/_2486_ ;
 wire \u_multiplier/_2487_ ;
 wire \u_multiplier/_2488_ ;
 wire \u_multiplier/_2489_ ;
 wire \u_multiplier/_2490_ ;
 wire \u_multiplier/_2491_ ;
 wire \u_multiplier/_2492_ ;
 wire \u_multiplier/_2493_ ;
 wire \u_multiplier/_2494_ ;
 wire \u_multiplier/_2495_ ;
 wire \u_multiplier/_2496_ ;
 wire \u_multiplier/_2497_ ;
 wire \u_multiplier/_2498_ ;
 wire \u_multiplier/_2499_ ;
 wire \u_multiplier/_2500_ ;
 wire \u_multiplier/_2501_ ;
 wire \u_multiplier/_2502_ ;
 wire \u_multiplier/_2503_ ;
 wire \u_multiplier/_2504_ ;
 wire \u_multiplier/_2505_ ;
 wire \u_multiplier/_2506_ ;
 wire \u_multiplier/_2507_ ;
 wire \u_multiplier/_2508_ ;
 wire \u_multiplier/_2509_ ;
 wire \u_multiplier/_2510_ ;
 wire \u_multiplier/_2511_ ;
 wire \u_multiplier/_2512_ ;
 wire \u_multiplier/_2513_ ;
 wire \u_multiplier/_2514_ ;
 wire \u_multiplier/_2515_ ;
 wire \u_multiplier/_2516_ ;
 wire \u_multiplier/_2517_ ;
 wire \u_multiplier/_2518_ ;
 wire \u_multiplier/_2519_ ;
 wire \u_multiplier/_2520_ ;
 wire \u_multiplier/_2521_ ;
 wire \u_multiplier/_2522_ ;
 wire \u_multiplier/_2523_ ;
 wire \u_multiplier/_2524_ ;
 wire \u_multiplier/_2525_ ;
 wire \u_multiplier/_2526_ ;
 wire \u_multiplier/_2527_ ;
 wire \u_multiplier/_2528_ ;
 wire \u_multiplier/_2529_ ;
 wire \u_multiplier/_2530_ ;
 wire \u_multiplier/_2531_ ;
 wire \u_multiplier/_2532_ ;
 wire \u_multiplier/_2533_ ;
 wire \u_multiplier/_2534_ ;
 wire \u_multiplier/_2535_ ;
 wire \u_multiplier/_2536_ ;
 wire \u_multiplier/_2537_ ;
 wire \u_multiplier/_2538_ ;
 wire \u_multiplier/_2539_ ;
 wire \u_multiplier/_2540_ ;
 wire \u_multiplier/_2541_ ;
 wire \u_multiplier/_2542_ ;
 wire \u_multiplier/_2543_ ;
 wire \u_multiplier/_2544_ ;
 wire \u_multiplier/_2545_ ;
 wire \u_multiplier/_2546_ ;
 wire \u_multiplier/_2547_ ;
 wire \u_multiplier/_2548_ ;
 wire \u_multiplier/_2549_ ;
 wire \u_multiplier/_2550_ ;
 wire \u_multiplier/_2551_ ;
 wire \u_multiplier/_2552_ ;
 wire \u_multiplier/_2553_ ;
 wire \u_multiplier/_2554_ ;
 wire \u_multiplier/_2555_ ;
 wire \u_multiplier/_2556_ ;
 wire \u_multiplier/_2557_ ;
 wire \u_multiplier/_2558_ ;
 wire \u_multiplier/_2559_ ;
 wire \u_multiplier/_2560_ ;
 wire \u_multiplier/_2561_ ;
 wire \u_multiplier/_2562_ ;
 wire \u_multiplier/_2563_ ;
 wire \u_multiplier/_2564_ ;
 wire \u_multiplier/_2565_ ;
 wire \u_multiplier/_2566_ ;
 wire \u_multiplier/_2567_ ;
 wire \u_multiplier/_2568_ ;
 wire \u_multiplier/_2569_ ;
 wire \u_multiplier/_2570_ ;
 wire \u_multiplier/_2571_ ;
 wire \u_multiplier/_2572_ ;
 wire \u_multiplier/_2573_ ;
 wire \u_multiplier/_2574_ ;
 wire \u_multiplier/_2575_ ;
 wire \u_multiplier/_2576_ ;
 wire \u_multiplier/_2577_ ;
 wire \u_multiplier/_2578_ ;
 wire \u_multiplier/_2579_ ;
 wire \u_multiplier/_2580_ ;
 wire \u_multiplier/_2581_ ;
 wire \u_multiplier/_2582_ ;
 wire \u_multiplier/_2583_ ;
 wire \u_multiplier/_2584_ ;
 wire \u_multiplier/_2585_ ;
 wire \u_multiplier/_2586_ ;
 wire \u_multiplier/_2587_ ;
 wire \u_multiplier/_2588_ ;
 wire \u_multiplier/_2589_ ;
 wire \u_multiplier/_2590_ ;
 wire \u_multiplier/_2591_ ;
 wire \u_multiplier/_2592_ ;
 wire \u_multiplier/_2593_ ;
 wire \u_multiplier/_2594_ ;
 wire \u_multiplier/_2595_ ;
 wire \u_multiplier/_2596_ ;
 wire \u_multiplier/_2597_ ;
 wire \u_multiplier/_2598_ ;
 wire \u_multiplier/_2599_ ;
 wire \u_multiplier/_2600_ ;
 wire \u_multiplier/_2601_ ;
 wire \u_multiplier/_2602_ ;
 wire \u_multiplier/_2603_ ;
 wire \u_multiplier/_2604_ ;
 wire \u_multiplier/_2605_ ;
 wire \u_multiplier/_2606_ ;
 wire \u_multiplier/_2607_ ;
 wire \u_multiplier/_2608_ ;
 wire \u_multiplier/_2609_ ;
 wire \u_multiplier/_2610_ ;
 wire \u_multiplier/_2611_ ;
 wire \u_multiplier/_2612_ ;
 wire \u_multiplier/_2613_ ;
 wire \u_multiplier/_2614_ ;
 wire \u_multiplier/_2615_ ;
 wire \u_multiplier/_2616_ ;
 wire \u_multiplier/_2617_ ;
 wire \u_multiplier/_2618_ ;
 wire \u_multiplier/_2619_ ;
 wire \u_multiplier/_2620_ ;
 wire \u_multiplier/_2621_ ;
 wire \u_multiplier/_2622_ ;
 wire \u_multiplier/_2623_ ;
 wire \u_multiplier/_2624_ ;
 wire \u_multiplier/_2625_ ;
 wire \u_multiplier/_2626_ ;
 wire \u_multiplier/_2627_ ;
 wire \u_multiplier/_2628_ ;
 wire \u_multiplier/_2629_ ;
 wire \u_multiplier/_2630_ ;
 wire \u_multiplier/_2631_ ;
 wire \u_multiplier/_2632_ ;
 wire \u_multiplier/_2633_ ;
 wire \u_multiplier/_2634_ ;
 wire \u_multiplier/_2635_ ;
 wire \u_multiplier/_2636_ ;
 wire \u_multiplier/_2637_ ;
 wire \u_multiplier/_2638_ ;
 wire \u_multiplier/_2639_ ;
 wire \u_multiplier/_2640_ ;
 wire \u_multiplier/_2641_ ;
 wire \u_multiplier/_2642_ ;
 wire \u_multiplier/_2643_ ;
 wire \u_multiplier/_2644_ ;
 wire \u_multiplier/_2645_ ;
 wire \u_multiplier/_2646_ ;
 wire \u_multiplier/_2647_ ;
 wire \u_multiplier/_2648_ ;
 wire \u_multiplier/_2649_ ;
 wire \u_multiplier/_2650_ ;
 wire \u_multiplier/_2651_ ;
 wire \u_multiplier/_2652_ ;
 wire \u_multiplier/_2653_ ;
 wire \u_multiplier/_2654_ ;
 wire \u_multiplier/_2655_ ;
 wire \u_multiplier/_2656_ ;
 wire \u_multiplier/_2657_ ;
 wire \u_multiplier/_2658_ ;
 wire \u_multiplier/_2659_ ;
 wire \u_multiplier/_2660_ ;
 wire \u_multiplier/_2661_ ;
 wire \u_multiplier/_2662_ ;
 wire \u_multiplier/_2663_ ;
 wire \u_multiplier/_2664_ ;
 wire \u_multiplier/_2665_ ;
 wire \u_multiplier/_2666_ ;
 wire \u_multiplier/_2667_ ;
 wire \u_multiplier/_2668_ ;
 wire \u_multiplier/_2669_ ;
 wire \u_multiplier/_2670_ ;
 wire \u_multiplier/_2671_ ;
 wire \u_multiplier/_2672_ ;
 wire \u_multiplier/_2673_ ;
 wire \u_multiplier/_2674_ ;
 wire \u_multiplier/_2675_ ;
 wire \u_multiplier/_2676_ ;
 wire \u_multiplier/_2677_ ;
 wire \u_multiplier/_2678_ ;
 wire \u_multiplier/_2679_ ;
 wire \u_multiplier/_2680_ ;
 wire \u_multiplier/_2681_ ;
 wire \u_multiplier/_2682_ ;
 wire \u_multiplier/_2683_ ;
 wire \u_multiplier/_2684_ ;
 wire \u_multiplier/_2685_ ;
 wire \u_multiplier/_2686_ ;
 wire \u_multiplier/_2687_ ;
 wire \u_multiplier/_2688_ ;
 wire \u_multiplier/_2689_ ;
 wire \u_multiplier/_2690_ ;
 wire \u_multiplier/_2691_ ;
 wire \u_multiplier/_2692_ ;
 wire \u_multiplier/_2693_ ;
 wire \u_multiplier/_2694_ ;
 wire \u_multiplier/_2695_ ;
 wire \u_multiplier/_2696_ ;
 wire \u_multiplier/_2697_ ;
 wire \u_multiplier/_2698_ ;
 wire \u_multiplier/_2699_ ;
 wire \u_multiplier/_2700_ ;
 wire \u_multiplier/_2701_ ;
 wire \u_multiplier/_2702_ ;
 wire \u_multiplier/_2703_ ;
 wire \u_multiplier/_2704_ ;
 wire \u_multiplier/_2705_ ;
 wire \u_multiplier/_2706_ ;
 wire \u_multiplier/_2707_ ;
 wire \u_multiplier/_2708_ ;
 wire \u_multiplier/_2709_ ;
 wire \u_multiplier/_2710_ ;
 wire \u_multiplier/_2711_ ;
 wire \u_multiplier/_2712_ ;
 wire \u_multiplier/_2713_ ;
 wire \u_multiplier/_2714_ ;
 wire \u_multiplier/_2715_ ;
 wire \u_multiplier/_2716_ ;
 wire \u_multiplier/_2717_ ;
 wire \u_multiplier/_2718_ ;
 wire \u_multiplier/_2719_ ;
 wire \u_multiplier/_2720_ ;
 wire \u_multiplier/_2721_ ;
 wire \u_multiplier/_2722_ ;
 wire \u_multiplier/_2723_ ;
 wire \u_multiplier/_2724_ ;
 wire \u_multiplier/_2725_ ;
 wire \u_multiplier/_2726_ ;
 wire \u_multiplier/_2727_ ;
 wire \u_multiplier/_2728_ ;
 wire \u_multiplier/_2729_ ;
 wire \u_multiplier/_2730_ ;
 wire \u_multiplier/_2731_ ;
 wire \u_multiplier/_2732_ ;
 wire \u_multiplier/_2733_ ;
 wire \u_multiplier/_2734_ ;
 wire \u_multiplier/_2735_ ;
 wire \u_multiplier/_2736_ ;
 wire \u_multiplier/_2737_ ;
 wire \u_multiplier/_2738_ ;
 wire \u_multiplier/_2739_ ;
 wire \u_multiplier/_2740_ ;
 wire \u_multiplier/_2741_ ;
 wire \u_multiplier/_2742_ ;
 wire \u_multiplier/_2743_ ;
 wire \u_multiplier/_2744_ ;
 wire \u_multiplier/_2745_ ;
 wire \u_multiplier/_2746_ ;
 wire \u_multiplier/_2747_ ;
 wire \u_multiplier/_2748_ ;
 wire \u_multiplier/_2749_ ;
 wire \u_multiplier/_2750_ ;
 wire \u_multiplier/_2751_ ;
 wire \u_multiplier/_2752_ ;
 wire \u_multiplier/_2753_ ;
 wire \u_multiplier/_2754_ ;
 wire \u_multiplier/_2755_ ;
 wire \u_multiplier/_2756_ ;
 wire \u_multiplier/_2757_ ;
 wire \u_multiplier/_2758_ ;
 wire \u_multiplier/_2759_ ;
 wire \u_multiplier/_2760_ ;
 wire \u_multiplier/_2761_ ;
 wire \u_multiplier/_2762_ ;
 wire \u_multiplier/_2763_ ;
 wire \u_multiplier/_2764_ ;
 wire \u_multiplier/_2765_ ;
 wire \u_multiplier/_2766_ ;
 wire \u_multiplier/_2767_ ;
 wire \u_multiplier/_2768_ ;
 wire \u_multiplier/_2769_ ;
 wire \u_multiplier/_2770_ ;
 wire \u_multiplier/_2771_ ;
 wire \u_multiplier/_2772_ ;
 wire \u_multiplier/_2773_ ;
 wire \u_multiplier/_2774_ ;
 wire \u_multiplier/_2775_ ;
 wire \u_multiplier/_2776_ ;
 wire \u_multiplier/_2777_ ;
 wire \u_multiplier/_2778_ ;
 wire \u_multiplier/_2779_ ;
 wire \u_multiplier/_2780_ ;
 wire \u_multiplier/_2781_ ;
 wire \u_multiplier/_2782_ ;
 wire \u_multiplier/_2783_ ;
 wire \u_multiplier/_2784_ ;
 wire \u_multiplier/_2785_ ;
 wire \u_multiplier/_2786_ ;
 wire \u_multiplier/_2787_ ;
 wire \u_multiplier/_2788_ ;
 wire \u_multiplier/_2789_ ;
 wire \u_multiplier/_2790_ ;
 wire \u_multiplier/_2791_ ;
 wire \u_multiplier/_2792_ ;
 wire \u_multiplier/_2793_ ;
 wire \u_multiplier/_2794_ ;
 wire \u_multiplier/_2795_ ;
 wire \u_multiplier/_2796_ ;
 wire \u_multiplier/_2797_ ;
 wire \u_multiplier/_2798_ ;
 wire \u_multiplier/_2799_ ;
 wire \u_multiplier/_2800_ ;
 wire \u_multiplier/_2801_ ;
 wire \u_multiplier/_2802_ ;
 wire \u_multiplier/_2803_ ;
 wire \u_multiplier/_2804_ ;
 wire \u_multiplier/_2805_ ;
 wire \u_multiplier/_2806_ ;
 wire \u_multiplier/_2807_ ;
 wire \u_multiplier/_2808_ ;
 wire \u_multiplier/_2809_ ;
 wire \u_multiplier/_2810_ ;
 wire \u_multiplier/_2811_ ;
 wire \u_multiplier/_2812_ ;
 wire \u_multiplier/_2813_ ;
 wire \u_multiplier/_2814_ ;
 wire \u_multiplier/_2815_ ;
 wire \u_multiplier/_2816_ ;
 wire \u_multiplier/_2817_ ;
 wire \u_multiplier/_2818_ ;
 wire \u_multiplier/_2819_ ;
 wire \u_multiplier/_2820_ ;
 wire \u_multiplier/_2821_ ;
 wire \u_multiplier/_2822_ ;
 wire \u_multiplier/_2823_ ;
 wire \u_multiplier/_2824_ ;
 wire \u_multiplier/_2825_ ;
 wire \u_multiplier/_2826_ ;
 wire \u_multiplier/_2827_ ;
 wire \u_multiplier/_2828_ ;
 wire \u_multiplier/_2829_ ;
 wire \u_multiplier/_2830_ ;
 wire \u_multiplier/_2831_ ;
 wire \u_multiplier/_2832_ ;
 wire \u_multiplier/_2833_ ;
 wire \u_multiplier/_2834_ ;
 wire \u_multiplier/_2835_ ;
 wire \u_multiplier/_2836_ ;
 wire \u_multiplier/_2837_ ;
 wire \u_multiplier/_2838_ ;
 wire \u_multiplier/_2839_ ;
 wire \u_multiplier/_2840_ ;
 wire \u_multiplier/_2841_ ;
 wire \u_multiplier/_2842_ ;
 wire \u_multiplier/_2843_ ;
 wire \u_multiplier/_2844_ ;
 wire \u_multiplier/_2845_ ;
 wire \u_multiplier/_2846_ ;
 wire \u_multiplier/_2847_ ;
 wire \u_multiplier/_2848_ ;
 wire \u_multiplier/_2849_ ;
 wire \u_multiplier/_2850_ ;
 wire \u_multiplier/_2851_ ;
 wire \u_multiplier/_2852_ ;
 wire \u_multiplier/_2853_ ;
 wire \u_multiplier/_2854_ ;
 wire \u_multiplier/_2855_ ;
 wire \u_multiplier/_2856_ ;
 wire \u_multiplier/_2857_ ;
 wire \u_multiplier/_2858_ ;
 wire \u_multiplier/_2859_ ;
 wire \u_multiplier/_2860_ ;
 wire \u_multiplier/_2861_ ;
 wire \u_multiplier/_2862_ ;
 wire \u_multiplier/_2863_ ;
 wire \u_multiplier/_2864_ ;
 wire \u_multiplier/_2865_ ;
 wire \u_multiplier/_2866_ ;
 wire \u_multiplier/_2867_ ;
 wire \u_multiplier/_2868_ ;
 wire \u_multiplier/_2869_ ;
 wire \u_multiplier/_2870_ ;
 wire \u_multiplier/_2871_ ;
 wire \u_multiplier/_2872_ ;
 wire \u_multiplier/_2873_ ;
 wire \u_multiplier/_2874_ ;
 wire \u_multiplier/_2875_ ;
 wire \u_multiplier/_2876_ ;
 wire \u_multiplier/_2877_ ;
 wire \u_multiplier/_2878_ ;
 wire \u_multiplier/_2879_ ;
 wire \u_multiplier/_2880_ ;
 wire \u_multiplier/_2881_ ;
 wire \u_multiplier/_2882_ ;
 wire \u_multiplier/_2883_ ;
 wire \u_multiplier/_2884_ ;
 wire \u_multiplier/_2885_ ;
 wire \u_multiplier/_2886_ ;
 wire \u_multiplier/_2887_ ;
 wire \u_multiplier/_2888_ ;
 wire \u_multiplier/_2889_ ;
 wire \u_multiplier/_2890_ ;
 wire \u_multiplier/_2891_ ;
 wire \u_multiplier/_2892_ ;
 wire \u_multiplier/_2893_ ;
 wire \u_multiplier/_2894_ ;
 wire \u_multiplier/_2895_ ;
 wire \u_multiplier/_2896_ ;
 wire \u_multiplier/_2897_ ;
 wire \u_multiplier/_2898_ ;
 wire \u_multiplier/_2899_ ;
 wire \u_multiplier/_2900_ ;
 wire \u_multiplier/_2901_ ;
 wire \u_multiplier/_2902_ ;
 wire \u_multiplier/_2903_ ;
 wire \u_multiplier/_2904_ ;
 wire \u_multiplier/_2905_ ;
 wire \u_multiplier/_2906_ ;
 wire \u_multiplier/_2907_ ;
 wire \u_multiplier/_2908_ ;
 wire \u_multiplier/_2909_ ;
 wire \u_multiplier/_2910_ ;
 wire \u_multiplier/_2911_ ;
 wire \u_multiplier/_2912_ ;
 wire \u_multiplier/_2913_ ;
 wire \u_multiplier/_2914_ ;
 wire \u_multiplier/_2915_ ;
 wire \u_multiplier/_2916_ ;
 wire \u_multiplier/_2917_ ;
 wire \u_multiplier/_2918_ ;
 wire \u_multiplier/_2919_ ;
 wire \u_multiplier/_2920_ ;
 wire \u_multiplier/_2921_ ;
 wire \u_multiplier/_2922_ ;
 wire \u_multiplier/_2923_ ;
 wire \u_multiplier/_2924_ ;
 wire \u_multiplier/_2925_ ;
 wire \u_multiplier/_2926_ ;
 wire \u_multiplier/_2927_ ;
 wire \u_multiplier/_2928_ ;
 wire \u_multiplier/_2929_ ;
 wire \u_multiplier/_2930_ ;
 wire \u_multiplier/_2931_ ;
 wire \u_multiplier/_2932_ ;
 wire \u_multiplier/_2933_ ;
 wire \u_multiplier/_2934_ ;
 wire \u_multiplier/_2935_ ;
 wire \u_multiplier/_2936_ ;
 wire \u_multiplier/_2937_ ;
 wire \u_multiplier/_2938_ ;
 wire \u_multiplier/_2939_ ;
 wire \u_multiplier/_2940_ ;
 wire \u_multiplier/_2941_ ;
 wire \u_multiplier/_2942_ ;
 wire \u_multiplier/_2943_ ;
 wire \u_multiplier/_2944_ ;
 wire \u_multiplier/_2945_ ;
 wire \u_multiplier/_2946_ ;
 wire \u_multiplier/_2947_ ;
 wire \u_multiplier/_2948_ ;
 wire \u_multiplier/_2949_ ;
 wire \u_multiplier/_2950_ ;
 wire \u_multiplier/_2951_ ;
 wire \u_multiplier/_2952_ ;
 wire \u_multiplier/_2953_ ;
 wire \u_multiplier/_2954_ ;
 wire \u_multiplier/_2955_ ;
 wire \u_multiplier/_2956_ ;
 wire \u_multiplier/_2957_ ;
 wire \u_multiplier/_2958_ ;
 wire \u_multiplier/_2959_ ;
 wire \u_multiplier/_2960_ ;
 wire \u_multiplier/_2961_ ;
 wire \u_multiplier/_2962_ ;
 wire \u_multiplier/_2963_ ;
 wire \u_multiplier/_2964_ ;
 wire \u_multiplier/_2965_ ;
 wire \u_multiplier/_2966_ ;
 wire \u_multiplier/_2967_ ;
 wire \u_multiplier/_2968_ ;
 wire \u_multiplier/_2969_ ;
 wire \u_multiplier/_2970_ ;
 wire \u_multiplier/_2971_ ;
 wire \u_multiplier/_2972_ ;
 wire \u_multiplier/_2973_ ;
 wire \u_multiplier/_2974_ ;
 wire \u_multiplier/_2975_ ;
 wire \u_multiplier/_2976_ ;
 wire \u_multiplier/_2977_ ;
 wire \u_multiplier/_2978_ ;
 wire \u_multiplier/_2979_ ;
 wire \u_multiplier/_2980_ ;
 wire \u_multiplier/_2981_ ;
 wire \u_multiplier/_2982_ ;
 wire \u_multiplier/_2983_ ;
 wire \u_multiplier/_2984_ ;
 wire \u_multiplier/_2985_ ;
 wire \u_multiplier/_2986_ ;
 wire \u_multiplier/_2987_ ;
 wire \u_multiplier/_2988_ ;
 wire \u_multiplier/_2989_ ;
 wire \u_multiplier/_2990_ ;
 wire \u_multiplier/_2991_ ;
 wire \u_multiplier/_2992_ ;
 wire \u_multiplier/_2993_ ;
 wire \u_multiplier/_2994_ ;
 wire \u_multiplier/_2995_ ;
 wire \u_multiplier/_2996_ ;
 wire \u_multiplier/_2997_ ;
 wire \u_multiplier/_2998_ ;
 wire \u_multiplier/_2999_ ;
 wire \u_multiplier/_3000_ ;
 wire \u_multiplier/_3001_ ;
 wire \u_multiplier/_3002_ ;
 wire \u_multiplier/_3003_ ;
 wire \u_multiplier/_3004_ ;
 wire \u_multiplier/_3005_ ;
 wire \u_multiplier/_3006_ ;
 wire \u_multiplier/_3007_ ;
 wire \u_multiplier/_3008_ ;
 wire \u_multiplier/_3009_ ;
 wire \u_multiplier/_3010_ ;
 wire \u_multiplier/_3011_ ;
 wire \u_multiplier/_3012_ ;
 wire \u_multiplier/_3013_ ;
 wire \u_multiplier/_3014_ ;
 wire \u_multiplier/_3015_ ;
 wire \u_multiplier/_3016_ ;
 wire \u_multiplier/_3017_ ;
 wire \u_multiplier/_3018_ ;
 wire \u_multiplier/_3019_ ;
 wire \u_multiplier/_3020_ ;
 wire \u_multiplier/_3021_ ;
 wire \u_multiplier/_3022_ ;
 wire \u_multiplier/_3023_ ;
 wire \u_multiplier/_3024_ ;
 wire \u_multiplier/_3025_ ;
 wire \u_multiplier/_3026_ ;
 wire \u_multiplier/_3027_ ;
 wire \u_multiplier/_3028_ ;
 wire \u_multiplier/_3029_ ;
 wire \u_multiplier/_3030_ ;
 wire \u_multiplier/_3031_ ;
 wire \u_multiplier/_3032_ ;
 wire \u_multiplier/_3033_ ;
 wire \u_multiplier/_3034_ ;
 wire \u_multiplier/_3035_ ;
 wire \u_multiplier/_3036_ ;
 wire \u_multiplier/_3037_ ;
 wire \u_multiplier/_3038_ ;
 wire \u_multiplier/_3039_ ;
 wire \u_multiplier/_3040_ ;
 wire \u_multiplier/_3041_ ;
 wire \u_multiplier/_3042_ ;
 wire \u_multiplier/_3043_ ;
 wire \u_multiplier/_3044_ ;
 wire \u_multiplier/_3045_ ;
 wire \u_multiplier/_3046_ ;
 wire \u_multiplier/_3047_ ;
 wire \u_multiplier/_3048_ ;
 wire \u_multiplier/_3049_ ;
 wire \u_multiplier/_3050_ ;
 wire \u_multiplier/_3051_ ;
 wire \u_multiplier/_3052_ ;
 wire \u_multiplier/_3053_ ;
 wire \u_multiplier/_3054_ ;
 wire \u_multiplier/_3055_ ;
 wire \u_multiplier/_3056_ ;
 wire \u_multiplier/_3057_ ;
 wire \u_multiplier/_3058_ ;
 wire \u_multiplier/_3059_ ;
 wire \u_multiplier/_3060_ ;
 wire \u_multiplier/_3061_ ;
 wire \u_multiplier/_3062_ ;
 wire \u_multiplier/_3063_ ;
 wire \u_multiplier/_3064_ ;
 wire \u_multiplier/_3065_ ;
 wire \u_multiplier/_3066_ ;
 wire \u_multiplier/_3067_ ;
 wire \u_multiplier/_3068_ ;
 wire \u_multiplier/_3069_ ;
 wire \u_multiplier/_3070_ ;
 wire \u_multiplier/_3071_ ;
 wire \u_multiplier/_3072_ ;
 wire \u_multiplier/_3073_ ;
 wire \u_multiplier/_3074_ ;
 wire \u_multiplier/_3075_ ;
 wire \u_multiplier/_3076_ ;
 wire \u_multiplier/_3077_ ;
 wire \u_multiplier/_3078_ ;
 wire \u_multiplier/_3079_ ;
 wire \u_multiplier/_3080_ ;
 wire \u_multiplier/_3081_ ;
 wire \u_multiplier/_3082_ ;
 wire \u_multiplier/_3083_ ;
 wire \u_multiplier/_3084_ ;
 wire \u_multiplier/_3085_ ;
 wire \u_multiplier/_3086_ ;
 wire \u_multiplier/_3087_ ;
 wire \u_multiplier/_3088_ ;
 wire \u_multiplier/_3089_ ;
 wire \u_multiplier/_3090_ ;
 wire \u_multiplier/_3091_ ;
 wire \u_multiplier/_3092_ ;
 wire \u_multiplier/_3093_ ;
 wire \u_multiplier/_3094_ ;
 wire \u_multiplier/_3095_ ;
 wire \u_multiplier/_3096_ ;
 wire \u_multiplier/_3097_ ;
 wire \u_multiplier/_3098_ ;
 wire \u_multiplier/_3099_ ;
 wire \u_multiplier/_3100_ ;
 wire \u_multiplier/_3101_ ;
 wire \u_multiplier/_3102_ ;
 wire \u_multiplier/_3103_ ;
 wire \u_multiplier/_3104_ ;
 wire \u_multiplier/_3105_ ;
 wire \u_multiplier/_3106_ ;
 wire \u_multiplier/_3107_ ;
 wire \u_multiplier/_3108_ ;
 wire \u_multiplier/_3109_ ;
 wire \u_multiplier/_3110_ ;
 wire \u_multiplier/_3111_ ;
 wire \u_multiplier/_3112_ ;
 wire \u_multiplier/_3113_ ;
 wire \u_multiplier/_3114_ ;
 wire \u_multiplier/_3115_ ;
 wire \u_multiplier/_3116_ ;
 wire \u_multiplier/_3117_ ;
 wire \u_multiplier/_3118_ ;
 wire \u_multiplier/_3119_ ;
 wire \u_multiplier/_3120_ ;
 wire \u_multiplier/_3121_ ;
 wire \u_multiplier/_3122_ ;
 wire \u_multiplier/_3123_ ;
 wire \u_multiplier/_3124_ ;
 wire \u_multiplier/_3125_ ;
 wire \u_multiplier/_3126_ ;
 wire \u_multiplier/_3127_ ;
 wire \u_multiplier/_3128_ ;
 wire \u_multiplier/_3129_ ;
 wire \u_multiplier/_3130_ ;
 wire \u_multiplier/_3131_ ;
 wire \u_multiplier/_3132_ ;
 wire \u_multiplier/_3133_ ;
 wire \u_multiplier/_3134_ ;
 wire \u_multiplier/_3135_ ;
 wire \u_multiplier/_3136_ ;
 wire \u_multiplier/_3137_ ;
 wire \u_multiplier/_3138_ ;
 wire \u_multiplier/_3139_ ;
 wire \u_multiplier/_3140_ ;
 wire \u_multiplier/_3141_ ;
 wire \u_multiplier/_3142_ ;
 wire \u_multiplier/_3143_ ;
 wire \u_multiplier/_3144_ ;
 wire \u_multiplier/_3145_ ;
 wire \u_multiplier/_3146_ ;
 wire \u_multiplier/_3147_ ;
 wire \u_multiplier/_3148_ ;
 wire \u_multiplier/_3149_ ;
 wire \u_multiplier/_3150_ ;
 wire \u_multiplier/_3151_ ;
 wire \u_multiplier/_3152_ ;
 wire \u_multiplier/_3153_ ;
 wire \u_multiplier/_3154_ ;
 wire \u_multiplier/_3155_ ;
 wire \u_multiplier/_3156_ ;
 wire \u_multiplier/_3157_ ;
 wire \u_multiplier/_3158_ ;
 wire \u_multiplier/_3159_ ;
 wire \u_multiplier/_3160_ ;
 wire \u_multiplier/_3161_ ;
 wire \u_multiplier/_3162_ ;
 wire \u_multiplier/_3163_ ;
 wire \u_multiplier/_3164_ ;
 wire \u_multiplier/_3165_ ;
 wire \u_multiplier/_3166_ ;
 wire \u_multiplier/_3167_ ;
 wire \u_multiplier/_3168_ ;
 wire \u_multiplier/_3169_ ;
 wire \u_multiplier/_3170_ ;
 wire \u_multiplier/_3171_ ;
 wire \u_multiplier/_3172_ ;
 wire \u_multiplier/_3173_ ;
 wire \u_multiplier/_3174_ ;
 wire \u_multiplier/_3175_ ;
 wire \u_multiplier/_3176_ ;
 wire \u_multiplier/_3177_ ;
 wire \u_multiplier/_3178_ ;
 wire \u_multiplier/_3179_ ;
 wire \u_multiplier/_3180_ ;
 wire \u_multiplier/_3181_ ;
 wire \u_multiplier/_3182_ ;
 wire \u_multiplier/_3183_ ;
 wire \u_multiplier/_3184_ ;
 wire \u_multiplier/_3185_ ;
 wire \u_multiplier/_3186_ ;
 wire \u_multiplier/_3187_ ;
 wire \u_multiplier/_3188_ ;
 wire \u_multiplier/_3189_ ;
 wire \u_multiplier/_3190_ ;
 wire \u_multiplier/_3191_ ;
 wire \u_multiplier/_3192_ ;
 wire \u_multiplier/_3193_ ;
 wire \u_multiplier/_3194_ ;
 wire \u_multiplier/_3195_ ;
 wire \u_multiplier/_3196_ ;
 wire \u_multiplier/_3197_ ;
 wire \u_multiplier/_3198_ ;
 wire \u_multiplier/_3199_ ;
 wire \u_multiplier/_3200_ ;
 wire \u_multiplier/_3201_ ;
 wire \u_multiplier/_3202_ ;
 wire \u_multiplier/_3203_ ;
 wire \u_multiplier/_3204_ ;
 wire \u_multiplier/_3205_ ;
 wire \u_multiplier/_3206_ ;
 wire \u_multiplier/_3207_ ;
 wire \u_multiplier/_3208_ ;
 wire \u_multiplier/_3209_ ;
 wire \u_multiplier/_3210_ ;
 wire \u_multiplier/_3211_ ;
 wire \u_multiplier/_3212_ ;
 wire \u_multiplier/_3213_ ;
 wire \u_multiplier/_3214_ ;
 wire \u_multiplier/_3215_ ;
 wire \u_multiplier/_3216_ ;
 wire \u_multiplier/_3217_ ;
 wire \u_multiplier/_3218_ ;
 wire \u_multiplier/_3219_ ;
 wire \u_multiplier/_3220_ ;
 wire \u_multiplier/_3221_ ;
 wire \u_multiplier/_3222_ ;
 wire \u_multiplier/_3223_ ;
 wire \u_multiplier/_3224_ ;
 wire \u_multiplier/_3225_ ;
 wire \u_multiplier/_3226_ ;
 wire \u_multiplier/_3227_ ;
 wire \u_multiplier/_3228_ ;
 wire \u_multiplier/_3229_ ;
 wire \u_multiplier/_3230_ ;
 wire \u_multiplier/_3231_ ;
 wire \u_multiplier/_3232_ ;
 wire \u_multiplier/_3233_ ;
 wire \u_multiplier/_3234_ ;
 wire \u_multiplier/_3235_ ;
 wire \u_multiplier/_3236_ ;
 wire \u_multiplier/_3237_ ;
 wire \u_multiplier/_3238_ ;
 wire \u_multiplier/_3239_ ;
 wire \u_multiplier/_3240_ ;
 wire \u_multiplier/_3241_ ;
 wire \u_multiplier/_3242_ ;
 wire \u_multiplier/_3243_ ;
 wire \u_multiplier/_3244_ ;
 wire \u_multiplier/_3245_ ;
 wire \u_multiplier/_3246_ ;
 wire \u_multiplier/_3247_ ;
 wire \u_multiplier/_3248_ ;
 wire \u_multiplier/_3249_ ;
 wire \u_multiplier/_3250_ ;
 wire \u_multiplier/_3251_ ;
 wire \u_multiplier/_3252_ ;
 wire \u_multiplier/_3253_ ;
 wire \u_multiplier/_3254_ ;
 wire \u_multiplier/_3255_ ;
 wire \u_multiplier/_3256_ ;
 wire \u_multiplier/_3257_ ;
 wire \u_multiplier/_3258_ ;
 wire \u_multiplier/_3259_ ;
 wire \u_multiplier/_3260_ ;
 wire \u_multiplier/_3261_ ;
 wire \u_multiplier/_3262_ ;
 wire \u_multiplier/_3263_ ;
 wire \u_multiplier/_3264_ ;
 wire \u_multiplier/_3265_ ;
 wire \u_multiplier/_3266_ ;
 wire \u_multiplier/_3267_ ;
 wire \u_multiplier/_3268_ ;
 wire \u_multiplier/_3269_ ;
 wire \u_multiplier/_3270_ ;
 wire \u_multiplier/_3271_ ;
 wire \u_multiplier/_3272_ ;
 wire \u_multiplier/_3273_ ;
 wire \u_multiplier/_3274_ ;
 wire \u_multiplier/_3275_ ;
 wire \u_multiplier/_3276_ ;
 wire \u_multiplier/_3277_ ;
 wire \u_multiplier/_3278_ ;
 wire \u_multiplier/_3279_ ;
 wire \u_multiplier/_3280_ ;
 wire \u_multiplier/_3281_ ;
 wire \u_multiplier/_3282_ ;
 wire \u_multiplier/_3283_ ;
 wire \u_multiplier/_3284_ ;
 wire \u_multiplier/_3285_ ;
 wire \u_multiplier/_3286_ ;
 wire \u_multiplier/_3287_ ;
 wire \u_multiplier/_3288_ ;
 wire \u_multiplier/_3289_ ;
 wire \u_multiplier/_3290_ ;
 wire \u_multiplier/_3291_ ;
 wire \u_multiplier/_3292_ ;
 wire \u_multiplier/_3293_ ;
 wire \u_multiplier/_3294_ ;
 wire \u_multiplier/_3295_ ;
 wire \u_multiplier/_3296_ ;
 wire \u_multiplier/_3297_ ;
 wire \u_multiplier/_3298_ ;
 wire \u_multiplier/_3299_ ;
 wire \u_multiplier/_3300_ ;
 wire \u_multiplier/_3301_ ;
 wire \u_multiplier/_3302_ ;
 wire \u_multiplier/_3303_ ;
 wire \u_multiplier/_3304_ ;
 wire \u_multiplier/_3305_ ;
 wire \u_multiplier/_3306_ ;
 wire \u_multiplier/_3307_ ;
 wire \u_multiplier/_3308_ ;
 wire \u_multiplier/_3309_ ;
 wire \u_multiplier/_3310_ ;
 wire \u_multiplier/_3311_ ;
 wire \u_multiplier/_3312_ ;
 wire \u_multiplier/_3313_ ;
 wire \u_multiplier/_3314_ ;
 wire \u_multiplier/_3315_ ;
 wire \u_multiplier/_3316_ ;
 wire \u_multiplier/_3317_ ;
 wire \u_multiplier/_3318_ ;
 wire \u_multiplier/_3319_ ;
 wire \u_multiplier/_3320_ ;
 wire \u_multiplier/_3321_ ;
 wire \u_multiplier/_3322_ ;
 wire \u_multiplier/_3323_ ;
 wire \u_multiplier/_3324_ ;
 wire \u_multiplier/_3325_ ;
 wire \u_multiplier/_3326_ ;
 wire \u_multiplier/_3327_ ;
 wire \u_multiplier/_3328_ ;
 wire \u_multiplier/_3329_ ;
 wire \u_multiplier/_3330_ ;
 wire \u_multiplier/_3331_ ;
 wire \u_multiplier/_3332_ ;
 wire \u_multiplier/_3333_ ;
 wire \u_multiplier/_3334_ ;
 wire \u_multiplier/_3335_ ;
 wire \u_multiplier/_3336_ ;
 wire \u_multiplier/_3337_ ;
 wire \u_multiplier/_3338_ ;
 wire \u_multiplier/_3339_ ;
 wire \u_multiplier/_3340_ ;
 wire \u_multiplier/_3341_ ;
 wire \u_multiplier/_3342_ ;
 wire \u_multiplier/_3343_ ;
 wire \u_multiplier/_3344_ ;
 wire \u_multiplier/_3345_ ;
 wire \u_multiplier/_3346_ ;
 wire \u_multiplier/_3347_ ;
 wire \u_multiplier/_3348_ ;
 wire \u_multiplier/_3349_ ;
 wire \u_multiplier/_3350_ ;
 wire \u_multiplier/_3351_ ;
 wire \u_multiplier/_3352_ ;
 wire \u_multiplier/_3353_ ;
 wire \u_multiplier/_3354_ ;
 wire \u_multiplier/_3355_ ;
 wire \u_multiplier/_3356_ ;
 wire \u_multiplier/_3357_ ;
 wire \u_multiplier/_3358_ ;
 wire \u_multiplier/_3359_ ;
 wire \u_multiplier/_3360_ ;
 wire \u_multiplier/_3361_ ;
 wire \u_multiplier/_3362_ ;
 wire \u_multiplier/_3363_ ;
 wire \u_multiplier/_3364_ ;
 wire \u_multiplier/_3365_ ;
 wire \u_multiplier/_3366_ ;
 wire \u_multiplier/_3367_ ;
 wire \u_multiplier/_3368_ ;
 wire \u_multiplier/_3369_ ;
 wire \u_multiplier/_3370_ ;
 wire \u_multiplier/_3371_ ;
 wire \u_multiplier/_3372_ ;
 wire \u_multiplier/_3373_ ;
 wire \u_multiplier/_3374_ ;
 wire \u_multiplier/_3375_ ;
 wire \u_multiplier/_3376_ ;
 wire \u_multiplier/_3377_ ;
 wire \u_multiplier/_3378_ ;
 wire \u_multiplier/_3379_ ;
 wire \u_multiplier/_3380_ ;
 wire \u_multiplier/_3381_ ;
 wire \u_multiplier/_3382_ ;
 wire \u_multiplier/_3383_ ;
 wire \u_multiplier/_3384_ ;
 wire \u_multiplier/_3385_ ;
 wire \u_multiplier/_3386_ ;
 wire \u_multiplier/_3387_ ;
 wire \u_multiplier/_3388_ ;
 wire \u_multiplier/_3389_ ;
 wire \u_multiplier/_3390_ ;
 wire \u_multiplier/_3391_ ;
 wire \u_multiplier/_3392_ ;
 wire \u_multiplier/_3393_ ;
 wire \u_multiplier/_3394_ ;
 wire \u_multiplier/_3395_ ;
 wire \u_multiplier/_3396_ ;
 wire \u_multiplier/_3397_ ;
 wire \u_multiplier/_3398_ ;
 wire \u_multiplier/_3399_ ;
 wire \u_multiplier/_3400_ ;
 wire \u_multiplier/_3401_ ;
 wire \u_multiplier/_3402_ ;
 wire \u_multiplier/_3403_ ;
 wire \u_multiplier/_3404_ ;
 wire \u_multiplier/_3405_ ;
 wire \u_multiplier/_3406_ ;
 wire \u_multiplier/_3407_ ;
 wire \u_multiplier/_3408_ ;
 wire \u_multiplier/_3409_ ;
 wire \u_multiplier/_3410_ ;
 wire \u_multiplier/_3411_ ;
 wire \u_multiplier/_3412_ ;
 wire \u_multiplier/_3413_ ;
 wire \u_multiplier/_3414_ ;
 wire \u_multiplier/_3415_ ;
 wire \u_multiplier/_3416_ ;
 wire \u_multiplier/_3417_ ;
 wire \u_multiplier/_3418_ ;
 wire \u_multiplier/_3419_ ;
 wire \u_multiplier/_3420_ ;
 wire \u_multiplier/_3421_ ;
 wire \u_multiplier/_3422_ ;
 wire \u_multiplier/_3423_ ;
 wire \u_multiplier/_3424_ ;
 wire \u_multiplier/_3425_ ;
 wire \u_multiplier/_3426_ ;
 wire \u_multiplier/_3427_ ;
 wire \u_multiplier/_3428_ ;
 wire \u_multiplier/_3429_ ;
 wire \u_multiplier/_3430_ ;
 wire \u_multiplier/_3431_ ;
 wire \u_multiplier/_3432_ ;
 wire \u_multiplier/_3433_ ;
 wire \u_multiplier/_3434_ ;
 wire \u_multiplier/_3435_ ;
 wire \u_multiplier/_3436_ ;
 wire \u_multiplier/_3437_ ;
 wire \u_multiplier/_3438_ ;
 wire \u_multiplier/_3439_ ;
 wire \u_multiplier/_3440_ ;
 wire \u_multiplier/_3441_ ;
 wire \u_multiplier/_3442_ ;
 wire \u_multiplier/_3443_ ;
 wire \u_multiplier/_3444_ ;
 wire \u_multiplier/_3445_ ;
 wire \u_multiplier/_3446_ ;
 wire \u_multiplier/_3447_ ;
 wire \u_multiplier/_3448_ ;
 wire \u_multiplier/_3449_ ;
 wire \u_multiplier/_3450_ ;
 wire \u_multiplier/_3451_ ;
 wire \u_multiplier/_3452_ ;
 wire \u_multiplier/_3453_ ;
 wire \u_multiplier/_3454_ ;
 wire \u_multiplier/_3455_ ;
 wire \u_multiplier/_3456_ ;
 wire \u_multiplier/_3457_ ;
 wire \u_multiplier/_3458_ ;
 wire \u_multiplier/_3459_ ;
 wire \u_multiplier/_3460_ ;
 wire \u_multiplier/_3461_ ;
 wire \u_multiplier/_3462_ ;
 wire \u_multiplier/_3463_ ;
 wire \u_multiplier/_3464_ ;
 wire \u_multiplier/_3465_ ;
 wire \u_multiplier/_3466_ ;
 wire \u_multiplier/_3467_ ;
 wire \u_multiplier/_3468_ ;
 wire \u_multiplier/_3469_ ;
 wire \u_multiplier/_3470_ ;
 wire \u_multiplier/_3471_ ;
 wire \u_multiplier/_3472_ ;
 wire \u_multiplier/_3473_ ;
 wire \u_multiplier/_3474_ ;
 wire \u_multiplier/_3475_ ;
 wire \u_multiplier/_3476_ ;
 wire \u_multiplier/_3477_ ;
 wire \u_multiplier/_3478_ ;
 wire \u_multiplier/_3479_ ;
 wire \u_multiplier/_3480_ ;
 wire \u_multiplier/_3481_ ;
 wire \u_multiplier/_3482_ ;
 wire \u_multiplier/_3483_ ;
 wire \u_multiplier/_3484_ ;
 wire \u_multiplier/_3485_ ;
 wire \u_multiplier/_3486_ ;
 wire \u_multiplier/_3487_ ;
 wire \u_multiplier/_3488_ ;
 wire \u_multiplier/_3489_ ;
 wire \u_multiplier/_3490_ ;
 wire \u_multiplier/_3491_ ;
 wire \u_multiplier/_3492_ ;
 wire \u_multiplier/_3493_ ;
 wire \u_multiplier/_3494_ ;
 wire \u_multiplier/_3495_ ;
 wire \u_multiplier/_3496_ ;
 wire \u_multiplier/_3497_ ;
 wire \u_multiplier/_3498_ ;
 wire \u_multiplier/_3499_ ;
 wire \u_multiplier/_3500_ ;
 wire \u_multiplier/_3501_ ;
 wire \u_multiplier/_3502_ ;
 wire \u_multiplier/_3503_ ;
 wire \u_multiplier/_3504_ ;
 wire \u_multiplier/_3505_ ;
 wire \u_multiplier/_3506_ ;
 wire \u_multiplier/_3507_ ;
 wire \u_multiplier/_3508_ ;
 wire \u_multiplier/_3509_ ;
 wire \u_multiplier/_3510_ ;
 wire \u_multiplier/_3511_ ;
 wire \u_multiplier/_3512_ ;
 wire \u_multiplier/_3513_ ;
 wire \u_multiplier/_3514_ ;
 wire \u_multiplier/_3515_ ;
 wire \u_multiplier/_3516_ ;
 wire \u_multiplier/_3517_ ;
 wire \u_multiplier/_3518_ ;
 wire \u_multiplier/_3519_ ;
 wire \u_multiplier/_3520_ ;
 wire \u_multiplier/_3521_ ;
 wire \u_multiplier/_3522_ ;
 wire \u_multiplier/_3523_ ;
 wire \u_multiplier/_3524_ ;
 wire \u_multiplier/_3525_ ;
 wire \u_multiplier/_3526_ ;
 wire \u_multiplier/_3527_ ;
 wire \u_multiplier/_3528_ ;
 wire \u_multiplier/_3529_ ;
 wire \u_multiplier/_3530_ ;
 wire \u_multiplier/_3531_ ;
 wire \u_multiplier/_3532_ ;
 wire \u_multiplier/_3533_ ;
 wire \u_multiplier/_3534_ ;
 wire \u_multiplier/_3535_ ;
 wire \u_multiplier/_3536_ ;
 wire \u_multiplier/_3537_ ;
 wire \u_multiplier/_3538_ ;
 wire \u_multiplier/_3539_ ;
 wire \u_multiplier/_3540_ ;
 wire \u_multiplier/_3541_ ;
 wire \u_multiplier/_3542_ ;
 wire \u_multiplier/_3543_ ;
 wire \u_multiplier/_3544_ ;
 wire \u_multiplier/_3545_ ;
 wire \u_multiplier/_3546_ ;
 wire \u_multiplier/_3547_ ;
 wire \u_multiplier/_3548_ ;
 wire \u_multiplier/_3549_ ;
 wire \u_multiplier/_3550_ ;
 wire \u_multiplier/_3551_ ;
 wire \u_multiplier/_3552_ ;
 wire \u_multiplier/_3553_ ;
 wire \u_multiplier/_3554_ ;
 wire \u_multiplier/_3555_ ;
 wire \u_multiplier/_3556_ ;
 wire \u_multiplier/_3557_ ;
 wire \u_multiplier/_3558_ ;
 wire \u_multiplier/_3559_ ;
 wire \u_multiplier/_3560_ ;
 wire \u_multiplier/_3561_ ;
 wire \u_multiplier/_3562_ ;
 wire \u_multiplier/_3563_ ;
 wire \u_multiplier/_3564_ ;
 wire \u_multiplier/_3565_ ;
 wire \u_multiplier/_3566_ ;
 wire \u_multiplier/_3567_ ;
 wire \u_multiplier/_3568_ ;
 wire \u_multiplier/_3569_ ;
 wire \u_multiplier/_3570_ ;
 wire \u_multiplier/_3571_ ;
 wire \u_multiplier/_3572_ ;
 wire \u_multiplier/_3573_ ;
 wire \u_multiplier/_3574_ ;
 wire \u_multiplier/_3575_ ;
 wire \u_multiplier/_3576_ ;
 wire \u_multiplier/_3577_ ;
 wire \u_multiplier/_3578_ ;
 wire \u_multiplier/_3579_ ;
 wire \u_multiplier/_3580_ ;
 wire \u_multiplier/_3581_ ;
 wire \u_multiplier/_3582_ ;
 wire \u_multiplier/_3583_ ;
 wire \u_multiplier/_3584_ ;
 wire \u_multiplier/_3585_ ;
 wire \u_multiplier/_3586_ ;
 wire \u_multiplier/_3587_ ;
 wire \u_multiplier/_3588_ ;
 wire \u_multiplier/_3589_ ;
 wire \u_multiplier/_3590_ ;
 wire \u_multiplier/_3591_ ;
 wire \u_multiplier/_3592_ ;
 wire \u_multiplier/_3593_ ;
 wire \u_multiplier/_3594_ ;
 wire \u_multiplier/_3595_ ;
 wire \u_multiplier/_3596_ ;
 wire \u_multiplier/_3597_ ;
 wire \u_multiplier/_3598_ ;
 wire \u_multiplier/_3599_ ;
 wire \u_multiplier/_3600_ ;
 wire \u_multiplier/_3601_ ;
 wire \u_multiplier/_3602_ ;
 wire \u_multiplier/_3603_ ;
 wire \u_multiplier/_3604_ ;
 wire \u_multiplier/_3605_ ;
 wire \u_multiplier/_3606_ ;
 wire \u_multiplier/_3607_ ;
 wire \u_multiplier/_3608_ ;
 wire \u_multiplier/_3609_ ;
 wire \u_multiplier/_3610_ ;
 wire \u_multiplier/_3611_ ;
 wire \u_multiplier/_3612_ ;
 wire \u_multiplier/_3613_ ;
 wire \u_multiplier/_3614_ ;
 wire \u_multiplier/_3615_ ;
 wire \u_multiplier/_3616_ ;
 wire \u_multiplier/_3617_ ;
 wire \u_multiplier/_3618_ ;
 wire \u_multiplier/_3619_ ;
 wire \u_multiplier/_3620_ ;
 wire \u_multiplier/_3621_ ;
 wire \u_multiplier/_3622_ ;
 wire \u_multiplier/_3623_ ;
 wire \u_multiplier/_3624_ ;
 wire \u_multiplier/_3625_ ;
 wire \u_multiplier/_3626_ ;
 wire \u_multiplier/_3627_ ;
 wire \u_multiplier/_3628_ ;
 wire \u_multiplier/_3629_ ;
 wire \u_multiplier/_3630_ ;
 wire \u_multiplier/_3631_ ;
 wire \u_multiplier/_3632_ ;
 wire \u_multiplier/_3633_ ;
 wire \u_multiplier/_3634_ ;
 wire \u_multiplier/_3635_ ;
 wire \u_multiplier/_3636_ ;
 wire \u_multiplier/_3637_ ;
 wire \u_multiplier/_3638_ ;
 wire \u_multiplier/_3639_ ;
 wire \u_multiplier/_3640_ ;
 wire \u_multiplier/_3641_ ;
 wire \u_multiplier/_3642_ ;
 wire \u_multiplier/_3643_ ;
 wire \u_multiplier/_3644_ ;
 wire \u_multiplier/_3645_ ;
 wire \u_multiplier/_3646_ ;
 wire \u_multiplier/_3647_ ;
 wire \u_multiplier/_3648_ ;
 wire \u_multiplier/_3649_ ;
 wire \u_multiplier/_3650_ ;
 wire \u_multiplier/_3651_ ;
 wire \u_multiplier/_3652_ ;
 wire \u_multiplier/_3653_ ;
 wire \u_multiplier/_3654_ ;
 wire \u_multiplier/_3655_ ;
 wire \u_multiplier/_3656_ ;
 wire \u_multiplier/_3657_ ;
 wire \u_multiplier/_3658_ ;
 wire \u_multiplier/_3659_ ;
 wire \u_multiplier/_3660_ ;
 wire \u_multiplier/_3661_ ;
 wire \u_multiplier/_3662_ ;
 wire \u_multiplier/_3663_ ;
 wire \u_multiplier/_3664_ ;
 wire \u_multiplier/_3665_ ;
 wire \u_multiplier/_3666_ ;
 wire \u_multiplier/_3667_ ;
 wire \u_multiplier/_3668_ ;
 wire \u_multiplier/_3669_ ;
 wire \u_multiplier/_3670_ ;
 wire \u_multiplier/_3671_ ;
 wire \u_multiplier/_3672_ ;
 wire \u_multiplier/_3673_ ;
 wire \u_multiplier/_3674_ ;
 wire \u_multiplier/_3675_ ;
 wire \u_multiplier/_3676_ ;
 wire \u_multiplier/_3677_ ;
 wire \u_multiplier/_3678_ ;
 wire \u_multiplier/_3679_ ;
 wire \u_multiplier/_3680_ ;
 wire \u_multiplier/_3681_ ;
 wire \u_multiplier/_3682_ ;
 wire \u_multiplier/_3683_ ;
 wire \u_multiplier/_3684_ ;
 wire \u_multiplier/_3685_ ;
 wire \u_multiplier/_3686_ ;
 wire \u_multiplier/_3687_ ;
 wire \u_multiplier/_3688_ ;
 wire \u_multiplier/_3689_ ;
 wire \u_multiplier/_3690_ ;
 wire \u_multiplier/_3691_ ;
 wire \u_multiplier/_3692_ ;
 wire \u_multiplier/_3693_ ;
 wire \u_multiplier/_3694_ ;
 wire \u_multiplier/_3695_ ;
 wire \u_multiplier/_3696_ ;
 wire \u_multiplier/_3697_ ;
 wire \u_multiplier/_3698_ ;
 wire \u_multiplier/_3699_ ;
 wire \u_multiplier/_3700_ ;
 wire \u_multiplier/_3701_ ;
 wire \u_multiplier/_3702_ ;
 wire \u_multiplier/_3703_ ;
 wire \u_multiplier/_3704_ ;
 wire \u_multiplier/_3705_ ;
 wire \u_multiplier/_3706_ ;
 wire \u_multiplier/_3707_ ;
 wire \u_multiplier/_3708_ ;
 wire \u_multiplier/_3709_ ;
 wire \u_multiplier/_3710_ ;
 wire \u_multiplier/_3711_ ;
 wire \u_multiplier/_3712_ ;
 wire \u_multiplier/_3713_ ;
 wire \u_multiplier/_3714_ ;
 wire \u_multiplier/_3715_ ;
 wire \u_multiplier/_3716_ ;
 wire \u_multiplier/_3717_ ;
 wire \u_multiplier/_3718_ ;
 wire \u_multiplier/_3719_ ;
 wire \u_multiplier/_3720_ ;
 wire \u_multiplier/_3721_ ;
 wire \u_multiplier/_3722_ ;
 wire \u_multiplier/_3723_ ;
 wire \u_multiplier/_3724_ ;
 wire \u_multiplier/_3725_ ;
 wire \u_multiplier/_3726_ ;
 wire \u_multiplier/_3727_ ;
 wire \u_multiplier/_3728_ ;
 wire \u_multiplier/_3729_ ;
 wire \u_multiplier/_3730_ ;
 wire \u_multiplier/_3731_ ;
 wire \u_multiplier/_3732_ ;
 wire \u_multiplier/_3733_ ;
 wire \u_multiplier/_3734_ ;
 wire \u_multiplier/_3735_ ;
 wire \u_multiplier/_3736_ ;
 wire \u_multiplier/_3737_ ;
 wire \u_multiplier/_3738_ ;
 wire \u_multiplier/_3739_ ;
 wire \u_multiplier/_3740_ ;
 wire \u_multiplier/_3741_ ;
 wire \u_multiplier/_3742_ ;
 wire \u_multiplier/_3743_ ;
 wire \u_multiplier/_3744_ ;
 wire \u_multiplier/_3745_ ;
 wire \u_multiplier/_3746_ ;
 wire \u_multiplier/_3747_ ;
 wire \u_multiplier/_3748_ ;
 wire \u_multiplier/_3749_ ;
 wire \u_multiplier/_3750_ ;
 wire \u_multiplier/_3751_ ;
 wire net125;
 wire \u_multiplier/zero_x ;
 wire \u_multiplier/zero_y ;
 wire \u_multiplier/LODx/_054_ ;
 wire \u_multiplier/LODx/_055_ ;
 wire \u_multiplier/LODx/_056_ ;
 wire \u_multiplier/LODx/_057_ ;
 wire \u_multiplier/LODx/_058_ ;
 wire \u_multiplier/LODx/_059_ ;
 wire \u_multiplier/LODx/_060_ ;
 wire \u_multiplier/LODx/_061_ ;
 wire \u_multiplier/LODx/_062_ ;
 wire \u_multiplier/LODx/_063_ ;
 wire \u_multiplier/LODx/_064_ ;
 wire \u_multiplier/LODx/_065_ ;
 wire \u_multiplier/LODx/_066_ ;
 wire \u_multiplier/LODx/_067_ ;
 wire \u_multiplier/LODx/_068_ ;
 wire \u_multiplier/LODx/_077_ ;
 wire \u_multiplier/LODx/_078_ ;
 wire \u_multiplier/LODx/_079_ ;
 wire \u_multiplier/LODx/_080_ ;
 wire \u_multiplier/LODx/_081_ ;
 wire \u_multiplier/LODx/_082_ ;
 wire \u_multiplier/LODx/_083_ ;
 wire \u_multiplier/LODx/_084_ ;
 wire \u_multiplier/LODx/lod4_0/_09_ ;
 wire \u_multiplier/LODx/lod4_0/_10_ ;
 wire \u_multiplier/LODx/lod4_0/_11_ ;
 wire \u_multiplier/LODx/lod4_1/_09_ ;
 wire \u_multiplier/LODx/lod4_1/_10_ ;
 wire \u_multiplier/LODx/lod4_1/_11_ ;
 wire \u_multiplier/LODx/lod4_2/_09_ ;
 wire \u_multiplier/LODx/lod4_2/_10_ ;
 wire \u_multiplier/LODx/lod4_2/_11_ ;
 wire \u_multiplier/LODx/lod4_3/_09_ ;
 wire \u_multiplier/LODx/lod4_3/_10_ ;
 wire \u_multiplier/LODx/lod4_3/_11_ ;
 wire \u_multiplier/LODx/lod4_4/_09_ ;
 wire \u_multiplier/LODx/lod4_4/_10_ ;
 wire \u_multiplier/LODx/lod4_4/_11_ ;
 wire \u_multiplier/LODx/lod4_5/_09_ ;
 wire \u_multiplier/LODx/lod4_5/_10_ ;
 wire \u_multiplier/LODx/lod4_5/_11_ ;
 wire \u_multiplier/LODx/lod4_6/_09_ ;
 wire \u_multiplier/LODx/lod4_6/_10_ ;
 wire \u_multiplier/LODx/lod4_6/_11_ ;
 wire \u_multiplier/LODx/lod4_7/_09_ ;
 wire \u_multiplier/LODx/lod4_7/_10_ ;
 wire \u_multiplier/LODx/lod4_7/_11_ ;
 wire \u_multiplier/LODx/lod4_middle_high/_09_ ;
 wire \u_multiplier/LODx/lod4_middle_high/_10_ ;
 wire \u_multiplier/LODx/lod4_middle_high/_11_ ;
 wire \u_multiplier/LODx/lod4_middle_low/_09_ ;
 wire \u_multiplier/LODx/lod4_middle_low/_10_ ;
 wire \u_multiplier/LODx/lod4_middle_low/_11_ ;
 wire \u_multiplier/LODy/_054_ ;
 wire \u_multiplier/LODy/_055_ ;
 wire \u_multiplier/LODy/_056_ ;
 wire \u_multiplier/LODy/_057_ ;
 wire \u_multiplier/LODy/_058_ ;
 wire \u_multiplier/LODy/_059_ ;
 wire \u_multiplier/LODy/_060_ ;
 wire \u_multiplier/LODy/_061_ ;
 wire \u_multiplier/LODy/_062_ ;
 wire \u_multiplier/LODy/_063_ ;
 wire \u_multiplier/LODy/_064_ ;
 wire \u_multiplier/LODy/_065_ ;
 wire \u_multiplier/LODy/_066_ ;
 wire \u_multiplier/LODy/_067_ ;
 wire \u_multiplier/LODy/_068_ ;
 wire \u_multiplier/LODy/_077_ ;
 wire \u_multiplier/LODy/_078_ ;
 wire \u_multiplier/LODy/_079_ ;
 wire \u_multiplier/LODy/_080_ ;
 wire \u_multiplier/LODy/_081_ ;
 wire \u_multiplier/LODy/_082_ ;
 wire \u_multiplier/LODy/_083_ ;
 wire \u_multiplier/LODy/_084_ ;
 wire \u_multiplier/LODy/lod4_0/_09_ ;
 wire \u_multiplier/LODy/lod4_0/_10_ ;
 wire \u_multiplier/LODy/lod4_0/_11_ ;
 wire \u_multiplier/LODy/lod4_1/_09_ ;
 wire \u_multiplier/LODy/lod4_1/_10_ ;
 wire \u_multiplier/LODy/lod4_1/_11_ ;
 wire \u_multiplier/LODy/lod4_2/_09_ ;
 wire \u_multiplier/LODy/lod4_2/_10_ ;
 wire \u_multiplier/LODy/lod4_2/_11_ ;
 wire \u_multiplier/LODy/lod4_3/_09_ ;
 wire \u_multiplier/LODy/lod4_3/_10_ ;
 wire \u_multiplier/LODy/lod4_3/_11_ ;
 wire \u_multiplier/LODy/lod4_4/_09_ ;
 wire \u_multiplier/LODy/lod4_4/_10_ ;
 wire \u_multiplier/LODy/lod4_4/_11_ ;
 wire \u_multiplier/LODy/lod4_5/_09_ ;
 wire \u_multiplier/LODy/lod4_5/_10_ ;
 wire \u_multiplier/LODy/lod4_5/_11_ ;
 wire \u_multiplier/LODy/lod4_6/_09_ ;
 wire \u_multiplier/LODy/lod4_6/_10_ ;
 wire \u_multiplier/LODy/lod4_6/_11_ ;
 wire \u_multiplier/LODy/lod4_7/_09_ ;
 wire \u_multiplier/LODy/lod4_7/_10_ ;
 wire \u_multiplier/LODy/lod4_7/_11_ ;
 wire \u_multiplier/LODy/lod4_middle_high/_09_ ;
 wire \u_multiplier/LODy/lod4_middle_high/_10_ ;
 wire \u_multiplier/LODy/lod4_middle_high/_11_ ;
 wire \u_multiplier/LODy/lod4_middle_low/_09_ ;
 wire \u_multiplier/LODy/lod4_middle_low/_10_ ;
 wire \u_multiplier/LODy/lod4_middle_low/_11_ ;
 wire \u_multiplier/NOD/_11_ ;
 wire \u_multiplier/NOD/_12_ ;
 wire \u_multiplier/NOD/_13_ ;
 wire net126;
 wire \u_multiplier/NOD/nod_basic_unit31/_5_ ;
 wire \u_multiplier/NOD/nod_cels[10].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[10].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[10].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[10].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[11].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[11].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[11].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[11].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[12].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[12].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[12].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[12].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[13].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[13].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[13].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[13].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[14].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[14].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[14].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[14].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[15].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[15].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[15].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[15].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[16].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[16].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[16].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[16].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[17].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[17].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[17].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[17].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[18].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[18].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[18].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[18].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[19].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[19].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[19].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[19].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[20].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[20].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[20].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[20].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[21].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[21].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[21].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[21].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[22].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[22].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[22].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[22].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[23].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[23].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[23].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[23].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[24].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[24].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[24].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[24].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[25].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[25].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[25].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[25].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[26].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[26].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[26].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[26].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[27].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[27].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[27].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[27].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[28].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[28].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[28].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[28].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[29].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[29].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[29].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[29].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[2].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[2].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[2].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[2].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[3].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[3].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[3].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[3].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[4].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[4].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[4].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[4].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[5].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[5].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[5].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[5].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[6].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[6].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[6].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[6].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[7].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[7].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[7].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[7].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[8].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[8].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[8].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[8].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[9].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[9].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[9].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[9].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/PE/code0/_31_ ;
 wire \u_multiplier/PE/code0/_32_ ;
 wire \u_multiplier/PE/code0/_33_ ;
 wire \u_multiplier/PE/code0/_34_ ;
 wire \u_multiplier/PE/code0/_35_ ;
 wire \u_multiplier/PE/code1/_31_ ;
 wire \u_multiplier/PE/code1/_32_ ;
 wire \u_multiplier/PE/code1/_33_ ;
 wire \u_multiplier/PE/code1/_34_ ;
 wire \u_multiplier/PE/code1/_35_ ;
 wire \u_multiplier/PE/code2/_31_ ;
 wire \u_multiplier/PE/code2/_32_ ;
 wire \u_multiplier/PE/code2/_33_ ;
 wire \u_multiplier/PE/code2/_34_ ;
 wire \u_multiplier/PE/code2/_35_ ;
 wire \u_multiplier/PE/code3/_31_ ;
 wire \u_multiplier/PE/code3/_32_ ;
 wire \u_multiplier/PE/code3/_33_ ;
 wire \u_multiplier/PE/code3/_34_ ;
 wire \u_multiplier/PE/code3/_35_ ;
 wire \u_multiplier/PE/code4/_31_ ;
 wire \u_multiplier/PE/code4/_32_ ;
 wire \u_multiplier/PE/code4/_33_ ;
 wire \u_multiplier/PE/code4/_34_ ;
 wire \u_multiplier/PE/code4/_35_ ;
 wire \u_multiplier/PEx/code0/_31_ ;
 wire \u_multiplier/PEx/code0/_32_ ;
 wire \u_multiplier/PEx/code0/_33_ ;
 wire \u_multiplier/PEx/code0/_34_ ;
 wire \u_multiplier/PEx/code0/_35_ ;
 wire \u_multiplier/PEx/code1/_31_ ;
 wire \u_multiplier/PEx/code1/_32_ ;
 wire \u_multiplier/PEx/code1/_33_ ;
 wire \u_multiplier/PEx/code1/_34_ ;
 wire \u_multiplier/PEx/code1/_35_ ;
 wire \u_multiplier/PEx/code2/_31_ ;
 wire \u_multiplier/PEx/code2/_32_ ;
 wire \u_multiplier/PEx/code2/_33_ ;
 wire \u_multiplier/PEx/code2/_34_ ;
 wire \u_multiplier/PEx/code2/_35_ ;
 wire \u_multiplier/PEx/code3/_31_ ;
 wire \u_multiplier/PEx/code3/_32_ ;
 wire \u_multiplier/PEx/code3/_33_ ;
 wire \u_multiplier/PEx/code3/_34_ ;
 wire \u_multiplier/PEx/code3/_35_ ;
 wire \u_multiplier/PEx/code4/_31_ ;
 wire \u_multiplier/PEx/code4/_32_ ;
 wire \u_multiplier/PEx/code4/_33_ ;
 wire \u_multiplier/PEx/code4/_34_ ;
 wire \u_multiplier/PEx/code4/_35_ ;
 wire \u_multiplier/PEy/code0/_31_ ;
 wire \u_multiplier/PEy/code0/_32_ ;
 wire \u_multiplier/PEy/code0/_33_ ;
 wire \u_multiplier/PEy/code0/_34_ ;
 wire \u_multiplier/PEy/code0/_35_ ;
 wire \u_multiplier/PEy/code1/_31_ ;
 wire \u_multiplier/PEy/code1/_32_ ;
 wire \u_multiplier/PEy/code1/_33_ ;
 wire \u_multiplier/PEy/code1/_34_ ;
 wire \u_multiplier/PEy/code1/_35_ ;
 wire \u_multiplier/PEy/code2/_31_ ;
 wire \u_multiplier/PEy/code2/_32_ ;
 wire \u_multiplier/PEy/code2/_33_ ;
 wire \u_multiplier/PEy/code2/_34_ ;
 wire \u_multiplier/PEy/code2/_35_ ;
 wire \u_multiplier/PEy/code3/_31_ ;
 wire \u_multiplier/PEy/code3/_32_ ;
 wire \u_multiplier/PEy/code3/_33_ ;
 wire \u_multiplier/PEy/code3/_34_ ;
 wire \u_multiplier/PEy/code3/_35_ ;
 wire \u_multiplier/PEy/code4/_31_ ;
 wire \u_multiplier/PEy/code4/_32_ ;
 wire \u_multiplier/PEy/code4/_33_ ;
 wire \u_multiplier/PEy/code4/_34_ ;
 wire \u_multiplier/PEy/code4/_35_ ;
 wire \u_multiplier/dec/_134_ ;
 wire \u_multiplier/dec/_135_ ;
 wire \u_multiplier/dec/_136_ ;
 wire \u_multiplier/dec/_137_ ;
 wire \u_multiplier/dec/_138_ ;
 wire \u_multiplier/dec/_139_ ;
 wire \u_multiplier/dec/_140_ ;
 wire \u_multiplier/dec/_141_ ;
 wire \u_multiplier/dec/_142_ ;
 wire \u_multiplier/dec/_143_ ;
 wire \u_multiplier/dec/_144_ ;
 wire \u_multiplier/dec/_145_ ;
 wire \u_multiplier/dec/_146_ ;
 wire \u_multiplier/dec/_147_ ;
 wire \u_multiplier/dec/_148_ ;
 wire \u_multiplier/dec/_149_ ;
 wire \u_multiplier/dec/_150_ ;
 wire \u_multiplier/dec/_151_ ;
 wire \u_multiplier/dec/_152_ ;
 wire \u_multiplier/dec/_153_ ;
 wire \u_multiplier/dec/_154_ ;
 wire \u_multiplier/dec/_155_ ;
 wire \u_multiplier/dec/_156_ ;
 wire \u_multiplier/dec/_157_ ;
 wire \u_multiplier/dec/_158_ ;
 wire \u_multiplier/dec/_159_ ;
 wire \u_multiplier/dec/_160_ ;
 wire \u_multiplier/dec/_161_ ;
 wire \u_multiplier/dec/_162_ ;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire valid_reg_out;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire clknet_0_clk;
 wire clknet_1_0_0_clk;
 wire clknet_1_1_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_4_0__leaf_clk;
 wire clknet_4_1__leaf_clk;
 wire clknet_4_2__leaf_clk;
 wire clknet_4_3__leaf_clk;
 wire clknet_4_4__leaf_clk;
 wire clknet_4_5__leaf_clk;
 wire clknet_4_6__leaf_clk;
 wire clknet_4_7__leaf_clk;
 wire clknet_4_8__leaf_clk;
 wire clknet_4_9__leaf_clk;
 wire clknet_4_10__leaf_clk;
 wire clknet_4_11__leaf_clk;
 wire clknet_4_12__leaf_clk;
 wire clknet_4_13__leaf_clk;
 wire clknet_4_14__leaf_clk;
 wire clknet_4_15__leaf_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire [31:0] _0683_;
 wire [5:0] addr_ptr;
 wire [2:0] curr_state;
 wire [24:0] data_in_reg;
 wire [5:0] init_count;
 wire [63:0] product;
 wire [31:0] sram_rdata;
 wire [31:0] sram_rdata_reg;
 wire [4:0] \u_multiplier/K ;
 wire [3:0] \u_multiplier/LODx/select_high ;
 wire [3:0] \u_multiplier/LODx/select_low ;
 wire [31:0] \u_multiplier/LODx/z ;
 wire [3:0] \u_multiplier/LODy/select_high ;
 wire [3:0] \u_multiplier/LODy/select_low ;
 wire [31:0] \u_multiplier/LODy/z ;
 wire [28:0] \u_multiplier/NOD/t_in ;
 wire [31:0] \u_multiplier/NOD_Q1 ;
 wire [4:0] \u_multiplier/code_x ;
 wire [4:0] \u_multiplier/code_y ;
 wire [63:0] \u_multiplier/dec_out ;
 wire [31:0] \u_multiplier/kx ;
 wire [31:0] \u_multiplier/ky ;

 INV_X2 _0684_ (.A(net58),
    .ZN(_0371_));
 INV_X2 _0685_ (.A(net57),
    .ZN(_0308_));
 INV_X1 _0686_ (.A(net12),
    .ZN(_0372_));
 INV_X1 _0687_ (.A(curr_state[2]),
    .ZN(_0373_));
 INV_X1 _0688_ (.A(init_count[4]),
    .ZN(_0374_));
 INV_X1 _0689_ (.A(net59),
    .ZN(_0375_));
 INV_X1 _0690_ (.A(addr_ptr[0]),
    .ZN(_0376_));
 INV_X1 _0691_ (.A(net147),
    .ZN(_0377_));
 AND3_X1 _0692_ (.A1(init_count[1]),
    .A2(init_count[0]),
    .A3(init_count[2]),
    .ZN(_0378_));
 AND4_X1 _0693_ (.A1(init_count[1]),
    .A2(init_count[0]),
    .A3(init_count[3]),
    .A4(init_count[2]),
    .ZN(_0379_));
 NAND4_X4 _0694_ (.A1(init_count[1]),
    .A2(init_count[0]),
    .A3(init_count[3]),
    .A4(init_count[2]),
    .ZN(_0380_));
 AND2_X1 _0695_ (.A1(init_count[5]),
    .A2(init_count[4]),
    .ZN(_0381_));
 NAND2_X1 _0696_ (.A1(init_count[5]),
    .A2(init_count[4]),
    .ZN(_0382_));
 NOR2_X1 _0697_ (.A1(_0380_),
    .A2(_0382_),
    .ZN(_0383_));
 AND2_X1 _0698_ (.A1(net58),
    .A2(net57),
    .ZN(_0384_));
 NAND2_X2 _0699_ (.A1(net58),
    .A2(net57),
    .ZN(_0385_));
 OR2_X1 _0700_ (.A1(net163),
    .A2(_0385_),
    .ZN(_0386_));
 NAND2_X2 _0701_ (.A1(net58),
    .A2(net205),
    .ZN(_0309_));
 NAND3_X1 _0702_ (.A1(net56),
    .A2(net12),
    .A3(_0384_),
    .ZN(_0387_));
 OAI221_X1 _0703_ (.A(_0387_),
    .B1(net164),
    .B2(_0383_),
    .C1(net57),
    .C2(_0309_),
    .ZN(_0307_));
 NOR2_X4 _0704_ (.A1(_0371_),
    .A2(_0375_),
    .ZN(_0304_));
 AND3_X1 _0705_ (.A1(net58),
    .A2(net57),
    .A3(curr_state[2]),
    .ZN(_0388_));
 NAND3_X1 _0706_ (.A1(_0379_),
    .A2(_0381_),
    .A3(_0388_),
    .ZN(_0389_));
 OAI21_X1 _0707_ (.A(_0389_),
    .B1(_0375_),
    .B2(_0371_),
    .ZN(_0306_));
 AOI22_X1 _0708_ (.A1(net58),
    .A2(net13),
    .B1(_0384_),
    .B2(net56),
    .ZN(_0305_));
 AND2_X1 _0709_ (.A1(net58),
    .A2(sram_rdata[0]),
    .ZN(_0272_));
 AND2_X1 _0710_ (.A1(net58),
    .A2(sram_rdata[1]),
    .ZN(_0283_));
 AND2_X1 _0711_ (.A1(net58),
    .A2(sram_rdata[2]),
    .ZN(_0294_));
 AND2_X1 _0712_ (.A1(net58),
    .A2(sram_rdata[3]),
    .ZN(_0297_));
 AND2_X1 _0713_ (.A1(net58),
    .A2(sram_rdata[4]),
    .ZN(_0298_));
 AND2_X1 _0714_ (.A1(net58),
    .A2(sram_rdata[5]),
    .ZN(_0299_));
 AND2_X1 _0715_ (.A1(net58),
    .A2(sram_rdata[6]),
    .ZN(_0300_));
 AND2_X1 _0716_ (.A1(net58),
    .A2(sram_rdata[7]),
    .ZN(_0301_));
 AND2_X1 _0717_ (.A1(net58),
    .A2(sram_rdata[8]),
    .ZN(_0302_));
 AND2_X1 _0718_ (.A1(net58),
    .A2(sram_rdata[9]),
    .ZN(_0303_));
 AND2_X1 _0719_ (.A1(net58),
    .A2(sram_rdata[10]),
    .ZN(_0273_));
 AND2_X1 _0720_ (.A1(net58),
    .A2(sram_rdata[11]),
    .ZN(_0274_));
 AND2_X1 _0721_ (.A1(net58),
    .A2(sram_rdata[12]),
    .ZN(_0275_));
 AND2_X1 _0722_ (.A1(net58),
    .A2(sram_rdata[13]),
    .ZN(_0276_));
 AND2_X1 _0723_ (.A1(net58),
    .A2(sram_rdata[14]),
    .ZN(_0277_));
 AND2_X1 _0724_ (.A1(net58),
    .A2(sram_rdata[15]),
    .ZN(_0278_));
 AND2_X1 _0725_ (.A1(net58),
    .A2(sram_rdata[16]),
    .ZN(_0279_));
 AND2_X1 _0726_ (.A1(net58),
    .A2(sram_rdata[17]),
    .ZN(_0280_));
 AND2_X1 _0727_ (.A1(net58),
    .A2(sram_rdata[18]),
    .ZN(_0281_));
 AND2_X1 _0728_ (.A1(net58),
    .A2(sram_rdata[19]),
    .ZN(_0282_));
 AND2_X1 _0729_ (.A1(net58),
    .A2(sram_rdata[20]),
    .ZN(_0284_));
 AND2_X1 _0730_ (.A1(net58),
    .A2(sram_rdata[21]),
    .ZN(_0285_));
 AND2_X1 _0731_ (.A1(net58),
    .A2(sram_rdata[22]),
    .ZN(_0286_));
 AND2_X1 _0732_ (.A1(net58),
    .A2(sram_rdata[23]),
    .ZN(_0287_));
 AND2_X1 _0733_ (.A1(net58),
    .A2(sram_rdata[24]),
    .ZN(_0288_));
 AND2_X1 _0734_ (.A1(net58),
    .A2(sram_rdata[25]),
    .ZN(_0289_));
 AND2_X1 _0735_ (.A1(net58),
    .A2(sram_rdata[26]),
    .ZN(_0290_));
 AND2_X1 _0736_ (.A1(net58),
    .A2(sram_rdata[27]),
    .ZN(_0291_));
 AND2_X1 _0737_ (.A1(net58),
    .A2(sram_rdata[28]),
    .ZN(_0292_));
 AND2_X1 _0738_ (.A1(net58),
    .A2(sram_rdata[29]),
    .ZN(_0293_));
 AND2_X1 _0739_ (.A1(net58),
    .A2(sram_rdata[30]),
    .ZN(_0295_));
 AND2_X1 _0740_ (.A1(net58),
    .A2(sram_rdata[31]),
    .ZN(_0296_));
 AND2_X1 _0741_ (.A1(product[0]),
    .A2(net23),
    .ZN(_0202_));
 AND2_X1 _0742_ (.A1(product[1]),
    .A2(net23),
    .ZN(_0213_));
 AND2_X1 _0743_ (.A1(product[2]),
    .A2(net22),
    .ZN(_0224_));
 AND2_X1 _0744_ (.A1(product[3]),
    .A2(net23),
    .ZN(_0235_));
 AND2_X1 _0745_ (.A1(product[4]),
    .A2(_0304_),
    .ZN(_0246_));
 AND2_X1 _0746_ (.A1(product[5]),
    .A2(net23),
    .ZN(_0257_));
 AND2_X1 _0747_ (.A1(product[6]),
    .A2(net22),
    .ZN(_0262_));
 AND2_X1 _0748_ (.A1(product[7]),
    .A2(net22),
    .ZN(_0263_));
 AND2_X1 _0749_ (.A1(product[8]),
    .A2(_0304_),
    .ZN(_0264_));
 AND2_X1 _0750_ (.A1(product[9]),
    .A2(_0304_),
    .ZN(_0265_));
 AND2_X1 _0751_ (.A1(product[10]),
    .A2(net23),
    .ZN(_0203_));
 AND2_X1 _0752_ (.A1(product[11]),
    .A2(net22),
    .ZN(_0204_));
 AND2_X1 _0753_ (.A1(product[12]),
    .A2(net22),
    .ZN(_0205_));
 AND2_X1 _0754_ (.A1(product[13]),
    .A2(net23),
    .ZN(_0206_));
 AND2_X1 _0755_ (.A1(product[14]),
    .A2(net22),
    .ZN(_0207_));
 AND2_X1 _0756_ (.A1(product[15]),
    .A2(net23),
    .ZN(_0208_));
 AND2_X1 _0757_ (.A1(product[16]),
    .A2(net23),
    .ZN(_0209_));
 AND2_X1 _0758_ (.A1(product[17]),
    .A2(net23),
    .ZN(_0210_));
 AND2_X1 _0759_ (.A1(product[18]),
    .A2(net22),
    .ZN(_0211_));
 AND2_X1 _0760_ (.A1(product[19]),
    .A2(net22),
    .ZN(_0212_));
 AND2_X1 _0761_ (.A1(product[20]),
    .A2(net23),
    .ZN(_0214_));
 AND2_X1 _0762_ (.A1(product[21]),
    .A2(net22),
    .ZN(_0215_));
 AND2_X1 _0763_ (.A1(product[22]),
    .A2(net22),
    .ZN(_0216_));
 AND2_X1 _0764_ (.A1(product[23]),
    .A2(_0304_),
    .ZN(_0217_));
 AND2_X1 _0765_ (.A1(product[24]),
    .A2(net23),
    .ZN(_0218_));
 AND2_X1 _0766_ (.A1(product[25]),
    .A2(_0304_),
    .ZN(_0219_));
 AND2_X1 _0767_ (.A1(product[26]),
    .A2(net22),
    .ZN(_0220_));
 AND2_X1 _0768_ (.A1(product[27]),
    .A2(net22),
    .ZN(_0221_));
 AND2_X1 _0769_ (.A1(product[28]),
    .A2(net22),
    .ZN(_0222_));
 AND2_X1 _0770_ (.A1(product[29]),
    .A2(net23),
    .ZN(_0223_));
 AND2_X1 _0771_ (.A1(product[30]),
    .A2(net22),
    .ZN(_0225_));
 AND2_X1 _0772_ (.A1(product[31]),
    .A2(net23),
    .ZN(_0226_));
 AND2_X1 _0773_ (.A1(product[32]),
    .A2(net23),
    .ZN(_0227_));
 AND2_X1 _0774_ (.A1(product[33]),
    .A2(net23),
    .ZN(_0228_));
 AND2_X1 _0775_ (.A1(product[34]),
    .A2(net22),
    .ZN(_0229_));
 AND2_X1 _0776_ (.A1(product[35]),
    .A2(net23),
    .ZN(_0230_));
 AND2_X1 _0777_ (.A1(product[36]),
    .A2(net23),
    .ZN(_0231_));
 AND2_X1 _0778_ (.A1(product[37]),
    .A2(net23),
    .ZN(_0232_));
 AND2_X1 _0779_ (.A1(product[38]),
    .A2(net23),
    .ZN(_0233_));
 AND2_X1 _0780_ (.A1(product[39]),
    .A2(_0304_),
    .ZN(_0234_));
 AND2_X1 _0781_ (.A1(product[40]),
    .A2(net23),
    .ZN(_0236_));
 AND2_X1 _0782_ (.A1(product[41]),
    .A2(net23),
    .ZN(_0237_));
 AND2_X1 _0783_ (.A1(product[42]),
    .A2(net23),
    .ZN(_0238_));
 AND2_X1 _0784_ (.A1(product[43]),
    .A2(_0304_),
    .ZN(_0239_));
 AND2_X1 _0785_ (.A1(product[44]),
    .A2(net22),
    .ZN(_0240_));
 AND2_X1 _0786_ (.A1(product[45]),
    .A2(net23),
    .ZN(_0241_));
 AND2_X1 _0787_ (.A1(product[46]),
    .A2(net23),
    .ZN(_0242_));
 AND2_X1 _0788_ (.A1(product[47]),
    .A2(net23),
    .ZN(_0243_));
 AND2_X1 _0789_ (.A1(product[48]),
    .A2(net22),
    .ZN(_0244_));
 AND2_X1 _0790_ (.A1(product[49]),
    .A2(net22),
    .ZN(_0245_));
 AND2_X1 _0791_ (.A1(product[50]),
    .A2(net23),
    .ZN(_0247_));
 AND2_X1 _0792_ (.A1(product[51]),
    .A2(net23),
    .ZN(_0248_));
 AND2_X1 _0793_ (.A1(product[52]),
    .A2(net23),
    .ZN(_0249_));
 AND2_X1 _0794_ (.A1(product[53]),
    .A2(net23),
    .ZN(_0250_));
 AND2_X1 _0795_ (.A1(product[54]),
    .A2(net22),
    .ZN(_0251_));
 AND2_X1 _0796_ (.A1(product[55]),
    .A2(net23),
    .ZN(_0252_));
 AND2_X1 _0797_ (.A1(product[56]),
    .A2(net23),
    .ZN(_0253_));
 AND2_X1 _0798_ (.A1(product[57]),
    .A2(net23),
    .ZN(_0254_));
 AND2_X1 _0799_ (.A1(product[58]),
    .A2(_0304_),
    .ZN(_0255_));
 AND2_X1 _0800_ (.A1(product[59]),
    .A2(net22),
    .ZN(_0256_));
 AND2_X1 _0801_ (.A1(product[60]),
    .A2(net23),
    .ZN(_0258_));
 AND2_X1 _0802_ (.A1(product[61]),
    .A2(net23),
    .ZN(_0259_));
 AND2_X1 _0803_ (.A1(product[62]),
    .A2(net23),
    .ZN(_0260_));
 AND2_X1 _0804_ (.A1(product[63]),
    .A2(net23),
    .ZN(_0261_));
 AND2_X1 _0805_ (.A1(net58),
    .A2(net24),
    .ZN(_0170_));
 AND2_X1 _0806_ (.A1(net58),
    .A2(net35),
    .ZN(_0181_));
 AND2_X1 _0807_ (.A1(net58),
    .A2(net46),
    .ZN(_0192_));
 AND2_X1 _0808_ (.A1(net58),
    .A2(net49),
    .ZN(_0195_));
 AND2_X1 _0809_ (.A1(net58),
    .A2(net50),
    .ZN(_0196_));
 AND2_X1 _0810_ (.A1(net58),
    .A2(net51),
    .ZN(_0197_));
 AND2_X1 _0811_ (.A1(net58),
    .A2(net52),
    .ZN(_0198_));
 AND2_X1 _0812_ (.A1(net58),
    .A2(net53),
    .ZN(_0199_));
 AND2_X1 _0813_ (.A1(net58),
    .A2(net54),
    .ZN(_0200_));
 AND2_X1 _0814_ (.A1(net58),
    .A2(net55),
    .ZN(_0201_));
 AND2_X1 _0815_ (.A1(net58),
    .A2(net25),
    .ZN(_0171_));
 AND2_X1 _0816_ (.A1(net58),
    .A2(net26),
    .ZN(_0172_));
 AND2_X1 _0817_ (.A1(net58),
    .A2(net27),
    .ZN(_0173_));
 AND2_X1 _0818_ (.A1(net58),
    .A2(net28),
    .ZN(_0174_));
 AND2_X1 _0819_ (.A1(net58),
    .A2(net29),
    .ZN(_0175_));
 AND2_X1 _0820_ (.A1(net58),
    .A2(net30),
    .ZN(_0176_));
 AND2_X1 _0821_ (.A1(net58),
    .A2(net31),
    .ZN(_0177_));
 AND2_X2 _0822_ (.A1(net58),
    .A2(net32),
    .ZN(_0178_));
 AND2_X1 _0823_ (.A1(net58),
    .A2(net33),
    .ZN(_0179_));
 AND2_X1 _0824_ (.A1(net58),
    .A2(net34),
    .ZN(_0180_));
 AND2_X1 _0825_ (.A1(net58),
    .A2(net36),
    .ZN(_0182_));
 AND2_X1 _0826_ (.A1(net58),
    .A2(net37),
    .ZN(_0183_));
 AND2_X1 _0827_ (.A1(net58),
    .A2(net38),
    .ZN(_0184_));
 AND2_X1 _0828_ (.A1(net58),
    .A2(net39),
    .ZN(_0185_));
 AND2_X1 _0829_ (.A1(net58),
    .A2(net40),
    .ZN(_0186_));
 AND2_X2 _0830_ (.A1(net58),
    .A2(net41),
    .ZN(_0187_));
 AND2_X2 _0831_ (.A1(net58),
    .A2(net42),
    .ZN(_0188_));
 AND2_X1 _0832_ (.A1(net58),
    .A2(net43),
    .ZN(_0189_));
 AND2_X1 _0833_ (.A1(net58),
    .A2(net44),
    .ZN(_0190_));
 AND2_X1 _0834_ (.A1(net58),
    .A2(net45),
    .ZN(_0191_));
 AND2_X1 _0835_ (.A1(net58),
    .A2(net47),
    .ZN(_0193_));
 AND2_X1 _0836_ (.A1(net58),
    .A2(net48),
    .ZN(_0194_));
 NAND2_X4 _0837_ (.A1(net58),
    .A2(_0308_),
    .ZN(_0390_));
 AND2_X1 _0838_ (.A1(_0389_),
    .A2(_0390_),
    .ZN(_0391_));
 AOI21_X2 _0839_ (.A(_0373_),
    .B1(_0379_),
    .B2(_0381_),
    .ZN(_0392_));
 OAI21_X1 _0840_ (.A(curr_state[2]),
    .B1(_0380_),
    .B2(_0382_),
    .ZN(_0393_));
 AOI22_X1 _0841_ (.A1(init_count[0]),
    .A2(net59),
    .B1(net167),
    .B2(_0392_),
    .ZN(_0394_));
 OAI22_X1 _0842_ (.A1(net168),
    .A2(_0391_),
    .B1(_0394_),
    .B2(_0385_),
    .ZN(_0266_));
 AND2_X1 _0843_ (.A1(net59),
    .A2(_0384_),
    .ZN(_0395_));
 NAND2_X1 _0844_ (.A1(init_count[1]),
    .A2(_0395_),
    .ZN(_0396_));
 XOR2_X1 _0845_ (.A(init_count[1]),
    .B(init_count[0]),
    .Z(_0397_));
 OAI21_X1 _0846_ (.A(_0388_),
    .B1(_0397_),
    .B2(_0383_),
    .ZN(_0398_));
 OAI211_X1 _0847_ (.A(_0396_),
    .B(_0398_),
    .C1(net180),
    .C2(_0390_),
    .ZN(_0267_));
 AOI21_X1 _0848_ (.A(init_count[2]),
    .B1(init_count[0]),
    .B2(init_count[1]),
    .ZN(_0399_));
 NAND2_X1 _0849_ (.A1(init_count[2]),
    .A2(_0395_),
    .ZN(_0400_));
 OAI22_X1 _0850_ (.A1(_0380_),
    .A2(_0382_),
    .B1(_0399_),
    .B2(_0378_),
    .ZN(_0401_));
 NAND2_X1 _0851_ (.A1(_0388_),
    .A2(_0401_),
    .ZN(_0402_));
 OAI211_X1 _0852_ (.A(_0400_),
    .B(_0402_),
    .C1(net177),
    .C2(_0390_),
    .ZN(_0268_));
 NAND2_X1 _0853_ (.A1(_0379_),
    .A2(_0382_),
    .ZN(_0403_));
 OAI211_X1 _0854_ (.A(_0388_),
    .B(_0403_),
    .C1(init_count[3]),
    .C2(_0378_),
    .ZN(_0404_));
 NAND2_X1 _0855_ (.A1(init_count[3]),
    .A2(_0395_),
    .ZN(_0405_));
 OAI211_X1 _0856_ (.A(_0404_),
    .B(_0405_),
    .C1(net174),
    .C2(_0390_),
    .ZN(_0269_));
 OR3_X1 _0857_ (.A1(init_count[5]),
    .A2(_0374_),
    .A3(_0380_),
    .ZN(_0406_));
 AOI21_X1 _0858_ (.A(_0373_),
    .B1(_0374_),
    .B2(_0380_),
    .ZN(_0407_));
 AOI22_X1 _0859_ (.A1(init_count[4]),
    .A2(net59),
    .B1(_0406_),
    .B2(_0407_),
    .ZN(_0408_));
 OAI22_X1 _0860_ (.A1(net10),
    .A2(_0390_),
    .B1(_0408_),
    .B2(_0385_),
    .ZN(_0270_));
 NAND2_X1 _0861_ (.A1(net224),
    .A2(_0395_),
    .ZN(_0409_));
 OAI21_X1 _0862_ (.A(net157),
    .B1(_0380_),
    .B2(net9),
    .ZN(_0410_));
 NAND2_X1 _0863_ (.A1(_0388_),
    .A2(_0410_),
    .ZN(_0411_));
 OAI211_X1 _0864_ (.A(_0409_),
    .B(_0411_),
    .C1(net158),
    .C2(_0390_),
    .ZN(_0271_));
 AOI22_X1 _0865_ (.A1(net59),
    .A2(_0376_),
    .B1(net160),
    .B2(_0392_),
    .ZN(_0412_));
 OAI22_X1 _0866_ (.A1(net161),
    .A2(_0390_),
    .B1(_0412_),
    .B2(_0385_),
    .ZN(_0164_));
 NAND2_X1 _0867_ (.A1(addr_ptr[0]),
    .A2(addr_ptr[1]),
    .ZN(_0413_));
 OR2_X1 _0868_ (.A1(addr_ptr[0]),
    .A2(addr_ptr[1]),
    .ZN(_0414_));
 OAI211_X1 _0869_ (.A(_0413_),
    .B(_0414_),
    .C1(net59),
    .C2(_0392_),
    .ZN(_0415_));
 OAI22_X1 _0870_ (.A1(net126),
    .A2(_0390_),
    .B1(_0415_),
    .B2(_0385_),
    .ZN(_0165_));
 NAND4_X2 _0871_ (.A1(addr_ptr[0]),
    .A2(addr_ptr[1]),
    .A3(addr_ptr[3]),
    .A4(addr_ptr[2]),
    .ZN(_0416_));
 NAND2_X1 _0872_ (.A1(addr_ptr[5]),
    .A2(addr_ptr[4]),
    .ZN(_0417_));
 OAI21_X1 _0873_ (.A(net59),
    .B1(_0416_),
    .B2(_0417_),
    .ZN(_0418_));
 AND2_X1 _0874_ (.A1(_0393_),
    .A2(_0418_),
    .ZN(_0419_));
 AOI21_X1 _0875_ (.A(_0385_),
    .B1(_0413_),
    .B2(net192),
    .ZN(_0420_));
 OAI21_X1 _0876_ (.A(_0420_),
    .B1(_0413_),
    .B2(net192),
    .ZN(_0421_));
 OAI22_X1 _0877_ (.A1(net193),
    .A2(_0390_),
    .B1(_0419_),
    .B2(_0421_),
    .ZN(_0166_));
 NOR3_X1 _0878_ (.A1(_0308_),
    .A2(net192),
    .A3(_0413_),
    .ZN(_0422_));
 OAI21_X1 _0879_ (.A(net58),
    .B1(_0377_),
    .B2(_0422_),
    .ZN(_0423_));
 AOI221_X1 _0880_ (.A(_0423_),
    .B1(_0422_),
    .B2(_0377_),
    .C1(net57),
    .C2(_0419_),
    .ZN(_0167_));
 NOR3_X1 _0881_ (.A1(_0308_),
    .A2(net153),
    .A3(_0416_),
    .ZN(_0424_));
 OAI21_X1 _0882_ (.A(net153),
    .B1(_0416_),
    .B2(_0308_),
    .ZN(_0425_));
 NAND2_X1 _0883_ (.A1(net58),
    .A2(net154),
    .ZN(_0426_));
 AOI211_X1 _0884_ (.A(_0424_),
    .B(_0426_),
    .C1(net57),
    .C2(_0419_),
    .ZN(_0168_));
 XOR2_X1 _0885_ (.A(net14),
    .B(_0424_),
    .Z(_0427_));
 AOI211_X1 _0886_ (.A(_0371_),
    .B(net15),
    .C1(_0419_),
    .C2(net57),
    .ZN(_0169_));
 DFF_X1 _0887_ (.D(_0202_),
    .CK(clknet_4_12__leaf_clk),
    .Q(net60),
    .QN(_0526_));
 DFF_X1 _0888_ (.D(_0213_),
    .CK(clknet_4_11__leaf_clk),
    .Q(net71),
    .QN(_0527_));
 DFF_X2 _0889_ (.D(_0224_),
    .CK(clknet_4_11__leaf_clk),
    .Q(net82),
    .QN(_0528_));
 DFF_X1 _0890_ (.D(_0235_),
    .CK(clknet_4_15__leaf_clk),
    .Q(net93),
    .QN(_0529_));
 DFF_X2 _0891_ (.D(_0246_),
    .CK(clknet_4_1__leaf_clk),
    .Q(net104),
    .QN(_0530_));
 DFF_X1 _0892_ (.D(_0257_),
    .CK(clknet_4_1__leaf_clk),
    .Q(net115),
    .QN(_0531_));
 DFF_X2 _0893_ (.D(_0262_),
    .CK(clknet_4_13__leaf_clk),
    .Q(net120),
    .QN(_0532_));
 DFF_X2 _0894_ (.D(_0263_),
    .CK(clknet_4_13__leaf_clk),
    .Q(net121),
    .QN(_0533_));
 DFF_X2 _0895_ (.D(_0264_),
    .CK(clknet_4_5__leaf_clk),
    .Q(net122),
    .QN(_0534_));
 DFF_X2 _0896_ (.D(_0265_),
    .CK(clknet_4_4__leaf_clk),
    .Q(net123),
    .QN(_0535_));
 DFF_X2 _0897_ (.D(_0203_),
    .CK(clknet_4_11__leaf_clk),
    .Q(net61),
    .QN(_0536_));
 DFF_X2 _0898_ (.D(_0204_),
    .CK(clknet_4_7__leaf_clk),
    .Q(net62),
    .QN(_0537_));
 DFF_X2 _0899_ (.D(_0205_),
    .CK(clknet_4_7__leaf_clk),
    .Q(net63),
    .QN(_0538_));
 DFF_X1 _0900_ (.D(_0206_),
    .CK(clknet_4_8__leaf_clk),
    .Q(net64),
    .QN(_0539_));
 DFF_X1 _0901_ (.D(_0207_),
    .CK(clknet_4_1__leaf_clk),
    .Q(net65),
    .QN(_0540_));
 DFF_X2 _0902_ (.D(_0208_),
    .CK(clknet_4_11__leaf_clk),
    .Q(net66),
    .QN(_0541_));
 DFF_X1 _0903_ (.D(_0209_),
    .CK(clknet_4_11__leaf_clk),
    .Q(net67),
    .QN(_0542_));
 DFF_X1 _0904_ (.D(_0210_),
    .CK(clknet_4_15__leaf_clk),
    .Q(net68),
    .QN(_0543_));
 DFF_X2 _0905_ (.D(_0211_),
    .CK(clknet_4_9__leaf_clk),
    .Q(net69),
    .QN(_0544_));
 DFF_X2 _0906_ (.D(_0212_),
    .CK(clknet_4_6__leaf_clk),
    .Q(net70),
    .QN(_0545_));
 DFF_X2 _0907_ (.D(_0214_),
    .CK(clknet_4_12__leaf_clk),
    .Q(net72),
    .QN(_0546_));
 DFF_X2 _0908_ (.D(_0215_),
    .CK(clknet_4_14__leaf_clk),
    .Q(net73),
    .QN(_0547_));
 DFF_X2 _0909_ (.D(_0216_),
    .CK(clknet_4_6__leaf_clk),
    .Q(net74),
    .QN(_0548_));
 DFF_X2 _0910_ (.D(_0217_),
    .CK(clknet_4_4__leaf_clk),
    .Q(net75),
    .QN(_0549_));
 DFF_X1 _0911_ (.D(_0218_),
    .CK(clknet_4_12__leaf_clk),
    .Q(net76),
    .QN(_0550_));
 DFF_X2 _0912_ (.D(_0219_),
    .CK(clknet_4_4__leaf_clk),
    .Q(net77),
    .QN(_0551_));
 DFF_X2 _0913_ (.D(_0220_),
    .CK(clknet_4_1__leaf_clk),
    .Q(net78),
    .QN(_0552_));
 DFF_X2 _0914_ (.D(_0221_),
    .CK(clknet_4_8__leaf_clk),
    .Q(net79),
    .QN(_0553_));
 DFF_X2 _0915_ (.D(_0222_),
    .CK(clknet_4_1__leaf_clk),
    .Q(net80),
    .QN(_0554_));
 DFF_X1 _0916_ (.D(_0223_),
    .CK(clknet_4_10__leaf_clk),
    .Q(net81),
    .QN(_0555_));
 DFF_X2 _0917_ (.D(_0225_),
    .CK(clknet_4_1__leaf_clk),
    .Q(net83),
    .QN(_0556_));
 DFF_X2 _0918_ (.D(_0226_),
    .CK(clknet_4_1__leaf_clk),
    .Q(net84),
    .QN(_0557_));
 DFF_X1 _0919_ (.D(_0227_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net85),
    .QN(_0558_));
 DFF_X1 _0920_ (.D(_0228_),
    .CK(clknet_4_10__leaf_clk),
    .Q(net86),
    .QN(_0559_));
 DFF_X1 _0921_ (.D(_0229_),
    .CK(clknet_4_15__leaf_clk),
    .Q(net87),
    .QN(_0560_));
 DFF_X1 _0922_ (.D(_0230_),
    .CK(clknet_4_12__leaf_clk),
    .Q(net88),
    .QN(_0561_));
 DFF_X2 _0923_ (.D(_0231_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net89),
    .QN(_0562_));
 DFF_X2 _0924_ (.D(_0232_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net90),
    .QN(_0563_));
 DFF_X1 _0925_ (.D(_0233_),
    .CK(clknet_4_10__leaf_clk),
    .Q(net91),
    .QN(_0564_));
 DFF_X2 _0926_ (.D(_0234_),
    .CK(clknet_4_4__leaf_clk),
    .Q(net92),
    .QN(_0565_));
 DFF_X2 _0927_ (.D(_0236_),
    .CK(clknet_4_10__leaf_clk),
    .Q(net94),
    .QN(_0566_));
 DFF_X1 _0928_ (.D(_0237_),
    .CK(clknet_4_11__leaf_clk),
    .Q(net95),
    .QN(_0567_));
 DFF_X2 _0929_ (.D(_0238_),
    .CK(clknet_4_10__leaf_clk),
    .Q(net96),
    .QN(_0568_));
 DFF_X2 _0930_ (.D(_0239_),
    .CK(clknet_4_1__leaf_clk),
    .Q(net97),
    .QN(_0569_));
 DFF_X2 _0931_ (.D(_0240_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net98),
    .QN(_0570_));
 DFF_X2 _0932_ (.D(_0241_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net99),
    .QN(_0571_));
 DFF_X1 _0933_ (.D(_0242_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net100),
    .QN(_0572_));
 DFF_X1 _0934_ (.D(_0243_),
    .CK(clknet_4_8__leaf_clk),
    .Q(net101),
    .QN(_0573_));
 DFF_X2 _0935_ (.D(_0244_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net102),
    .QN(_0574_));
 DFF_X2 _0936_ (.D(_0245_),
    .CK(clknet_4_1__leaf_clk),
    .Q(net103),
    .QN(_0575_));
 DFF_X2 _0937_ (.D(_0247_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net105),
    .QN(_0576_));
 DFF_X1 _0938_ (.D(_0248_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net106),
    .QN(_0577_));
 DFF_X1 _0939_ (.D(_0249_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net107),
    .QN(_0578_));
 DFF_X2 _0940_ (.D(_0250_),
    .CK(clknet_4_10__leaf_clk),
    .Q(net108),
    .QN(_0579_));
 DFF_X2 _0941_ (.D(_0251_),
    .CK(clknet_4_9__leaf_clk),
    .Q(net109),
    .QN(_0580_));
 DFF_X1 _0942_ (.D(_0252_),
    .CK(clknet_4_2__leaf_clk),
    .Q(net110),
    .QN(_0581_));
 DFF_X2 _0943_ (.D(_0253_),
    .CK(clknet_4_10__leaf_clk),
    .Q(net111),
    .QN(_0582_));
 DFF_X1 _0944_ (.D(_0254_),
    .CK(clknet_4_10__leaf_clk),
    .Q(net112),
    .QN(_0583_));
 DFF_X2 _0945_ (.D(_0255_),
    .CK(clknet_4_4__leaf_clk),
    .Q(net113),
    .QN(_0584_));
 DFF_X2 _0946_ (.D(_0256_),
    .CK(clknet_4_15__leaf_clk),
    .Q(net114),
    .QN(_0585_));
 DFF_X1 _0947_ (.D(_0258_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net116),
    .QN(_0586_));
 DFF_X2 _0948_ (.D(_0259_),
    .CK(clknet_4_7__leaf_clk),
    .Q(net117),
    .QN(_0587_));
 DFF_X2 _0949_ (.D(_0260_),
    .CK(clknet_4_10__leaf_clk),
    .Q(net118),
    .QN(_0588_));
 DFF_X1 _0950_ (.D(_0261_),
    .CK(clknet_4_2__leaf_clk),
    .Q(net119),
    .QN(_0589_));
 DFF_X1 _0951_ (.D(_0305_),
    .CK(clknet_4_5__leaf_clk),
    .Q(curr_state[0]),
    .QN(_0590_));
 DFF_X2 _0952_ (.D(_0306_),
    .CK(clknet_4_5__leaf_clk),
    .Q(net59),
    .QN(_0591_));
 DFF_X2 _0953_ (.D(net165),
    .CK(clknet_4_5__leaf_clk),
    .Q(curr_state[2]),
    .QN(_0592_));
 DFF_X2 _0954_ (.D(_0170_),
    .CK(clknet_4_9__leaf_clk),
    .Q(data_in_reg[0]),
    .QN(_0593_));
 DFF_X2 _0955_ (.D(_0181_),
    .CK(clknet_4_7__leaf_clk),
    .Q(data_in_reg[1]),
    .QN(_0594_));
 DFF_X2 _0956_ (.D(_0192_),
    .CK(clknet_4_13__leaf_clk),
    .Q(data_in_reg[2]),
    .QN(_0595_));
 DFF_X2 _0957_ (.D(_0195_),
    .CK(clknet_4_8__leaf_clk),
    .Q(\u_multiplier/LODx/z [3]),
    .QN(_0596_));
 DFF_X2 _0958_ (.D(_0196_),
    .CK(clknet_4_6__leaf_clk),
    .Q(data_in_reg[4]),
    .QN(_0597_));
 DFF_X2 _0959_ (.D(_0197_),
    .CK(clknet_4_14__leaf_clk),
    .Q(data_in_reg[5]),
    .QN(_0598_));
 DFF_X2 _0960_ (.D(_0198_),
    .CK(clknet_4_2__leaf_clk),
    .Q(data_in_reg[6]),
    .QN(_0599_));
 DFF_X2 _0961_ (.D(_0199_),
    .CK(clknet_4_1__leaf_clk),
    .Q(\u_multiplier/LODx/z [7]),
    .QN(_0600_));
 DFF_X2 _0962_ (.D(_0200_),
    .CK(clknet_4_14__leaf_clk),
    .Q(data_in_reg[8]),
    .QN(_0601_));
 DFF_X2 _0963_ (.D(_0201_),
    .CK(clknet_4_3__leaf_clk),
    .Q(data_in_reg[9]),
    .QN(_0602_));
 DFF_X2 _0964_ (.D(_0171_),
    .CK(clknet_4_11__leaf_clk),
    .Q(data_in_reg[10]),
    .QN(_0603_));
 DFF_X2 _0965_ (.D(_0172_),
    .CK(clknet_4_1__leaf_clk),
    .Q(\u_multiplier/LODx/z [11]),
    .QN(_0604_));
 DFF_X2 _0966_ (.D(_0173_),
    .CK(clknet_4_13__leaf_clk),
    .Q(data_in_reg[12]),
    .QN(_0605_));
 DFF_X2 _0967_ (.D(_0174_),
    .CK(clknet_4_7__leaf_clk),
    .Q(data_in_reg[13]),
    .QN(_0606_));
 DFF_X2 _0968_ (.D(_0175_),
    .CK(clknet_4_12__leaf_clk),
    .Q(data_in_reg[14]),
    .QN(_0607_));
 DFF_X2 _0969_ (.D(_0176_),
    .CK(clknet_4_10__leaf_clk),
    .Q(\u_multiplier/LODx/z [15]),
    .QN(_0608_));
 DFF_X2 _0970_ (.D(_0177_),
    .CK(clknet_4_1__leaf_clk),
    .Q(data_in_reg[16]),
    .QN(_0609_));
 DFF_X2 _0971_ (.D(_0178_),
    .CK(clknet_4_8__leaf_clk),
    .Q(data_in_reg[17]),
    .QN(_0610_));
 DFF_X2 _0972_ (.D(_0179_),
    .CK(clknet_4_7__leaf_clk),
    .Q(data_in_reg[18]),
    .QN(_0611_));
 DFF_X2 _0973_ (.D(_0180_),
    .CK(clknet_4_9__leaf_clk),
    .Q(\u_multiplier/LODx/z [19]),
    .QN(_0612_));
 DFF_X2 _0974_ (.D(_0182_),
    .CK(clknet_4_8__leaf_clk),
    .Q(data_in_reg[20]),
    .QN(_0613_));
 DFF_X2 _0975_ (.D(_0183_),
    .CK(clknet_4_9__leaf_clk),
    .Q(data_in_reg[21]),
    .QN(_0614_));
 DFF_X2 _0976_ (.D(_0184_),
    .CK(clknet_4_12__leaf_clk),
    .Q(data_in_reg[22]),
    .QN(_0615_));
 DFF_X2 _0977_ (.D(_0185_),
    .CK(clknet_4_9__leaf_clk),
    .Q(\u_multiplier/LODx/z [23]),
    .QN(_0616_));
 DFF_X2 _0978_ (.D(_0186_),
    .CK(clknet_4_13__leaf_clk),
    .Q(data_in_reg[24]),
    .QN(_0617_));
 DFF_X2 _0979_ (.D(_0187_),
    .CK(clknet_4_11__leaf_clk),
    .Q(_0683_[25]),
    .QN(_0618_));
 DFF_X2 _0980_ (.D(_0188_),
    .CK(clknet_4_13__leaf_clk),
    .Q(_0683_[26]),
    .QN(_0619_));
 DFF_X2 _0981_ (.D(_0189_),
    .CK(clknet_4_13__leaf_clk),
    .Q(\u_multiplier/LODx/z [27]),
    .QN(_0620_));
 DFF_X2 _0982_ (.D(_0190_),
    .CK(clknet_4_10__leaf_clk),
    .Q(_0683_[28]),
    .QN(_0621_));
 DFF_X2 _0983_ (.D(_0191_),
    .CK(clknet_4_10__leaf_clk),
    .Q(_0683_[29]),
    .QN(_0622_));
 DFF_X2 _0984_ (.D(_0193_),
    .CK(clknet_4_1__leaf_clk),
    .Q(_0683_[30]),
    .QN(_0623_));
 DFF_X2 _0985_ (.D(_0194_),
    .CK(clknet_4_14__leaf_clk),
    .Q(\u_multiplier/LODx/z [31]),
    .QN(_0624_));
 DFF_X2 _0986_ (.D(_0272_),
    .CK(clknet_4_6__leaf_clk),
    .Q(sram_rdata_reg[0]),
    .QN(_0625_));
 DFF_X2 _0987_ (.D(_0283_),
    .CK(clknet_4_6__leaf_clk),
    .Q(sram_rdata_reg[1]),
    .QN(_0626_));
 DFF_X2 _0988_ (.D(_0294_),
    .CK(clknet_4_6__leaf_clk),
    .Q(sram_rdata_reg[2]),
    .QN(_0627_));
 DFF_X2 _0989_ (.D(_0297_),
    .CK(clknet_4_6__leaf_clk),
    .Q(\u_multiplier/LODy/z [3]),
    .QN(_0628_));
 DFF_X2 _0990_ (.D(_0298_),
    .CK(clknet_4_6__leaf_clk),
    .Q(sram_rdata_reg[4]),
    .QN(_0629_));
 DFF_X2 _0991_ (.D(_0299_),
    .CK(clknet_4_3__leaf_clk),
    .Q(sram_rdata_reg[5]),
    .QN(_0630_));
 DFF_X2 _0992_ (.D(_0300_),
    .CK(clknet_4_3__leaf_clk),
    .Q(sram_rdata_reg[6]),
    .QN(_0631_));
 DFF_X2 _0993_ (.D(_0301_),
    .CK(clknet_4_3__leaf_clk),
    .Q(\u_multiplier/LODy/z [7]),
    .QN(_0632_));
 DFF_X2 _0994_ (.D(_0302_),
    .CK(clknet_4_3__leaf_clk),
    .Q(sram_rdata_reg[8]),
    .QN(_0633_));
 DFF_X2 _0995_ (.D(_0303_),
    .CK(clknet_4_3__leaf_clk),
    .Q(sram_rdata_reg[9]),
    .QN(_0634_));
 DFF_X2 _0996_ (.D(_0273_),
    .CK(clknet_4_3__leaf_clk),
    .Q(sram_rdata_reg[10]),
    .QN(_0635_));
 DFF_X2 _0997_ (.D(_0274_),
    .CK(clknet_4_3__leaf_clk),
    .Q(\u_multiplier/LODy/z [11]),
    .QN(_0636_));
 DFF_X2 _0998_ (.D(_0275_),
    .CK(clknet_4_2__leaf_clk),
    .Q(sram_rdata_reg[12]),
    .QN(_0637_));
 DFF_X2 _0999_ (.D(_0276_),
    .CK(clknet_4_3__leaf_clk),
    .Q(sram_rdata_reg[13]),
    .QN(_0638_));
 DFF_X2 _1000_ (.D(_0277_),
    .CK(clknet_4_2__leaf_clk),
    .Q(sram_rdata_reg[14]),
    .QN(_0639_));
 DFF_X2 _1001_ (.D(_0278_),
    .CK(clknet_4_2__leaf_clk),
    .Q(\u_multiplier/LODy/z [15]),
    .QN(_0640_));
 DFF_X2 _1002_ (.D(_0279_),
    .CK(clknet_4_3__leaf_clk),
    .Q(sram_rdata_reg[16]),
    .QN(_0641_));
 DFF_X2 _1003_ (.D(_0280_),
    .CK(clknet_4_2__leaf_clk),
    .Q(sram_rdata_reg[17]),
    .QN(_0642_));
 DFF_X2 _1004_ (.D(_0281_),
    .CK(clknet_4_2__leaf_clk),
    .Q(sram_rdata_reg[18]),
    .QN(_0643_));
 DFF_X2 _1005_ (.D(_0282_),
    .CK(clknet_4_2__leaf_clk),
    .Q(\u_multiplier/LODy/z [19]),
    .QN(_0644_));
 DFF_X2 _1006_ (.D(_0284_),
    .CK(clknet_4_2__leaf_clk),
    .Q(sram_rdata_reg[20]),
    .QN(_0645_));
 DFF_X2 _1007_ (.D(_0285_),
    .CK(clknet_4_2__leaf_clk),
    .Q(sram_rdata_reg[21]),
    .QN(_0646_));
 DFF_X2 _1008_ (.D(_0286_),
    .CK(clknet_4_3__leaf_clk),
    .Q(sram_rdata_reg[22]),
    .QN(_0647_));
 DFF_X2 _1009_ (.D(_0287_),
    .CK(clknet_4_2__leaf_clk),
    .Q(\u_multiplier/LODy/z [23]),
    .QN(_0648_));
 DFF_X2 _1010_ (.D(_0288_),
    .CK(clknet_4_3__leaf_clk),
    .Q(sram_rdata_reg[24]),
    .QN(_0649_));
 DFF_X2 _1011_ (.D(_0289_),
    .CK(clknet_4_3__leaf_clk),
    .Q(sram_rdata_reg[25]),
    .QN(_0650_));
 DFF_X2 _1012_ (.D(_0290_),
    .CK(clknet_4_3__leaf_clk),
    .Q(sram_rdata_reg[26]),
    .QN(_0651_));
 DFF_X2 _1013_ (.D(_0291_),
    .CK(clknet_4_3__leaf_clk),
    .Q(\u_multiplier/LODy/z [27]),
    .QN(_0652_));
 DFF_X2 _1014_ (.D(_0292_),
    .CK(clknet_4_9__leaf_clk),
    .Q(sram_rdata_reg[28]),
    .QN(_0653_));
 DFF_X2 _1015_ (.D(_0293_),
    .CK(clknet_4_3__leaf_clk),
    .Q(sram_rdata_reg[29]),
    .QN(_0654_));
 DFF_X2 _1016_ (.D(_0295_),
    .CK(clknet_4_9__leaf_clk),
    .Q(sram_rdata_reg[30]),
    .QN(_0655_));
 DFF_X2 _1017_ (.D(_0296_),
    .CK(clknet_4_9__leaf_clk),
    .Q(\u_multiplier/LODy/z [31]),
    .QN(_0656_));
 DFF_X1 _1018_ (.D(net22),
    .CK(clknet_4_15__leaf_clk),
    .Q(net124),
    .QN(_0657_));
 DFF_X2 _1019_ (.D(net162),
    .CK(clknet_4_5__leaf_clk),
    .Q(addr_ptr[0]),
    .QN(_0658_));
 DFF_X1 _1020_ (.D(net127),
    .CK(clknet_4_4__leaf_clk),
    .Q(addr_ptr[1]),
    .QN(_0659_));
 DFF_X1 _1021_ (.D(_0166_),
    .CK(clknet_4_4__leaf_clk),
    .Q(addr_ptr[2]),
    .QN(_0660_));
 DFF_X1 _1022_ (.D(_0167_),
    .CK(clknet_4_5__leaf_clk),
    .Q(addr_ptr[3]),
    .QN(_0661_));
 DFF_X1 _1023_ (.D(_0168_),
    .CK(clknet_4_5__leaf_clk),
    .Q(addr_ptr[4]),
    .QN(_0662_));
 DFF_X1 _1024_ (.D(_0169_),
    .CK(clknet_4_5__leaf_clk),
    .Q(addr_ptr[5]),
    .QN(_0663_));
 DFF_X2 _1025_ (.D(net169),
    .CK(clknet_4_4__leaf_clk),
    .Q(init_count[0]),
    .QN(_0664_));
 DFF_X2 _1026_ (.D(net181),
    .CK(clknet_4_5__leaf_clk),
    .Q(init_count[1]),
    .QN(_0665_));
 DFF_X2 _1027_ (.D(net178),
    .CK(clknet_4_5__leaf_clk),
    .Q(init_count[2]),
    .QN(_0666_));
 DFF_X2 _1028_ (.D(net175),
    .CK(clknet_4_4__leaf_clk),
    .Q(init_count[3]),
    .QN(_0667_));
 DFF_X1 _1029_ (.D(net11),
    .CK(clknet_4_5__leaf_clk),
    .Q(init_count[4]),
    .QN(_0668_));
 DFF_X1 _1030_ (.D(net159),
    .CK(clknet_4_5__leaf_clk),
    .Q(init_count[5]),
    .QN(_0669_));
 SRAM_6T_CORE_64x32_MC_TB sram_inst (.ce_in(_0308_),
    .we_in(_0309_),
    .clk(clknet_4_7__leaf_clk),
    .addr_in({net190,
    net185,
    net197,
    net195,
    net139,
    net141}),
    .rd_out({sram_rdata[31],
    sram_rdata[30],
    sram_rdata[29],
    sram_rdata[28],
    sram_rdata[27],
    sram_rdata[26],
    sram_rdata[25],
    sram_rdata[24],
    sram_rdata[23],
    sram_rdata[22],
    sram_rdata[21],
    sram_rdata[20],
    sram_rdata[19],
    sram_rdata[18],
    sram_rdata[17],
    sram_rdata[16],
    sram_rdata[15],
    sram_rdata[14],
    sram_rdata[13],
    sram_rdata[12],
    sram_rdata[11],
    sram_rdata[10],
    sram_rdata[9],
    sram_rdata[8],
    sram_rdata[7],
    sram_rdata[6],
    sram_rdata[5],
    sram_rdata[4],
    sram_rdata[3],
    sram_rdata[2],
    sram_rdata[1],
    sram_rdata[0]}),
    .wd_in({net144,
    net206,
    net171,
    net149,
    net1,
    net148,
    net145,
    net199,
    net150,
    net4,
    net146,
    net142,
    net16,
    net166,
    net172,
    net191,
    net188,
    net3,
    net170,
    net151,
    net183,
    net187,
    net152,
    net5,
    net156,
    net182,
    net8,
    net2,
    net186,
    net6,
    net7,
    net155}));
 AND2_X1 \u_multiplier/LODx/Inst_MUX214_0/_09_  (.A1(\u_multiplier/LODx/z [1]),
    .A2(\u_multiplier/LODx/_061_ ),
    .ZN(\u_multiplier/kx [1]));
 AND2_X1 \u_multiplier/LODx/Inst_MUX214_0/_10_  (.A1(\u_multiplier/LODx/_061_ ),
    .A2(\u_multiplier/LODx/z [0]),
    .ZN(\u_multiplier/kx [0]));
 AND2_X1 \u_multiplier/LODx/Inst_MUX214_0/_11_  (.A1(\u_multiplier/LODx/_061_ ),
    .A2(\u_multiplier/LODx/z [3]),
    .ZN(\u_multiplier/kx [3]));
 AND2_X1 \u_multiplier/LODx/Inst_MUX214_0/_12_  (.A1(\u_multiplier/LODx/_061_ ),
    .A2(\u_multiplier/LODx/z [2]),
    .ZN(\u_multiplier/kx [2]));
 AND2_X1 \u_multiplier/LODx/Inst_MUX214_1/_09_  (.A1(\u_multiplier/LODx/z [5]),
    .A2(\u_multiplier/LODx/_062_ ),
    .ZN(\u_multiplier/kx [5]));
 AND2_X1 \u_multiplier/LODx/Inst_MUX214_1/_10_  (.A1(\u_multiplier/LODx/_062_ ),
    .A2(\u_multiplier/LODx/z [4]),
    .ZN(\u_multiplier/kx [4]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_1/_11_  (.A1(\u_multiplier/LODx/_062_ ),
    .A2(\u_multiplier/LODx/z [7]),
    .ZN(\u_multiplier/kx [7]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_1/_12_  (.A1(\u_multiplier/LODx/_062_ ),
    .A2(\u_multiplier/LODx/z [6]),
    .ZN(\u_multiplier/kx [6]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_2/_09_  (.A1(\u_multiplier/LODx/z [9]),
    .A2(\u_multiplier/LODx/_063_ ),
    .ZN(\u_multiplier/kx [9]));
 AND2_X1 \u_multiplier/LODx/Inst_MUX214_2/_10_  (.A1(\u_multiplier/LODx/_063_ ),
    .A2(\u_multiplier/LODx/z [8]),
    .ZN(\u_multiplier/kx [8]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_2/_11_  (.A1(\u_multiplier/LODx/_063_ ),
    .A2(\u_multiplier/LODx/z [11]),
    .ZN(\u_multiplier/kx [11]));
 AND2_X1 \u_multiplier/LODx/Inst_MUX214_2/_12_  (.A1(\u_multiplier/LODx/_063_ ),
    .A2(\u_multiplier/LODx/z [10]),
    .ZN(\u_multiplier/kx [10]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_3/_09_  (.A1(\u_multiplier/LODx/z [13]),
    .A2(\u_multiplier/LODx/_064_ ),
    .ZN(\u_multiplier/kx [13]));
 AND2_X1 \u_multiplier/LODx/Inst_MUX214_3/_10_  (.A1(\u_multiplier/LODx/_064_ ),
    .A2(\u_multiplier/LODx/z [12]),
    .ZN(\u_multiplier/kx [12]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_3/_11_  (.A1(\u_multiplier/LODx/_064_ ),
    .A2(\u_multiplier/LODx/z [15]),
    .ZN(\u_multiplier/kx [15]));
 AND2_X1 \u_multiplier/LODx/Inst_MUX214_3/_12_  (.A1(\u_multiplier/LODx/_064_ ),
    .A2(\u_multiplier/LODx/z [14]),
    .ZN(\u_multiplier/kx [14]));
 AND2_X1 \u_multiplier/LODx/Inst_MUX214_4/_09_  (.A1(\u_multiplier/LODx/z [17]),
    .A2(\u_multiplier/LODx/_065_ ),
    .ZN(\u_multiplier/kx [17]));
 AND2_X1 \u_multiplier/LODx/Inst_MUX214_4/_10_  (.A1(\u_multiplier/LODx/_065_ ),
    .A2(\u_multiplier/LODx/z [16]),
    .ZN(\u_multiplier/kx [16]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_4/_11_  (.A1(\u_multiplier/LODx/_065_ ),
    .A2(\u_multiplier/LODx/z [19]),
    .ZN(\u_multiplier/kx [19]));
 AND2_X1 \u_multiplier/LODx/Inst_MUX214_4/_12_  (.A1(\u_multiplier/LODx/_065_ ),
    .A2(\u_multiplier/LODx/z [18]),
    .ZN(\u_multiplier/kx [18]));
 AND2_X1 \u_multiplier/LODx/Inst_MUX214_5/_09_  (.A1(\u_multiplier/LODx/z [21]),
    .A2(\u_multiplier/LODx/_066_ ),
    .ZN(\u_multiplier/kx [21]));
 AND2_X1 \u_multiplier/LODx/Inst_MUX214_5/_10_  (.A1(\u_multiplier/LODx/_066_ ),
    .A2(\u_multiplier/LODx/z [20]),
    .ZN(\u_multiplier/kx [20]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_5/_11_  (.A1(\u_multiplier/LODx/_066_ ),
    .A2(\u_multiplier/LODx/z [23]),
    .ZN(\u_multiplier/kx [23]));
 AND2_X1 \u_multiplier/LODx/Inst_MUX214_5/_12_  (.A1(\u_multiplier/LODx/_066_ ),
    .A2(\u_multiplier/LODx/z [22]),
    .ZN(\u_multiplier/kx [22]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_6/_09_  (.A1(\u_multiplier/LODx/z [25]),
    .A2(\u_multiplier/LODx/_067_ ),
    .ZN(\u_multiplier/kx [25]));
 AND2_X1 \u_multiplier/LODx/Inst_MUX214_6/_10_  (.A1(\u_multiplier/LODx/_067_ ),
    .A2(\u_multiplier/LODx/z [24]),
    .ZN(\u_multiplier/kx [24]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_6/_11_  (.A1(\u_multiplier/LODx/_067_ ),
    .A2(\u_multiplier/LODx/z [27]),
    .ZN(\u_multiplier/kx [27]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_6/_12_  (.A1(\u_multiplier/LODx/_067_ ),
    .A2(\u_multiplier/LODx/z [26]),
    .ZN(\u_multiplier/kx [26]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_7/_09_  (.A1(\u_multiplier/LODx/z [29]),
    .A2(\u_multiplier/LODx/_068_ ),
    .ZN(\u_multiplier/kx [29]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_7/_10_  (.A1(\u_multiplier/LODx/_068_ ),
    .A2(\u_multiplier/LODx/z [28]),
    .ZN(\u_multiplier/kx [28]));
 AND2_X1 \u_multiplier/LODx/Inst_MUX214_7/_11_  (.A1(\u_multiplier/LODx/_068_ ),
    .A2(\u_multiplier/LODx/z [31]),
    .ZN(\u_multiplier/kx [31]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_7/_12_  (.A1(\u_multiplier/LODx/_068_ ),
    .A2(\u_multiplier/LODx/z [30]),
    .ZN(\u_multiplier/kx [30]));
 NOR4_X2 \u_multiplier/LODx/_086_  (.A1(_0683_[30]),
    .A2(\u_multiplier/LODx/z [31]),
    .A3(_0683_[28]),
    .A4(_0683_[29]),
    .ZN(\u_multiplier/LODx/_054_ ));
 INV_X1 \u_multiplier/LODx/_087_  (.A(\u_multiplier/LODx/_054_ ),
    .ZN(\u_multiplier/LODx/select_high [3]));
 NOR4_X4 \u_multiplier/LODx/_088_  (.A1(_0683_[26]),
    .A2(\u_multiplier/LODx/z [27]),
    .A3(data_in_reg[24]),
    .A4(_0683_[25]),
    .ZN(\u_multiplier/LODx/_055_ ));
 INV_X1 \u_multiplier/LODx/_089_  (.A(\u_multiplier/LODx/_055_ ),
    .ZN(\u_multiplier/LODx/_083_ ));
 OR4_X2 \u_multiplier/LODx/_090_  (.A1(data_in_reg[14]),
    .A2(\u_multiplier/LODx/z [15]),
    .A3(data_in_reg[12]),
    .A4(data_in_reg[13]),
    .ZN(\u_multiplier/LODx/select_low [3]));
 OR4_X2 \u_multiplier/LODx/_091_  (.A1(data_in_reg[10]),
    .A2(\u_multiplier/LODx/z [11]),
    .A3(data_in_reg[8]),
    .A4(data_in_reg[9]),
    .ZN(\u_multiplier/LODx/_079_ ));
 OR4_X1 \u_multiplier/LODx/_092_  (.A1(data_in_reg[6]),
    .A2(\u_multiplier/LODx/z [7]),
    .A3(data_in_reg[4]),
    .A4(data_in_reg[5]),
    .ZN(\u_multiplier/LODx/_078_ ));
 OR4_X1 \u_multiplier/LODx/_093_  (.A1(data_in_reg[2]),
    .A2(\u_multiplier/LODx/z [3]),
    .A3(data_in_reg[0]),
    .A4(data_in_reg[1]),
    .ZN(\u_multiplier/LODx/_077_ ));
 NOR4_X4 \u_multiplier/LODx/_094_  (.A1(data_in_reg[22]),
    .A2(\u_multiplier/LODx/z [23]),
    .A3(data_in_reg[20]),
    .A4(data_in_reg[21]),
    .ZN(\u_multiplier/LODx/_056_ ));
 INV_X1 \u_multiplier/LODx/_095_  (.A(\u_multiplier/LODx/_056_ ),
    .ZN(\u_multiplier/LODx/_082_ ));
 NOR4_X4 \u_multiplier/LODx/_096_  (.A1(data_in_reg[18]),
    .A2(\u_multiplier/LODx/z [19]),
    .A3(data_in_reg[16]),
    .A4(data_in_reg[17]),
    .ZN(\u_multiplier/LODx/_057_ ));
 INV_X1 \u_multiplier/LODx/_097_  (.A(\u_multiplier/LODx/_057_ ),
    .ZN(\u_multiplier/LODx/_081_ ));
 AND4_X1 \u_multiplier/LODx/_098_  (.A1(\u_multiplier/LODx/_054_ ),
    .A2(\u_multiplier/LODx/_055_ ),
    .A3(\u_multiplier/LODx/_056_ ),
    .A4(\u_multiplier/LODx/_057_ ),
    .ZN(\u_multiplier/LODx/_058_ ));
 NAND4_X2 \u_multiplier/LODx/_099_  (.A1(\u_multiplier/LODx/_054_ ),
    .A2(\u_multiplier/LODx/_055_ ),
    .A3(\u_multiplier/LODx/_056_ ),
    .A4(\u_multiplier/LODx/_057_ ),
    .ZN(\u_multiplier/LODx/_059_ ));
 AND2_X1 \u_multiplier/LODx/_100_  (.A1(\u_multiplier/LODx/select_high [0]),
    .A2(\u_multiplier/LODx/_059_ ),
    .ZN(\u_multiplier/LODx/_065_ ));
 AND2_X1 \u_multiplier/LODx/_101_  (.A1(\u_multiplier/LODx/select_high [1]),
    .A2(\u_multiplier/LODx/_059_ ),
    .ZN(\u_multiplier/LODx/_066_ ));
 AND2_X1 \u_multiplier/LODx/_102_  (.A1(\u_multiplier/LODx/select_high [2]),
    .A2(\u_multiplier/LODx/_059_ ),
    .ZN(\u_multiplier/LODx/_067_ ));
 AND2_X1 \u_multiplier/LODx/_103_  (.A1(\u_multiplier/LODx/select_high [3]),
    .A2(\u_multiplier/LODx/_059_ ),
    .ZN(\u_multiplier/LODx/_068_ ));
 AND2_X1 \u_multiplier/LODx/_104_  (.A1(\u_multiplier/LODx/select_low [0]),
    .A2(\u_multiplier/LODx/_058_ ),
    .ZN(\u_multiplier/LODx/_061_ ));
 AND2_X1 \u_multiplier/LODx/_105_  (.A1(\u_multiplier/LODx/select_low [1]),
    .A2(\u_multiplier/LODx/_058_ ),
    .ZN(\u_multiplier/LODx/_062_ ));
 AND2_X1 \u_multiplier/LODx/_106_  (.A1(\u_multiplier/LODx/select_low [2]),
    .A2(\u_multiplier/LODx/_058_ ),
    .ZN(\u_multiplier/LODx/_063_ ));
 AND2_X1 \u_multiplier/LODx/_107_  (.A1(\u_multiplier/LODx/select_low [3]),
    .A2(\u_multiplier/LODx/_058_ ),
    .ZN(\u_multiplier/LODx/_064_ ));
 NOR4_X1 \u_multiplier/LODx/_108_  (.A1(\u_multiplier/LODx/select_low [3]),
    .A2(\u_multiplier/LODx/_079_ ),
    .A3(\u_multiplier/LODx/_078_ ),
    .A4(\u_multiplier/LODx/_077_ ),
    .ZN(\u_multiplier/LODx/_060_ ));
 AND2_X1 \u_multiplier/LODx/_109_  (.A1(\u_multiplier/LODx/_058_ ),
    .A2(\u_multiplier/LODx/_060_ ),
    .ZN(\u_multiplier/zero_x ));
 INV_X1 \u_multiplier/LODx/lod4_0/_12_  (.A(data_in_reg[2]),
    .ZN(\u_multiplier/LODx/lod4_0/_10_ ));
 INV_X1 \u_multiplier/LODx/lod4_0/_13_  (.A(data_in_reg[1]),
    .ZN(\u_multiplier/LODx/lod4_0/_11_ ));
 INV_X1 \u_multiplier/LODx/lod4_0/_14_  (.A(data_in_reg[0]),
    .ZN(\u_multiplier/LODx/lod4_0/_09_ ));
 NOR2_X1 \u_multiplier/LODx/lod4_0/_15_  (.A1(\u_multiplier/LODx/lod4_0/_10_ ),
    .A2(\u_multiplier/LODx/z [3]),
    .ZN(\u_multiplier/LODx/z [2]));
 NOR3_X1 \u_multiplier/LODx/lod4_0/_16_  (.A1(data_in_reg[2]),
    .A2(\u_multiplier/LODx/z [3]),
    .A3(\u_multiplier/LODx/lod4_0/_11_ ),
    .ZN(\u_multiplier/LODx/z [1]));
 NOR4_X1 \u_multiplier/LODx/lod4_0/_17_  (.A1(data_in_reg[2]),
    .A2(\u_multiplier/LODx/z [3]),
    .A3(data_in_reg[1]),
    .A4(\u_multiplier/LODx/lod4_0/_09_ ),
    .ZN(\u_multiplier/LODx/z [0]));
 INV_X1 \u_multiplier/LODx/lod4_1/_12_  (.A(data_in_reg[6]),
    .ZN(\u_multiplier/LODx/lod4_1/_10_ ));
 INV_X1 \u_multiplier/LODx/lod4_1/_13_  (.A(data_in_reg[5]),
    .ZN(\u_multiplier/LODx/lod4_1/_11_ ));
 INV_X1 \u_multiplier/LODx/lod4_1/_14_  (.A(data_in_reg[4]),
    .ZN(\u_multiplier/LODx/lod4_1/_09_ ));
 NOR2_X1 \u_multiplier/LODx/lod4_1/_15_  (.A1(\u_multiplier/LODx/lod4_1/_10_ ),
    .A2(\u_multiplier/LODx/z [7]),
    .ZN(\u_multiplier/LODx/z [6]));
 NOR3_X1 \u_multiplier/LODx/lod4_1/_16_  (.A1(data_in_reg[6]),
    .A2(\u_multiplier/LODx/z [7]),
    .A3(\u_multiplier/LODx/lod4_1/_11_ ),
    .ZN(\u_multiplier/LODx/z [5]));
 NOR4_X1 \u_multiplier/LODx/lod4_1/_17_  (.A1(data_in_reg[6]),
    .A2(\u_multiplier/LODx/z [7]),
    .A3(data_in_reg[5]),
    .A4(\u_multiplier/LODx/lod4_1/_09_ ),
    .ZN(\u_multiplier/LODx/z [4]));
 INV_X1 \u_multiplier/LODx/lod4_2/_12_  (.A(data_in_reg[10]),
    .ZN(\u_multiplier/LODx/lod4_2/_10_ ));
 INV_X1 \u_multiplier/LODx/lod4_2/_13_  (.A(data_in_reg[9]),
    .ZN(\u_multiplier/LODx/lod4_2/_11_ ));
 INV_X1 \u_multiplier/LODx/lod4_2/_14_  (.A(data_in_reg[8]),
    .ZN(\u_multiplier/LODx/lod4_2/_09_ ));
 NOR2_X1 \u_multiplier/LODx/lod4_2/_15_  (.A1(\u_multiplier/LODx/lod4_2/_10_ ),
    .A2(\u_multiplier/LODx/z [11]),
    .ZN(\u_multiplier/LODx/z [10]));
 NOR3_X1 \u_multiplier/LODx/lod4_2/_16_  (.A1(data_in_reg[10]),
    .A2(\u_multiplier/LODx/z [11]),
    .A3(\u_multiplier/LODx/lod4_2/_11_ ),
    .ZN(\u_multiplier/LODx/z [9]));
 NOR4_X1 \u_multiplier/LODx/lod4_2/_17_  (.A1(data_in_reg[10]),
    .A2(\u_multiplier/LODx/z [11]),
    .A3(data_in_reg[9]),
    .A4(\u_multiplier/LODx/lod4_2/_09_ ),
    .ZN(\u_multiplier/LODx/z [8]));
 INV_X1 \u_multiplier/LODx/lod4_3/_12_  (.A(data_in_reg[14]),
    .ZN(\u_multiplier/LODx/lod4_3/_10_ ));
 INV_X1 \u_multiplier/LODx/lod4_3/_13_  (.A(data_in_reg[13]),
    .ZN(\u_multiplier/LODx/lod4_3/_11_ ));
 INV_X1 \u_multiplier/LODx/lod4_3/_14_  (.A(data_in_reg[12]),
    .ZN(\u_multiplier/LODx/lod4_3/_09_ ));
 NOR2_X1 \u_multiplier/LODx/lod4_3/_15_  (.A1(\u_multiplier/LODx/lod4_3/_10_ ),
    .A2(\u_multiplier/LODx/z [15]),
    .ZN(\u_multiplier/LODx/z [14]));
 NOR3_X1 \u_multiplier/LODx/lod4_3/_16_  (.A1(data_in_reg[14]),
    .A2(\u_multiplier/LODx/z [15]),
    .A3(\u_multiplier/LODx/lod4_3/_11_ ),
    .ZN(\u_multiplier/LODx/z [13]));
 NOR4_X1 \u_multiplier/LODx/lod4_3/_17_  (.A1(data_in_reg[14]),
    .A2(\u_multiplier/LODx/z [15]),
    .A3(data_in_reg[13]),
    .A4(\u_multiplier/LODx/lod4_3/_09_ ),
    .ZN(\u_multiplier/LODx/z [12]));
 INV_X1 \u_multiplier/LODx/lod4_4/_12_  (.A(data_in_reg[18]),
    .ZN(\u_multiplier/LODx/lod4_4/_10_ ));
 INV_X1 \u_multiplier/LODx/lod4_4/_13_  (.A(data_in_reg[17]),
    .ZN(\u_multiplier/LODx/lod4_4/_11_ ));
 INV_X1 \u_multiplier/LODx/lod4_4/_14_  (.A(data_in_reg[16]),
    .ZN(\u_multiplier/LODx/lod4_4/_09_ ));
 NOR2_X1 \u_multiplier/LODx/lod4_4/_15_  (.A1(\u_multiplier/LODx/lod4_4/_10_ ),
    .A2(\u_multiplier/LODx/z [19]),
    .ZN(\u_multiplier/LODx/z [18]));
 NOR3_X1 \u_multiplier/LODx/lod4_4/_16_  (.A1(data_in_reg[18]),
    .A2(\u_multiplier/LODx/z [19]),
    .A3(\u_multiplier/LODx/lod4_4/_11_ ),
    .ZN(\u_multiplier/LODx/z [17]));
 NOR4_X1 \u_multiplier/LODx/lod4_4/_17_  (.A1(data_in_reg[18]),
    .A2(\u_multiplier/LODx/z [19]),
    .A3(data_in_reg[17]),
    .A4(\u_multiplier/LODx/lod4_4/_09_ ),
    .ZN(\u_multiplier/LODx/z [16]));
 INV_X1 \u_multiplier/LODx/lod4_5/_12_  (.A(data_in_reg[22]),
    .ZN(\u_multiplier/LODx/lod4_5/_10_ ));
 INV_X1 \u_multiplier/LODx/lod4_5/_13_  (.A(data_in_reg[21]),
    .ZN(\u_multiplier/LODx/lod4_5/_11_ ));
 INV_X1 \u_multiplier/LODx/lod4_5/_14_  (.A(data_in_reg[20]),
    .ZN(\u_multiplier/LODx/lod4_5/_09_ ));
 NOR2_X1 \u_multiplier/LODx/lod4_5/_15_  (.A1(\u_multiplier/LODx/lod4_5/_10_ ),
    .A2(\u_multiplier/LODx/z [23]),
    .ZN(\u_multiplier/LODx/z [22]));
 NOR3_X1 \u_multiplier/LODx/lod4_5/_16_  (.A1(data_in_reg[22]),
    .A2(\u_multiplier/LODx/z [23]),
    .A3(\u_multiplier/LODx/lod4_5/_11_ ),
    .ZN(\u_multiplier/LODx/z [21]));
 NOR4_X1 \u_multiplier/LODx/lod4_5/_17_  (.A1(data_in_reg[22]),
    .A2(\u_multiplier/LODx/z [23]),
    .A3(data_in_reg[21]),
    .A4(\u_multiplier/LODx/lod4_5/_09_ ),
    .ZN(\u_multiplier/LODx/z [20]));
 INV_X1 \u_multiplier/LODx/lod4_6/_12_  (.A(_0683_[26]),
    .ZN(\u_multiplier/LODx/lod4_6/_10_ ));
 INV_X1 \u_multiplier/LODx/lod4_6/_13_  (.A(_0683_[25]),
    .ZN(\u_multiplier/LODx/lod4_6/_11_ ));
 INV_X1 \u_multiplier/LODx/lod4_6/_14_  (.A(data_in_reg[24]),
    .ZN(\u_multiplier/LODx/lod4_6/_09_ ));
 NOR2_X1 \u_multiplier/LODx/lod4_6/_15_  (.A1(\u_multiplier/LODx/lod4_6/_10_ ),
    .A2(\u_multiplier/LODx/z [27]),
    .ZN(\u_multiplier/LODx/z [26]));
 NOR3_X1 \u_multiplier/LODx/lod4_6/_16_  (.A1(_0683_[26]),
    .A2(\u_multiplier/LODx/z [27]),
    .A3(\u_multiplier/LODx/lod4_6/_11_ ),
    .ZN(\u_multiplier/LODx/z [25]));
 NOR4_X1 \u_multiplier/LODx/lod4_6/_17_  (.A1(_0683_[26]),
    .A2(\u_multiplier/LODx/z [27]),
    .A3(_0683_[25]),
    .A4(\u_multiplier/LODx/lod4_6/_09_ ),
    .ZN(\u_multiplier/LODx/z [24]));
 INV_X1 \u_multiplier/LODx/lod4_7/_12_  (.A(_0683_[30]),
    .ZN(\u_multiplier/LODx/lod4_7/_10_ ));
 INV_X1 \u_multiplier/LODx/lod4_7/_13_  (.A(_0683_[29]),
    .ZN(\u_multiplier/LODx/lod4_7/_11_ ));
 INV_X1 \u_multiplier/LODx/lod4_7/_14_  (.A(_0683_[28]),
    .ZN(\u_multiplier/LODx/lod4_7/_09_ ));
 NOR2_X1 \u_multiplier/LODx/lod4_7/_15_  (.A1(\u_multiplier/LODx/lod4_7/_10_ ),
    .A2(\u_multiplier/LODx/z [31]),
    .ZN(\u_multiplier/LODx/z [30]));
 NOR3_X1 \u_multiplier/LODx/lod4_7/_16_  (.A1(_0683_[30]),
    .A2(\u_multiplier/LODx/z [31]),
    .A3(\u_multiplier/LODx/lod4_7/_11_ ),
    .ZN(\u_multiplier/LODx/z [29]));
 NOR4_X1 \u_multiplier/LODx/lod4_7/_17_  (.A1(_0683_[30]),
    .A2(\u_multiplier/LODx/z [31]),
    .A3(_0683_[29]),
    .A4(\u_multiplier/LODx/lod4_7/_09_ ),
    .ZN(\u_multiplier/LODx/z [28]));
 INV_X1 \u_multiplier/LODx/lod4_middle_high/_12_  (.A(\u_multiplier/LODx/_083_ ),
    .ZN(\u_multiplier/LODx/lod4_middle_high/_10_ ));
 INV_X1 \u_multiplier/LODx/lod4_middle_high/_13_  (.A(\u_multiplier/LODx/_082_ ),
    .ZN(\u_multiplier/LODx/lod4_middle_high/_11_ ));
 INV_X1 \u_multiplier/LODx/lod4_middle_high/_14_  (.A(\u_multiplier/LODx/_081_ ),
    .ZN(\u_multiplier/LODx/lod4_middle_high/_09_ ));
 NOR2_X1 \u_multiplier/LODx/lod4_middle_high/_15_  (.A1(\u_multiplier/LODx/lod4_middle_high/_10_ ),
    .A2(\u_multiplier/LODx/select_high [3]),
    .ZN(\u_multiplier/LODx/select_high [2]));
 NOR3_X1 \u_multiplier/LODx/lod4_middle_high/_16_  (.A1(\u_multiplier/LODx/_083_ ),
    .A2(\u_multiplier/LODx/select_high [3]),
    .A3(\u_multiplier/LODx/lod4_middle_high/_11_ ),
    .ZN(\u_multiplier/LODx/select_high [1]));
 NOR4_X1 \u_multiplier/LODx/lod4_middle_high/_17_  (.A1(\u_multiplier/LODx/_083_ ),
    .A2(\u_multiplier/LODx/select_high [3]),
    .A3(\u_multiplier/LODx/_082_ ),
    .A4(\u_multiplier/LODx/lod4_middle_high/_09_ ),
    .ZN(\u_multiplier/LODx/select_high [0]));
 INV_X1 \u_multiplier/LODx/lod4_middle_low/_12_  (.A(\u_multiplier/LODx/_079_ ),
    .ZN(\u_multiplier/LODx/lod4_middle_low/_10_ ));
 INV_X1 \u_multiplier/LODx/lod4_middle_low/_13_  (.A(\u_multiplier/LODx/_078_ ),
    .ZN(\u_multiplier/LODx/lod4_middle_low/_11_ ));
 INV_X1 \u_multiplier/LODx/lod4_middle_low/_14_  (.A(\u_multiplier/LODx/_077_ ),
    .ZN(\u_multiplier/LODx/lod4_middle_low/_09_ ));
 NOR2_X1 \u_multiplier/LODx/lod4_middle_low/_15_  (.A1(\u_multiplier/LODx/lod4_middle_low/_10_ ),
    .A2(\u_multiplier/LODx/select_low [3]),
    .ZN(\u_multiplier/LODx/select_low [2]));
 NOR3_X1 \u_multiplier/LODx/lod4_middle_low/_16_  (.A1(\u_multiplier/LODx/_079_ ),
    .A2(\u_multiplier/LODx/select_low [3]),
    .A3(\u_multiplier/LODx/lod4_middle_low/_11_ ),
    .ZN(\u_multiplier/LODx/select_low [1]));
 NOR4_X1 \u_multiplier/LODx/lod4_middle_low/_17_  (.A1(\u_multiplier/LODx/_079_ ),
    .A2(\u_multiplier/LODx/select_low [3]),
    .A3(\u_multiplier/LODx/_078_ ),
    .A4(\u_multiplier/LODx/lod4_middle_low/_09_ ),
    .ZN(\u_multiplier/LODx/select_low [0]));
 AND2_X1 \u_multiplier/LODy/Inst_MUX214_0/_09_  (.A1(\u_multiplier/LODy/z [1]),
    .A2(\u_multiplier/LODy/_061_ ),
    .ZN(\u_multiplier/ky [1]));
 AND2_X1 \u_multiplier/LODy/Inst_MUX214_0/_10_  (.A1(\u_multiplier/LODy/_061_ ),
    .A2(\u_multiplier/LODy/z [0]),
    .ZN(\u_multiplier/ky [0]));
 AND2_X1 \u_multiplier/LODy/Inst_MUX214_0/_11_  (.A1(\u_multiplier/LODy/_061_ ),
    .A2(\u_multiplier/LODy/z [3]),
    .ZN(\u_multiplier/ky [3]));
 AND2_X1 \u_multiplier/LODy/Inst_MUX214_0/_12_  (.A1(\u_multiplier/LODy/_061_ ),
    .A2(\u_multiplier/LODy/z [2]),
    .ZN(\u_multiplier/ky [2]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_1/_09_  (.A1(\u_multiplier/LODy/z [5]),
    .A2(\u_multiplier/LODy/_062_ ),
    .ZN(\u_multiplier/ky [5]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_1/_10_  (.A1(\u_multiplier/LODy/_062_ ),
    .A2(\u_multiplier/LODy/z [4]),
    .ZN(\u_multiplier/ky [4]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_1/_11_  (.A1(\u_multiplier/LODy/_062_ ),
    .A2(\u_multiplier/LODy/z [7]),
    .ZN(\u_multiplier/ky [7]));
 AND2_X1 \u_multiplier/LODy/Inst_MUX214_1/_12_  (.A1(\u_multiplier/LODy/_062_ ),
    .A2(\u_multiplier/LODy/z [6]),
    .ZN(\u_multiplier/ky [6]));
 AND2_X1 \u_multiplier/LODy/Inst_MUX214_2/_09_  (.A1(\u_multiplier/LODy/z [9]),
    .A2(\u_multiplier/LODy/_063_ ),
    .ZN(\u_multiplier/ky [9]));
 AND2_X1 \u_multiplier/LODy/Inst_MUX214_2/_10_  (.A1(\u_multiplier/LODy/_063_ ),
    .A2(\u_multiplier/LODy/z [8]),
    .ZN(\u_multiplier/ky [8]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_2/_11_  (.A1(\u_multiplier/LODy/_063_ ),
    .A2(\u_multiplier/LODy/z [11]),
    .ZN(\u_multiplier/ky [11]));
 AND2_X1 \u_multiplier/LODy/Inst_MUX214_2/_12_  (.A1(\u_multiplier/LODy/_063_ ),
    .A2(\u_multiplier/LODy/z [10]),
    .ZN(\u_multiplier/ky [10]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_3/_09_  (.A1(\u_multiplier/LODy/z [13]),
    .A2(\u_multiplier/LODy/_064_ ),
    .ZN(\u_multiplier/ky [13]));
 AND2_X1 \u_multiplier/LODy/Inst_MUX214_3/_10_  (.A1(\u_multiplier/LODy/_064_ ),
    .A2(\u_multiplier/LODy/z [12]),
    .ZN(\u_multiplier/ky [12]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_3/_11_  (.A1(\u_multiplier/LODy/_064_ ),
    .A2(\u_multiplier/LODy/z [15]),
    .ZN(\u_multiplier/ky [15]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_3/_12_  (.A1(\u_multiplier/LODy/_064_ ),
    .A2(\u_multiplier/LODy/z [14]),
    .ZN(\u_multiplier/ky [14]));
 AND2_X1 \u_multiplier/LODy/Inst_MUX214_4/_09_  (.A1(\u_multiplier/LODy/z [17]),
    .A2(\u_multiplier/LODy/_065_ ),
    .ZN(\u_multiplier/ky [17]));
 AND2_X1 \u_multiplier/LODy/Inst_MUX214_4/_10_  (.A1(\u_multiplier/LODy/_065_ ),
    .A2(\u_multiplier/LODy/z [16]),
    .ZN(\u_multiplier/ky [16]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_4/_11_  (.A1(\u_multiplier/LODy/_065_ ),
    .A2(\u_multiplier/LODy/z [19]),
    .ZN(\u_multiplier/ky [19]));
 AND2_X1 \u_multiplier/LODy/Inst_MUX214_4/_12_  (.A1(\u_multiplier/LODy/_065_ ),
    .A2(\u_multiplier/LODy/z [18]),
    .ZN(\u_multiplier/ky [18]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_5/_09_  (.A1(\u_multiplier/LODy/z [21]),
    .A2(\u_multiplier/LODy/_066_ ),
    .ZN(\u_multiplier/ky [21]));
 AND2_X1 \u_multiplier/LODy/Inst_MUX214_5/_10_  (.A1(\u_multiplier/LODy/_066_ ),
    .A2(\u_multiplier/LODy/z [20]),
    .ZN(\u_multiplier/ky [20]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_5/_11_  (.A1(\u_multiplier/LODy/_066_ ),
    .A2(\u_multiplier/LODy/z [23]),
    .ZN(\u_multiplier/ky [23]));
 AND2_X1 \u_multiplier/LODy/Inst_MUX214_5/_12_  (.A1(\u_multiplier/LODy/_066_ ),
    .A2(\u_multiplier/LODy/z [22]),
    .ZN(\u_multiplier/ky [22]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_6/_09_  (.A1(\u_multiplier/LODy/z [25]),
    .A2(\u_multiplier/LODy/_067_ ),
    .ZN(\u_multiplier/ky [25]));
 AND2_X1 \u_multiplier/LODy/Inst_MUX214_6/_10_  (.A1(\u_multiplier/LODy/_067_ ),
    .A2(\u_multiplier/LODy/z [24]),
    .ZN(\u_multiplier/ky [24]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_6/_11_  (.A1(\u_multiplier/LODy/_067_ ),
    .A2(\u_multiplier/LODy/z [27]),
    .ZN(\u_multiplier/ky [27]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_6/_12_  (.A1(\u_multiplier/LODy/_067_ ),
    .A2(\u_multiplier/LODy/z [26]),
    .ZN(\u_multiplier/ky [26]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_7/_09_  (.A1(\u_multiplier/LODy/z [29]),
    .A2(\u_multiplier/LODy/_068_ ),
    .ZN(\u_multiplier/ky [29]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_7/_10_  (.A1(\u_multiplier/LODy/_068_ ),
    .A2(\u_multiplier/LODy/z [28]),
    .ZN(\u_multiplier/ky [28]));
 AND2_X1 \u_multiplier/LODy/Inst_MUX214_7/_11_  (.A1(\u_multiplier/LODy/_068_ ),
    .A2(\u_multiplier/LODy/z [31]),
    .ZN(\u_multiplier/ky [31]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_7/_12_  (.A1(\u_multiplier/LODy/_068_ ),
    .A2(\u_multiplier/LODy/z [30]),
    .ZN(\u_multiplier/ky [30]));
 NOR4_X4 \u_multiplier/LODy/_086_  (.A1(sram_rdata_reg[30]),
    .A2(\u_multiplier/LODy/z [31]),
    .A3(sram_rdata_reg[28]),
    .A4(sram_rdata_reg[29]),
    .ZN(\u_multiplier/LODy/_054_ ));
 INV_X1 \u_multiplier/LODy/_087_  (.A(\u_multiplier/LODy/_054_ ),
    .ZN(\u_multiplier/LODy/select_high [3]));
 NOR4_X2 \u_multiplier/LODy/_088_  (.A1(sram_rdata_reg[26]),
    .A2(\u_multiplier/LODy/z [27]),
    .A3(sram_rdata_reg[24]),
    .A4(sram_rdata_reg[25]),
    .ZN(\u_multiplier/LODy/_055_ ));
 INV_X1 \u_multiplier/LODy/_089_  (.A(\u_multiplier/LODy/_055_ ),
    .ZN(\u_multiplier/LODy/_083_ ));
 OR4_X2 \u_multiplier/LODy/_090_  (.A1(sram_rdata_reg[14]),
    .A2(\u_multiplier/LODy/z [15]),
    .A3(sram_rdata_reg[12]),
    .A4(sram_rdata_reg[13]),
    .ZN(\u_multiplier/LODy/select_low [3]));
 OR4_X2 \u_multiplier/LODy/_091_  (.A1(sram_rdata_reg[10]),
    .A2(\u_multiplier/LODy/z [11]),
    .A3(sram_rdata_reg[8]),
    .A4(sram_rdata_reg[9]),
    .ZN(\u_multiplier/LODy/_079_ ));
 OR4_X1 \u_multiplier/LODy/_092_  (.A1(sram_rdata_reg[6]),
    .A2(\u_multiplier/LODy/z [7]),
    .A3(sram_rdata_reg[4]),
    .A4(sram_rdata_reg[5]),
    .ZN(\u_multiplier/LODy/_078_ ));
 OR4_X1 \u_multiplier/LODy/_093_  (.A1(sram_rdata_reg[2]),
    .A2(\u_multiplier/LODy/z [3]),
    .A3(sram_rdata_reg[0]),
    .A4(sram_rdata_reg[1]),
    .ZN(\u_multiplier/LODy/_077_ ));
 NOR4_X4 \u_multiplier/LODy/_094_  (.A1(sram_rdata_reg[22]),
    .A2(\u_multiplier/LODy/z [23]),
    .A3(sram_rdata_reg[20]),
    .A4(sram_rdata_reg[21]),
    .ZN(\u_multiplier/LODy/_056_ ));
 INV_X1 \u_multiplier/LODy/_095_  (.A(\u_multiplier/LODy/_056_ ),
    .ZN(\u_multiplier/LODy/_082_ ));
 NOR4_X4 \u_multiplier/LODy/_096_  (.A1(sram_rdata_reg[18]),
    .A2(\u_multiplier/LODy/z [19]),
    .A3(sram_rdata_reg[16]),
    .A4(sram_rdata_reg[17]),
    .ZN(\u_multiplier/LODy/_057_ ));
 INV_X1 \u_multiplier/LODy/_097_  (.A(\u_multiplier/LODy/_057_ ),
    .ZN(\u_multiplier/LODy/_081_ ));
 AND4_X1 \u_multiplier/LODy/_098_  (.A1(\u_multiplier/LODy/_054_ ),
    .A2(\u_multiplier/LODy/_055_ ),
    .A3(\u_multiplier/LODy/_056_ ),
    .A4(\u_multiplier/LODy/_057_ ),
    .ZN(\u_multiplier/LODy/_058_ ));
 NAND4_X2 \u_multiplier/LODy/_099_  (.A1(\u_multiplier/LODy/_054_ ),
    .A2(\u_multiplier/LODy/_055_ ),
    .A3(\u_multiplier/LODy/_056_ ),
    .A4(\u_multiplier/LODy/_057_ ),
    .ZN(\u_multiplier/LODy/_059_ ));
 AND2_X1 \u_multiplier/LODy/_100_  (.A1(\u_multiplier/LODy/select_high [0]),
    .A2(\u_multiplier/LODy/_059_ ),
    .ZN(\u_multiplier/LODy/_065_ ));
 AND2_X1 \u_multiplier/LODy/_101_  (.A1(\u_multiplier/LODy/select_high [1]),
    .A2(\u_multiplier/LODy/_059_ ),
    .ZN(\u_multiplier/LODy/_066_ ));
 AND2_X1 \u_multiplier/LODy/_102_  (.A1(\u_multiplier/LODy/select_high [2]),
    .A2(\u_multiplier/LODy/_059_ ),
    .ZN(\u_multiplier/LODy/_067_ ));
 AND2_X1 \u_multiplier/LODy/_103_  (.A1(\u_multiplier/LODy/select_high [3]),
    .A2(\u_multiplier/LODy/_059_ ),
    .ZN(\u_multiplier/LODy/_068_ ));
 AND2_X1 \u_multiplier/LODy/_104_  (.A1(\u_multiplier/LODy/select_low [0]),
    .A2(\u_multiplier/LODy/_058_ ),
    .ZN(\u_multiplier/LODy/_061_ ));
 AND2_X1 \u_multiplier/LODy/_105_  (.A1(\u_multiplier/LODy/select_low [1]),
    .A2(\u_multiplier/LODy/_058_ ),
    .ZN(\u_multiplier/LODy/_062_ ));
 AND2_X1 \u_multiplier/LODy/_106_  (.A1(\u_multiplier/LODy/select_low [2]),
    .A2(\u_multiplier/LODy/_058_ ),
    .ZN(\u_multiplier/LODy/_063_ ));
 AND2_X1 \u_multiplier/LODy/_107_  (.A1(\u_multiplier/LODy/select_low [3]),
    .A2(\u_multiplier/LODy/_058_ ),
    .ZN(\u_multiplier/LODy/_064_ ));
 NOR4_X1 \u_multiplier/LODy/_108_  (.A1(\u_multiplier/LODy/select_low [3]),
    .A2(\u_multiplier/LODy/_079_ ),
    .A3(\u_multiplier/LODy/_078_ ),
    .A4(\u_multiplier/LODy/_077_ ),
    .ZN(\u_multiplier/LODy/_060_ ));
 AND2_X2 \u_multiplier/LODy/_109_  (.A1(\u_multiplier/LODy/_058_ ),
    .A2(\u_multiplier/LODy/_060_ ),
    .ZN(\u_multiplier/zero_y ));
 INV_X1 \u_multiplier/LODy/lod4_0/_12_  (.A(sram_rdata_reg[2]),
    .ZN(\u_multiplier/LODy/lod4_0/_10_ ));
 INV_X1 \u_multiplier/LODy/lod4_0/_13_  (.A(sram_rdata_reg[1]),
    .ZN(\u_multiplier/LODy/lod4_0/_11_ ));
 INV_X1 \u_multiplier/LODy/lod4_0/_14_  (.A(sram_rdata_reg[0]),
    .ZN(\u_multiplier/LODy/lod4_0/_09_ ));
 NOR2_X1 \u_multiplier/LODy/lod4_0/_15_  (.A1(\u_multiplier/LODy/lod4_0/_10_ ),
    .A2(\u_multiplier/LODy/z [3]),
    .ZN(\u_multiplier/LODy/z [2]));
 NOR3_X1 \u_multiplier/LODy/lod4_0/_16_  (.A1(sram_rdata_reg[2]),
    .A2(\u_multiplier/LODy/z [3]),
    .A3(\u_multiplier/LODy/lod4_0/_11_ ),
    .ZN(\u_multiplier/LODy/z [1]));
 NOR4_X1 \u_multiplier/LODy/lod4_0/_17_  (.A1(sram_rdata_reg[2]),
    .A2(\u_multiplier/LODy/z [3]),
    .A3(sram_rdata_reg[1]),
    .A4(\u_multiplier/LODy/lod4_0/_09_ ),
    .ZN(\u_multiplier/LODy/z [0]));
 INV_X1 \u_multiplier/LODy/lod4_1/_12_  (.A(sram_rdata_reg[6]),
    .ZN(\u_multiplier/LODy/lod4_1/_10_ ));
 INV_X1 \u_multiplier/LODy/lod4_1/_13_  (.A(sram_rdata_reg[5]),
    .ZN(\u_multiplier/LODy/lod4_1/_11_ ));
 INV_X1 \u_multiplier/LODy/lod4_1/_14_  (.A(sram_rdata_reg[4]),
    .ZN(\u_multiplier/LODy/lod4_1/_09_ ));
 NOR2_X1 \u_multiplier/LODy/lod4_1/_15_  (.A1(\u_multiplier/LODy/lod4_1/_10_ ),
    .A2(\u_multiplier/LODy/z [7]),
    .ZN(\u_multiplier/LODy/z [6]));
 NOR3_X1 \u_multiplier/LODy/lod4_1/_16_  (.A1(sram_rdata_reg[6]),
    .A2(\u_multiplier/LODy/z [7]),
    .A3(\u_multiplier/LODy/lod4_1/_11_ ),
    .ZN(\u_multiplier/LODy/z [5]));
 NOR4_X1 \u_multiplier/LODy/lod4_1/_17_  (.A1(sram_rdata_reg[6]),
    .A2(\u_multiplier/LODy/z [7]),
    .A3(sram_rdata_reg[5]),
    .A4(\u_multiplier/LODy/lod4_1/_09_ ),
    .ZN(\u_multiplier/LODy/z [4]));
 INV_X1 \u_multiplier/LODy/lod4_2/_12_  (.A(sram_rdata_reg[10]),
    .ZN(\u_multiplier/LODy/lod4_2/_10_ ));
 INV_X1 \u_multiplier/LODy/lod4_2/_13_  (.A(sram_rdata_reg[9]),
    .ZN(\u_multiplier/LODy/lod4_2/_11_ ));
 INV_X1 \u_multiplier/LODy/lod4_2/_14_  (.A(sram_rdata_reg[8]),
    .ZN(\u_multiplier/LODy/lod4_2/_09_ ));
 NOR2_X1 \u_multiplier/LODy/lod4_2/_15_  (.A1(\u_multiplier/LODy/lod4_2/_10_ ),
    .A2(\u_multiplier/LODy/z [11]),
    .ZN(\u_multiplier/LODy/z [10]));
 NOR3_X1 \u_multiplier/LODy/lod4_2/_16_  (.A1(sram_rdata_reg[10]),
    .A2(\u_multiplier/LODy/z [11]),
    .A3(\u_multiplier/LODy/lod4_2/_11_ ),
    .ZN(\u_multiplier/LODy/z [9]));
 NOR4_X1 \u_multiplier/LODy/lod4_2/_17_  (.A1(sram_rdata_reg[10]),
    .A2(\u_multiplier/LODy/z [11]),
    .A3(sram_rdata_reg[9]),
    .A4(\u_multiplier/LODy/lod4_2/_09_ ),
    .ZN(\u_multiplier/LODy/z [8]));
 INV_X1 \u_multiplier/LODy/lod4_3/_12_  (.A(sram_rdata_reg[14]),
    .ZN(\u_multiplier/LODy/lod4_3/_10_ ));
 INV_X1 \u_multiplier/LODy/lod4_3/_13_  (.A(sram_rdata_reg[13]),
    .ZN(\u_multiplier/LODy/lod4_3/_11_ ));
 INV_X1 \u_multiplier/LODy/lod4_3/_14_  (.A(sram_rdata_reg[12]),
    .ZN(\u_multiplier/LODy/lod4_3/_09_ ));
 NOR2_X1 \u_multiplier/LODy/lod4_3/_15_  (.A1(\u_multiplier/LODy/lod4_3/_10_ ),
    .A2(\u_multiplier/LODy/z [15]),
    .ZN(\u_multiplier/LODy/z [14]));
 NOR3_X1 \u_multiplier/LODy/lod4_3/_16_  (.A1(sram_rdata_reg[14]),
    .A2(\u_multiplier/LODy/z [15]),
    .A3(\u_multiplier/LODy/lod4_3/_11_ ),
    .ZN(\u_multiplier/LODy/z [13]));
 NOR4_X1 \u_multiplier/LODy/lod4_3/_17_  (.A1(sram_rdata_reg[14]),
    .A2(\u_multiplier/LODy/z [15]),
    .A3(sram_rdata_reg[13]),
    .A4(\u_multiplier/LODy/lod4_3/_09_ ),
    .ZN(\u_multiplier/LODy/z [12]));
 INV_X1 \u_multiplier/LODy/lod4_4/_12_  (.A(sram_rdata_reg[18]),
    .ZN(\u_multiplier/LODy/lod4_4/_10_ ));
 INV_X1 \u_multiplier/LODy/lod4_4/_13_  (.A(sram_rdata_reg[17]),
    .ZN(\u_multiplier/LODy/lod4_4/_11_ ));
 INV_X1 \u_multiplier/LODy/lod4_4/_14_  (.A(sram_rdata_reg[16]),
    .ZN(\u_multiplier/LODy/lod4_4/_09_ ));
 NOR2_X1 \u_multiplier/LODy/lod4_4/_15_  (.A1(\u_multiplier/LODy/lod4_4/_10_ ),
    .A2(\u_multiplier/LODy/z [19]),
    .ZN(\u_multiplier/LODy/z [18]));
 NOR3_X1 \u_multiplier/LODy/lod4_4/_16_  (.A1(sram_rdata_reg[18]),
    .A2(\u_multiplier/LODy/z [19]),
    .A3(\u_multiplier/LODy/lod4_4/_11_ ),
    .ZN(\u_multiplier/LODy/z [17]));
 NOR4_X1 \u_multiplier/LODy/lod4_4/_17_  (.A1(sram_rdata_reg[18]),
    .A2(\u_multiplier/LODy/z [19]),
    .A3(sram_rdata_reg[17]),
    .A4(\u_multiplier/LODy/lod4_4/_09_ ),
    .ZN(\u_multiplier/LODy/z [16]));
 INV_X1 \u_multiplier/LODy/lod4_5/_12_  (.A(sram_rdata_reg[22]),
    .ZN(\u_multiplier/LODy/lod4_5/_10_ ));
 INV_X1 \u_multiplier/LODy/lod4_5/_13_  (.A(sram_rdata_reg[21]),
    .ZN(\u_multiplier/LODy/lod4_5/_11_ ));
 INV_X1 \u_multiplier/LODy/lod4_5/_14_  (.A(sram_rdata_reg[20]),
    .ZN(\u_multiplier/LODy/lod4_5/_09_ ));
 NOR2_X1 \u_multiplier/LODy/lod4_5/_15_  (.A1(\u_multiplier/LODy/lod4_5/_10_ ),
    .A2(\u_multiplier/LODy/z [23]),
    .ZN(\u_multiplier/LODy/z [22]));
 NOR3_X1 \u_multiplier/LODy/lod4_5/_16_  (.A1(sram_rdata_reg[22]),
    .A2(\u_multiplier/LODy/z [23]),
    .A3(\u_multiplier/LODy/lod4_5/_11_ ),
    .ZN(\u_multiplier/LODy/z [21]));
 NOR4_X1 \u_multiplier/LODy/lod4_5/_17_  (.A1(sram_rdata_reg[22]),
    .A2(\u_multiplier/LODy/z [23]),
    .A3(sram_rdata_reg[21]),
    .A4(\u_multiplier/LODy/lod4_5/_09_ ),
    .ZN(\u_multiplier/LODy/z [20]));
 INV_X1 \u_multiplier/LODy/lod4_6/_12_  (.A(sram_rdata_reg[26]),
    .ZN(\u_multiplier/LODy/lod4_6/_10_ ));
 INV_X1 \u_multiplier/LODy/lod4_6/_13_  (.A(sram_rdata_reg[25]),
    .ZN(\u_multiplier/LODy/lod4_6/_11_ ));
 INV_X1 \u_multiplier/LODy/lod4_6/_14_  (.A(sram_rdata_reg[24]),
    .ZN(\u_multiplier/LODy/lod4_6/_09_ ));
 NOR2_X1 \u_multiplier/LODy/lod4_6/_15_  (.A1(\u_multiplier/LODy/lod4_6/_10_ ),
    .A2(\u_multiplier/LODy/z [27]),
    .ZN(\u_multiplier/LODy/z [26]));
 NOR3_X1 \u_multiplier/LODy/lod4_6/_16_  (.A1(sram_rdata_reg[26]),
    .A2(\u_multiplier/LODy/z [27]),
    .A3(\u_multiplier/LODy/lod4_6/_11_ ),
    .ZN(\u_multiplier/LODy/z [25]));
 NOR4_X1 \u_multiplier/LODy/lod4_6/_17_  (.A1(sram_rdata_reg[26]),
    .A2(\u_multiplier/LODy/z [27]),
    .A3(sram_rdata_reg[25]),
    .A4(\u_multiplier/LODy/lod4_6/_09_ ),
    .ZN(\u_multiplier/LODy/z [24]));
 INV_X1 \u_multiplier/LODy/lod4_7/_12_  (.A(sram_rdata_reg[30]),
    .ZN(\u_multiplier/LODy/lod4_7/_10_ ));
 INV_X1 \u_multiplier/LODy/lod4_7/_13_  (.A(sram_rdata_reg[29]),
    .ZN(\u_multiplier/LODy/lod4_7/_11_ ));
 INV_X1 \u_multiplier/LODy/lod4_7/_14_  (.A(sram_rdata_reg[28]),
    .ZN(\u_multiplier/LODy/lod4_7/_09_ ));
 NOR2_X1 \u_multiplier/LODy/lod4_7/_15_  (.A1(\u_multiplier/LODy/lod4_7/_10_ ),
    .A2(\u_multiplier/LODy/z [31]),
    .ZN(\u_multiplier/LODy/z [30]));
 NOR3_X1 \u_multiplier/LODy/lod4_7/_16_  (.A1(sram_rdata_reg[30]),
    .A2(\u_multiplier/LODy/z [31]),
    .A3(\u_multiplier/LODy/lod4_7/_11_ ),
    .ZN(\u_multiplier/LODy/z [29]));
 NOR4_X1 \u_multiplier/LODy/lod4_7/_17_  (.A1(sram_rdata_reg[30]),
    .A2(\u_multiplier/LODy/z [31]),
    .A3(sram_rdata_reg[29]),
    .A4(\u_multiplier/LODy/lod4_7/_09_ ),
    .ZN(\u_multiplier/LODy/z [28]));
 INV_X1 \u_multiplier/LODy/lod4_middle_high/_12_  (.A(\u_multiplier/LODy/_083_ ),
    .ZN(\u_multiplier/LODy/lod4_middle_high/_10_ ));
 INV_X1 \u_multiplier/LODy/lod4_middle_high/_13_  (.A(\u_multiplier/LODy/_082_ ),
    .ZN(\u_multiplier/LODy/lod4_middle_high/_11_ ));
 INV_X1 \u_multiplier/LODy/lod4_middle_high/_14_  (.A(\u_multiplier/LODy/_081_ ),
    .ZN(\u_multiplier/LODy/lod4_middle_high/_09_ ));
 NOR2_X1 \u_multiplier/LODy/lod4_middle_high/_15_  (.A1(\u_multiplier/LODy/lod4_middle_high/_10_ ),
    .A2(\u_multiplier/LODy/select_high [3]),
    .ZN(\u_multiplier/LODy/select_high [2]));
 NOR3_X1 \u_multiplier/LODy/lod4_middle_high/_16_  (.A1(\u_multiplier/LODy/_083_ ),
    .A2(\u_multiplier/LODy/select_high [3]),
    .A3(\u_multiplier/LODy/lod4_middle_high/_11_ ),
    .ZN(\u_multiplier/LODy/select_high [1]));
 NOR4_X1 \u_multiplier/LODy/lod4_middle_high/_17_  (.A1(\u_multiplier/LODy/_083_ ),
    .A2(\u_multiplier/LODy/select_high [3]),
    .A3(\u_multiplier/LODy/_082_ ),
    .A4(\u_multiplier/LODy/lod4_middle_high/_09_ ),
    .ZN(\u_multiplier/LODy/select_high [0]));
 INV_X1 \u_multiplier/LODy/lod4_middle_low/_12_  (.A(\u_multiplier/LODy/_079_ ),
    .ZN(\u_multiplier/LODy/lod4_middle_low/_10_ ));
 INV_X1 \u_multiplier/LODy/lod4_middle_low/_13_  (.A(\u_multiplier/LODy/_078_ ),
    .ZN(\u_multiplier/LODy/lod4_middle_low/_11_ ));
 INV_X1 \u_multiplier/LODy/lod4_middle_low/_14_  (.A(\u_multiplier/LODy/_077_ ),
    .ZN(\u_multiplier/LODy/lod4_middle_low/_09_ ));
 NOR2_X1 \u_multiplier/LODy/lod4_middle_low/_15_  (.A1(\u_multiplier/LODy/lod4_middle_low/_10_ ),
    .A2(\u_multiplier/LODy/select_low [3]),
    .ZN(\u_multiplier/LODy/select_low [2]));
 NOR3_X1 \u_multiplier/LODy/lod4_middle_low/_16_  (.A1(\u_multiplier/LODy/_079_ ),
    .A2(\u_multiplier/LODy/select_low [3]),
    .A3(\u_multiplier/LODy/lod4_middle_low/_11_ ),
    .ZN(\u_multiplier/LODy/select_low [1]));
 NOR4_X1 \u_multiplier/LODy/lod4_middle_low/_17_  (.A1(\u_multiplier/LODy/_079_ ),
    .A2(\u_multiplier/LODy/select_low [3]),
    .A3(\u_multiplier/LODy/_078_ ),
    .A4(\u_multiplier/LODy/lod4_middle_low/_09_ ),
    .ZN(\u_multiplier/LODy/select_low [0]));
 INV_X1 \u_multiplier/NOD/_15_  (.A(\u_multiplier/NOD/t_in [1]),
    .ZN(\u_multiplier/NOD/_11_ ));
 INV_X1 \u_multiplier/NOD/_16_  (.A(\u_multiplier/_1841_ ),
    .ZN(\u_multiplier/NOD/_12_ ));
 INV_X1 \u_multiplier/NOD/_17_  (.A(\u_multiplier/_1830_ ),
    .ZN(\u_multiplier/NOD/_13_ ));
 AND2_X1 \u_multiplier/NOD/_18_  (.A1(\u_multiplier/_1851_ ),
    .A2(\u_multiplier/_1853_ ),
    .ZN(\u_multiplier/NOD_Q1 [31]));
 NOR4_X1 \u_multiplier/NOD/_19_  (.A1(\u_multiplier/_1852_ ),
    .A2(\u_multiplier/NOD/_11_ ),
    .A3(\u_multiplier/NOD/_12_ ),
    .A4(\u_multiplier/_1830_ ),
    .ZN(\u_multiplier/NOD_Q1 [1]));
 NOR4_X1 \u_multiplier/NOD/_20_  (.A1(\u_multiplier/_1852_ ),
    .A2(\u_multiplier/NOD/_11_ ),
    .A3(\u_multiplier/_1841_ ),
    .A4(\u_multiplier/NOD/_13_ ),
    .ZN(\u_multiplier/NOD_Q1 [0]));
 AOI21_X1 \u_multiplier/NOD/nod_basic_unit31/_7_  (.A(\u_multiplier/_1853_ ),
    .B1(\u_multiplier/_1850_ ),
    .B2(\u_multiplier/_1851_ ),
    .ZN(\u_multiplier/NOD/nod_basic_unit31/_5_ ));
 AOI21_X2 \u_multiplier/NOD/nod_basic_unit31/_8_  (.A(\u_multiplier/NOD/nod_basic_unit31/_5_ ),
    .B1(\u_multiplier/_1853_ ),
    .B2(\u_multiplier/_1851_ ),
    .ZN(\u_multiplier/NOD_Q1 [30]));
 INV_X1 \u_multiplier/NOD/nod_cels[10].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [10]),
    .ZN(\u_multiplier/NOD/nod_cels[10].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[10].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[10].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[10].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[10].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[10].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1832_ ),
    .ZN(\u_multiplier/NOD/t_in [9]));
 NOR3_X1 \u_multiplier/NOD/nod_cels[10].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[10].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1832_ ),
    .A3(\u_multiplier/NOD/nod_cels[10].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [10]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[10].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1831_ ),
    .B1(\u_multiplier/_1859_ ),
    .B2(\u_multiplier/_1860_ ),
    .ZN(\u_multiplier/NOD/nod_cels[10].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[10].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[10].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1831_ ),
    .B2(\u_multiplier/_1860_ ),
    .ZN(\u_multiplier/NOD/nod_cels[10].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[11].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [11]),
    .ZN(\u_multiplier/NOD/nod_cels[11].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[11].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[11].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[11].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[11].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[11].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1833_ ),
    .ZN(\u_multiplier/NOD/t_in [10]));
 NOR3_X2 \u_multiplier/NOD/nod_cels[11].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[11].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1833_ ),
    .A3(\u_multiplier/NOD/nod_cels[11].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [11]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[11].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1832_ ),
    .B1(\u_multiplier/_1860_ ),
    .B2(\u_multiplier/_1831_ ),
    .ZN(\u_multiplier/NOD/nod_cels[11].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[11].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[11].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1832_ ),
    .B2(\u_multiplier/_1831_ ),
    .ZN(\u_multiplier/NOD/nod_cels[11].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[12].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [12]),
    .ZN(\u_multiplier/NOD/nod_cels[12].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[12].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[12].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[12].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[12].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[12].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1834_ ),
    .ZN(\u_multiplier/NOD/t_in [11]));
 NOR3_X1 \u_multiplier/NOD/nod_cels[12].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[12].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1834_ ),
    .A3(\u_multiplier/NOD/nod_cels[12].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [12]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[12].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1833_ ),
    .B1(\u_multiplier/_1831_ ),
    .B2(\u_multiplier/_1832_ ),
    .ZN(\u_multiplier/NOD/nod_cels[12].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[12].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[12].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1833_ ),
    .B2(\u_multiplier/_1832_ ),
    .ZN(\u_multiplier/NOD/nod_cels[12].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[13].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [13]),
    .ZN(\u_multiplier/NOD/nod_cels[13].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[13].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[13].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[13].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[13].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[13].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1835_ ),
    .ZN(\u_multiplier/NOD/t_in [12]));
 NOR3_X2 \u_multiplier/NOD/nod_cels[13].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[13].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1835_ ),
    .A3(\u_multiplier/NOD/nod_cels[13].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [13]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[13].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1834_ ),
    .B1(\u_multiplier/_1832_ ),
    .B2(\u_multiplier/_1833_ ),
    .ZN(\u_multiplier/NOD/nod_cels[13].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[13].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[13].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1834_ ),
    .B2(\u_multiplier/_1833_ ),
    .ZN(\u_multiplier/NOD/nod_cels[13].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[14].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [14]),
    .ZN(\u_multiplier/NOD/nod_cels[14].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[14].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[14].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[14].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[14].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[14].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1836_ ),
    .ZN(\u_multiplier/NOD/t_in [13]));
 NOR3_X2 \u_multiplier/NOD/nod_cels[14].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[14].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1836_ ),
    .A3(\u_multiplier/NOD/nod_cels[14].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [14]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[14].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1835_ ),
    .B1(\u_multiplier/_1833_ ),
    .B2(\u_multiplier/_1834_ ),
    .ZN(\u_multiplier/NOD/nod_cels[14].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[14].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[14].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1835_ ),
    .B2(\u_multiplier/_1834_ ),
    .ZN(\u_multiplier/NOD/nod_cels[14].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[15].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [15]),
    .ZN(\u_multiplier/NOD/nod_cels[15].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[15].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[15].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[15].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[15].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[15].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1837_ ),
    .ZN(\u_multiplier/NOD/t_in [14]));
 NOR3_X2 \u_multiplier/NOD/nod_cels[15].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[15].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1837_ ),
    .A3(\u_multiplier/NOD/nod_cels[15].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [15]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[15].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1836_ ),
    .B1(\u_multiplier/_1834_ ),
    .B2(\u_multiplier/_1835_ ),
    .ZN(\u_multiplier/NOD/nod_cels[15].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[15].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[15].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1836_ ),
    .B2(\u_multiplier/_1835_ ),
    .ZN(\u_multiplier/NOD/nod_cels[15].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[16].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [16]),
    .ZN(\u_multiplier/NOD/nod_cels[16].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[16].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[16].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[16].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[16].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[16].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1838_ ),
    .ZN(\u_multiplier/NOD/t_in [15]));
 NOR3_X1 \u_multiplier/NOD/nod_cels[16].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[16].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1838_ ),
    .A3(\u_multiplier/NOD/nod_cels[16].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [16]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[16].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1837_ ),
    .B1(\u_multiplier/_1835_ ),
    .B2(\u_multiplier/_1836_ ),
    .ZN(\u_multiplier/NOD/nod_cels[16].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[16].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[16].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1837_ ),
    .B2(\u_multiplier/_1836_ ),
    .ZN(\u_multiplier/NOD/nod_cels[16].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[17].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [17]),
    .ZN(\u_multiplier/NOD/nod_cels[17].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[17].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[17].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[17].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[17].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[17].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1839_ ),
    .ZN(\u_multiplier/NOD/t_in [16]));
 NOR3_X1 \u_multiplier/NOD/nod_cels[17].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[17].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1839_ ),
    .A3(\u_multiplier/NOD/nod_cels[17].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [17]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[17].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1838_ ),
    .B1(\u_multiplier/_1836_ ),
    .B2(\u_multiplier/_1837_ ),
    .ZN(\u_multiplier/NOD/nod_cels[17].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[17].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[17].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1838_ ),
    .B2(\u_multiplier/_1837_ ),
    .ZN(\u_multiplier/NOD/nod_cels[17].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[18].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [18]),
    .ZN(\u_multiplier/NOD/nod_cels[18].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[18].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[18].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[18].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[18].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[18].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1840_ ),
    .ZN(\u_multiplier/NOD/t_in [17]));
 NOR3_X1 \u_multiplier/NOD/nod_cels[18].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[18].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1840_ ),
    .A3(\u_multiplier/NOD/nod_cels[18].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [18]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[18].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1839_ ),
    .B1(\u_multiplier/_1837_ ),
    .B2(\u_multiplier/_1838_ ),
    .ZN(\u_multiplier/NOD/nod_cels[18].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[18].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[18].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1839_ ),
    .B2(\u_multiplier/_1838_ ),
    .ZN(\u_multiplier/NOD/nod_cels[18].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[19].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [19]),
    .ZN(\u_multiplier/NOD/nod_cels[19].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[19].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[19].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[19].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[19].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[19].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1842_ ),
    .ZN(\u_multiplier/NOD/t_in [18]));
 NOR3_X2 \u_multiplier/NOD/nod_cels[19].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[19].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1842_ ),
    .A3(\u_multiplier/NOD/nod_cels[19].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [19]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[19].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1840_ ),
    .B1(\u_multiplier/_1838_ ),
    .B2(\u_multiplier/_1839_ ),
    .ZN(\u_multiplier/NOD/nod_cels[19].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[19].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[19].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1840_ ),
    .B2(\u_multiplier/_1839_ ),
    .ZN(\u_multiplier/NOD/nod_cels[19].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[20].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [20]),
    .ZN(\u_multiplier/NOD/nod_cels[20].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[20].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[20].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[20].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[20].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[20].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1843_ ),
    .ZN(\u_multiplier/NOD/t_in [19]));
 NOR3_X1 \u_multiplier/NOD/nod_cels[20].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[20].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1843_ ),
    .A3(\u_multiplier/NOD/nod_cels[20].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [20]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[20].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1842_ ),
    .B1(\u_multiplier/_1839_ ),
    .B2(\u_multiplier/_1840_ ),
    .ZN(\u_multiplier/NOD/nod_cels[20].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[20].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[20].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1842_ ),
    .B2(\u_multiplier/_1840_ ),
    .ZN(\u_multiplier/NOD/nod_cels[20].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[21].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [21]),
    .ZN(\u_multiplier/NOD/nod_cels[21].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[21].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[21].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[21].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[21].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[21].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1844_ ),
    .ZN(\u_multiplier/NOD/t_in [20]));
 NOR3_X2 \u_multiplier/NOD/nod_cels[21].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[21].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1844_ ),
    .A3(\u_multiplier/NOD/nod_cels[21].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [21]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[21].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1843_ ),
    .B1(\u_multiplier/_1840_ ),
    .B2(\u_multiplier/_1842_ ),
    .ZN(\u_multiplier/NOD/nod_cels[21].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[21].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[21].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1843_ ),
    .B2(\u_multiplier/_1842_ ),
    .ZN(\u_multiplier/NOD/nod_cels[21].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[22].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [22]),
    .ZN(\u_multiplier/NOD/nod_cels[22].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[22].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[22].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[22].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[22].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[22].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1845_ ),
    .ZN(\u_multiplier/NOD/t_in [21]));
 NOR3_X2 \u_multiplier/NOD/nod_cels[22].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[22].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1845_ ),
    .A3(\u_multiplier/NOD/nod_cels[22].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [22]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[22].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1844_ ),
    .B1(\u_multiplier/_1842_ ),
    .B2(\u_multiplier/_1843_ ),
    .ZN(\u_multiplier/NOD/nod_cels[22].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[22].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[22].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1844_ ),
    .B2(\u_multiplier/_1843_ ),
    .ZN(\u_multiplier/NOD/nod_cels[22].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[23].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [23]),
    .ZN(\u_multiplier/NOD/nod_cels[23].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[23].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[23].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[23].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[23].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[23].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1846_ ),
    .ZN(\u_multiplier/NOD/t_in [22]));
 NOR3_X2 \u_multiplier/NOD/nod_cels[23].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[23].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1846_ ),
    .A3(\u_multiplier/NOD/nod_cels[23].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [23]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[23].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1845_ ),
    .B1(\u_multiplier/_1843_ ),
    .B2(\u_multiplier/_1844_ ),
    .ZN(\u_multiplier/NOD/nod_cels[23].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[23].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[23].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1845_ ),
    .B2(\u_multiplier/_1844_ ),
    .ZN(\u_multiplier/NOD/nod_cels[23].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[24].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [24]),
    .ZN(\u_multiplier/NOD/nod_cels[24].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[24].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[24].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[24].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[24].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[24].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1847_ ),
    .ZN(\u_multiplier/NOD/t_in [23]));
 NOR3_X2 \u_multiplier/NOD/nod_cels[24].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[24].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1847_ ),
    .A3(\u_multiplier/NOD/nod_cels[24].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [24]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[24].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1846_ ),
    .B1(\u_multiplier/_1844_ ),
    .B2(\u_multiplier/_1845_ ),
    .ZN(\u_multiplier/NOD/nod_cels[24].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[24].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[24].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1846_ ),
    .B2(\u_multiplier/_1845_ ),
    .ZN(\u_multiplier/NOD/nod_cels[24].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[25].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [25]),
    .ZN(\u_multiplier/NOD/nod_cels[25].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[25].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[25].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[25].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[25].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[25].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1848_ ),
    .ZN(\u_multiplier/NOD/t_in [24]));
 NOR3_X2 \u_multiplier/NOD/nod_cels[25].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[25].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1848_ ),
    .A3(\u_multiplier/NOD/nod_cels[25].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [25]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[25].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1847_ ),
    .B1(\u_multiplier/_1845_ ),
    .B2(\u_multiplier/_1846_ ),
    .ZN(\u_multiplier/NOD/nod_cels[25].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[25].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[25].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1847_ ),
    .B2(\u_multiplier/_1846_ ),
    .ZN(\u_multiplier/NOD/nod_cels[25].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[26].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [26]),
    .ZN(\u_multiplier/NOD/nod_cels[26].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[26].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[26].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[26].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[26].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[26].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1849_ ),
    .ZN(\u_multiplier/NOD/t_in [25]));
 NOR3_X2 \u_multiplier/NOD/nod_cels[26].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[26].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1849_ ),
    .A3(\u_multiplier/NOD/nod_cels[26].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [26]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[26].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1848_ ),
    .B1(\u_multiplier/_1846_ ),
    .B2(\u_multiplier/_1847_ ),
    .ZN(\u_multiplier/NOD/nod_cels[26].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[26].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[26].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1848_ ),
    .B2(\u_multiplier/_1847_ ),
    .ZN(\u_multiplier/NOD/nod_cels[26].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[27].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [27]),
    .ZN(\u_multiplier/NOD/nod_cels[27].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[27].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[27].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[27].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[27].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[27].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1850_ ),
    .ZN(\u_multiplier/NOD/t_in [26]));
 NOR3_X2 \u_multiplier/NOD/nod_cels[27].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[27].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1850_ ),
    .A3(\u_multiplier/NOD/nod_cels[27].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [27]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[27].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1849_ ),
    .B1(\u_multiplier/_1847_ ),
    .B2(\u_multiplier/_1848_ ),
    .ZN(\u_multiplier/NOD/nod_cels[27].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[27].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[27].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1849_ ),
    .B2(\u_multiplier/_1848_ ),
    .ZN(\u_multiplier/NOD/nod_cels[27].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[28].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [28]),
    .ZN(\u_multiplier/NOD/nod_cels[28].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[28].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[28].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[28].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[28].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[28].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1851_ ),
    .ZN(\u_multiplier/NOD/t_in [27]));
 NOR3_X4 \u_multiplier/NOD/nod_cels[28].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[28].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1851_ ),
    .A3(\u_multiplier/NOD/nod_cels[28].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [28]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[28].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1850_ ),
    .B1(\u_multiplier/_1848_ ),
    .B2(\u_multiplier/_1849_ ),
    .ZN(\u_multiplier/NOD/nod_cels[28].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[28].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[28].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1850_ ),
    .B2(\u_multiplier/_1849_ ),
    .ZN(\u_multiplier/NOD/nod_cels[28].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[29].Nod_bits/_07_  (.A(net125),
    .ZN(\u_multiplier/NOD/nod_cels[29].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[29].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[29].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[29].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[29].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[29].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1853_ ),
    .ZN(\u_multiplier/NOD/t_in [28]));
 NOR3_X2 \u_multiplier/NOD/nod_cels[29].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[29].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1853_ ),
    .A3(\u_multiplier/NOD/nod_cels[29].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [29]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[29].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1851_ ),
    .B1(\u_multiplier/_1849_ ),
    .B2(\u_multiplier/_1850_ ),
    .ZN(\u_multiplier/NOD/nod_cels[29].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[29].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[29].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1851_ ),
    .B2(\u_multiplier/_1850_ ),
    .ZN(\u_multiplier/NOD/nod_cels[29].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[2].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [2]),
    .ZN(\u_multiplier/NOD/nod_cels[2].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[2].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[2].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[2].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[2].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[2].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1854_ ),
    .ZN(\u_multiplier/NOD/t_in [1]));
 NOR3_X1 \u_multiplier/NOD/nod_cels[2].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[2].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1854_ ),
    .A3(\u_multiplier/NOD/nod_cels[2].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [2]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[2].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1852_ ),
    .B1(\u_multiplier/_1830_ ),
    .B2(\u_multiplier/_1841_ ),
    .ZN(\u_multiplier/NOD/nod_cels[2].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[2].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[2].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1852_ ),
    .B2(\u_multiplier/_1841_ ),
    .ZN(\u_multiplier/NOD/nod_cels[2].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[3].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [3]),
    .ZN(\u_multiplier/NOD/nod_cels[3].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[3].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[3].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[3].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[3].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[3].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1855_ ),
    .ZN(\u_multiplier/NOD/t_in [2]));
 NOR3_X2 \u_multiplier/NOD/nod_cels[3].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[3].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1855_ ),
    .A3(\u_multiplier/NOD/nod_cels[3].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [3]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[3].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1854_ ),
    .B1(\u_multiplier/_1841_ ),
    .B2(\u_multiplier/_1852_ ),
    .ZN(\u_multiplier/NOD/nod_cels[3].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[3].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[3].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1854_ ),
    .B2(\u_multiplier/_1852_ ),
    .ZN(\u_multiplier/NOD/nod_cels[3].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[4].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [4]),
    .ZN(\u_multiplier/NOD/nod_cels[4].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[4].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[4].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[4].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[4].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[4].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1856_ ),
    .ZN(\u_multiplier/NOD/t_in [3]));
 NOR3_X1 \u_multiplier/NOD/nod_cels[4].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[4].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1856_ ),
    .A3(\u_multiplier/NOD/nod_cels[4].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [4]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[4].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1855_ ),
    .B1(\u_multiplier/_1852_ ),
    .B2(\u_multiplier/_1854_ ),
    .ZN(\u_multiplier/NOD/nod_cels[4].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[4].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[4].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1855_ ),
    .B2(\u_multiplier/_1854_ ),
    .ZN(\u_multiplier/NOD/nod_cels[4].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[5].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [5]),
    .ZN(\u_multiplier/NOD/nod_cels[5].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[5].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[5].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[5].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[5].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[5].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1857_ ),
    .ZN(\u_multiplier/NOD/t_in [4]));
 NOR3_X1 \u_multiplier/NOD/nod_cels[5].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[5].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1857_ ),
    .A3(\u_multiplier/NOD/nod_cels[5].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [5]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[5].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1856_ ),
    .B1(\u_multiplier/_1854_ ),
    .B2(\u_multiplier/_1855_ ),
    .ZN(\u_multiplier/NOD/nod_cels[5].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[5].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[5].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1856_ ),
    .B2(\u_multiplier/_1855_ ),
    .ZN(\u_multiplier/NOD/nod_cels[5].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[6].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [6]),
    .ZN(\u_multiplier/NOD/nod_cels[6].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[6].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[6].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[6].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[6].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[6].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1858_ ),
    .ZN(\u_multiplier/NOD/t_in [5]));
 NOR3_X1 \u_multiplier/NOD/nod_cels[6].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[6].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1858_ ),
    .A3(\u_multiplier/NOD/nod_cels[6].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [6]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[6].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1857_ ),
    .B1(\u_multiplier/_1855_ ),
    .B2(\u_multiplier/_1856_ ),
    .ZN(\u_multiplier/NOD/nod_cels[6].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[6].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[6].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1857_ ),
    .B2(\u_multiplier/_1856_ ),
    .ZN(\u_multiplier/NOD/nod_cels[6].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[7].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [7]),
    .ZN(\u_multiplier/NOD/nod_cels[7].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[7].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[7].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[7].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[7].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[7].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1859_ ),
    .ZN(\u_multiplier/NOD/t_in [6]));
 NOR3_X4 \u_multiplier/NOD/nod_cels[7].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[7].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1859_ ),
    .A3(\u_multiplier/NOD/nod_cels[7].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [7]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[7].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1858_ ),
    .B1(\u_multiplier/_1856_ ),
    .B2(\u_multiplier/_1857_ ),
    .ZN(\u_multiplier/NOD/nod_cels[7].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[7].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[7].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1858_ ),
    .B2(\u_multiplier/_1857_ ),
    .ZN(\u_multiplier/NOD/nod_cels[7].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[8].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [8]),
    .ZN(\u_multiplier/NOD/nod_cels[8].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[8].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[8].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[8].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[8].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[8].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1860_ ),
    .ZN(\u_multiplier/NOD/t_in [7]));
 NOR3_X1 \u_multiplier/NOD/nod_cels[8].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[8].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1860_ ),
    .A3(\u_multiplier/NOD/nod_cels[8].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [8]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[8].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1859_ ),
    .B1(\u_multiplier/_1857_ ),
    .B2(\u_multiplier/_1858_ ),
    .ZN(\u_multiplier/NOD/nod_cels[8].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[8].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[8].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1859_ ),
    .B2(\u_multiplier/_1858_ ),
    .ZN(\u_multiplier/NOD/nod_cels[8].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[9].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [9]),
    .ZN(\u_multiplier/NOD/nod_cels[9].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[9].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[9].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[9].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[9].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[9].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1831_ ),
    .ZN(\u_multiplier/NOD/t_in [8]));
 NOR3_X1 \u_multiplier/NOD/nod_cels[9].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[9].Nod_bits/_02_ ),
    .A2(\u_multiplier/_1831_ ),
    .A3(\u_multiplier/NOD/nod_cels[9].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [9]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[9].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_1860_ ),
    .B1(\u_multiplier/_1858_ ),
    .B2(\u_multiplier/_1859_ ),
    .ZN(\u_multiplier/NOD/nod_cels[9].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[9].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[9].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_1860_ ),
    .B2(\u_multiplier/_1859_ ),
    .ZN(\u_multiplier/NOD/nod_cels[9].Nod_bits/tmp1 ));
 NOR3_X1 \u_multiplier/PE/code0/_36_  (.A1(\u_multiplier/NOD_Q1 [17]),
    .A2(\u_multiplier/NOD_Q1 [9]),
    .A3(\u_multiplier/NOD_Q1 [23]),
    .ZN(\u_multiplier/PE/code0/_31_ ));
 NOR3_X1 \u_multiplier/PE/code0/_37_  (.A1(\u_multiplier/NOD_Q1 [3]),
    .A2(\u_multiplier/NOD_Q1 [27]),
    .A3(\u_multiplier/NOD_Q1 [15]),
    .ZN(\u_multiplier/PE/code0/_32_ ));
 NOR4_X1 \u_multiplier/PE/code0/_38_  (.A1(\u_multiplier/NOD_Q1 [5]),
    .A2(\u_multiplier/NOD_Q1 [29]),
    .A3(\u_multiplier/NOD_Q1 [19]),
    .A4(\u_multiplier/NOD_Q1 [11]),
    .ZN(\u_multiplier/PE/code0/_33_ ));
 NOR4_X1 \u_multiplier/PE/code0/_39_  (.A1(\u_multiplier/NOD_Q1 [1]),
    .A2(\u_multiplier/NOD_Q1 [21]),
    .A3(\u_multiplier/NOD_Q1 [13]),
    .A4(\u_multiplier/NOD_Q1 [31]),
    .ZN(\u_multiplier/PE/code0/_34_ ));
 NAND4_X1 \u_multiplier/PE/code0/_40_  (.A1(\u_multiplier/PE/code0/_31_ ),
    .A2(\u_multiplier/PE/code0/_32_ ),
    .A3(\u_multiplier/PE/code0/_33_ ),
    .A4(\u_multiplier/PE/code0/_34_ ),
    .ZN(\u_multiplier/PE/code0/_35_ ));
 OR3_X4 \u_multiplier/PE/code0/_41_  (.A1(\u_multiplier/NOD_Q1 [25]),
    .A2(\u_multiplier/NOD_Q1 [7]),
    .A3(\u_multiplier/PE/code0/_35_ ),
    .ZN(\u_multiplier/K [0]));
 NOR3_X1 \u_multiplier/PE/code1/_36_  (.A1(\u_multiplier/NOD_Q1 [18]),
    .A2(\u_multiplier/NOD_Q1 [10]),
    .A3(\u_multiplier/NOD_Q1 [23]),
    .ZN(\u_multiplier/PE/code1/_31_ ));
 NOR3_X1 \u_multiplier/PE/code1/_37_  (.A1(\u_multiplier/NOD_Q1 [3]),
    .A2(\u_multiplier/NOD_Q1 [27]),
    .A3(\u_multiplier/NOD_Q1 [15]),
    .ZN(\u_multiplier/PE/code1/_32_ ));
 NOR4_X1 \u_multiplier/PE/code1/_38_  (.A1(\u_multiplier/NOD_Q1 [6]),
    .A2(\u_multiplier/NOD_Q1 [30]),
    .A3(\u_multiplier/NOD_Q1 [19]),
    .A4(\u_multiplier/NOD_Q1 [11]),
    .ZN(\u_multiplier/PE/code1/_33_ ));
 NOR4_X1 \u_multiplier/PE/code1/_39_  (.A1(\u_multiplier/NOD_Q1 [2]),
    .A2(\u_multiplier/NOD_Q1 [22]),
    .A3(\u_multiplier/NOD_Q1 [14]),
    .A4(\u_multiplier/NOD_Q1 [31]),
    .ZN(\u_multiplier/PE/code1/_34_ ));
 NAND4_X1 \u_multiplier/PE/code1/_40_  (.A1(\u_multiplier/PE/code1/_31_ ),
    .A2(\u_multiplier/PE/code1/_32_ ),
    .A3(\u_multiplier/PE/code1/_33_ ),
    .A4(\u_multiplier/PE/code1/_34_ ),
    .ZN(\u_multiplier/PE/code1/_35_ ));
 OR3_X4 \u_multiplier/PE/code1/_41_  (.A1(\u_multiplier/NOD_Q1 [26]),
    .A2(\u_multiplier/NOD_Q1 [7]),
    .A3(\u_multiplier/PE/code1/_35_ ),
    .ZN(\u_multiplier/K [1]));
 NOR3_X1 \u_multiplier/PE/code2/_36_  (.A1(\u_multiplier/NOD_Q1 [20]),
    .A2(\u_multiplier/NOD_Q1 [12]),
    .A3(\u_multiplier/NOD_Q1 [23]),
    .ZN(\u_multiplier/PE/code2/_31_ ));
 NOR3_X1 \u_multiplier/PE/code2/_37_  (.A1(\u_multiplier/NOD_Q1 [5]),
    .A2(\u_multiplier/NOD_Q1 [29]),
    .A3(\u_multiplier/NOD_Q1 [15]),
    .ZN(\u_multiplier/PE/code2/_32_ ));
 NOR4_X1 \u_multiplier/PE/code2/_38_  (.A1(\u_multiplier/NOD_Q1 [6]),
    .A2(\u_multiplier/NOD_Q1 [30]),
    .A3(\u_multiplier/NOD_Q1 [21]),
    .A4(\u_multiplier/NOD_Q1 [13]),
    .ZN(\u_multiplier/PE/code2/_33_ ));
 NOR4_X1 \u_multiplier/PE/code2/_39_  (.A1(\u_multiplier/NOD_Q1 [4]),
    .A2(\u_multiplier/NOD_Q1 [22]),
    .A3(\u_multiplier/NOD_Q1 [14]),
    .A4(\u_multiplier/NOD_Q1 [31]),
    .ZN(\u_multiplier/PE/code2/_34_ ));
 NAND4_X1 \u_multiplier/PE/code2/_40_  (.A1(\u_multiplier/PE/code2/_31_ ),
    .A2(\u_multiplier/PE/code2/_32_ ),
    .A3(\u_multiplier/PE/code2/_33_ ),
    .A4(\u_multiplier/PE/code2/_34_ ),
    .ZN(\u_multiplier/PE/code2/_35_ ));
 OR3_X4 \u_multiplier/PE/code2/_41_  (.A1(\u_multiplier/NOD_Q1 [28]),
    .A2(\u_multiplier/NOD_Q1 [7]),
    .A3(\u_multiplier/PE/code2/_35_ ),
    .ZN(\u_multiplier/K [2]));
 NOR3_X1 \u_multiplier/PE/code3/_36_  (.A1(\u_multiplier/NOD_Q1 [24]),
    .A2(\u_multiplier/NOD_Q1 [12]),
    .A3(\u_multiplier/NOD_Q1 [27]),
    .ZN(\u_multiplier/PE/code3/_31_ ));
 NOR3_X1 \u_multiplier/PE/code3/_37_  (.A1(\u_multiplier/NOD_Q1 [9]),
    .A2(\u_multiplier/NOD_Q1 [29]),
    .A3(\u_multiplier/NOD_Q1 [15]),
    .ZN(\u_multiplier/PE/code3/_32_ ));
 NOR4_X1 \u_multiplier/PE/code3/_38_  (.A1(\u_multiplier/NOD_Q1 [10]),
    .A2(\u_multiplier/NOD_Q1 [30]),
    .A3(\u_multiplier/NOD_Q1 [25]),
    .A4(\u_multiplier/NOD_Q1 [13]),
    .ZN(\u_multiplier/PE/code3/_33_ ));
 NOR4_X1 \u_multiplier/PE/code3/_39_  (.A1(\u_multiplier/NOD_Q1 [8]),
    .A2(\u_multiplier/NOD_Q1 [26]),
    .A3(\u_multiplier/NOD_Q1 [14]),
    .A4(\u_multiplier/NOD_Q1 [31]),
    .ZN(\u_multiplier/PE/code3/_34_ ));
 NAND4_X1 \u_multiplier/PE/code3/_40_  (.A1(\u_multiplier/PE/code3/_31_ ),
    .A2(\u_multiplier/PE/code3/_32_ ),
    .A3(\u_multiplier/PE/code3/_33_ ),
    .A4(\u_multiplier/PE/code3/_34_ ),
    .ZN(\u_multiplier/PE/code3/_35_ ));
 OR3_X4 \u_multiplier/PE/code3/_41_  (.A1(\u_multiplier/NOD_Q1 [28]),
    .A2(\u_multiplier/NOD_Q1 [11]),
    .A3(\u_multiplier/PE/code3/_35_ ),
    .ZN(\u_multiplier/K [3]));
 NOR3_X1 \u_multiplier/PE/code4/_36_  (.A1(\u_multiplier/NOD_Q1 [24]),
    .A2(\u_multiplier/NOD_Q1 [20]),
    .A3(\u_multiplier/NOD_Q1 [27]),
    .ZN(\u_multiplier/PE/code4/_31_ ));
 NOR3_X1 \u_multiplier/PE/code4/_37_  (.A1(\u_multiplier/NOD_Q1 [17]),
    .A2(\u_multiplier/NOD_Q1 [29]),
    .A3(\u_multiplier/NOD_Q1 [23]),
    .ZN(\u_multiplier/PE/code4/_32_ ));
 NOR4_X1 \u_multiplier/PE/code4/_38_  (.A1(\u_multiplier/NOD_Q1 [18]),
    .A2(\u_multiplier/NOD_Q1 [30]),
    .A3(\u_multiplier/NOD_Q1 [25]),
    .A4(\u_multiplier/NOD_Q1 [21]),
    .ZN(\u_multiplier/PE/code4/_33_ ));
 NOR4_X1 \u_multiplier/PE/code4/_39_  (.A1(\u_multiplier/NOD_Q1 [16]),
    .A2(\u_multiplier/NOD_Q1 [26]),
    .A3(\u_multiplier/NOD_Q1 [22]),
    .A4(\u_multiplier/NOD_Q1 [31]),
    .ZN(\u_multiplier/PE/code4/_34_ ));
 NAND4_X1 \u_multiplier/PE/code4/_40_  (.A1(\u_multiplier/PE/code4/_31_ ),
    .A2(\u_multiplier/PE/code4/_32_ ),
    .A3(\u_multiplier/PE/code4/_33_ ),
    .A4(\u_multiplier/PE/code4/_34_ ),
    .ZN(\u_multiplier/PE/code4/_35_ ));
 OR3_X4 \u_multiplier/PE/code4/_41_  (.A1(\u_multiplier/NOD_Q1 [28]),
    .A2(\u_multiplier/NOD_Q1 [19]),
    .A3(\u_multiplier/PE/code4/_35_ ),
    .ZN(\u_multiplier/K [4]));
 NOR3_X1 \u_multiplier/PEx/code0/_36_  (.A1(\u_multiplier/kx [17]),
    .A2(\u_multiplier/kx [9]),
    .A3(\u_multiplier/kx [23]),
    .ZN(\u_multiplier/PEx/code0/_31_ ));
 NOR3_X1 \u_multiplier/PEx/code0/_37_  (.A1(\u_multiplier/kx [3]),
    .A2(\u_multiplier/kx [27]),
    .A3(\u_multiplier/kx [15]),
    .ZN(\u_multiplier/PEx/code0/_32_ ));
 NOR4_X1 \u_multiplier/PEx/code0/_38_  (.A1(\u_multiplier/kx [5]),
    .A2(\u_multiplier/kx [29]),
    .A3(\u_multiplier/kx [19]),
    .A4(\u_multiplier/kx [11]),
    .ZN(\u_multiplier/PEx/code0/_33_ ));
 NOR4_X1 \u_multiplier/PEx/code0/_39_  (.A1(\u_multiplier/kx [1]),
    .A2(\u_multiplier/kx [21]),
    .A3(\u_multiplier/kx [13]),
    .A4(\u_multiplier/kx [31]),
    .ZN(\u_multiplier/PEx/code0/_34_ ));
 NAND4_X1 \u_multiplier/PEx/code0/_40_  (.A1(\u_multiplier/PEx/code0/_31_ ),
    .A2(\u_multiplier/PEx/code0/_32_ ),
    .A3(\u_multiplier/PEx/code0/_33_ ),
    .A4(\u_multiplier/PEx/code0/_34_ ),
    .ZN(\u_multiplier/PEx/code0/_35_ ));
 OR3_X4 \u_multiplier/PEx/code0/_41_  (.A1(\u_multiplier/kx [25]),
    .A2(\u_multiplier/kx [7]),
    .A3(\u_multiplier/PEx/code0/_35_ ),
    .ZN(\u_multiplier/code_x [0]));
 NOR3_X1 \u_multiplier/PEx/code1/_36_  (.A1(\u_multiplier/kx [18]),
    .A2(\u_multiplier/kx [10]),
    .A3(\u_multiplier/kx [23]),
    .ZN(\u_multiplier/PEx/code1/_31_ ));
 NOR3_X1 \u_multiplier/PEx/code1/_37_  (.A1(\u_multiplier/kx [3]),
    .A2(\u_multiplier/kx [27]),
    .A3(\u_multiplier/kx [15]),
    .ZN(\u_multiplier/PEx/code1/_32_ ));
 NOR4_X1 \u_multiplier/PEx/code1/_38_  (.A1(\u_multiplier/kx [6]),
    .A2(\u_multiplier/kx [30]),
    .A3(\u_multiplier/kx [19]),
    .A4(\u_multiplier/kx [11]),
    .ZN(\u_multiplier/PEx/code1/_33_ ));
 NOR4_X1 \u_multiplier/PEx/code1/_39_  (.A1(\u_multiplier/kx [2]),
    .A2(\u_multiplier/kx [22]),
    .A3(\u_multiplier/kx [14]),
    .A4(\u_multiplier/kx [31]),
    .ZN(\u_multiplier/PEx/code1/_34_ ));
 NAND4_X1 \u_multiplier/PEx/code1/_40_  (.A1(\u_multiplier/PEx/code1/_31_ ),
    .A2(\u_multiplier/PEx/code1/_32_ ),
    .A3(\u_multiplier/PEx/code1/_33_ ),
    .A4(\u_multiplier/PEx/code1/_34_ ),
    .ZN(\u_multiplier/PEx/code1/_35_ ));
 OR3_X4 \u_multiplier/PEx/code1/_41_  (.A1(\u_multiplier/kx [26]),
    .A2(\u_multiplier/kx [7]),
    .A3(\u_multiplier/PEx/code1/_35_ ),
    .ZN(\u_multiplier/code_x [1]));
 NOR3_X1 \u_multiplier/PEx/code2/_36_  (.A1(\u_multiplier/kx [20]),
    .A2(\u_multiplier/kx [12]),
    .A3(\u_multiplier/kx [23]),
    .ZN(\u_multiplier/PEx/code2/_31_ ));
 NOR3_X1 \u_multiplier/PEx/code2/_37_  (.A1(\u_multiplier/kx [5]),
    .A2(\u_multiplier/kx [29]),
    .A3(\u_multiplier/kx [15]),
    .ZN(\u_multiplier/PEx/code2/_32_ ));
 NOR4_X1 \u_multiplier/PEx/code2/_38_  (.A1(\u_multiplier/kx [6]),
    .A2(\u_multiplier/kx [30]),
    .A3(\u_multiplier/kx [21]),
    .A4(\u_multiplier/kx [13]),
    .ZN(\u_multiplier/PEx/code2/_33_ ));
 NOR4_X1 \u_multiplier/PEx/code2/_39_  (.A1(\u_multiplier/kx [4]),
    .A2(\u_multiplier/kx [22]),
    .A3(\u_multiplier/kx [14]),
    .A4(\u_multiplier/kx [31]),
    .ZN(\u_multiplier/PEx/code2/_34_ ));
 NAND4_X1 \u_multiplier/PEx/code2/_40_  (.A1(\u_multiplier/PEx/code2/_31_ ),
    .A2(\u_multiplier/PEx/code2/_32_ ),
    .A3(\u_multiplier/PEx/code2/_33_ ),
    .A4(\u_multiplier/PEx/code2/_34_ ),
    .ZN(\u_multiplier/PEx/code2/_35_ ));
 OR3_X4 \u_multiplier/PEx/code2/_41_  (.A1(\u_multiplier/kx [28]),
    .A2(\u_multiplier/kx [7]),
    .A3(\u_multiplier/PEx/code2/_35_ ),
    .ZN(\u_multiplier/code_x [2]));
 NOR3_X1 \u_multiplier/PEx/code3/_36_  (.A1(\u_multiplier/kx [24]),
    .A2(\u_multiplier/kx [12]),
    .A3(\u_multiplier/kx [27]),
    .ZN(\u_multiplier/PEx/code3/_31_ ));
 NOR3_X1 \u_multiplier/PEx/code3/_37_  (.A1(\u_multiplier/kx [9]),
    .A2(\u_multiplier/kx [29]),
    .A3(\u_multiplier/kx [15]),
    .ZN(\u_multiplier/PEx/code3/_32_ ));
 NOR4_X1 \u_multiplier/PEx/code3/_38_  (.A1(\u_multiplier/kx [10]),
    .A2(\u_multiplier/kx [30]),
    .A3(\u_multiplier/kx [25]),
    .A4(\u_multiplier/kx [13]),
    .ZN(\u_multiplier/PEx/code3/_33_ ));
 NOR4_X1 \u_multiplier/PEx/code3/_39_  (.A1(\u_multiplier/kx [8]),
    .A2(\u_multiplier/kx [26]),
    .A3(\u_multiplier/kx [14]),
    .A4(\u_multiplier/kx [31]),
    .ZN(\u_multiplier/PEx/code3/_34_ ));
 NAND4_X1 \u_multiplier/PEx/code3/_40_  (.A1(\u_multiplier/PEx/code3/_31_ ),
    .A2(\u_multiplier/PEx/code3/_32_ ),
    .A3(\u_multiplier/PEx/code3/_33_ ),
    .A4(\u_multiplier/PEx/code3/_34_ ),
    .ZN(\u_multiplier/PEx/code3/_35_ ));
 OR3_X4 \u_multiplier/PEx/code3/_41_  (.A1(\u_multiplier/kx [28]),
    .A2(\u_multiplier/kx [11]),
    .A3(\u_multiplier/PEx/code3/_35_ ),
    .ZN(\u_multiplier/code_x [3]));
 NOR3_X1 \u_multiplier/PEx/code4/_36_  (.A1(\u_multiplier/kx [24]),
    .A2(\u_multiplier/kx [20]),
    .A3(\u_multiplier/kx [27]),
    .ZN(\u_multiplier/PEx/code4/_31_ ));
 NOR3_X1 \u_multiplier/PEx/code4/_37_  (.A1(\u_multiplier/kx [17]),
    .A2(\u_multiplier/kx [29]),
    .A3(\u_multiplier/kx [23]),
    .ZN(\u_multiplier/PEx/code4/_32_ ));
 NOR4_X1 \u_multiplier/PEx/code4/_38_  (.A1(\u_multiplier/kx [18]),
    .A2(\u_multiplier/kx [30]),
    .A3(\u_multiplier/kx [25]),
    .A4(\u_multiplier/kx [21]),
    .ZN(\u_multiplier/PEx/code4/_33_ ));
 NOR4_X1 \u_multiplier/PEx/code4/_39_  (.A1(\u_multiplier/kx [16]),
    .A2(\u_multiplier/kx [26]),
    .A3(\u_multiplier/kx [22]),
    .A4(\u_multiplier/kx [31]),
    .ZN(\u_multiplier/PEx/code4/_34_ ));
 NAND4_X1 \u_multiplier/PEx/code4/_40_  (.A1(\u_multiplier/PEx/code4/_31_ ),
    .A2(\u_multiplier/PEx/code4/_32_ ),
    .A3(\u_multiplier/PEx/code4/_33_ ),
    .A4(\u_multiplier/PEx/code4/_34_ ),
    .ZN(\u_multiplier/PEx/code4/_35_ ));
 OR3_X4 \u_multiplier/PEx/code4/_41_  (.A1(\u_multiplier/kx [28]),
    .A2(\u_multiplier/kx [19]),
    .A3(\u_multiplier/PEx/code4/_35_ ),
    .ZN(\u_multiplier/code_x [4]));
 NOR3_X1 \u_multiplier/PEy/code0/_36_  (.A1(\u_multiplier/ky [17]),
    .A2(\u_multiplier/ky [9]),
    .A3(\u_multiplier/ky [23]),
    .ZN(\u_multiplier/PEy/code0/_31_ ));
 NOR3_X1 \u_multiplier/PEy/code0/_37_  (.A1(\u_multiplier/ky [3]),
    .A2(\u_multiplier/ky [27]),
    .A3(\u_multiplier/ky [15]),
    .ZN(\u_multiplier/PEy/code0/_32_ ));
 NOR4_X1 \u_multiplier/PEy/code0/_38_  (.A1(\u_multiplier/ky [5]),
    .A2(\u_multiplier/ky [29]),
    .A3(\u_multiplier/ky [19]),
    .A4(\u_multiplier/ky [11]),
    .ZN(\u_multiplier/PEy/code0/_33_ ));
 NOR4_X1 \u_multiplier/PEy/code0/_39_  (.A1(\u_multiplier/ky [1]),
    .A2(\u_multiplier/ky [21]),
    .A3(\u_multiplier/ky [13]),
    .A4(\u_multiplier/ky [31]),
    .ZN(\u_multiplier/PEy/code0/_34_ ));
 NAND4_X1 \u_multiplier/PEy/code0/_40_  (.A1(\u_multiplier/PEy/code0/_31_ ),
    .A2(\u_multiplier/PEy/code0/_32_ ),
    .A3(\u_multiplier/PEy/code0/_33_ ),
    .A4(\u_multiplier/PEy/code0/_34_ ),
    .ZN(\u_multiplier/PEy/code0/_35_ ));
 OR3_X4 \u_multiplier/PEy/code0/_41_  (.A1(\u_multiplier/ky [25]),
    .A2(\u_multiplier/ky [7]),
    .A3(\u_multiplier/PEy/code0/_35_ ),
    .ZN(\u_multiplier/code_y [0]));
 NOR3_X1 \u_multiplier/PEy/code1/_36_  (.A1(\u_multiplier/ky [18]),
    .A2(\u_multiplier/ky [10]),
    .A3(\u_multiplier/ky [23]),
    .ZN(\u_multiplier/PEy/code1/_31_ ));
 NOR3_X1 \u_multiplier/PEy/code1/_37_  (.A1(\u_multiplier/ky [3]),
    .A2(\u_multiplier/ky [27]),
    .A3(\u_multiplier/ky [15]),
    .ZN(\u_multiplier/PEy/code1/_32_ ));
 NOR4_X1 \u_multiplier/PEy/code1/_38_  (.A1(\u_multiplier/ky [6]),
    .A2(\u_multiplier/ky [30]),
    .A3(\u_multiplier/ky [19]),
    .A4(\u_multiplier/ky [11]),
    .ZN(\u_multiplier/PEy/code1/_33_ ));
 NOR4_X1 \u_multiplier/PEy/code1/_39_  (.A1(\u_multiplier/ky [2]),
    .A2(\u_multiplier/ky [22]),
    .A3(\u_multiplier/ky [14]),
    .A4(\u_multiplier/ky [31]),
    .ZN(\u_multiplier/PEy/code1/_34_ ));
 NAND4_X1 \u_multiplier/PEy/code1/_40_  (.A1(\u_multiplier/PEy/code1/_31_ ),
    .A2(\u_multiplier/PEy/code1/_32_ ),
    .A3(\u_multiplier/PEy/code1/_33_ ),
    .A4(\u_multiplier/PEy/code1/_34_ ),
    .ZN(\u_multiplier/PEy/code1/_35_ ));
 OR3_X4 \u_multiplier/PEy/code1/_41_  (.A1(\u_multiplier/ky [26]),
    .A2(\u_multiplier/ky [7]),
    .A3(\u_multiplier/PEy/code1/_35_ ),
    .ZN(\u_multiplier/code_y [1]));
 NOR3_X1 \u_multiplier/PEy/code2/_36_  (.A1(\u_multiplier/ky [20]),
    .A2(\u_multiplier/ky [12]),
    .A3(\u_multiplier/ky [23]),
    .ZN(\u_multiplier/PEy/code2/_31_ ));
 NOR3_X1 \u_multiplier/PEy/code2/_37_  (.A1(\u_multiplier/ky [5]),
    .A2(\u_multiplier/ky [29]),
    .A3(\u_multiplier/ky [15]),
    .ZN(\u_multiplier/PEy/code2/_32_ ));
 NOR4_X1 \u_multiplier/PEy/code2/_38_  (.A1(\u_multiplier/ky [6]),
    .A2(\u_multiplier/ky [30]),
    .A3(\u_multiplier/ky [21]),
    .A4(\u_multiplier/ky [13]),
    .ZN(\u_multiplier/PEy/code2/_33_ ));
 NOR4_X1 \u_multiplier/PEy/code2/_39_  (.A1(\u_multiplier/ky [4]),
    .A2(\u_multiplier/ky [22]),
    .A3(\u_multiplier/ky [14]),
    .A4(\u_multiplier/ky [31]),
    .ZN(\u_multiplier/PEy/code2/_34_ ));
 NAND4_X1 \u_multiplier/PEy/code2/_40_  (.A1(\u_multiplier/PEy/code2/_31_ ),
    .A2(\u_multiplier/PEy/code2/_32_ ),
    .A3(\u_multiplier/PEy/code2/_33_ ),
    .A4(\u_multiplier/PEy/code2/_34_ ),
    .ZN(\u_multiplier/PEy/code2/_35_ ));
 OR3_X4 \u_multiplier/PEy/code2/_41_  (.A1(\u_multiplier/ky [28]),
    .A2(\u_multiplier/ky [7]),
    .A3(\u_multiplier/PEy/code2/_35_ ),
    .ZN(\u_multiplier/code_y [2]));
 NOR3_X1 \u_multiplier/PEy/code3/_36_  (.A1(\u_multiplier/ky [24]),
    .A2(\u_multiplier/ky [12]),
    .A3(\u_multiplier/ky [27]),
    .ZN(\u_multiplier/PEy/code3/_31_ ));
 NOR3_X1 \u_multiplier/PEy/code3/_37_  (.A1(\u_multiplier/ky [9]),
    .A2(\u_multiplier/ky [29]),
    .A3(\u_multiplier/ky [15]),
    .ZN(\u_multiplier/PEy/code3/_32_ ));
 NOR4_X1 \u_multiplier/PEy/code3/_38_  (.A1(\u_multiplier/ky [10]),
    .A2(\u_multiplier/ky [30]),
    .A3(\u_multiplier/ky [25]),
    .A4(\u_multiplier/ky [13]),
    .ZN(\u_multiplier/PEy/code3/_33_ ));
 NOR4_X1 \u_multiplier/PEy/code3/_39_  (.A1(\u_multiplier/ky [8]),
    .A2(\u_multiplier/ky [26]),
    .A3(\u_multiplier/ky [14]),
    .A4(\u_multiplier/ky [31]),
    .ZN(\u_multiplier/PEy/code3/_34_ ));
 NAND4_X1 \u_multiplier/PEy/code3/_40_  (.A1(\u_multiplier/PEy/code3/_31_ ),
    .A2(\u_multiplier/PEy/code3/_32_ ),
    .A3(\u_multiplier/PEy/code3/_33_ ),
    .A4(\u_multiplier/PEy/code3/_34_ ),
    .ZN(\u_multiplier/PEy/code3/_35_ ));
 OR3_X4 \u_multiplier/PEy/code3/_41_  (.A1(\u_multiplier/ky [28]),
    .A2(\u_multiplier/ky [11]),
    .A3(\u_multiplier/PEy/code3/_35_ ),
    .ZN(\u_multiplier/code_y [3]));
 NOR3_X1 \u_multiplier/PEy/code4/_36_  (.A1(\u_multiplier/ky [24]),
    .A2(\u_multiplier/ky [20]),
    .A3(\u_multiplier/ky [27]),
    .ZN(\u_multiplier/PEy/code4/_31_ ));
 NOR3_X1 \u_multiplier/PEy/code4/_37_  (.A1(\u_multiplier/ky [17]),
    .A2(\u_multiplier/ky [29]),
    .A3(\u_multiplier/ky [23]),
    .ZN(\u_multiplier/PEy/code4/_32_ ));
 NOR4_X1 \u_multiplier/PEy/code4/_38_  (.A1(\u_multiplier/ky [18]),
    .A2(\u_multiplier/ky [30]),
    .A3(\u_multiplier/ky [25]),
    .A4(\u_multiplier/ky [21]),
    .ZN(\u_multiplier/PEy/code4/_33_ ));
 NOR4_X1 \u_multiplier/PEy/code4/_39_  (.A1(\u_multiplier/ky [16]),
    .A2(\u_multiplier/ky [26]),
    .A3(\u_multiplier/ky [22]),
    .A4(\u_multiplier/ky [31]),
    .ZN(\u_multiplier/PEy/code4/_34_ ));
 NAND4_X1 \u_multiplier/PEy/code4/_40_  (.A1(\u_multiplier/PEy/code4/_31_ ),
    .A2(\u_multiplier/PEy/code4/_32_ ),
    .A3(\u_multiplier/PEy/code4/_33_ ),
    .A4(\u_multiplier/PEy/code4/_34_ ),
    .ZN(\u_multiplier/PEy/code4/_35_ ));
 OR3_X4 \u_multiplier/PEy/code4/_41_  (.A1(\u_multiplier/ky [28]),
    .A2(\u_multiplier/ky [19]),
    .A3(\u_multiplier/PEy/code4/_35_ ),
    .ZN(\u_multiplier/code_y [4]));
 INV_X4 \u_multiplier/_3880_  (.A(\u_multiplier/code_y [0]),
    .ZN(\u_multiplier/_3105_ ));
 INV_X16 \u_multiplier/_3881_  (.A(\u_multiplier/code_y [2]),
    .ZN(\u_multiplier/_3106_ ));
 INV_X16 \u_multiplier/_3882_  (.A(\u_multiplier/code_y [3]),
    .ZN(\u_multiplier/_3107_ ));
 INV_X8 \u_multiplier/_3883_  (.A(\u_multiplier/code_y [4]),
    .ZN(\u_multiplier/_3108_ ));
 INV_X8 \u_multiplier/_3884_  (.A(\u_multiplier/code_x [4]),
    .ZN(\u_multiplier/_3109_ ));
 INV_X8 \u_multiplier/_3885_  (.A(\u_multiplier/code_x [2]),
    .ZN(\u_multiplier/_3110_ ));
 INV_X16 \u_multiplier/_3886_  (.A(\u_multiplier/code_x [3]),
    .ZN(\u_multiplier/_3111_ ));
 INV_X8 \u_multiplier/_3887_  (.A(\u_multiplier/K [2]),
    .ZN(\u_multiplier/_3112_ ));
 INV_X8 \u_multiplier/_3888_  (.A(\u_multiplier/K [0]),
    .ZN(\u_multiplier/_3113_ ));
 INV_X8 \u_multiplier/_3889_  (.A(\u_multiplier/K [1]),
    .ZN(\u_multiplier/_3114_ ));
 INV_X16 \u_multiplier/_3890_  (.A(\u_multiplier/K [3]),
    .ZN(\u_multiplier/_3115_ ));
 INV_X16 \u_multiplier/_3891_  (.A(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_3116_ ));
 INV_X1 \u_multiplier/_3892_  (.A(\u_multiplier/dec_out [9]),
    .ZN(\u_multiplier/_3117_ ));
 INV_X1 \u_multiplier/_3893_  (.A(\u_multiplier/dec_out [14]),
    .ZN(\u_multiplier/_3118_ ));
 INV_X1 \u_multiplier/_3894_  (.A(\u_multiplier/dec_out [16]),
    .ZN(\u_multiplier/_3119_ ));
 INV_X1 \u_multiplier/_3895_  (.A(\u_multiplier/dec_out [18]),
    .ZN(\u_multiplier/_3120_ ));
 INV_X1 \u_multiplier/_3896_  (.A(\u_multiplier/dec_out [54]),
    .ZN(\u_multiplier/_3121_ ));
 INV_X1 \u_multiplier/_3897_  (.A(\u_multiplier/dec_out [55]),
    .ZN(\u_multiplier/_3122_ ));
 INV_X1 \u_multiplier/_3898_  (.A(\u_multiplier/dec_out [56]),
    .ZN(\u_multiplier/_3123_ ));
 INV_X1 \u_multiplier/_3899_  (.A(\u_multiplier/dec_out [57]),
    .ZN(\u_multiplier/_3124_ ));
 INV_X1 \u_multiplier/_3900_  (.A(\u_multiplier/dec_out [61]),
    .ZN(\u_multiplier/_3125_ ));
 INV_X1 \u_multiplier/_3901_  (.A(\u_multiplier/dec_out [62]),
    .ZN(\u_multiplier/_3126_ ));
 XNOR2_X2 \u_multiplier/_3902_  (.A(\u_multiplier/ky [0]),
    .B(sram_rdata_reg[0]),
    .ZN(\u_multiplier/_3127_ ));
 XOR2_X2 \u_multiplier/_3903_  (.A(\u_multiplier/ky [0]),
    .B(sram_rdata_reg[0]),
    .Z(\u_multiplier/_3128_ ));
 XOR2_X2 \u_multiplier/_3904_  (.A(\u_multiplier/kx [30]),
    .B(_0683_[30]),
    .Z(\u_multiplier/_3129_ ));
 XNOR2_X2 \u_multiplier/_3905_  (.A(\u_multiplier/kx [30]),
    .B(_0683_[30]),
    .ZN(\u_multiplier/_3130_ ));
 XOR2_X2 \u_multiplier/_3906_  (.A(\u_multiplier/ky [30]),
    .B(sram_rdata_reg[30]),
    .Z(\u_multiplier/_3131_ ));
 NOR2_X1 \u_multiplier/_3907_  (.A1(\u_multiplier/_3130_ ),
    .A2(\u_multiplier/_3131_ ),
    .ZN(\u_multiplier/_3132_ ));
 XOR2_X2 \u_multiplier/_3908_  (.A(\u_multiplier/ky [6]),
    .B(sram_rdata_reg[6]),
    .Z(\u_multiplier/_3133_ ));
 XNOR2_X1 \u_multiplier/_3909_  (.A(\u_multiplier/kx [6]),
    .B(data_in_reg[6]),
    .ZN(\u_multiplier/_3134_ ));
 XOR2_X2 \u_multiplier/_3910_  (.A(\u_multiplier/kx [6]),
    .B(data_in_reg[6]),
    .Z(\u_multiplier/_3135_ ));
 NOR2_X1 \u_multiplier/_3911_  (.A1(\u_multiplier/_3133_ ),
    .A2(\u_multiplier/_3134_ ),
    .ZN(\u_multiplier/_3136_ ));
 XOR2_X2 \u_multiplier/_3912_  (.A(\u_multiplier/ky [5]),
    .B(sram_rdata_reg[5]),
    .Z(\u_multiplier/_3137_ ));
 XNOR2_X2 \u_multiplier/_3913_  (.A(\u_multiplier/ky [5]),
    .B(sram_rdata_reg[5]),
    .ZN(\u_multiplier/_3138_ ));
 XOR2_X2 \u_multiplier/_3914_  (.A(\u_multiplier/kx [5]),
    .B(data_in_reg[5]),
    .Z(\u_multiplier/_3139_ ));
 OR2_X1 \u_multiplier/_3915_  (.A1(\u_multiplier/_3138_ ),
    .A2(\u_multiplier/_3139_ ),
    .ZN(\u_multiplier/_3140_ ));
 XOR2_X2 \u_multiplier/_3916_  (.A(\u_multiplier/ky [1]),
    .B(sram_rdata_reg[1]),
    .Z(\u_multiplier/_3141_ ));
 XNOR2_X1 \u_multiplier/_3917_  (.A(\u_multiplier/ky [1]),
    .B(sram_rdata_reg[1]),
    .ZN(\u_multiplier/_3142_ ));
 XNOR2_X2 \u_multiplier/_3918_  (.A(\u_multiplier/kx [1]),
    .B(data_in_reg[1]),
    .ZN(\u_multiplier/_3143_ ));
 XOR2_X1 \u_multiplier/_3919_  (.A(\u_multiplier/kx [1]),
    .B(data_in_reg[1]),
    .Z(\u_multiplier/_3144_ ));
 XNOR2_X2 \u_multiplier/_3920_  (.A(\u_multiplier/kx [0]),
    .B(data_in_reg[0]),
    .ZN(\u_multiplier/_3145_ ));
 XOR2_X2 \u_multiplier/_3921_  (.A(\u_multiplier/kx [0]),
    .B(data_in_reg[0]),
    .Z(\u_multiplier/_3146_ ));
 OAI22_X1 \u_multiplier/_3922_  (.A1(\u_multiplier/_3141_ ),
    .A2(\u_multiplier/_3143_ ),
    .B1(\u_multiplier/_3145_ ),
    .B2(\u_multiplier/_3128_ ),
    .ZN(\u_multiplier/_3147_ ));
 XOR2_X2 \u_multiplier/_3923_  (.A(\u_multiplier/ky [2]),
    .B(sram_rdata_reg[2]),
    .Z(\u_multiplier/_3148_ ));
 XNOR2_X1 \u_multiplier/_3924_  (.A(\u_multiplier/ky [2]),
    .B(sram_rdata_reg[2]),
    .ZN(\u_multiplier/_3149_ ));
 XNOR2_X2 \u_multiplier/_3925_  (.A(\u_multiplier/kx [2]),
    .B(data_in_reg[2]),
    .ZN(\u_multiplier/_3150_ ));
 XOR2_X1 \u_multiplier/_3926_  (.A(\u_multiplier/kx [2]),
    .B(data_in_reg[2]),
    .Z(\u_multiplier/_3151_ ));
 AOI22_X1 \u_multiplier/_3927_  (.A1(\u_multiplier/_3141_ ),
    .A2(\u_multiplier/_3143_ ),
    .B1(\u_multiplier/_3148_ ),
    .B2(\u_multiplier/_3150_ ),
    .ZN(\u_multiplier/_3152_ ));
 XOR2_X2 \u_multiplier/_3928_  (.A(\u_multiplier/ky [3]),
    .B(\u_multiplier/LODy/z [3]),
    .Z(\u_multiplier/_3153_ ));
 XNOR2_X1 \u_multiplier/_3929_  (.A(\u_multiplier/ky [3]),
    .B(\u_multiplier/LODy/z [3]),
    .ZN(\u_multiplier/_3154_ ));
 XNOR2_X2 \u_multiplier/_3930_  (.A(\u_multiplier/kx [3]),
    .B(\u_multiplier/LODx/z [3]),
    .ZN(\u_multiplier/_3155_ ));
 OAI22_X1 \u_multiplier/_3931_  (.A1(\u_multiplier/_3148_ ),
    .A2(\u_multiplier/_3150_ ),
    .B1(\u_multiplier/_3153_ ),
    .B2(\u_multiplier/_3155_ ),
    .ZN(\u_multiplier/_3156_ ));
 AOI21_X1 \u_multiplier/_3932_  (.A(\u_multiplier/_3156_ ),
    .B1(\u_multiplier/_3152_ ),
    .B2(\u_multiplier/_3147_ ),
    .ZN(\u_multiplier/_3157_ ));
 XOR2_X2 \u_multiplier/_3933_  (.A(\u_multiplier/ky [4]),
    .B(sram_rdata_reg[4]),
    .Z(\u_multiplier/_3158_ ));
 XNOR2_X2 \u_multiplier/_3934_  (.A(\u_multiplier/ky [4]),
    .B(sram_rdata_reg[4]),
    .ZN(\u_multiplier/_3159_ ));
 XNOR2_X1 \u_multiplier/_3935_  (.A(\u_multiplier/kx [4]),
    .B(data_in_reg[4]),
    .ZN(\u_multiplier/_3160_ ));
 XOR2_X2 \u_multiplier/_3936_  (.A(\u_multiplier/kx [4]),
    .B(data_in_reg[4]),
    .Z(\u_multiplier/_3161_ ));
 NAND2_X1 \u_multiplier/_3937_  (.A1(\u_multiplier/_3153_ ),
    .A2(\u_multiplier/_3155_ ),
    .ZN(\u_multiplier/_3162_ ));
 OAI21_X1 \u_multiplier/_3938_  (.A(\u_multiplier/_3162_ ),
    .B1(\u_multiplier/_3161_ ),
    .B2(\u_multiplier/_3159_ ),
    .ZN(\u_multiplier/_3163_ ));
 AOI22_X1 \u_multiplier/_3939_  (.A1(\u_multiplier/_3138_ ),
    .A2(\u_multiplier/_3139_ ),
    .B1(\u_multiplier/_3159_ ),
    .B2(\u_multiplier/_3161_ ),
    .ZN(\u_multiplier/_3164_ ));
 OAI21_X1 \u_multiplier/_3940_  (.A(\u_multiplier/_3164_ ),
    .B1(\u_multiplier/_3163_ ),
    .B2(\u_multiplier/_3157_ ),
    .ZN(\u_multiplier/_3165_ ));
 AOI21_X1 \u_multiplier/_3941_  (.A(\u_multiplier/_3136_ ),
    .B1(\u_multiplier/_3140_ ),
    .B2(\u_multiplier/_3165_ ),
    .ZN(\u_multiplier/_3166_ ));
 XOR2_X2 \u_multiplier/_3942_  (.A(\u_multiplier/ky [7]),
    .B(\u_multiplier/LODy/z [7]),
    .Z(\u_multiplier/_3167_ ));
 XNOR2_X2 \u_multiplier/_3943_  (.A(\u_multiplier/ky [7]),
    .B(\u_multiplier/LODy/z [7]),
    .ZN(\u_multiplier/_3168_ ));
 XOR2_X2 \u_multiplier/_3944_  (.A(\u_multiplier/kx [7]),
    .B(\u_multiplier/LODx/z [7]),
    .Z(\u_multiplier/_3169_ ));
 NAND2_X1 \u_multiplier/_3945_  (.A1(\u_multiplier/_3133_ ),
    .A2(\u_multiplier/_3134_ ),
    .ZN(\u_multiplier/_3170_ ));
 OAI21_X1 \u_multiplier/_3946_  (.A(\u_multiplier/_3170_ ),
    .B1(\u_multiplier/_3169_ ),
    .B2(\u_multiplier/_3168_ ),
    .ZN(\u_multiplier/_3171_ ));
 XOR2_X2 \u_multiplier/_3947_  (.A(\u_multiplier/ky [10]),
    .B(sram_rdata_reg[10]),
    .Z(\u_multiplier/_3172_ ));
 INV_X1 \u_multiplier/_3948_  (.A(\u_multiplier/_3172_ ),
    .ZN(\u_multiplier/_3173_ ));
 XOR2_X2 \u_multiplier/_3949_  (.A(\u_multiplier/kx [10]),
    .B(data_in_reg[10]),
    .Z(\u_multiplier/_3174_ ));
 XOR2_X2 \u_multiplier/_3950_  (.A(\u_multiplier/ky [11]),
    .B(\u_multiplier/LODy/z [11]),
    .Z(\u_multiplier/_3175_ ));
 XNOR2_X2 \u_multiplier/_3951_  (.A(\u_multiplier/ky [11]),
    .B(\u_multiplier/LODy/z [11]),
    .ZN(\u_multiplier/_3176_ ));
 XOR2_X2 \u_multiplier/_3952_  (.A(\u_multiplier/kx [11]),
    .B(\u_multiplier/LODx/z [11]),
    .Z(\u_multiplier/_3177_ ));
 NOR2_X1 \u_multiplier/_3953_  (.A1(\u_multiplier/_3176_ ),
    .A2(\u_multiplier/_3177_ ),
    .ZN(\u_multiplier/_3178_ ));
 AND2_X1 \u_multiplier/_3954_  (.A1(\u_multiplier/_3176_ ),
    .A2(\u_multiplier/_3177_ ),
    .ZN(\u_multiplier/_3179_ ));
 XOR2_X1 \u_multiplier/_3955_  (.A(\u_multiplier/_3172_ ),
    .B(\u_multiplier/_3174_ ),
    .Z(\u_multiplier/_3180_ ));
 OR3_X1 \u_multiplier/_3956_  (.A1(\u_multiplier/_3178_ ),
    .A2(\u_multiplier/_3179_ ),
    .A3(\u_multiplier/_3180_ ),
    .ZN(\u_multiplier/_3181_ ));
 XOR2_X2 \u_multiplier/_3957_  (.A(\u_multiplier/ky [8]),
    .B(sram_rdata_reg[8]),
    .Z(\u_multiplier/_3182_ ));
 INV_X1 \u_multiplier/_3958_  (.A(\u_multiplier/_3182_ ),
    .ZN(\u_multiplier/_3183_ ));
 XOR2_X2 \u_multiplier/_3959_  (.A(\u_multiplier/kx [8]),
    .B(data_in_reg[8]),
    .Z(\u_multiplier/_3184_ ));
 NAND2_X1 \u_multiplier/_3960_  (.A1(\u_multiplier/_3168_ ),
    .A2(\u_multiplier/_3169_ ),
    .ZN(\u_multiplier/_3185_ ));
 XOR2_X2 \u_multiplier/_3961_  (.A(\u_multiplier/ky [9]),
    .B(sram_rdata_reg[9]),
    .Z(\u_multiplier/_3186_ ));
 XNOR2_X1 \u_multiplier/_3962_  (.A(\u_multiplier/kx [9]),
    .B(data_in_reg[9]),
    .ZN(\u_multiplier/_3187_ ));
 XOR2_X2 \u_multiplier/_3963_  (.A(\u_multiplier/kx [9]),
    .B(data_in_reg[9]),
    .Z(\u_multiplier/_3188_ ));
 NAND2_X1 \u_multiplier/_3964_  (.A1(\u_multiplier/_3186_ ),
    .A2(\u_multiplier/_3187_ ),
    .ZN(\u_multiplier/_3189_ ));
 OR2_X1 \u_multiplier/_3965_  (.A1(\u_multiplier/_3186_ ),
    .A2(\u_multiplier/_3187_ ),
    .ZN(\u_multiplier/_3190_ ));
 XOR2_X1 \u_multiplier/_3966_  (.A(\u_multiplier/_3182_ ),
    .B(\u_multiplier/_3184_ ),
    .Z(\u_multiplier/_3191_ ));
 NAND3_X1 \u_multiplier/_3967_  (.A1(\u_multiplier/_3185_ ),
    .A2(\u_multiplier/_3189_ ),
    .A3(\u_multiplier/_3190_ ),
    .ZN(\u_multiplier/_3192_ ));
 NOR3_X1 \u_multiplier/_3968_  (.A1(\u_multiplier/_3181_ ),
    .A2(\u_multiplier/_3191_ ),
    .A3(\u_multiplier/_3192_ ),
    .ZN(\u_multiplier/_3193_ ));
 OAI21_X1 \u_multiplier/_3969_  (.A(\u_multiplier/_3193_ ),
    .B1(\u_multiplier/_3171_ ),
    .B2(\u_multiplier/_3166_ ),
    .ZN(\u_multiplier/_3194_ ));
 OAI21_X1 \u_multiplier/_3970_  (.A(\u_multiplier/_3189_ ),
    .B1(\u_multiplier/_3184_ ),
    .B2(\u_multiplier/_3183_ ),
    .ZN(\u_multiplier/_3195_ ));
 NAND2_X1 \u_multiplier/_3971_  (.A1(\u_multiplier/_3190_ ),
    .A2(\u_multiplier/_3195_ ),
    .ZN(\u_multiplier/_3196_ ));
 NOR2_X1 \u_multiplier/_3972_  (.A1(\u_multiplier/_3181_ ),
    .A2(\u_multiplier/_3196_ ),
    .ZN(\u_multiplier/_3197_ ));
 NOR3_X1 \u_multiplier/_3973_  (.A1(\u_multiplier/_3173_ ),
    .A2(\u_multiplier/_3174_ ),
    .A3(\u_multiplier/_3179_ ),
    .ZN(\u_multiplier/_3198_ ));
 NOR3_X1 \u_multiplier/_3974_  (.A1(\u_multiplier/_3178_ ),
    .A2(\u_multiplier/_3197_ ),
    .A3(\u_multiplier/_3198_ ),
    .ZN(\u_multiplier/_3199_ ));
 XOR2_X2 \u_multiplier/_3975_  (.A(\u_multiplier/ky [14]),
    .B(sram_rdata_reg[14]),
    .Z(\u_multiplier/_3200_ ));
 XNOR2_X2 \u_multiplier/_3976_  (.A(\u_multiplier/ky [14]),
    .B(sram_rdata_reg[14]),
    .ZN(\u_multiplier/_3201_ ));
 XOR2_X2 \u_multiplier/_3977_  (.A(\u_multiplier/kx [14]),
    .B(data_in_reg[14]),
    .Z(\u_multiplier/_3202_ ));
 OR2_X1 \u_multiplier/_3978_  (.A1(\u_multiplier/_3201_ ),
    .A2(\u_multiplier/_3202_ ),
    .ZN(\u_multiplier/_3203_ ));
 XOR2_X2 \u_multiplier/_3979_  (.A(\u_multiplier/ky [15]),
    .B(\u_multiplier/LODy/z [15]),
    .Z(\u_multiplier/_3204_ ));
 XNOR2_X1 \u_multiplier/_3980_  (.A(\u_multiplier/kx [15]),
    .B(\u_multiplier/LODx/z [15]),
    .ZN(\u_multiplier/_3205_ ));
 XOR2_X2 \u_multiplier/_3981_  (.A(\u_multiplier/kx [15]),
    .B(\u_multiplier/LODx/z [15]),
    .Z(\u_multiplier/_3206_ ));
 NAND2_X1 \u_multiplier/_3982_  (.A1(\u_multiplier/_3204_ ),
    .A2(\u_multiplier/_3205_ ),
    .ZN(\u_multiplier/_3207_ ));
 NOR2_X1 \u_multiplier/_3983_  (.A1(\u_multiplier/_3204_ ),
    .A2(\u_multiplier/_3205_ ),
    .ZN(\u_multiplier/_3208_ ));
 AOI21_X1 \u_multiplier/_3984_  (.A(\u_multiplier/_3208_ ),
    .B1(\u_multiplier/_3202_ ),
    .B2(\u_multiplier/_3201_ ),
    .ZN(\u_multiplier/_3209_ ));
 AND3_X1 \u_multiplier/_3985_  (.A1(\u_multiplier/_3203_ ),
    .A2(\u_multiplier/_3207_ ),
    .A3(\u_multiplier/_3209_ ),
    .ZN(\u_multiplier/_3210_ ));
 XOR2_X2 \u_multiplier/_3986_  (.A(\u_multiplier/ky [13]),
    .B(sram_rdata_reg[13]),
    .Z(\u_multiplier/_3211_ ));
 XNOR2_X1 \u_multiplier/_3987_  (.A(\u_multiplier/kx [13]),
    .B(data_in_reg[13]),
    .ZN(\u_multiplier/_3212_ ));
 XOR2_X2 \u_multiplier/_3988_  (.A(\u_multiplier/kx [13]),
    .B(data_in_reg[13]),
    .Z(\u_multiplier/_3213_ ));
 NAND2_X1 \u_multiplier/_3989_  (.A1(\u_multiplier/_3211_ ),
    .A2(\u_multiplier/_3212_ ),
    .ZN(\u_multiplier/_3214_ ));
 XOR2_X2 \u_multiplier/_3990_  (.A(\u_multiplier/ky [12]),
    .B(sram_rdata_reg[12]),
    .Z(\u_multiplier/_3215_ ));
 XOR2_X2 \u_multiplier/_3991_  (.A(\u_multiplier/kx [12]),
    .B(data_in_reg[12]),
    .Z(\u_multiplier/_3216_ ));
 INV_X1 \u_multiplier/_3992_  (.A(\u_multiplier/_3216_ ),
    .ZN(\u_multiplier/_3217_ ));
 NAND2_X1 \u_multiplier/_3993_  (.A1(\u_multiplier/_3215_ ),
    .A2(\u_multiplier/_3217_ ),
    .ZN(\u_multiplier/_3218_ ));
 NAND2_X1 \u_multiplier/_3994_  (.A1(\u_multiplier/_3214_ ),
    .A2(\u_multiplier/_3218_ ),
    .ZN(\u_multiplier/_3219_ ));
 OR2_X1 \u_multiplier/_3995_  (.A1(\u_multiplier/_3211_ ),
    .A2(\u_multiplier/_3212_ ),
    .ZN(\u_multiplier/_3220_ ));
 XNOR2_X1 \u_multiplier/_3996_  (.A(\u_multiplier/_3215_ ),
    .B(\u_multiplier/_3216_ ),
    .ZN(\u_multiplier/_3221_ ));
 NAND4_X1 \u_multiplier/_3997_  (.A1(\u_multiplier/_3210_ ),
    .A2(\u_multiplier/_3214_ ),
    .A3(\u_multiplier/_3220_ ),
    .A4(\u_multiplier/_3221_ ),
    .ZN(\u_multiplier/_3222_ ));
 AOI21_X1 \u_multiplier/_3998_  (.A(\u_multiplier/_3222_ ),
    .B1(\u_multiplier/_3199_ ),
    .B2(\u_multiplier/_3194_ ),
    .ZN(\u_multiplier/_3223_ ));
 NAND3_X1 \u_multiplier/_3999_  (.A1(\u_multiplier/_3210_ ),
    .A2(\u_multiplier/_3219_ ),
    .A3(\u_multiplier/_3220_ ),
    .ZN(\u_multiplier/_3224_ ));
 OAI211_X1 \u_multiplier/_4000_  (.A(\u_multiplier/_3207_ ),
    .B(\u_multiplier/_3224_ ),
    .C1(\u_multiplier/_3208_ ),
    .C2(\u_multiplier/_3203_ ),
    .ZN(\u_multiplier/_3225_ ));
 XOR2_X2 \u_multiplier/_4001_  (.A(\u_multiplier/ky [22]),
    .B(sram_rdata_reg[22]),
    .Z(\u_multiplier/_3226_ ));
 XOR2_X2 \u_multiplier/_4002_  (.A(\u_multiplier/kx [22]),
    .B(data_in_reg[22]),
    .Z(\u_multiplier/_3227_ ));
 INV_X1 \u_multiplier/_4003_  (.A(\u_multiplier/_3227_ ),
    .ZN(\u_multiplier/_3228_ ));
 XOR2_X2 \u_multiplier/_4004_  (.A(\u_multiplier/kx [23]),
    .B(\u_multiplier/LODx/z [23]),
    .Z(\u_multiplier/_3229_ ));
 XNOR2_X2 \u_multiplier/_4005_  (.A(\u_multiplier/ky [23]),
    .B(\u_multiplier/LODy/z [23]),
    .ZN(\u_multiplier/_3230_ ));
 XOR2_X2 \u_multiplier/_4006_  (.A(\u_multiplier/ky [23]),
    .B(\u_multiplier/LODy/z [23]),
    .Z(\u_multiplier/_3231_ ));
 NOR2_X1 \u_multiplier/_4007_  (.A1(\u_multiplier/_3229_ ),
    .A2(\u_multiplier/_3230_ ),
    .ZN(\u_multiplier/_3232_ ));
 NAND2_X1 \u_multiplier/_4008_  (.A1(\u_multiplier/_3229_ ),
    .A2(\u_multiplier/_3230_ ),
    .ZN(\u_multiplier/_3233_ ));
 OAI21_X1 \u_multiplier/_4009_  (.A(\u_multiplier/_3233_ ),
    .B1(\u_multiplier/_3228_ ),
    .B2(\u_multiplier/_3226_ ),
    .ZN(\u_multiplier/_3234_ ));
 AOI211_X2 \u_multiplier/_4010_  (.A(\u_multiplier/_3232_ ),
    .B(\u_multiplier/_3234_ ),
    .C1(\u_multiplier/_3226_ ),
    .C2(\u_multiplier/_3228_ ),
    .ZN(\u_multiplier/_3235_ ));
 XOR2_X2 \u_multiplier/_4011_  (.A(\u_multiplier/kx [21]),
    .B(data_in_reg[21]),
    .Z(\u_multiplier/_3236_ ));
 XNOR2_X2 \u_multiplier/_4012_  (.A(\u_multiplier/ky [21]),
    .B(sram_rdata_reg[21]),
    .ZN(\u_multiplier/_3237_ ));
 XOR2_X2 \u_multiplier/_4013_  (.A(\u_multiplier/ky [21]),
    .B(sram_rdata_reg[21]),
    .Z(\u_multiplier/_3238_ ));
 NAND2_X1 \u_multiplier/_4014_  (.A1(\u_multiplier/_3236_ ),
    .A2(\u_multiplier/_3237_ ),
    .ZN(\u_multiplier/_3239_ ));
 XOR2_X2 \u_multiplier/_4015_  (.A(\u_multiplier/kx [20]),
    .B(data_in_reg[20]),
    .Z(\u_multiplier/_3240_ ));
 XOR2_X2 \u_multiplier/_4016_  (.A(\u_multiplier/ky [20]),
    .B(sram_rdata_reg[20]),
    .Z(\u_multiplier/_3241_ ));
 INV_X1 \u_multiplier/_4017_  (.A(\u_multiplier/_3241_ ),
    .ZN(\u_multiplier/_3242_ ));
 OR2_X1 \u_multiplier/_4018_  (.A1(\u_multiplier/_3236_ ),
    .A2(\u_multiplier/_3237_ ),
    .ZN(\u_multiplier/_3243_ ));
 XNOR2_X1 \u_multiplier/_4019_  (.A(\u_multiplier/_3240_ ),
    .B(\u_multiplier/_3241_ ),
    .ZN(\u_multiplier/_3244_ ));
 NAND4_X1 \u_multiplier/_4020_  (.A1(\u_multiplier/_3235_ ),
    .A2(\u_multiplier/_3239_ ),
    .A3(\u_multiplier/_3243_ ),
    .A4(\u_multiplier/_3244_ ),
    .ZN(\u_multiplier/_3245_ ));
 XOR2_X2 \u_multiplier/_4021_  (.A(\u_multiplier/kx [19]),
    .B(\u_multiplier/LODx/z [19]),
    .Z(\u_multiplier/_3246_ ));
 XNOR2_X2 \u_multiplier/_4022_  (.A(\u_multiplier/ky [19]),
    .B(\u_multiplier/LODy/z [19]),
    .ZN(\u_multiplier/_3247_ ));
 XOR2_X2 \u_multiplier/_4023_  (.A(\u_multiplier/ky [19]),
    .B(\u_multiplier/LODy/z [19]),
    .Z(\u_multiplier/_3248_ ));
 NOR2_X1 \u_multiplier/_4024_  (.A1(\u_multiplier/_3246_ ),
    .A2(\u_multiplier/_3247_ ),
    .ZN(\u_multiplier/_3249_ ));
 XOR2_X2 \u_multiplier/_4025_  (.A(\u_multiplier/ky [18]),
    .B(sram_rdata_reg[18]),
    .Z(\u_multiplier/_3250_ ));
 INV_X1 \u_multiplier/_4026_  (.A(\u_multiplier/_3250_ ),
    .ZN(\u_multiplier/_3251_ ));
 XOR2_X2 \u_multiplier/_4027_  (.A(\u_multiplier/kx [18]),
    .B(data_in_reg[18]),
    .Z(\u_multiplier/_3252_ ));
 XNOR2_X1 \u_multiplier/_4028_  (.A(\u_multiplier/_3246_ ),
    .B(\u_multiplier/_3247_ ),
    .ZN(\u_multiplier/_3253_ ));
 AOI21_X1 \u_multiplier/_4029_  (.A(\u_multiplier/_3253_ ),
    .B1(\u_multiplier/_3252_ ),
    .B2(\u_multiplier/_3251_ ),
    .ZN(\u_multiplier/_3254_ ));
 XOR2_X2 \u_multiplier/_4030_  (.A(\u_multiplier/kx [17]),
    .B(data_in_reg[17]),
    .Z(\u_multiplier/_3255_ ));
 XNOR2_X1 \u_multiplier/_4031_  (.A(\u_multiplier/kx [17]),
    .B(data_in_reg[17]),
    .ZN(\u_multiplier/_3256_ ));
 XOR2_X2 \u_multiplier/_4032_  (.A(\u_multiplier/ky [17]),
    .B(sram_rdata_reg[17]),
    .Z(\u_multiplier/_3257_ ));
 NOR2_X1 \u_multiplier/_4033_  (.A1(\u_multiplier/_3256_ ),
    .A2(\u_multiplier/_3257_ ),
    .ZN(\u_multiplier/_3258_ ));
 OAI21_X1 \u_multiplier/_4034_  (.A(\u_multiplier/_3254_ ),
    .B1(\u_multiplier/_3252_ ),
    .B2(\u_multiplier/_3251_ ),
    .ZN(\u_multiplier/_3259_ ));
 XNOR2_X1 \u_multiplier/_4035_  (.A(\u_multiplier/kx [16]),
    .B(data_in_reg[16]),
    .ZN(\u_multiplier/_3260_ ));
 XOR2_X2 \u_multiplier/_4036_  (.A(\u_multiplier/kx [16]),
    .B(data_in_reg[16]),
    .Z(\u_multiplier/_3261_ ));
 XOR2_X2 \u_multiplier/_4037_  (.A(\u_multiplier/ky [16]),
    .B(sram_rdata_reg[16]),
    .Z(\u_multiplier/_3262_ ));
 AOI22_X1 \u_multiplier/_4038_  (.A1(\u_multiplier/_3256_ ),
    .A2(\u_multiplier/_3257_ ),
    .B1(\u_multiplier/_3260_ ),
    .B2(\u_multiplier/_3262_ ),
    .ZN(\u_multiplier/_3263_ ));
 OAI21_X1 \u_multiplier/_4039_  (.A(\u_multiplier/_3263_ ),
    .B1(\u_multiplier/_3262_ ),
    .B2(\u_multiplier/_3260_ ),
    .ZN(\u_multiplier/_3264_ ));
 NOR4_X1 \u_multiplier/_4040_  (.A1(\u_multiplier/_3245_ ),
    .A2(\u_multiplier/_3258_ ),
    .A3(\u_multiplier/_3259_ ),
    .A4(\u_multiplier/_3264_ ),
    .ZN(\u_multiplier/_3265_ ));
 OAI21_X1 \u_multiplier/_4041_  (.A(\u_multiplier/_3265_ ),
    .B1(\u_multiplier/_3225_ ),
    .B2(\u_multiplier/_3223_ ),
    .ZN(\u_multiplier/_3266_ ));
 OAI21_X1 \u_multiplier/_4042_  (.A(\u_multiplier/_3243_ ),
    .B1(\u_multiplier/_3242_ ),
    .B2(\u_multiplier/_3240_ ),
    .ZN(\u_multiplier/_3267_ ));
 NAND3_X1 \u_multiplier/_4043_  (.A1(\u_multiplier/_3235_ ),
    .A2(\u_multiplier/_3239_ ),
    .A3(\u_multiplier/_3267_ ),
    .ZN(\u_multiplier/_3268_ ));
 NAND3_X1 \u_multiplier/_4044_  (.A1(\u_multiplier/_3226_ ),
    .A2(\u_multiplier/_3228_ ),
    .A3(\u_multiplier/_3233_ ),
    .ZN(\u_multiplier/_3269_ ));
 OAI211_X1 \u_multiplier/_4045_  (.A(\u_multiplier/_3268_ ),
    .B(\u_multiplier/_3269_ ),
    .C1(\u_multiplier/_3229_ ),
    .C2(\u_multiplier/_3230_ ),
    .ZN(\u_multiplier/_3270_ ));
 AOI211_X1 \u_multiplier/_4046_  (.A(\u_multiplier/_3251_ ),
    .B(\u_multiplier/_3252_ ),
    .C1(\u_multiplier/_3246_ ),
    .C2(\u_multiplier/_3247_ ),
    .ZN(\u_multiplier/_3271_ ));
 NOR2_X1 \u_multiplier/_4047_  (.A1(\u_multiplier/_3249_ ),
    .A2(\u_multiplier/_3271_ ),
    .ZN(\u_multiplier/_3272_ ));
 OR3_X1 \u_multiplier/_4048_  (.A1(\u_multiplier/_3258_ ),
    .A2(\u_multiplier/_3259_ ),
    .A3(\u_multiplier/_3263_ ),
    .ZN(\u_multiplier/_3273_ ));
 AOI21_X1 \u_multiplier/_4049_  (.A(\u_multiplier/_3245_ ),
    .B1(\u_multiplier/_3272_ ),
    .B2(\u_multiplier/_3273_ ),
    .ZN(\u_multiplier/_3274_ ));
 NOR2_X1 \u_multiplier/_4050_  (.A1(\u_multiplier/_3270_ ),
    .A2(\u_multiplier/_3274_ ),
    .ZN(\u_multiplier/_3275_ ));
 XOR2_X2 \u_multiplier/_4051_  (.A(\u_multiplier/kx [26]),
    .B(_0683_[26]),
    .Z(\u_multiplier/_3276_ ));
 XOR2_X2 \u_multiplier/_4052_  (.A(\u_multiplier/ky [26]),
    .B(sram_rdata_reg[26]),
    .Z(\u_multiplier/_3277_ ));
 XNOR2_X2 \u_multiplier/_4053_  (.A(\u_multiplier/ky [26]),
    .B(sram_rdata_reg[26]),
    .ZN(\u_multiplier/_3278_ ));
 OR2_X1 \u_multiplier/_4054_  (.A1(\u_multiplier/_3276_ ),
    .A2(\u_multiplier/_3278_ ),
    .ZN(\u_multiplier/_3279_ ));
 XOR2_X2 \u_multiplier/_4055_  (.A(\u_multiplier/kx [27]),
    .B(\u_multiplier/LODx/z [27]),
    .Z(\u_multiplier/_3280_ ));
 XNOR2_X1 \u_multiplier/_4056_  (.A(\u_multiplier/kx [27]),
    .B(\u_multiplier/LODx/z [27]),
    .ZN(\u_multiplier/_3281_ ));
 XOR2_X2 \u_multiplier/_4057_  (.A(\u_multiplier/ky [27]),
    .B(\u_multiplier/LODy/z [27]),
    .Z(\u_multiplier/_3282_ ));
 NAND2_X1 \u_multiplier/_4058_  (.A1(\u_multiplier/_3281_ ),
    .A2(\u_multiplier/_3282_ ),
    .ZN(\u_multiplier/_3283_ ));
 NOR2_X1 \u_multiplier/_4059_  (.A1(\u_multiplier/_3281_ ),
    .A2(\u_multiplier/_3282_ ),
    .ZN(\u_multiplier/_3284_ ));
 AOI21_X1 \u_multiplier/_4060_  (.A(\u_multiplier/_3284_ ),
    .B1(\u_multiplier/_3278_ ),
    .B2(\u_multiplier/_3276_ ),
    .ZN(\u_multiplier/_3285_ ));
 AND3_X1 \u_multiplier/_4061_  (.A1(\u_multiplier/_3279_ ),
    .A2(\u_multiplier/_3283_ ),
    .A3(\u_multiplier/_3285_ ),
    .ZN(\u_multiplier/_3286_ ));
 XOR2_X2 \u_multiplier/_4062_  (.A(\u_multiplier/kx [25]),
    .B(_0683_[25]),
    .Z(\u_multiplier/_3287_ ));
 XNOR2_X2 \u_multiplier/_4063_  (.A(\u_multiplier/ky [25]),
    .B(sram_rdata_reg[25]),
    .ZN(\u_multiplier/_3288_ ));
 XOR2_X2 \u_multiplier/_4064_  (.A(\u_multiplier/ky [25]),
    .B(sram_rdata_reg[25]),
    .Z(\u_multiplier/_3289_ ));
 OR2_X1 \u_multiplier/_4065_  (.A1(\u_multiplier/_3287_ ),
    .A2(\u_multiplier/_3288_ ),
    .ZN(\u_multiplier/_3290_ ));
 XOR2_X2 \u_multiplier/_4066_  (.A(\u_multiplier/kx [24]),
    .B(data_in_reg[24]),
    .Z(\u_multiplier/_3291_ ));
 XOR2_X2 \u_multiplier/_4067_  (.A(\u_multiplier/ky [24]),
    .B(sram_rdata_reg[24]),
    .Z(\u_multiplier/_3292_ ));
 INV_X1 \u_multiplier/_4068_  (.A(\u_multiplier/_3292_ ),
    .ZN(\u_multiplier/_3293_ ));
 NAND2_X1 \u_multiplier/_4069_  (.A1(\u_multiplier/_3287_ ),
    .A2(\u_multiplier/_3288_ ),
    .ZN(\u_multiplier/_3294_ ));
 XNOR2_X1 \u_multiplier/_4070_  (.A(\u_multiplier/_3291_ ),
    .B(\u_multiplier/_3292_ ),
    .ZN(\u_multiplier/_3295_ ));
 NAND4_X1 \u_multiplier/_4071_  (.A1(\u_multiplier/_3286_ ),
    .A2(\u_multiplier/_3290_ ),
    .A3(\u_multiplier/_3294_ ),
    .A4(\u_multiplier/_3295_ ),
    .ZN(\u_multiplier/_3296_ ));
 AOI21_X1 \u_multiplier/_4072_  (.A(\u_multiplier/_3296_ ),
    .B1(\u_multiplier/_3275_ ),
    .B2(\u_multiplier/_3266_ ),
    .ZN(\u_multiplier/_3297_ ));
 OAI21_X1 \u_multiplier/_4073_  (.A(\u_multiplier/_3290_ ),
    .B1(\u_multiplier/_3291_ ),
    .B2(\u_multiplier/_3293_ ),
    .ZN(\u_multiplier/_3298_ ));
 NAND3_X1 \u_multiplier/_4074_  (.A1(\u_multiplier/_3286_ ),
    .A2(\u_multiplier/_3294_ ),
    .A3(\u_multiplier/_3298_ ),
    .ZN(\u_multiplier/_3299_ ));
 OAI211_X1 \u_multiplier/_4075_  (.A(\u_multiplier/_3283_ ),
    .B(\u_multiplier/_3299_ ),
    .C1(\u_multiplier/_3284_ ),
    .C2(\u_multiplier/_3279_ ),
    .ZN(\u_multiplier/_3300_ ));
 XOR2_X2 \u_multiplier/_4076_  (.A(\u_multiplier/kx [29]),
    .B(_0683_[29]),
    .Z(\u_multiplier/_3301_ ));
 INV_X1 \u_multiplier/_4077_  (.A(\u_multiplier/_3301_ ),
    .ZN(\u_multiplier/_3302_ ));
 XOR2_X2 \u_multiplier/_4078_  (.A(\u_multiplier/ky [29]),
    .B(sram_rdata_reg[29]),
    .Z(\u_multiplier/_3303_ ));
 INV_X1 \u_multiplier/_4079_  (.A(\u_multiplier/_3303_ ),
    .ZN(\u_multiplier/_3304_ ));
 XNOR2_X1 \u_multiplier/_4080_  (.A(\u_multiplier/_3301_ ),
    .B(\u_multiplier/_3303_ ),
    .ZN(\u_multiplier/_3305_ ));
 XOR2_X2 \u_multiplier/_4081_  (.A(\u_multiplier/kx [28]),
    .B(_0683_[28]),
    .Z(\u_multiplier/_3306_ ));
 XOR2_X2 \u_multiplier/_4082_  (.A(\u_multiplier/ky [28]),
    .B(sram_rdata_reg[28]),
    .Z(\u_multiplier/_3307_ ));
 INV_X1 \u_multiplier/_4083_  (.A(\u_multiplier/_3307_ ),
    .ZN(\u_multiplier/_3308_ ));
 XNOR2_X1 \u_multiplier/_4084_  (.A(\u_multiplier/_3306_ ),
    .B(\u_multiplier/_3307_ ),
    .ZN(\u_multiplier/_3309_ ));
 OAI211_X2 \u_multiplier/_4085_  (.A(\u_multiplier/_3305_ ),
    .B(\u_multiplier/_3309_ ),
    .C1(\u_multiplier/_3297_ ),
    .C2(\u_multiplier/_3300_ ),
    .ZN(\u_multiplier/_3310_ ));
 AOI211_X2 \u_multiplier/_4086_  (.A(\u_multiplier/_3306_ ),
    .B(\u_multiplier/_3308_ ),
    .C1(\u_multiplier/_3301_ ),
    .C2(\u_multiplier/_3304_ ),
    .ZN(\u_multiplier/_3311_ ));
 AOI221_X2 \u_multiplier/_4087_  (.A(\u_multiplier/_3311_ ),
    .B1(\u_multiplier/_3303_ ),
    .B2(\u_multiplier/_3302_ ),
    .C1(\u_multiplier/_3130_ ),
    .C2(\u_multiplier/_3131_ ),
    .ZN(\u_multiplier/_3312_ ));
 AOI21_X4 \u_multiplier/_4088_  (.A(\u_multiplier/_3132_ ),
    .B1(\u_multiplier/_3310_ ),
    .B2(\u_multiplier/_3312_ ),
    .ZN(\u_multiplier/_3313_ ));
 MUX2_X1 \u_multiplier/_4089_  (.A(\u_multiplier/_3145_ ),
    .B(\u_multiplier/_3127_ ),
    .S(net17),
    .Z(\u_multiplier/_3314_ ));
 INV_X1 \u_multiplier/_4090_  (.A(\u_multiplier/_3314_ ),
    .ZN(\u_multiplier/_1830_ ));
 MUX2_X2 \u_multiplier/_4091_  (.A(\u_multiplier/_3144_ ),
    .B(\u_multiplier/_3141_ ),
    .S(net17),
    .Z(\u_multiplier/_1841_ ));
 MUX2_X2 \u_multiplier/_4092_  (.A(\u_multiplier/_3151_ ),
    .B(\u_multiplier/_3148_ ),
    .S(net17),
    .Z(\u_multiplier/_1852_ ));
 NAND2_X1 \u_multiplier/_4093_  (.A1(\u_multiplier/_3153_ ),
    .A2(net17),
    .ZN(\u_multiplier/_3315_ ));
 OAI21_X4 \u_multiplier/_4094_  (.A(\u_multiplier/_3315_ ),
    .B1(net17),
    .B2(\u_multiplier/_3155_ ),
    .ZN(\u_multiplier/_1854_ ));
 MUX2_X2 \u_multiplier/_4095_  (.A(\u_multiplier/_3161_ ),
    .B(\u_multiplier/_3158_ ),
    .S(net17),
    .Z(\u_multiplier/_1855_ ));
 MUX2_X2 \u_multiplier/_4096_  (.A(\u_multiplier/_3139_ ),
    .B(\u_multiplier/_3137_ ),
    .S(net17),
    .Z(\u_multiplier/_1856_ ));
 MUX2_X2 \u_multiplier/_4097_  (.A(\u_multiplier/_3135_ ),
    .B(\u_multiplier/_3133_ ),
    .S(net17),
    .Z(\u_multiplier/_1857_ ));
 MUX2_X2 \u_multiplier/_4098_  (.A(\u_multiplier/_3169_ ),
    .B(\u_multiplier/_3167_ ),
    .S(net17),
    .Z(\u_multiplier/_1858_ ));
 MUX2_X2 \u_multiplier/_4099_  (.A(\u_multiplier/_3184_ ),
    .B(\u_multiplier/_3182_ ),
    .S(net17),
    .Z(\u_multiplier/_1859_ ));
 MUX2_X2 \u_multiplier/_4100_  (.A(\u_multiplier/_3188_ ),
    .B(\u_multiplier/_3186_ ),
    .S(net17),
    .Z(\u_multiplier/_1860_ ));
 MUX2_X2 \u_multiplier/_4101_  (.A(\u_multiplier/_3174_ ),
    .B(\u_multiplier/_3172_ ),
    .S(net17),
    .Z(\u_multiplier/_1831_ ));
 MUX2_X2 \u_multiplier/_4102_  (.A(\u_multiplier/_3177_ ),
    .B(\u_multiplier/_3175_ ),
    .S(net17),
    .Z(\u_multiplier/_1832_ ));
 MUX2_X2 \u_multiplier/_4103_  (.A(\u_multiplier/_3216_ ),
    .B(\u_multiplier/_3215_ ),
    .S(net17),
    .Z(\u_multiplier/_1833_ ));
 MUX2_X2 \u_multiplier/_4104_  (.A(\u_multiplier/_3213_ ),
    .B(\u_multiplier/_3211_ ),
    .S(net17),
    .Z(\u_multiplier/_1834_ ));
 MUX2_X2 \u_multiplier/_4105_  (.A(\u_multiplier/_3202_ ),
    .B(\u_multiplier/_3200_ ),
    .S(net17),
    .Z(\u_multiplier/_1835_ ));
 MUX2_X2 \u_multiplier/_4106_  (.A(\u_multiplier/_3206_ ),
    .B(\u_multiplier/_3204_ ),
    .S(net17),
    .Z(\u_multiplier/_1836_ ));
 MUX2_X2 \u_multiplier/_4107_  (.A(\u_multiplier/_3261_ ),
    .B(\u_multiplier/_3262_ ),
    .S(net17),
    .Z(\u_multiplier/_1837_ ));
 MUX2_X2 \u_multiplier/_4108_  (.A(\u_multiplier/_3255_ ),
    .B(\u_multiplier/_3257_ ),
    .S(\u_multiplier/_3313_ ),
    .Z(\u_multiplier/_1838_ ));
 MUX2_X2 \u_multiplier/_4109_  (.A(\u_multiplier/_3252_ ),
    .B(\u_multiplier/_3250_ ),
    .S(\u_multiplier/_3313_ ),
    .Z(\u_multiplier/_1839_ ));
 MUX2_X2 \u_multiplier/_4110_  (.A(\u_multiplier/_3246_ ),
    .B(\u_multiplier/_3248_ ),
    .S(\u_multiplier/_3313_ ),
    .Z(\u_multiplier/_1840_ ));
 MUX2_X2 \u_multiplier/_4111_  (.A(\u_multiplier/_3240_ ),
    .B(\u_multiplier/_3241_ ),
    .S(\u_multiplier/_3313_ ),
    .Z(\u_multiplier/_1842_ ));
 MUX2_X2 \u_multiplier/_4112_  (.A(\u_multiplier/_3236_ ),
    .B(\u_multiplier/_3238_ ),
    .S(\u_multiplier/_3313_ ),
    .Z(\u_multiplier/_1843_ ));
 MUX2_X2 \u_multiplier/_4113_  (.A(\u_multiplier/_3227_ ),
    .B(\u_multiplier/_3226_ ),
    .S(\u_multiplier/_3313_ ),
    .Z(\u_multiplier/_1844_ ));
 MUX2_X2 \u_multiplier/_4114_  (.A(\u_multiplier/_3229_ ),
    .B(\u_multiplier/_3231_ ),
    .S(\u_multiplier/_3313_ ),
    .Z(\u_multiplier/_1845_ ));
 MUX2_X2 \u_multiplier/_4115_  (.A(\u_multiplier/_3291_ ),
    .B(\u_multiplier/_3292_ ),
    .S(\u_multiplier/_3313_ ),
    .Z(\u_multiplier/_1846_ ));
 MUX2_X2 \u_multiplier/_4116_  (.A(\u_multiplier/_3287_ ),
    .B(\u_multiplier/_3289_ ),
    .S(\u_multiplier/_3313_ ),
    .Z(\u_multiplier/_1847_ ));
 MUX2_X2 \u_multiplier/_4117_  (.A(\u_multiplier/_3276_ ),
    .B(\u_multiplier/_3277_ ),
    .S(\u_multiplier/_3313_ ),
    .Z(\u_multiplier/_1848_ ));
 MUX2_X2 \u_multiplier/_4118_  (.A(\u_multiplier/_3280_ ),
    .B(\u_multiplier/_3282_ ),
    .S(\u_multiplier/_3313_ ),
    .Z(\u_multiplier/_1849_ ));
 MUX2_X2 \u_multiplier/_4119_  (.A(\u_multiplier/_3306_ ),
    .B(\u_multiplier/_3307_ ),
    .S(\u_multiplier/_3313_ ),
    .Z(\u_multiplier/_1850_ ));
 MUX2_X2 \u_multiplier/_4120_  (.A(\u_multiplier/_3301_ ),
    .B(\u_multiplier/_3303_ ),
    .S(\u_multiplier/_3313_ ),
    .Z(\u_multiplier/_1851_ ));
 OR2_X2 \u_multiplier/_4121_  (.A1(\u_multiplier/_3129_ ),
    .A2(\u_multiplier/_3131_ ),
    .ZN(\u_multiplier/_1853_ ));
 MUX2_X1 \u_multiplier/_4122_  (.A(\u_multiplier/_3128_ ),
    .B(\u_multiplier/_3146_ ),
    .S(net17),
    .Z(\u_multiplier/_3316_ ));
 MUX2_X1 \u_multiplier/_4123_  (.A(\u_multiplier/_3127_ ),
    .B(\u_multiplier/_3145_ ),
    .S(net17),
    .Z(\u_multiplier/_3317_ ));
 NAND2_X1 \u_multiplier/_4124_  (.A1(\u_multiplier/_3113_ ),
    .A2(\u_multiplier/_3316_ ),
    .ZN(\u_multiplier/_3318_ ));
 NAND3_X2 \u_multiplier/_4125_  (.A1(\u_multiplier/_3113_ ),
    .A2(\u_multiplier/_3114_ ),
    .A3(\u_multiplier/_3316_ ),
    .ZN(\u_multiplier/_3319_ ));
 NOR2_X1 \u_multiplier/_4126_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/_3319_ ),
    .ZN(\u_multiplier/_3320_ ));
 NOR3_X2 \u_multiplier/_4127_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/K [3]),
    .A3(\u_multiplier/_3319_ ),
    .ZN(\u_multiplier/_3321_ ));
 AOI21_X4 \u_multiplier/_4128_  (.A(\u_multiplier/dec_out [0]),
    .B1(\u_multiplier/_3321_ ),
    .B2(\u_multiplier/_3116_ ),
    .ZN(\u_multiplier/_3322_ ));
 NOR2_X1 \u_multiplier/_4129_  (.A1(\u_multiplier/code_x [0]),
    .A2(\u_multiplier/_3127_ ),
    .ZN(\u_multiplier/_3323_ ));
 NOR3_X1 \u_multiplier/_4130_  (.A1(\u_multiplier/code_x [0]),
    .A2(\u_multiplier/code_x [1]),
    .A3(\u_multiplier/_3127_ ),
    .ZN(\u_multiplier/_3324_ ));
 AND2_X1 \u_multiplier/_4131_  (.A1(\u_multiplier/_3110_ ),
    .A2(\u_multiplier/_3324_ ),
    .ZN(\u_multiplier/_3325_ ));
 NAND2_X2 \u_multiplier/_4132_  (.A1(\u_multiplier/_3111_ ),
    .A2(\u_multiplier/_3325_ ),
    .ZN(\u_multiplier/_3326_ ));
 NAND2_X2 \u_multiplier/_4133_  (.A1(\u_multiplier/_3105_ ),
    .A2(\u_multiplier/_3146_ ),
    .ZN(\u_multiplier/_3327_ ));
 NOR3_X4 \u_multiplier/_4134_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/code_y [2]),
    .A3(\u_multiplier/_3327_ ),
    .ZN(\u_multiplier/_3328_ ));
 NAND2_X2 \u_multiplier/_4135_  (.A1(\u_multiplier/_3107_ ),
    .A2(\u_multiplier/_3328_ ),
    .ZN(\u_multiplier/_3329_ ));
 OAI22_X2 \u_multiplier/_4136_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_3326_ ),
    .B1(\u_multiplier/_3329_ ),
    .B2(\u_multiplier/code_y [4]),
    .ZN(\u_multiplier/_3330_ ));
 OR4_X4 \u_multiplier/_4137_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/code_x [4]),
    .A3(\u_multiplier/_3326_ ),
    .A4(\u_multiplier/_3329_ ),
    .ZN(\u_multiplier/_3331_ ));
 NAND2_X4 \u_multiplier/_4138_  (.A1(\u_multiplier/_3330_ ),
    .A2(\u_multiplier/_3331_ ),
    .ZN(\u_multiplier/_3332_ ));
 NOR2_X4 \u_multiplier/_4139_  (.A1(\u_multiplier/zero_y ),
    .A2(\u_multiplier/zero_x ),
    .ZN(\u_multiplier/_3333_ ));
 OR2_X4 \u_multiplier/_4140_  (.A1(\u_multiplier/zero_y ),
    .A2(\u_multiplier/zero_x ),
    .ZN(\u_multiplier/_3334_ ));
 OAI21_X2 \u_multiplier/_4141_  (.A(\u_multiplier/_3333_ ),
    .B1(\u_multiplier/_3332_ ),
    .B2(\u_multiplier/_3322_ ),
    .ZN(\u_multiplier/_3335_ ));
 AOI21_X4 \u_multiplier/_4142_  (.A(\u_multiplier/_3335_ ),
    .B1(\u_multiplier/_3332_ ),
    .B2(\u_multiplier/_3322_ ),
    .ZN(product[0]));
 OAI21_X4 \u_multiplier/_4143_  (.A(\u_multiplier/_3331_ ),
    .B1(\u_multiplier/_3332_ ),
    .B2(\u_multiplier/_3322_ ),
    .ZN(\u_multiplier/_3336_ ));
 MUX2_X1 \u_multiplier/_4144_  (.A(\u_multiplier/_3142_ ),
    .B(\u_multiplier/_3143_ ),
    .S(net17),
    .Z(\u_multiplier/_3337_ ));
 MUX2_X2 \u_multiplier/_4145_  (.A(\u_multiplier/_3317_ ),
    .B(\u_multiplier/_3337_ ),
    .S(\u_multiplier/_3113_ ),
    .Z(\u_multiplier/_3338_ ));
 OR2_X1 \u_multiplier/_4146_  (.A1(\u_multiplier/K [1]),
    .A2(\u_multiplier/_3338_ ),
    .ZN(\u_multiplier/_3339_ ));
 NOR2_X1 \u_multiplier/_4147_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/_3339_ ),
    .ZN(\u_multiplier/_3340_ ));
 NOR4_X4 \u_multiplier/_4148_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/K [1]),
    .A3(\u_multiplier/K [3]),
    .A4(\u_multiplier/_3338_ ),
    .ZN(\u_multiplier/_3341_ ));
 AOI21_X4 \u_multiplier/_4149_  (.A(\u_multiplier/dec_out [1]),
    .B1(\u_multiplier/_3341_ ),
    .B2(\u_multiplier/_3116_ ),
    .ZN(\u_multiplier/_3342_ ));
 MUX2_X1 \u_multiplier/_4150_  (.A(\u_multiplier/_3142_ ),
    .B(\u_multiplier/_3127_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_3343_ ));
 OR2_X1 \u_multiplier/_4151_  (.A1(\u_multiplier/code_x [1]),
    .A2(\u_multiplier/_3343_ ),
    .ZN(\u_multiplier/_3344_ ));
 NOR2_X2 \u_multiplier/_4152_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_3344_ ),
    .ZN(\u_multiplier/_3345_ ));
 NAND2_X1 \u_multiplier/_4153_  (.A1(\u_multiplier/_3111_ ),
    .A2(\u_multiplier/_3345_ ),
    .ZN(\u_multiplier/_3346_ ));
 MUX2_X1 \u_multiplier/_4154_  (.A(\u_multiplier/_3143_ ),
    .B(\u_multiplier/_3145_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_3347_ ));
 OR2_X1 \u_multiplier/_4155_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_3347_ ),
    .ZN(\u_multiplier/_3348_ ));
 OR2_X1 \u_multiplier/_4156_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_3348_ ),
    .ZN(\u_multiplier/_3349_ ));
 OR2_X1 \u_multiplier/_4157_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_3349_ ),
    .ZN(\u_multiplier/_3350_ ));
 OAI22_X1 \u_multiplier/_4158_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_3346_ ),
    .B1(\u_multiplier/_3350_ ),
    .B2(\u_multiplier/code_y [4]),
    .ZN(\u_multiplier/_3351_ ));
 OR4_X1 \u_multiplier/_4159_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/code_x [4]),
    .A3(\u_multiplier/_3346_ ),
    .A4(\u_multiplier/_3350_ ),
    .ZN(\u_multiplier/_3352_ ));
 NAND2_X1 \u_multiplier/_4160_  (.A1(\u_multiplier/_3351_ ),
    .A2(\u_multiplier/_3352_ ),
    .ZN(\u_multiplier/_3353_ ));
 XOR2_X2 \u_multiplier/_4161_  (.A(\u_multiplier/_3342_ ),
    .B(\u_multiplier/_3353_ ),
    .Z(\u_multiplier/_3354_ ));
 NAND2_X2 \u_multiplier/_4162_  (.A1(\u_multiplier/_3336_ ),
    .A2(\u_multiplier/_3354_ ),
    .ZN(\u_multiplier/_3355_ ));
 OAI21_X2 \u_multiplier/_4163_  (.A(net21),
    .B1(\u_multiplier/_3336_ ),
    .B2(\u_multiplier/_3354_ ),
    .ZN(\u_multiplier/_3356_ ));
 AOI21_X4 \u_multiplier/_4164_  (.A(\u_multiplier/_3356_ ),
    .B1(\u_multiplier/_3354_ ),
    .B2(\u_multiplier/_3336_ ),
    .ZN(product[1]));
 OAI21_X2 \u_multiplier/_4165_  (.A(\u_multiplier/_3352_ ),
    .B1(\u_multiplier/_3353_ ),
    .B2(\u_multiplier/_3342_ ),
    .ZN(\u_multiplier/_3357_ ));
 MUX2_X1 \u_multiplier/_4166_  (.A(\u_multiplier/_3149_ ),
    .B(\u_multiplier/_3150_ ),
    .S(net17),
    .Z(\u_multiplier/_3358_ ));
 MUX2_X1 \u_multiplier/_4167_  (.A(\u_multiplier/_3337_ ),
    .B(\u_multiplier/_3358_ ),
    .S(\u_multiplier/_3113_ ),
    .Z(\u_multiplier/_3359_ ));
 MUX2_X2 \u_multiplier/_4168_  (.A(\u_multiplier/_3318_ ),
    .B(\u_multiplier/_3359_ ),
    .S(\u_multiplier/_3114_ ),
    .Z(\u_multiplier/_3360_ ));
 NOR2_X1 \u_multiplier/_4169_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/_3360_ ),
    .ZN(\u_multiplier/_3361_ ));
 NOR4_X2 \u_multiplier/_4170_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/K [3]),
    .A3(\u_multiplier/K [4]),
    .A4(\u_multiplier/_3360_ ),
    .ZN(\u_multiplier/_3362_ ));
 MUX2_X1 \u_multiplier/_4171_  (.A(\u_multiplier/_3148_ ),
    .B(\u_multiplier/_3141_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_3363_ ));
 MUX2_X1 \u_multiplier/_4172_  (.A(\u_multiplier/_3363_ ),
    .B(\u_multiplier/_3323_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_3364_ ));
 NAND2_X1 \u_multiplier/_4173_  (.A1(\u_multiplier/_3110_ ),
    .A2(\u_multiplier/_3364_ ),
    .ZN(\u_multiplier/_3365_ ));
 NAND3_X1 \u_multiplier/_4174_  (.A1(\u_multiplier/_3110_ ),
    .A2(\u_multiplier/_3111_ ),
    .A3(\u_multiplier/_3364_ ),
    .ZN(\u_multiplier/_3366_ ));
 MUX2_X1 \u_multiplier/_4175_  (.A(\u_multiplier/_3144_ ),
    .B(\u_multiplier/_3151_ ),
    .S(\u_multiplier/_3105_ ),
    .Z(\u_multiplier/_3367_ ));
 NOR2_X1 \u_multiplier/_4176_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_3367_ ),
    .ZN(\u_multiplier/_3368_ ));
 AOI21_X2 \u_multiplier/_4177_  (.A(\u_multiplier/_3368_ ),
    .B1(\u_multiplier/_3327_ ),
    .B2(\u_multiplier/code_y [1]),
    .ZN(\u_multiplier/_3369_ ));
 NAND2_X1 \u_multiplier/_4178_  (.A1(\u_multiplier/_3106_ ),
    .A2(\u_multiplier/_3369_ ),
    .ZN(\u_multiplier/_3370_ ));
 NAND3_X1 \u_multiplier/_4179_  (.A1(\u_multiplier/_3106_ ),
    .A2(\u_multiplier/_3107_ ),
    .A3(\u_multiplier/_3369_ ),
    .ZN(\u_multiplier/_3371_ ));
 OAI22_X1 \u_multiplier/_4180_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_3366_ ),
    .B1(\u_multiplier/_3371_ ),
    .B2(\u_multiplier/code_y [4]),
    .ZN(\u_multiplier/_3372_ ));
 OR4_X1 \u_multiplier/_4181_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/code_x [4]),
    .A3(\u_multiplier/_3366_ ),
    .A4(\u_multiplier/_3371_ ),
    .ZN(\u_multiplier/_3373_ ));
 NAND2_X1 \u_multiplier/_4182_  (.A1(\u_multiplier/_3372_ ),
    .A2(\u_multiplier/_3373_ ),
    .ZN(\u_multiplier/_3374_ ));
 INV_X1 \u_multiplier/_4183_  (.A(\u_multiplier/_3374_ ),
    .ZN(\u_multiplier/_3375_ ));
 OAI21_X2 \u_multiplier/_4184_  (.A(\u_multiplier/_3375_ ),
    .B1(\u_multiplier/_3362_ ),
    .B2(\u_multiplier/dec_out [2]),
    .ZN(\u_multiplier/_3376_ ));
 OR3_X2 \u_multiplier/_4185_  (.A1(\u_multiplier/dec_out [2]),
    .A2(\u_multiplier/_3362_ ),
    .A3(\u_multiplier/_3375_ ),
    .ZN(\u_multiplier/_3377_ ));
 AND3_X1 \u_multiplier/_4186_  (.A1(\u_multiplier/_3357_ ),
    .A2(\u_multiplier/_3376_ ),
    .A3(\u_multiplier/_3377_ ),
    .ZN(\u_multiplier/_3378_ ));
 NAND3_X1 \u_multiplier/_4187_  (.A1(\u_multiplier/_3357_ ),
    .A2(\u_multiplier/_3376_ ),
    .A3(\u_multiplier/_3377_ ),
    .ZN(\u_multiplier/_3379_ ));
 AOI21_X2 \u_multiplier/_4188_  (.A(\u_multiplier/_3357_ ),
    .B1(\u_multiplier/_3376_ ),
    .B2(\u_multiplier/_3377_ ),
    .ZN(\u_multiplier/_3380_ ));
 NOR3_X2 \u_multiplier/_4189_  (.A1(\u_multiplier/_3355_ ),
    .A2(\u_multiplier/_3378_ ),
    .A3(\u_multiplier/_3380_ ),
    .ZN(\u_multiplier/_3381_ ));
 OAI21_X1 \u_multiplier/_4190_  (.A(\u_multiplier/_3355_ ),
    .B1(\u_multiplier/_3378_ ),
    .B2(\u_multiplier/_3380_ ),
    .ZN(\u_multiplier/_3382_ ));
 INV_X1 \u_multiplier/_4191_  (.A(\u_multiplier/_3382_ ),
    .ZN(\u_multiplier/_3383_ ));
 NOR3_X2 \u_multiplier/_4192_  (.A1(\u_multiplier/_3334_ ),
    .A2(\u_multiplier/_3381_ ),
    .A3(\u_multiplier/_3383_ ),
    .ZN(product[2]));
 NOR2_X1 \u_multiplier/_4193_  (.A1(\u_multiplier/_3378_ ),
    .A2(\u_multiplier/_3381_ ),
    .ZN(\u_multiplier/_3384_ ));
 OAI21_X2 \u_multiplier/_4194_  (.A(\u_multiplier/_3379_ ),
    .B1(\u_multiplier/_3380_ ),
    .B2(\u_multiplier/_3355_ ),
    .ZN(\u_multiplier/_3385_ ));
 NAND2_X1 \u_multiplier/_4195_  (.A1(\u_multiplier/_3373_ ),
    .A2(\u_multiplier/_3376_ ),
    .ZN(\u_multiplier/_3386_ ));
 MUX2_X1 \u_multiplier/_4196_  (.A(\u_multiplier/_3154_ ),
    .B(\u_multiplier/_3155_ ),
    .S(net17),
    .Z(\u_multiplier/_3387_ ));
 MUX2_X1 \u_multiplier/_4197_  (.A(\u_multiplier/_3358_ ),
    .B(\u_multiplier/_3387_ ),
    .S(\u_multiplier/_3113_ ),
    .Z(\u_multiplier/_3388_ ));
 MUX2_X2 \u_multiplier/_4198_  (.A(\u_multiplier/_3338_ ),
    .B(\u_multiplier/_3388_ ),
    .S(\u_multiplier/_3114_ ),
    .Z(\u_multiplier/_3389_ ));
 NOR2_X1 \u_multiplier/_4199_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/_3389_ ),
    .ZN(\u_multiplier/_3390_ ));
 NOR3_X4 \u_multiplier/_4200_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/K [3]),
    .A3(\u_multiplier/_3389_ ),
    .ZN(\u_multiplier/_3391_ ));
 AOI21_X4 \u_multiplier/_4201_  (.A(\u_multiplier/dec_out [3]),
    .B1(\u_multiplier/_3391_ ),
    .B2(\u_multiplier/_3116_ ),
    .ZN(\u_multiplier/_3392_ ));
 MUX2_X1 \u_multiplier/_4202_  (.A(\u_multiplier/_3154_ ),
    .B(\u_multiplier/_3149_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_3393_ ));
 MUX2_X1 \u_multiplier/_4203_  (.A(\u_multiplier/_3393_ ),
    .B(\u_multiplier/_3343_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_3394_ ));
 OR2_X1 \u_multiplier/_4204_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_3394_ ),
    .ZN(\u_multiplier/_3395_ ));
 OR2_X1 \u_multiplier/_4205_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_3395_ ),
    .ZN(\u_multiplier/_3396_ ));
 MUX2_X1 \u_multiplier/_4206_  (.A(\u_multiplier/_3150_ ),
    .B(\u_multiplier/_3155_ ),
    .S(\u_multiplier/_3105_ ),
    .Z(\u_multiplier/_3397_ ));
 MUX2_X1 \u_multiplier/_4207_  (.A(\u_multiplier/_3397_ ),
    .B(\u_multiplier/_3347_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_3398_ ));
 OR2_X1 \u_multiplier/_4208_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_3398_ ),
    .ZN(\u_multiplier/_3399_ ));
 OR2_X1 \u_multiplier/_4209_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_3399_ ),
    .ZN(\u_multiplier/_3400_ ));
 OAI22_X1 \u_multiplier/_4210_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_3396_ ),
    .B1(\u_multiplier/_3400_ ),
    .B2(\u_multiplier/code_y [4]),
    .ZN(\u_multiplier/_3401_ ));
 OR4_X1 \u_multiplier/_4211_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/code_x [4]),
    .A3(\u_multiplier/_3396_ ),
    .A4(\u_multiplier/_3400_ ),
    .ZN(\u_multiplier/_3402_ ));
 NAND2_X1 \u_multiplier/_4212_  (.A1(\u_multiplier/_3401_ ),
    .A2(\u_multiplier/_3402_ ),
    .ZN(\u_multiplier/_3403_ ));
 XOR2_X2 \u_multiplier/_4213_  (.A(\u_multiplier/_3392_ ),
    .B(\u_multiplier/_3403_ ),
    .Z(\u_multiplier/_3404_ ));
 AND2_X1 \u_multiplier/_4214_  (.A1(\u_multiplier/_3386_ ),
    .A2(\u_multiplier/_3404_ ),
    .ZN(\u_multiplier/_3405_ ));
 OR2_X1 \u_multiplier/_4215_  (.A1(\u_multiplier/_3386_ ),
    .A2(\u_multiplier/_3404_ ),
    .ZN(\u_multiplier/_3406_ ));
 XNOR2_X2 \u_multiplier/_4216_  (.A(\u_multiplier/_3386_ ),
    .B(\u_multiplier/_3404_ ),
    .ZN(\u_multiplier/_3407_ ));
 AOI21_X1 \u_multiplier/_4217_  (.A(\u_multiplier/_3334_ ),
    .B1(\u_multiplier/_3384_ ),
    .B2(\u_multiplier/_3407_ ),
    .ZN(\u_multiplier/_3408_ ));
 OAI21_X2 \u_multiplier/_4218_  (.A(\u_multiplier/_3408_ ),
    .B1(\u_multiplier/_3407_ ),
    .B2(\u_multiplier/_3384_ ),
    .ZN(\u_multiplier/_3409_ ));
 INV_X1 \u_multiplier/_4219_  (.A(\u_multiplier/_3409_ ),
    .ZN(product[3]));
 AOI21_X4 \u_multiplier/_4220_  (.A(\u_multiplier/_3405_ ),
    .B1(\u_multiplier/_3406_ ),
    .B2(\u_multiplier/_3385_ ),
    .ZN(\u_multiplier/_3410_ ));
 OAI21_X2 \u_multiplier/_4221_  (.A(\u_multiplier/_3402_ ),
    .B1(\u_multiplier/_3403_ ),
    .B2(\u_multiplier/_3392_ ),
    .ZN(\u_multiplier/_3411_ ));
 MUX2_X1 \u_multiplier/_4222_  (.A(\u_multiplier/_3159_ ),
    .B(\u_multiplier/_3160_ ),
    .S(net17),
    .Z(\u_multiplier/_3412_ ));
 MUX2_X1 \u_multiplier/_4223_  (.A(\u_multiplier/_3387_ ),
    .B(\u_multiplier/_3412_ ),
    .S(\u_multiplier/_3113_ ),
    .Z(\u_multiplier/_3413_ ));
 MUX2_X1 \u_multiplier/_4224_  (.A(\u_multiplier/_3359_ ),
    .B(\u_multiplier/_3413_ ),
    .S(\u_multiplier/_3114_ ),
    .Z(\u_multiplier/_3414_ ));
 MUX2_X1 \u_multiplier/_4225_  (.A(\u_multiplier/_3319_ ),
    .B(\u_multiplier/_3414_ ),
    .S(\u_multiplier/_3112_ ),
    .Z(\u_multiplier/_3415_ ));
 NOR2_X2 \u_multiplier/_4226_  (.A1(\u_multiplier/K [3]),
    .A2(\u_multiplier/_3415_ ),
    .ZN(\u_multiplier/_3416_ ));
 AOI21_X4 \u_multiplier/_4227_  (.A(\u_multiplier/dec_out [4]),
    .B1(\u_multiplier/_3416_ ),
    .B2(\u_multiplier/_3116_ ),
    .ZN(\u_multiplier/_3417_ ));
 MUX2_X1 \u_multiplier/_4228_  (.A(\u_multiplier/_3158_ ),
    .B(\u_multiplier/_3153_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_3418_ ));
 INV_X1 \u_multiplier/_4229_  (.A(\u_multiplier/_3418_ ),
    .ZN(\u_multiplier/_3419_ ));
 MUX2_X1 \u_multiplier/_4230_  (.A(\u_multiplier/_3418_ ),
    .B(\u_multiplier/_3363_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_3420_ ));
 MUX2_X1 \u_multiplier/_4231_  (.A(\u_multiplier/_3324_ ),
    .B(\u_multiplier/_3420_ ),
    .S(\u_multiplier/_3110_ ),
    .Z(\u_multiplier/_3421_ ));
 NAND2_X1 \u_multiplier/_4232_  (.A1(\u_multiplier/_3111_ ),
    .A2(\u_multiplier/_3421_ ),
    .ZN(\u_multiplier/_3422_ ));
 NOR2_X1 \u_multiplier/_4233_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_3422_ ),
    .ZN(\u_multiplier/_3423_ ));
 MUX2_X1 \u_multiplier/_4234_  (.A(\u_multiplier/_3155_ ),
    .B(\u_multiplier/_3160_ ),
    .S(\u_multiplier/_3105_ ),
    .Z(\u_multiplier/_3424_ ));
 NAND2_X1 \u_multiplier/_4235_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_3367_ ),
    .ZN(\u_multiplier/_3425_ ));
 OAI21_X1 \u_multiplier/_4236_  (.A(\u_multiplier/code_y [2]),
    .B1(\u_multiplier/_3327_ ),
    .B2(\u_multiplier/code_y [1]),
    .ZN(\u_multiplier/_3426_ ));
 OAI211_X1 \u_multiplier/_4237_  (.A(\u_multiplier/_3106_ ),
    .B(\u_multiplier/_3425_ ),
    .C1(\u_multiplier/_3424_ ),
    .C2(\u_multiplier/code_y [1]),
    .ZN(\u_multiplier/_3427_ ));
 AND2_X1 \u_multiplier/_4238_  (.A1(\u_multiplier/_3426_ ),
    .A2(\u_multiplier/_3427_ ),
    .ZN(\u_multiplier/_3428_ ));
 NAND2_X1 \u_multiplier/_4239_  (.A1(\u_multiplier/_3107_ ),
    .A2(\u_multiplier/_3428_ ),
    .ZN(\u_multiplier/_3429_ ));
 NOR2_X1 \u_multiplier/_4240_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_3429_ ),
    .ZN(\u_multiplier/_3430_ ));
 AND2_X1 \u_multiplier/_4241_  (.A1(\u_multiplier/_3423_ ),
    .A2(\u_multiplier/_3430_ ),
    .ZN(\u_multiplier/_3431_ ));
 XNOR2_X2 \u_multiplier/_4242_  (.A(\u_multiplier/_3423_ ),
    .B(\u_multiplier/_3430_ ),
    .ZN(\u_multiplier/_3432_ ));
 NOR2_X1 \u_multiplier/_4243_  (.A1(\u_multiplier/_3417_ ),
    .A2(\u_multiplier/_3432_ ),
    .ZN(\u_multiplier/_3433_ ));
 XOR2_X2 \u_multiplier/_4244_  (.A(\u_multiplier/_3417_ ),
    .B(\u_multiplier/_3432_ ),
    .Z(\u_multiplier/_3434_ ));
 NAND2_X1 \u_multiplier/_4245_  (.A1(\u_multiplier/_3411_ ),
    .A2(\u_multiplier/_3434_ ),
    .ZN(\u_multiplier/_3435_ ));
 XNOR2_X2 \u_multiplier/_4246_  (.A(\u_multiplier/_3411_ ),
    .B(\u_multiplier/_3434_ ),
    .ZN(\u_multiplier/_3436_ ));
 AOI21_X1 \u_multiplier/_4247_  (.A(\u_multiplier/_3334_ ),
    .B1(\u_multiplier/_3410_ ),
    .B2(\u_multiplier/_3436_ ),
    .ZN(\u_multiplier/_3437_ ));
 OAI21_X2 \u_multiplier/_4248_  (.A(\u_multiplier/_3437_ ),
    .B1(\u_multiplier/_3436_ ),
    .B2(\u_multiplier/_3410_ ),
    .ZN(\u_multiplier/_3438_ ));
 INV_X1 \u_multiplier/_4249_  (.A(\u_multiplier/_3438_ ),
    .ZN(product[4]));
 OAI21_X4 \u_multiplier/_4250_  (.A(\u_multiplier/_3435_ ),
    .B1(\u_multiplier/_3436_ ),
    .B2(\u_multiplier/_3410_ ),
    .ZN(\u_multiplier/_3439_ ));
 OR2_X1 \u_multiplier/_4251_  (.A1(\u_multiplier/_3431_ ),
    .A2(\u_multiplier/_3433_ ),
    .ZN(\u_multiplier/_3440_ ));
 MUX2_X1 \u_multiplier/_4252_  (.A(\u_multiplier/_3137_ ),
    .B(\u_multiplier/_3139_ ),
    .S(net17),
    .Z(\u_multiplier/_3441_ ));
 NAND2_X1 \u_multiplier/_4253_  (.A1(\u_multiplier/_3113_ ),
    .A2(\u_multiplier/_3441_ ),
    .ZN(\u_multiplier/_3442_ ));
 OAI21_X1 \u_multiplier/_4254_  (.A(\u_multiplier/_3442_ ),
    .B1(\u_multiplier/_3412_ ),
    .B2(\u_multiplier/_3113_ ),
    .ZN(\u_multiplier/_3443_ ));
 NOR2_X1 \u_multiplier/_4255_  (.A1(\u_multiplier/_3114_ ),
    .A2(\u_multiplier/_3388_ ),
    .ZN(\u_multiplier/_3444_ ));
 AOI21_X1 \u_multiplier/_4256_  (.A(\u_multiplier/_3444_ ),
    .B1(\u_multiplier/_3443_ ),
    .B2(\u_multiplier/_3114_ ),
    .ZN(\u_multiplier/_3445_ ));
 MUX2_X1 \u_multiplier/_4257_  (.A(\u_multiplier/_3339_ ),
    .B(\u_multiplier/_3445_ ),
    .S(\u_multiplier/_3112_ ),
    .Z(\u_multiplier/_3446_ ));
 NOR2_X2 \u_multiplier/_4258_  (.A1(\u_multiplier/K [3]),
    .A2(\u_multiplier/_3446_ ),
    .ZN(\u_multiplier/_3447_ ));
 AOI21_X2 \u_multiplier/_4259_  (.A(\u_multiplier/dec_out [5]),
    .B1(\u_multiplier/_3447_ ),
    .B2(\u_multiplier/_3116_ ),
    .ZN(\u_multiplier/_3448_ ));
 MUX2_X1 \u_multiplier/_4260_  (.A(\u_multiplier/_3137_ ),
    .B(\u_multiplier/_3158_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_3449_ ));
 NOR2_X1 \u_multiplier/_4261_  (.A1(\u_multiplier/code_x [1]),
    .A2(\u_multiplier/_3449_ ),
    .ZN(\u_multiplier/_3450_ ));
 AOI21_X1 \u_multiplier/_4262_  (.A(\u_multiplier/_3450_ ),
    .B1(\u_multiplier/_3393_ ),
    .B2(\u_multiplier/code_x [1]),
    .ZN(\u_multiplier/_3451_ ));
 NOR2_X1 \u_multiplier/_4263_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_3451_ ),
    .ZN(\u_multiplier/_3452_ ));
 AOI21_X2 \u_multiplier/_4264_  (.A(\u_multiplier/_3452_ ),
    .B1(\u_multiplier/_3344_ ),
    .B2(\u_multiplier/code_x [2]),
    .ZN(\u_multiplier/_3453_ ));
 NAND2_X1 \u_multiplier/_4265_  (.A1(\u_multiplier/_3111_ ),
    .A2(\u_multiplier/_3453_ ),
    .ZN(\u_multiplier/_3454_ ));
 NOR2_X1 \u_multiplier/_4266_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_3454_ ),
    .ZN(\u_multiplier/_3455_ ));
 MUX2_X1 \u_multiplier/_4267_  (.A(\u_multiplier/_3139_ ),
    .B(\u_multiplier/_3161_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_3456_ ));
 INV_X1 \u_multiplier/_4268_  (.A(\u_multiplier/_3456_ ),
    .ZN(\u_multiplier/_3457_ ));
 NOR2_X1 \u_multiplier/_4269_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_3456_ ),
    .ZN(\u_multiplier/_3458_ ));
 AOI21_X1 \u_multiplier/_4270_  (.A(\u_multiplier/_3458_ ),
    .B1(\u_multiplier/_3397_ ),
    .B2(\u_multiplier/code_y [1]),
    .ZN(\u_multiplier/_3459_ ));
 NAND2_X1 \u_multiplier/_4271_  (.A1(\u_multiplier/_3106_ ),
    .A2(\u_multiplier/_3459_ ),
    .ZN(\u_multiplier/_3460_ ));
 OAI21_X2 \u_multiplier/_4272_  (.A(\u_multiplier/_3460_ ),
    .B1(\u_multiplier/_3348_ ),
    .B2(\u_multiplier/_3106_ ),
    .ZN(\u_multiplier/_3461_ ));
 NAND2_X1 \u_multiplier/_4273_  (.A1(\u_multiplier/_3107_ ),
    .A2(\u_multiplier/_3461_ ),
    .ZN(\u_multiplier/_3462_ ));
 NOR2_X1 \u_multiplier/_4274_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_3462_ ),
    .ZN(\u_multiplier/_3463_ ));
 AND2_X1 \u_multiplier/_4275_  (.A1(\u_multiplier/_3455_ ),
    .A2(\u_multiplier/_3463_ ),
    .ZN(\u_multiplier/_3464_ ));
 XNOR2_X2 \u_multiplier/_4276_  (.A(\u_multiplier/_3455_ ),
    .B(\u_multiplier/_3463_ ),
    .ZN(\u_multiplier/_3465_ ));
 NOR2_X1 \u_multiplier/_4277_  (.A1(\u_multiplier/_3448_ ),
    .A2(\u_multiplier/_3465_ ),
    .ZN(\u_multiplier/_3466_ ));
 XOR2_X2 \u_multiplier/_4278_  (.A(\u_multiplier/_3448_ ),
    .B(\u_multiplier/_3465_ ),
    .Z(\u_multiplier/_3467_ ));
 AND2_X1 \u_multiplier/_4279_  (.A1(\u_multiplier/_3440_ ),
    .A2(\u_multiplier/_3467_ ),
    .ZN(\u_multiplier/_3468_ ));
 XOR2_X2 \u_multiplier/_4280_  (.A(\u_multiplier/_3440_ ),
    .B(\u_multiplier/_3467_ ),
    .Z(\u_multiplier/_3469_ ));
 OAI21_X1 \u_multiplier/_4281_  (.A(net21),
    .B1(\u_multiplier/_3439_ ),
    .B2(\u_multiplier/_3469_ ),
    .ZN(\u_multiplier/_3470_ ));
 AOI21_X2 \u_multiplier/_4282_  (.A(\u_multiplier/_3470_ ),
    .B1(\u_multiplier/_3469_ ),
    .B2(\u_multiplier/_3439_ ),
    .ZN(product[5]));
 AOI21_X4 \u_multiplier/_4283_  (.A(\u_multiplier/_3468_ ),
    .B1(\u_multiplier/_3469_ ),
    .B2(\u_multiplier/_3439_ ),
    .ZN(\u_multiplier/_3471_ ));
 NOR2_X1 \u_multiplier/_4284_  (.A1(\u_multiplier/_3464_ ),
    .A2(\u_multiplier/_3466_ ),
    .ZN(\u_multiplier/_3472_ ));
 MUX2_X1 \u_multiplier/_4285_  (.A(\u_multiplier/_3133_ ),
    .B(\u_multiplier/_3135_ ),
    .S(net17),
    .Z(\u_multiplier/_3473_ ));
 MUX2_X1 \u_multiplier/_4286_  (.A(\u_multiplier/_3441_ ),
    .B(\u_multiplier/_3473_ ),
    .S(\u_multiplier/_3113_ ),
    .Z(\u_multiplier/_3474_ ));
 NAND2_X1 \u_multiplier/_4287_  (.A1(\u_multiplier/_3114_ ),
    .A2(\u_multiplier/_3474_ ),
    .ZN(\u_multiplier/_3475_ ));
 OAI21_X1 \u_multiplier/_4288_  (.A(\u_multiplier/_3475_ ),
    .B1(\u_multiplier/_3413_ ),
    .B2(\u_multiplier/_3114_ ),
    .ZN(\u_multiplier/_3476_ ));
 NOR2_X1 \u_multiplier/_4289_  (.A1(\u_multiplier/_3112_ ),
    .A2(\u_multiplier/_3360_ ),
    .ZN(\u_multiplier/_3477_ ));
 AOI21_X2 \u_multiplier/_4290_  (.A(\u_multiplier/_3477_ ),
    .B1(\u_multiplier/_3476_ ),
    .B2(\u_multiplier/_3112_ ),
    .ZN(\u_multiplier/_3478_ ));
 NOR2_X2 \u_multiplier/_4291_  (.A1(\u_multiplier/K [3]),
    .A2(\u_multiplier/_3478_ ),
    .ZN(\u_multiplier/_3479_ ));
 AOI21_X2 \u_multiplier/_4292_  (.A(\u_multiplier/dec_out [6]),
    .B1(\u_multiplier/_3479_ ),
    .B2(\u_multiplier/_3116_ ),
    .ZN(\u_multiplier/_3480_ ));
 MUX2_X1 \u_multiplier/_4293_  (.A(\u_multiplier/_3133_ ),
    .B(\u_multiplier/_3137_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_3481_ ));
 NAND2_X1 \u_multiplier/_4294_  (.A1(\u_multiplier/code_x [1]),
    .A2(\u_multiplier/_3419_ ),
    .ZN(\u_multiplier/_3482_ ));
 OAI21_X1 \u_multiplier/_4295_  (.A(\u_multiplier/_3482_ ),
    .B1(\u_multiplier/_3481_ ),
    .B2(\u_multiplier/code_x [1]),
    .ZN(\u_multiplier/_3483_ ));
 NAND2_X1 \u_multiplier/_4296_  (.A1(\u_multiplier/_3110_ ),
    .A2(\u_multiplier/_3483_ ),
    .ZN(\u_multiplier/_3484_ ));
 OAI21_X1 \u_multiplier/_4297_  (.A(\u_multiplier/_3484_ ),
    .B1(\u_multiplier/_3364_ ),
    .B2(\u_multiplier/_3110_ ),
    .ZN(\u_multiplier/_3485_ ));
 OR2_X1 \u_multiplier/_4298_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_3485_ ),
    .ZN(\u_multiplier/_3486_ ));
 NOR2_X1 \u_multiplier/_4299_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_3486_ ),
    .ZN(\u_multiplier/_3487_ ));
 MUX2_X1 \u_multiplier/_4300_  (.A(\u_multiplier/_3135_ ),
    .B(\u_multiplier/_3139_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_3488_ ));
 NAND2_X1 \u_multiplier/_4301_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_3424_ ),
    .ZN(\u_multiplier/_3489_ ));
 OAI21_X1 \u_multiplier/_4302_  (.A(\u_multiplier/_3489_ ),
    .B1(\u_multiplier/_3488_ ),
    .B2(\u_multiplier/code_y [1]),
    .ZN(\u_multiplier/_3490_ ));
 NAND2_X1 \u_multiplier/_4303_  (.A1(\u_multiplier/_3106_ ),
    .A2(\u_multiplier/_3490_ ),
    .ZN(\u_multiplier/_3491_ ));
 OAI21_X1 \u_multiplier/_4304_  (.A(\u_multiplier/_3491_ ),
    .B1(\u_multiplier/_3369_ ),
    .B2(\u_multiplier/_3106_ ),
    .ZN(\u_multiplier/_3492_ ));
 OR2_X1 \u_multiplier/_4305_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_3492_ ),
    .ZN(\u_multiplier/_3493_ ));
 NOR2_X1 \u_multiplier/_4306_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_3493_ ),
    .ZN(\u_multiplier/_3494_ ));
 AND2_X1 \u_multiplier/_4307_  (.A1(\u_multiplier/_3487_ ),
    .A2(\u_multiplier/_3494_ ),
    .ZN(\u_multiplier/_3495_ ));
 XNOR2_X2 \u_multiplier/_4308_  (.A(\u_multiplier/_3487_ ),
    .B(\u_multiplier/_3494_ ),
    .ZN(\u_multiplier/_3496_ ));
 NOR2_X1 \u_multiplier/_4309_  (.A1(\u_multiplier/_3480_ ),
    .A2(\u_multiplier/_3496_ ),
    .ZN(\u_multiplier/_3497_ ));
 XOR2_X2 \u_multiplier/_4310_  (.A(\u_multiplier/_3480_ ),
    .B(\u_multiplier/_3496_ ),
    .Z(\u_multiplier/_3498_ ));
 OAI21_X2 \u_multiplier/_4311_  (.A(\u_multiplier/_3498_ ),
    .B1(\u_multiplier/_3466_ ),
    .B2(\u_multiplier/_3464_ ),
    .ZN(\u_multiplier/_3499_ ));
 XOR2_X2 \u_multiplier/_4312_  (.A(\u_multiplier/_3472_ ),
    .B(\u_multiplier/_3498_ ),
    .Z(\u_multiplier/_3500_ ));
 AOI21_X2 \u_multiplier/_4313_  (.A(\u_multiplier/_3334_ ),
    .B1(\u_multiplier/_3471_ ),
    .B2(\u_multiplier/_3500_ ),
    .ZN(\u_multiplier/_3501_ ));
 OAI21_X4 \u_multiplier/_4314_  (.A(\u_multiplier/_3501_ ),
    .B1(\u_multiplier/_3500_ ),
    .B2(\u_multiplier/_3471_ ),
    .ZN(\u_multiplier/_3502_ ));
 INV_X1 \u_multiplier/_4315_  (.A(\u_multiplier/_3502_ ),
    .ZN(product[6]));
 OAI21_X4 \u_multiplier/_4316_  (.A(\u_multiplier/_3499_ ),
    .B1(\u_multiplier/_3500_ ),
    .B2(\u_multiplier/_3471_ ),
    .ZN(\u_multiplier/_3503_ ));
 MUX2_X1 \u_multiplier/_4317_  (.A(\u_multiplier/_3167_ ),
    .B(\u_multiplier/_3169_ ),
    .S(net17),
    .Z(\u_multiplier/_3504_ ));
 AND2_X1 \u_multiplier/_4318_  (.A1(\u_multiplier/_3113_ ),
    .A2(\u_multiplier/_3504_ ),
    .ZN(\u_multiplier/_3505_ ));
 AOI21_X1 \u_multiplier/_4319_  (.A(\u_multiplier/_3505_ ),
    .B1(\u_multiplier/_3473_ ),
    .B2(\u_multiplier/K [0]),
    .ZN(\u_multiplier/_3506_ ));
 NOR2_X1 \u_multiplier/_4320_  (.A1(\u_multiplier/K [1]),
    .A2(\u_multiplier/_3506_ ),
    .ZN(\u_multiplier/_3507_ ));
 AOI21_X1 \u_multiplier/_4321_  (.A(\u_multiplier/_3507_ ),
    .B1(\u_multiplier/_3443_ ),
    .B2(\u_multiplier/K [1]),
    .ZN(\u_multiplier/_3508_ ));
 MUX2_X2 \u_multiplier/_4322_  (.A(\u_multiplier/_3389_ ),
    .B(\u_multiplier/_3508_ ),
    .S(\u_multiplier/_3112_ ),
    .Z(\u_multiplier/_3509_ ));
 NOR2_X4 \u_multiplier/_4323_  (.A1(\u_multiplier/K [3]),
    .A2(\u_multiplier/_3509_ ),
    .ZN(\u_multiplier/_3510_ ));
 AOI21_X4 \u_multiplier/_4324_  (.A(\u_multiplier/dec_out [7]),
    .B1(\u_multiplier/_3510_ ),
    .B2(\u_multiplier/_3116_ ),
    .ZN(\u_multiplier/_3511_ ));
 MUX2_X1 \u_multiplier/_4325_  (.A(\u_multiplier/_3167_ ),
    .B(\u_multiplier/_3133_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_3512_ ));
 MUX2_X1 \u_multiplier/_4326_  (.A(\u_multiplier/_3512_ ),
    .B(\u_multiplier/_3449_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_3513_ ));
 NAND2_X1 \u_multiplier/_4327_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_3394_ ),
    .ZN(\u_multiplier/_3514_ ));
 OAI21_X2 \u_multiplier/_4328_  (.A(\u_multiplier/_3514_ ),
    .B1(\u_multiplier/_3513_ ),
    .B2(\u_multiplier/code_x [2]),
    .ZN(\u_multiplier/_3515_ ));
 OR2_X1 \u_multiplier/_4329_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_3515_ ),
    .ZN(\u_multiplier/_3516_ ));
 MUX2_X1 \u_multiplier/_4330_  (.A(\u_multiplier/_3135_ ),
    .B(\u_multiplier/_3169_ ),
    .S(\u_multiplier/_3105_ ),
    .Z(\u_multiplier/_3517_ ));
 NAND2_X1 \u_multiplier/_4331_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_3457_ ),
    .ZN(\u_multiplier/_3518_ ));
 OAI21_X1 \u_multiplier/_4332_  (.A(\u_multiplier/_3518_ ),
    .B1(\u_multiplier/_3517_ ),
    .B2(\u_multiplier/code_y [1]),
    .ZN(\u_multiplier/_3519_ ));
 MUX2_X1 \u_multiplier/_4333_  (.A(\u_multiplier/_3398_ ),
    .B(\u_multiplier/_3519_ ),
    .S(\u_multiplier/_3106_ ),
    .Z(\u_multiplier/_3520_ ));
 OR2_X2 \u_multiplier/_4334_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_3520_ ),
    .ZN(\u_multiplier/_3521_ ));
 OAI22_X1 \u_multiplier/_4335_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_3516_ ),
    .B1(\u_multiplier/_3521_ ),
    .B2(\u_multiplier/code_y [4]),
    .ZN(\u_multiplier/_3522_ ));
 OR4_X1 \u_multiplier/_4336_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/code_x [4]),
    .A3(\u_multiplier/_3516_ ),
    .A4(\u_multiplier/_3521_ ),
    .ZN(\u_multiplier/_3523_ ));
 NAND2_X1 \u_multiplier/_4337_  (.A1(\u_multiplier/_3522_ ),
    .A2(\u_multiplier/_3523_ ),
    .ZN(\u_multiplier/_3524_ ));
 XOR2_X2 \u_multiplier/_4338_  (.A(\u_multiplier/_3511_ ),
    .B(\u_multiplier/_3524_ ),
    .Z(\u_multiplier/_3525_ ));
 OAI21_X2 \u_multiplier/_4339_  (.A(\u_multiplier/_3525_ ),
    .B1(\u_multiplier/_3497_ ),
    .B2(\u_multiplier/_3495_ ),
    .ZN(\u_multiplier/_3526_ ));
 OR3_X1 \u_multiplier/_4340_  (.A1(\u_multiplier/_3495_ ),
    .A2(\u_multiplier/_3497_ ),
    .A3(\u_multiplier/_3525_ ),
    .ZN(\u_multiplier/_3527_ ));
 AND2_X2 \u_multiplier/_4341_  (.A1(\u_multiplier/_3526_ ),
    .A2(\u_multiplier/_3527_ ),
    .ZN(\u_multiplier/_3528_ ));
 NAND2_X2 \u_multiplier/_4342_  (.A1(\u_multiplier/_3503_ ),
    .A2(\u_multiplier/_3528_ ),
    .ZN(\u_multiplier/_3529_ ));
 OAI21_X2 \u_multiplier/_4343_  (.A(net21),
    .B1(\u_multiplier/_3503_ ),
    .B2(\u_multiplier/_3528_ ),
    .ZN(\u_multiplier/_3530_ ));
 AOI21_X4 \u_multiplier/_4344_  (.A(\u_multiplier/_3530_ ),
    .B1(\u_multiplier/_3528_ ),
    .B2(\u_multiplier/_3503_ ),
    .ZN(product[7]));
 NAND2_X2 \u_multiplier/_4345_  (.A1(\u_multiplier/_3526_ ),
    .A2(\u_multiplier/_3529_ ),
    .ZN(\u_multiplier/_3531_ ));
 OAI21_X2 \u_multiplier/_4346_  (.A(\u_multiplier/_3523_ ),
    .B1(\u_multiplier/_3524_ ),
    .B2(\u_multiplier/_3511_ ),
    .ZN(\u_multiplier/_3532_ ));
 MUX2_X1 \u_multiplier/_4347_  (.A(\u_multiplier/_3182_ ),
    .B(\u_multiplier/_3184_ ),
    .S(net17),
    .Z(\u_multiplier/_3533_ ));
 MUX2_X1 \u_multiplier/_4348_  (.A(\u_multiplier/_3504_ ),
    .B(\u_multiplier/_3533_ ),
    .S(\u_multiplier/_3113_ ),
    .Z(\u_multiplier/_3534_ ));
 MUX2_X1 \u_multiplier/_4349_  (.A(\u_multiplier/_3474_ ),
    .B(\u_multiplier/_3534_ ),
    .S(\u_multiplier/_3114_ ),
    .Z(\u_multiplier/_3535_ ));
 NAND2_X1 \u_multiplier/_4350_  (.A1(\u_multiplier/_3112_ ),
    .A2(\u_multiplier/_3535_ ),
    .ZN(\u_multiplier/_3536_ ));
 OAI21_X1 \u_multiplier/_4351_  (.A(\u_multiplier/_3536_ ),
    .B1(\u_multiplier/_3414_ ),
    .B2(\u_multiplier/_3112_ ),
    .ZN(\u_multiplier/_3537_ ));
 MUX2_X2 \u_multiplier/_4352_  (.A(\u_multiplier/_3320_ ),
    .B(\u_multiplier/_3537_ ),
    .S(\u_multiplier/_3115_ ),
    .Z(\u_multiplier/_3538_ ));
 AOI21_X4 \u_multiplier/_4353_  (.A(\u_multiplier/dec_out [8]),
    .B1(\u_multiplier/_3538_ ),
    .B2(\u_multiplier/_3116_ ),
    .ZN(\u_multiplier/_3539_ ));
 MUX2_X1 \u_multiplier/_4354_  (.A(\u_multiplier/_3182_ ),
    .B(\u_multiplier/_3167_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_3540_ ));
 MUX2_X1 \u_multiplier/_4355_  (.A(\u_multiplier/_3540_ ),
    .B(\u_multiplier/_3481_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_3541_ ));
 OR2_X1 \u_multiplier/_4356_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_3541_ ),
    .ZN(\u_multiplier/_3542_ ));
 OAI21_X1 \u_multiplier/_4357_  (.A(\u_multiplier/_3542_ ),
    .B1(\u_multiplier/_3420_ ),
    .B2(\u_multiplier/_3110_ ),
    .ZN(\u_multiplier/_3543_ ));
 NAND2_X1 \u_multiplier/_4358_  (.A1(\u_multiplier/_3111_ ),
    .A2(\u_multiplier/_3543_ ),
    .ZN(\u_multiplier/_3544_ ));
 OAI21_X2 \u_multiplier/_4359_  (.A(\u_multiplier/_3544_ ),
    .B1(\u_multiplier/_3325_ ),
    .B2(\u_multiplier/_3111_ ),
    .ZN(\u_multiplier/_3545_ ));
 NOR2_X2 \u_multiplier/_4360_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_3545_ ),
    .ZN(\u_multiplier/_3546_ ));
 MUX2_X1 \u_multiplier/_4361_  (.A(\u_multiplier/_3169_ ),
    .B(\u_multiplier/_3184_ ),
    .S(\u_multiplier/_3105_ ),
    .Z(\u_multiplier/_3547_ ));
 MUX2_X1 \u_multiplier/_4362_  (.A(\u_multiplier/_3547_ ),
    .B(\u_multiplier/_3488_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_3548_ ));
 OAI211_X1 \u_multiplier/_4363_  (.A(\u_multiplier/code_y [2]),
    .B(\u_multiplier/_3425_ ),
    .C1(\u_multiplier/_3424_ ),
    .C2(\u_multiplier/code_y [1]),
    .ZN(\u_multiplier/_3549_ ));
 OAI21_X1 \u_multiplier/_4364_  (.A(\u_multiplier/_3549_ ),
    .B1(\u_multiplier/_3548_ ),
    .B2(\u_multiplier/code_y [2]),
    .ZN(\u_multiplier/_3550_ ));
 NOR2_X1 \u_multiplier/_4365_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_3550_ ),
    .ZN(\u_multiplier/_3551_ ));
 AOI21_X4 \u_multiplier/_4366_  (.A(\u_multiplier/_3551_ ),
    .B1(\u_multiplier/_3328_ ),
    .B2(\u_multiplier/code_y [3]),
    .ZN(\u_multiplier/_3552_ ));
 NOR2_X2 \u_multiplier/_4367_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_3552_ ),
    .ZN(\u_multiplier/_3553_ ));
 NOR2_X1 \u_multiplier/_4368_  (.A1(\u_multiplier/_3546_ ),
    .A2(\u_multiplier/_3553_ ),
    .ZN(\u_multiplier/_3554_ ));
 NAND2_X1 \u_multiplier/_4369_  (.A1(\u_multiplier/_3546_ ),
    .A2(\u_multiplier/_3553_ ),
    .ZN(\u_multiplier/_3555_ ));
 XOR2_X2 \u_multiplier/_4370_  (.A(\u_multiplier/_3546_ ),
    .B(\u_multiplier/_3553_ ),
    .Z(\u_multiplier/_3556_ ));
 XNOR2_X2 \u_multiplier/_4371_  (.A(\u_multiplier/_3539_ ),
    .B(\u_multiplier/_3556_ ),
    .ZN(\u_multiplier/_3557_ ));
 NAND2_X1 \u_multiplier/_4372_  (.A1(\u_multiplier/_3532_ ),
    .A2(\u_multiplier/_3557_ ),
    .ZN(\u_multiplier/_3558_ ));
 XOR2_X2 \u_multiplier/_4373_  (.A(\u_multiplier/_3532_ ),
    .B(\u_multiplier/_3557_ ),
    .Z(\u_multiplier/_3559_ ));
 INV_X1 \u_multiplier/_4374_  (.A(\u_multiplier/_3559_ ),
    .ZN(\u_multiplier/_3560_ ));
 OAI21_X2 \u_multiplier/_4375_  (.A(net21),
    .B1(\u_multiplier/_3531_ ),
    .B2(\u_multiplier/_3559_ ),
    .ZN(\u_multiplier/_3561_ ));
 AOI21_X4 \u_multiplier/_4376_  (.A(\u_multiplier/_3561_ ),
    .B1(\u_multiplier/_3559_ ),
    .B2(\u_multiplier/_3531_ ),
    .ZN(product[8]));
 OAI21_X2 \u_multiplier/_4377_  (.A(\u_multiplier/_3555_ ),
    .B1(\u_multiplier/_3554_ ),
    .B2(\u_multiplier/_3539_ ),
    .ZN(\u_multiplier/_3562_ ));
 MUX2_X1 \u_multiplier/_4378_  (.A(\u_multiplier/_3186_ ),
    .B(\u_multiplier/_3188_ ),
    .S(net17),
    .Z(\u_multiplier/_3563_ ));
 AND2_X1 \u_multiplier/_4379_  (.A1(\u_multiplier/_3113_ ),
    .A2(\u_multiplier/_3563_ ),
    .ZN(\u_multiplier/_3564_ ));
 AOI21_X1 \u_multiplier/_4380_  (.A(\u_multiplier/_3564_ ),
    .B1(\u_multiplier/_3533_ ),
    .B2(\u_multiplier/K [0]),
    .ZN(\u_multiplier/_3565_ ));
 MUX2_X1 \u_multiplier/_4381_  (.A(\u_multiplier/_3506_ ),
    .B(\u_multiplier/_3565_ ),
    .S(\u_multiplier/_3114_ ),
    .Z(\u_multiplier/_3566_ ));
 MUX2_X1 \u_multiplier/_4382_  (.A(\u_multiplier/_3445_ ),
    .B(\u_multiplier/_3566_ ),
    .S(\u_multiplier/_3112_ ),
    .Z(\u_multiplier/_3567_ ));
 NOR2_X1 \u_multiplier/_4383_  (.A1(\u_multiplier/K [3]),
    .A2(\u_multiplier/_3567_ ),
    .ZN(\u_multiplier/_3568_ ));
 AOI21_X4 \u_multiplier/_4384_  (.A(\u_multiplier/_3568_ ),
    .B1(\u_multiplier/_3340_ ),
    .B2(\u_multiplier/K [3]),
    .ZN(\u_multiplier/_3569_ ));
 OAI21_X2 \u_multiplier/_4385_  (.A(\u_multiplier/_3117_ ),
    .B1(\u_multiplier/_3569_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_3570_ ));
 MUX2_X1 \u_multiplier/_4386_  (.A(\u_multiplier/_3186_ ),
    .B(\u_multiplier/_3182_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_3571_ ));
 MUX2_X1 \u_multiplier/_4387_  (.A(\u_multiplier/_3571_ ),
    .B(\u_multiplier/_3512_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_3572_ ));
 OR2_X1 \u_multiplier/_4388_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_3572_ ),
    .ZN(\u_multiplier/_3573_ ));
 OAI21_X1 \u_multiplier/_4389_  (.A(\u_multiplier/_3573_ ),
    .B1(\u_multiplier/_3451_ ),
    .B2(\u_multiplier/_3110_ ),
    .ZN(\u_multiplier/_3574_ ));
 NAND2_X1 \u_multiplier/_4390_  (.A1(\u_multiplier/_3111_ ),
    .A2(\u_multiplier/_3574_ ),
    .ZN(\u_multiplier/_3575_ ));
 OAI21_X2 \u_multiplier/_4391_  (.A(\u_multiplier/_3575_ ),
    .B1(\u_multiplier/_3345_ ),
    .B2(\u_multiplier/_3111_ ),
    .ZN(\u_multiplier/_3576_ ));
 OR2_X1 \u_multiplier/_4392_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_3576_ ),
    .ZN(\u_multiplier/_3577_ ));
 MUX2_X1 \u_multiplier/_4393_  (.A(\u_multiplier/_3184_ ),
    .B(\u_multiplier/_3188_ ),
    .S(\u_multiplier/_3105_ ),
    .Z(\u_multiplier/_3578_ ));
 MUX2_X1 \u_multiplier/_4394_  (.A(\u_multiplier/_3578_ ),
    .B(\u_multiplier/_3517_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_3579_ ));
 OR2_X1 \u_multiplier/_4395_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_3579_ ),
    .ZN(\u_multiplier/_3580_ ));
 OAI21_X1 \u_multiplier/_4396_  (.A(\u_multiplier/_3580_ ),
    .B1(\u_multiplier/_3459_ ),
    .B2(\u_multiplier/_3106_ ),
    .ZN(\u_multiplier/_3581_ ));
 MUX2_X2 \u_multiplier/_4397_  (.A(\u_multiplier/_3349_ ),
    .B(\u_multiplier/_3581_ ),
    .S(\u_multiplier/_3107_ ),
    .Z(\u_multiplier/_3582_ ));
 OR2_X1 \u_multiplier/_4398_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_3582_ ),
    .ZN(\u_multiplier/_3583_ ));
 XOR2_X2 \u_multiplier/_4399_  (.A(\u_multiplier/_3577_ ),
    .B(\u_multiplier/_3583_ ),
    .Z(\u_multiplier/_3584_ ));
 NAND2_X1 \u_multiplier/_4400_  (.A1(\u_multiplier/_3570_ ),
    .A2(\u_multiplier/_3584_ ),
    .ZN(\u_multiplier/_3585_ ));
 XOR2_X2 \u_multiplier/_4401_  (.A(\u_multiplier/_3570_ ),
    .B(\u_multiplier/_3584_ ),
    .Z(\u_multiplier/_3586_ ));
 NAND2_X1 \u_multiplier/_4402_  (.A1(\u_multiplier/_3562_ ),
    .A2(\u_multiplier/_3586_ ),
    .ZN(\u_multiplier/_3587_ ));
 XNOR2_X2 \u_multiplier/_4403_  (.A(\u_multiplier/_3562_ ),
    .B(\u_multiplier/_3586_ ),
    .ZN(\u_multiplier/_3588_ ));
 NAND2_X1 \u_multiplier/_4404_  (.A1(\u_multiplier/_3558_ ),
    .A2(\u_multiplier/_3588_ ),
    .ZN(\u_multiplier/_3589_ ));
 AOI21_X1 \u_multiplier/_4405_  (.A(\u_multiplier/_3589_ ),
    .B1(\u_multiplier/_3559_ ),
    .B2(\u_multiplier/_3531_ ),
    .ZN(\u_multiplier/_3590_ ));
 AOI211_X2 \u_multiplier/_4406_  (.A(\u_multiplier/_3560_ ),
    .B(\u_multiplier/_3588_ ),
    .C1(\u_multiplier/_3526_ ),
    .C2(\u_multiplier/_3529_ ),
    .ZN(\u_multiplier/_3591_ ));
 NOR2_X1 \u_multiplier/_4407_  (.A1(\u_multiplier/_3558_ ),
    .A2(\u_multiplier/_3588_ ),
    .ZN(\u_multiplier/_3592_ ));
 NOR4_X2 \u_multiplier/_4408_  (.A1(\u_multiplier/_3334_ ),
    .A2(\u_multiplier/_3590_ ),
    .A3(\u_multiplier/_3591_ ),
    .A4(\u_multiplier/_3592_ ),
    .ZN(product[9]));
 OAI21_X2 \u_multiplier/_4409_  (.A(\u_multiplier/_3587_ ),
    .B1(\u_multiplier/_3588_ ),
    .B2(\u_multiplier/_3558_ ),
    .ZN(\u_multiplier/_3593_ ));
 OR2_X1 \u_multiplier/_4410_  (.A1(\u_multiplier/_3591_ ),
    .A2(\u_multiplier/_3593_ ),
    .ZN(\u_multiplier/_3594_ ));
 OAI21_X2 \u_multiplier/_4411_  (.A(\u_multiplier/_3585_ ),
    .B1(\u_multiplier/_3583_ ),
    .B2(\u_multiplier/_3577_ ),
    .ZN(\u_multiplier/_3595_ ));
 MUX2_X1 \u_multiplier/_4412_  (.A(\u_multiplier/_3172_ ),
    .B(\u_multiplier/_3174_ ),
    .S(net17),
    .Z(\u_multiplier/_3596_ ));
 MUX2_X1 \u_multiplier/_4413_  (.A(\u_multiplier/_3563_ ),
    .B(\u_multiplier/_3596_ ),
    .S(\u_multiplier/_3113_ ),
    .Z(\u_multiplier/_3597_ ));
 MUX2_X1 \u_multiplier/_4414_  (.A(\u_multiplier/_3534_ ),
    .B(\u_multiplier/_3597_ ),
    .S(\u_multiplier/_3114_ ),
    .Z(\u_multiplier/_3598_ ));
 MUX2_X1 \u_multiplier/_4415_  (.A(\u_multiplier/_3476_ ),
    .B(\u_multiplier/_3598_ ),
    .S(\u_multiplier/_3112_ ),
    .Z(\u_multiplier/_3599_ ));
 MUX2_X2 \u_multiplier/_4416_  (.A(\u_multiplier/_3361_ ),
    .B(\u_multiplier/_3599_ ),
    .S(\u_multiplier/_3115_ ),
    .Z(\u_multiplier/_3600_ ));
 AOI21_X4 \u_multiplier/_4417_  (.A(\u_multiplier/dec_out [10]),
    .B1(\u_multiplier/_3600_ ),
    .B2(\u_multiplier/_3116_ ),
    .ZN(\u_multiplier/_3601_ ));
 MUX2_X1 \u_multiplier/_4418_  (.A(\u_multiplier/_3172_ ),
    .B(\u_multiplier/_3186_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_3602_ ));
 MUX2_X1 \u_multiplier/_4419_  (.A(\u_multiplier/_3602_ ),
    .B(\u_multiplier/_3540_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_3603_ ));
 NAND2_X1 \u_multiplier/_4420_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_3483_ ),
    .ZN(\u_multiplier/_3604_ ));
 OAI21_X1 \u_multiplier/_4421_  (.A(\u_multiplier/_3604_ ),
    .B1(\u_multiplier/_3603_ ),
    .B2(\u_multiplier/code_x [2]),
    .ZN(\u_multiplier/_3605_ ));
 MUX2_X1 \u_multiplier/_4422_  (.A(\u_multiplier/_3365_ ),
    .B(\u_multiplier/_3605_ ),
    .S(\u_multiplier/_3111_ ),
    .Z(\u_multiplier/_3606_ ));
 MUX2_X1 \u_multiplier/_4423_  (.A(\u_multiplier/_3174_ ),
    .B(\u_multiplier/_3188_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_3607_ ));
 MUX2_X1 \u_multiplier/_4424_  (.A(\u_multiplier/_3607_ ),
    .B(\u_multiplier/_3547_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_3608_ ));
 NAND2_X1 \u_multiplier/_4425_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_3490_ ),
    .ZN(\u_multiplier/_3609_ ));
 OAI21_X1 \u_multiplier/_4426_  (.A(\u_multiplier/_3609_ ),
    .B1(\u_multiplier/_3608_ ),
    .B2(\u_multiplier/code_y [2]),
    .ZN(\u_multiplier/_3610_ ));
 MUX2_X2 \u_multiplier/_4427_  (.A(\u_multiplier/_3370_ ),
    .B(\u_multiplier/_3610_ ),
    .S(\u_multiplier/_3107_ ),
    .Z(\u_multiplier/_3611_ ));
 OAI22_X1 \u_multiplier/_4428_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_3606_ ),
    .B1(\u_multiplier/_3611_ ),
    .B2(\u_multiplier/code_y [4]),
    .ZN(\u_multiplier/_3612_ ));
 OR4_X1 \u_multiplier/_4429_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/code_x [4]),
    .A3(\u_multiplier/_3606_ ),
    .A4(\u_multiplier/_3611_ ),
    .ZN(\u_multiplier/_3613_ ));
 AND2_X1 \u_multiplier/_4430_  (.A1(\u_multiplier/_3612_ ),
    .A2(\u_multiplier/_3613_ ),
    .ZN(\u_multiplier/_3614_ ));
 INV_X1 \u_multiplier/_4431_  (.A(\u_multiplier/_3614_ ),
    .ZN(\u_multiplier/_3615_ ));
 XNOR2_X2 \u_multiplier/_4432_  (.A(\u_multiplier/_3601_ ),
    .B(\u_multiplier/_3614_ ),
    .ZN(\u_multiplier/_3616_ ));
 AND2_X1 \u_multiplier/_4433_  (.A1(\u_multiplier/_3595_ ),
    .A2(\u_multiplier/_3616_ ),
    .ZN(\u_multiplier/_3617_ ));
 XOR2_X2 \u_multiplier/_4434_  (.A(\u_multiplier/_3595_ ),
    .B(\u_multiplier/_3616_ ),
    .Z(\u_multiplier/_3618_ ));
 AND2_X1 \u_multiplier/_4435_  (.A1(\u_multiplier/_3594_ ),
    .A2(\u_multiplier/_3618_ ),
    .ZN(\u_multiplier/_3619_ ));
 NOR3_X2 \u_multiplier/_4436_  (.A1(\u_multiplier/_3591_ ),
    .A2(\u_multiplier/_3593_ ),
    .A3(\u_multiplier/_3618_ ),
    .ZN(\u_multiplier/_3620_ ));
 NOR3_X4 \u_multiplier/_4437_  (.A1(\u_multiplier/_3334_ ),
    .A2(\u_multiplier/_3619_ ),
    .A3(\u_multiplier/_3620_ ),
    .ZN(product[10]));
 OAI21_X2 \u_multiplier/_4438_  (.A(\u_multiplier/_3613_ ),
    .B1(\u_multiplier/_3615_ ),
    .B2(\u_multiplier/_3601_ ),
    .ZN(\u_multiplier/_3621_ ));
 MUX2_X1 \u_multiplier/_4439_  (.A(\u_multiplier/_3175_ ),
    .B(\u_multiplier/_3177_ ),
    .S(net17),
    .Z(\u_multiplier/_3622_ ));
 MUX2_X1 \u_multiplier/_4440_  (.A(\u_multiplier/_3596_ ),
    .B(\u_multiplier/_3622_ ),
    .S(\u_multiplier/_3113_ ),
    .Z(\u_multiplier/_3623_ ));
 NAND2_X1 \u_multiplier/_4441_  (.A1(\u_multiplier/_3114_ ),
    .A2(\u_multiplier/_3623_ ),
    .ZN(\u_multiplier/_3624_ ));
 OAI21_X1 \u_multiplier/_4442_  (.A(\u_multiplier/_3624_ ),
    .B1(\u_multiplier/_3565_ ),
    .B2(\u_multiplier/_3114_ ),
    .ZN(\u_multiplier/_3625_ ));
 NAND2_X1 \u_multiplier/_4443_  (.A1(\u_multiplier/_3112_ ),
    .A2(\u_multiplier/_3625_ ),
    .ZN(\u_multiplier/_3626_ ));
 OAI21_X1 \u_multiplier/_4444_  (.A(\u_multiplier/_3626_ ),
    .B1(\u_multiplier/_3508_ ),
    .B2(\u_multiplier/_3112_ ),
    .ZN(\u_multiplier/_3627_ ));
 MUX2_X2 \u_multiplier/_4445_  (.A(\u_multiplier/_3390_ ),
    .B(\u_multiplier/_3627_ ),
    .S(\u_multiplier/_3115_ ),
    .Z(\u_multiplier/_3628_ ));
 AOI21_X2 \u_multiplier/_4446_  (.A(\u_multiplier/dec_out [11]),
    .B1(\u_multiplier/_3628_ ),
    .B2(\u_multiplier/_3116_ ),
    .ZN(\u_multiplier/_3629_ ));
 MUX2_X1 \u_multiplier/_4447_  (.A(\u_multiplier/_3175_ ),
    .B(\u_multiplier/_3172_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_3630_ ));
 MUX2_X1 \u_multiplier/_4448_  (.A(\u_multiplier/_3630_ ),
    .B(\u_multiplier/_3571_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_3631_ ));
 MUX2_X1 \u_multiplier/_4449_  (.A(\u_multiplier/_3513_ ),
    .B(\u_multiplier/_3631_ ),
    .S(\u_multiplier/_3110_ ),
    .Z(\u_multiplier/_3632_ ));
 NAND2_X1 \u_multiplier/_4450_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_3395_ ),
    .ZN(\u_multiplier/_3633_ ));
 OAI21_X2 \u_multiplier/_4451_  (.A(\u_multiplier/_3633_ ),
    .B1(\u_multiplier/_3632_ ),
    .B2(\u_multiplier/code_x [3]),
    .ZN(\u_multiplier/_3634_ ));
 OR2_X1 \u_multiplier/_4452_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_3634_ ),
    .ZN(\u_multiplier/_3635_ ));
 MUX2_X1 \u_multiplier/_4453_  (.A(\u_multiplier/_3174_ ),
    .B(\u_multiplier/_3177_ ),
    .S(\u_multiplier/_3105_ ),
    .Z(\u_multiplier/_3636_ ));
 MUX2_X1 \u_multiplier/_4454_  (.A(\u_multiplier/_3636_ ),
    .B(\u_multiplier/_3578_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_3637_ ));
 NAND2_X1 \u_multiplier/_4455_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_3519_ ),
    .ZN(\u_multiplier/_3638_ ));
 OAI21_X1 \u_multiplier/_4456_  (.A(\u_multiplier/_3638_ ),
    .B1(\u_multiplier/_3637_ ),
    .B2(\u_multiplier/code_y [2]),
    .ZN(\u_multiplier/_3639_ ));
 MUX2_X2 \u_multiplier/_4457_  (.A(\u_multiplier/_3399_ ),
    .B(\u_multiplier/_3639_ ),
    .S(\u_multiplier/_3107_ ),
    .Z(\u_multiplier/_3640_ ));
 OAI21_X1 \u_multiplier/_4458_  (.A(\u_multiplier/_3635_ ),
    .B1(\u_multiplier/_3640_ ),
    .B2(\u_multiplier/code_y [4]),
    .ZN(\u_multiplier/_3641_ ));
 OR3_X1 \u_multiplier/_4459_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_3635_ ),
    .A3(\u_multiplier/_3640_ ),
    .ZN(\u_multiplier/_3642_ ));
 AND2_X1 \u_multiplier/_4460_  (.A1(\u_multiplier/_3641_ ),
    .A2(\u_multiplier/_3642_ ),
    .ZN(\u_multiplier/_3643_ ));
 INV_X1 \u_multiplier/_4461_  (.A(\u_multiplier/_3643_ ),
    .ZN(\u_multiplier/_3644_ ));
 XNOR2_X2 \u_multiplier/_4462_  (.A(\u_multiplier/_3629_ ),
    .B(\u_multiplier/_3643_ ),
    .ZN(\u_multiplier/_3645_ ));
 XOR2_X2 \u_multiplier/_4463_  (.A(\u_multiplier/_3621_ ),
    .B(\u_multiplier/_3645_ ),
    .Z(\u_multiplier/_3646_ ));
 OR3_X1 \u_multiplier/_4464_  (.A1(\u_multiplier/_3617_ ),
    .A2(\u_multiplier/_3619_ ),
    .A3(\u_multiplier/_3646_ ),
    .ZN(\u_multiplier/_3647_ ));
 OAI211_X4 \u_multiplier/_4465_  (.A(\u_multiplier/_3618_ ),
    .B(\u_multiplier/_3646_ ),
    .C1(\u_multiplier/_3591_ ),
    .C2(\u_multiplier/_3593_ ),
    .ZN(\u_multiplier/_3648_ ));
 NAND2_X1 \u_multiplier/_4466_  (.A1(\u_multiplier/_3617_ ),
    .A2(\u_multiplier/_3646_ ),
    .ZN(\u_multiplier/_3649_ ));
 INV_X1 \u_multiplier/_4467_  (.A(\u_multiplier/_3649_ ),
    .ZN(\u_multiplier/_3650_ ));
 AND4_X1 \u_multiplier/_4468_  (.A1(net21),
    .A2(\u_multiplier/_3647_ ),
    .A3(\u_multiplier/_3648_ ),
    .A4(\u_multiplier/_3649_ ),
    .ZN(product[11]));
 AOI21_X2 \u_multiplier/_4469_  (.A(\u_multiplier/_3650_ ),
    .B1(\u_multiplier/_3645_ ),
    .B2(\u_multiplier/_3621_ ),
    .ZN(\u_multiplier/_3651_ ));
 NAND2_X1 \u_multiplier/_4470_  (.A1(\u_multiplier/_3648_ ),
    .A2(\u_multiplier/_3651_ ),
    .ZN(\u_multiplier/_3652_ ));
 OAI21_X1 \u_multiplier/_4471_  (.A(\u_multiplier/_3642_ ),
    .B1(\u_multiplier/_3644_ ),
    .B2(\u_multiplier/_3629_ ),
    .ZN(\u_multiplier/_3653_ ));
 MUX2_X1 \u_multiplier/_4472_  (.A(\u_multiplier/_3215_ ),
    .B(\u_multiplier/_3216_ ),
    .S(net17),
    .Z(\u_multiplier/_3654_ ));
 MUX2_X1 \u_multiplier/_4473_  (.A(\u_multiplier/_3622_ ),
    .B(\u_multiplier/_3654_ ),
    .S(\u_multiplier/_3113_ ),
    .Z(\u_multiplier/_3655_ ));
 MUX2_X1 \u_multiplier/_4474_  (.A(\u_multiplier/_3597_ ),
    .B(\u_multiplier/_3655_ ),
    .S(\u_multiplier/_3114_ ),
    .Z(\u_multiplier/_3656_ ));
 MUX2_X2 \u_multiplier/_4475_  (.A(\u_multiplier/_3535_ ),
    .B(\u_multiplier/_3656_ ),
    .S(\u_multiplier/_3112_ ),
    .Z(\u_multiplier/_3657_ ));
 NOR2_X1 \u_multiplier/_4476_  (.A1(\u_multiplier/_3115_ ),
    .A2(\u_multiplier/_3415_ ),
    .ZN(\u_multiplier/_3658_ ));
 AOI21_X4 \u_multiplier/_4477_  (.A(\u_multiplier/_3658_ ),
    .B1(\u_multiplier/_3657_ ),
    .B2(\u_multiplier/_3115_ ),
    .ZN(\u_multiplier/_3659_ ));
 NOR2_X1 \u_multiplier/_4478_  (.A1(\u_multiplier/K [4]),
    .A2(\u_multiplier/_3659_ ),
    .ZN(\u_multiplier/_3660_ ));
 NOR2_X1 \u_multiplier/_4479_  (.A1(\u_multiplier/dec_out [12]),
    .A2(\u_multiplier/_3660_ ),
    .ZN(\u_multiplier/_3661_ ));
 MUX2_X1 \u_multiplier/_4480_  (.A(\u_multiplier/_3215_ ),
    .B(\u_multiplier/_3175_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_3662_ ));
 MUX2_X1 \u_multiplier/_4481_  (.A(\u_multiplier/_3662_ ),
    .B(\u_multiplier/_3602_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_3663_ ));
 OR2_X1 \u_multiplier/_4482_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_3663_ ),
    .ZN(\u_multiplier/_3664_ ));
 OAI21_X1 \u_multiplier/_4483_  (.A(\u_multiplier/_3664_ ),
    .B1(\u_multiplier/_3541_ ),
    .B2(\u_multiplier/_3110_ ),
    .ZN(\u_multiplier/_3665_ ));
 NAND2_X1 \u_multiplier/_4484_  (.A1(\u_multiplier/_3111_ ),
    .A2(\u_multiplier/_3665_ ),
    .ZN(\u_multiplier/_3666_ ));
 OAI21_X2 \u_multiplier/_4485_  (.A(\u_multiplier/_3666_ ),
    .B1(\u_multiplier/_3421_ ),
    .B2(\u_multiplier/_3111_ ),
    .ZN(\u_multiplier/_3667_ ));
 OR2_X1 \u_multiplier/_4486_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_3667_ ),
    .ZN(\u_multiplier/_3668_ ));
 MUX2_X1 \u_multiplier/_4487_  (.A(\u_multiplier/_3177_ ),
    .B(\u_multiplier/_3216_ ),
    .S(\u_multiplier/_3105_ ),
    .Z(\u_multiplier/_3669_ ));
 MUX2_X1 \u_multiplier/_4488_  (.A(\u_multiplier/_3669_ ),
    .B(\u_multiplier/_3607_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_3670_ ));
 OR2_X1 \u_multiplier/_4489_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_3670_ ),
    .ZN(\u_multiplier/_3671_ ));
 OAI21_X1 \u_multiplier/_4490_  (.A(\u_multiplier/_3671_ ),
    .B1(\u_multiplier/_3548_ ),
    .B2(\u_multiplier/_3106_ ),
    .ZN(\u_multiplier/_3672_ ));
 NOR2_X1 \u_multiplier/_4491_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_3672_ ),
    .ZN(\u_multiplier/_3673_ ));
 AOI21_X4 \u_multiplier/_4492_  (.A(\u_multiplier/_3673_ ),
    .B1(\u_multiplier/_3428_ ),
    .B2(\u_multiplier/code_y [3]),
    .ZN(\u_multiplier/_3674_ ));
 OR2_X1 \u_multiplier/_4493_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_3674_ ),
    .ZN(\u_multiplier/_3675_ ));
 XOR2_X2 \u_multiplier/_4494_  (.A(\u_multiplier/_3668_ ),
    .B(\u_multiplier/_3675_ ),
    .Z(\u_multiplier/_3676_ ));
 OAI21_X1 \u_multiplier/_4495_  (.A(\u_multiplier/_3676_ ),
    .B1(\u_multiplier/_3660_ ),
    .B2(\u_multiplier/dec_out [12]),
    .ZN(\u_multiplier/_3677_ ));
 XNOR2_X2 \u_multiplier/_4496_  (.A(\u_multiplier/_3661_ ),
    .B(\u_multiplier/_3676_ ),
    .ZN(\u_multiplier/_3678_ ));
 AND2_X1 \u_multiplier/_4497_  (.A1(\u_multiplier/_3653_ ),
    .A2(\u_multiplier/_3678_ ),
    .ZN(\u_multiplier/_3679_ ));
 XOR2_X2 \u_multiplier/_4498_  (.A(\u_multiplier/_3653_ ),
    .B(\u_multiplier/_3678_ ),
    .Z(\u_multiplier/_3680_ ));
 INV_X1 \u_multiplier/_4499_  (.A(\u_multiplier/_3680_ ),
    .ZN(\u_multiplier/_3681_ ));
 AOI21_X2 \u_multiplier/_4500_  (.A(\u_multiplier/_3681_ ),
    .B1(\u_multiplier/_3651_ ),
    .B2(\u_multiplier/_3648_ ),
    .ZN(\u_multiplier/_3682_ ));
 OAI21_X1 \u_multiplier/_4501_  (.A(net21),
    .B1(\u_multiplier/_3652_ ),
    .B2(\u_multiplier/_3680_ ),
    .ZN(\u_multiplier/_3683_ ));
 NOR2_X1 \u_multiplier/_4502_  (.A1(\u_multiplier/_3682_ ),
    .A2(\u_multiplier/_3683_ ),
    .ZN(product[12]));
 OAI21_X2 \u_multiplier/_4503_  (.A(\u_multiplier/_3677_ ),
    .B1(\u_multiplier/_3675_ ),
    .B2(\u_multiplier/_3668_ ),
    .ZN(\u_multiplier/_3684_ ));
 MUX2_X1 \u_multiplier/_4504_  (.A(\u_multiplier/_3211_ ),
    .B(\u_multiplier/_3213_ ),
    .S(net17),
    .Z(\u_multiplier/_3685_ ));
 MUX2_X1 \u_multiplier/_4505_  (.A(\u_multiplier/_3654_ ),
    .B(\u_multiplier/_3685_ ),
    .S(\u_multiplier/_3113_ ),
    .Z(\u_multiplier/_3686_ ));
 MUX2_X1 \u_multiplier/_4506_  (.A(\u_multiplier/_3623_ ),
    .B(\u_multiplier/_3686_ ),
    .S(\u_multiplier/_3114_ ),
    .Z(\u_multiplier/_3687_ ));
 NAND2_X1 \u_multiplier/_4507_  (.A1(\u_multiplier/_3112_ ),
    .A2(\u_multiplier/_3687_ ),
    .ZN(\u_multiplier/_3688_ ));
 OAI21_X2 \u_multiplier/_4508_  (.A(\u_multiplier/_3688_ ),
    .B1(\u_multiplier/_3566_ ),
    .B2(\u_multiplier/_3112_ ),
    .ZN(\u_multiplier/_3689_ ));
 NOR2_X1 \u_multiplier/_4509_  (.A1(\u_multiplier/_3115_ ),
    .A2(\u_multiplier/_3446_ ),
    .ZN(\u_multiplier/_3690_ ));
 AOI21_X4 \u_multiplier/_4510_  (.A(\u_multiplier/_3690_ ),
    .B1(\u_multiplier/_3689_ ),
    .B2(\u_multiplier/_3115_ ),
    .ZN(\u_multiplier/_3691_ ));
 NOR2_X1 \u_multiplier/_4511_  (.A1(\u_multiplier/K [4]),
    .A2(\u_multiplier/_3691_ ),
    .ZN(\u_multiplier/_3692_ ));
 NOR2_X2 \u_multiplier/_4512_  (.A1(\u_multiplier/dec_out [13]),
    .A2(\u_multiplier/_3692_ ),
    .ZN(\u_multiplier/_3693_ ));
 INV_X1 \u_multiplier/_4513_  (.A(\u_multiplier/_3693_ ),
    .ZN(\u_multiplier/_3694_ ));
 MUX2_X1 \u_multiplier/_4514_  (.A(\u_multiplier/_3211_ ),
    .B(\u_multiplier/_3215_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_3695_ ));
 MUX2_X1 \u_multiplier/_4515_  (.A(\u_multiplier/_3695_ ),
    .B(\u_multiplier/_3630_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_3696_ ));
 OR2_X1 \u_multiplier/_4516_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_3696_ ),
    .ZN(\u_multiplier/_3697_ ));
 OAI21_X1 \u_multiplier/_4517_  (.A(\u_multiplier/_3697_ ),
    .B1(\u_multiplier/_3572_ ),
    .B2(\u_multiplier/_3110_ ),
    .ZN(\u_multiplier/_3698_ ));
 NAND2_X1 \u_multiplier/_4518_  (.A1(\u_multiplier/_3111_ ),
    .A2(\u_multiplier/_3698_ ),
    .ZN(\u_multiplier/_3699_ ));
 OAI21_X2 \u_multiplier/_4519_  (.A(\u_multiplier/_3699_ ),
    .B1(\u_multiplier/_3453_ ),
    .B2(\u_multiplier/_3111_ ),
    .ZN(\u_multiplier/_3700_ ));
 OR2_X1 \u_multiplier/_4520_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_3700_ ),
    .ZN(\u_multiplier/_3701_ ));
 MUX2_X1 \u_multiplier/_4521_  (.A(\u_multiplier/_3213_ ),
    .B(\u_multiplier/_3216_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_3702_ ));
 MUX2_X1 \u_multiplier/_4522_  (.A(\u_multiplier/_3702_ ),
    .B(\u_multiplier/_3636_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_3703_ ));
 OR2_X1 \u_multiplier/_4523_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_3703_ ),
    .ZN(\u_multiplier/_3704_ ));
 OAI21_X1 \u_multiplier/_4524_  (.A(\u_multiplier/_3704_ ),
    .B1(\u_multiplier/_3579_ ),
    .B2(\u_multiplier/_3106_ ),
    .ZN(\u_multiplier/_3705_ ));
 NOR2_X1 \u_multiplier/_4525_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_3705_ ),
    .ZN(\u_multiplier/_3706_ ));
 AOI21_X4 \u_multiplier/_4526_  (.A(\u_multiplier/_3706_ ),
    .B1(\u_multiplier/_3461_ ),
    .B2(\u_multiplier/code_y [3]),
    .ZN(\u_multiplier/_3707_ ));
 NOR2_X1 \u_multiplier/_4527_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_3707_ ),
    .ZN(\u_multiplier/_3708_ ));
 NOR3_X1 \u_multiplier/_4528_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_3701_ ),
    .A3(\u_multiplier/_3707_ ),
    .ZN(\u_multiplier/_3709_ ));
 XNOR2_X2 \u_multiplier/_4529_  (.A(\u_multiplier/_3701_ ),
    .B(\u_multiplier/_3708_ ),
    .ZN(\u_multiplier/_3710_ ));
 XNOR2_X2 \u_multiplier/_4530_  (.A(\u_multiplier/_3693_ ),
    .B(\u_multiplier/_3710_ ),
    .ZN(\u_multiplier/_3711_ ));
 AND2_X1 \u_multiplier/_4531_  (.A1(\u_multiplier/_3684_ ),
    .A2(\u_multiplier/_3711_ ),
    .ZN(\u_multiplier/_3712_ ));
 XOR2_X2 \u_multiplier/_4532_  (.A(\u_multiplier/_3684_ ),
    .B(\u_multiplier/_3711_ ),
    .Z(\u_multiplier/_3713_ ));
 INV_X1 \u_multiplier/_4533_  (.A(\u_multiplier/_3713_ ),
    .ZN(\u_multiplier/_3714_ ));
 NOR3_X2 \u_multiplier/_4534_  (.A1(\u_multiplier/_3679_ ),
    .A2(\u_multiplier/_3682_ ),
    .A3(\u_multiplier/_3713_ ),
    .ZN(\u_multiplier/_3715_ ));
 AOI211_X2 \u_multiplier/_4535_  (.A(\u_multiplier/_3681_ ),
    .B(\u_multiplier/_3714_ ),
    .C1(\u_multiplier/_3648_ ),
    .C2(\u_multiplier/_3651_ ),
    .ZN(\u_multiplier/_3716_ ));
 AND2_X1 \u_multiplier/_4536_  (.A1(\u_multiplier/_3679_ ),
    .A2(\u_multiplier/_3713_ ),
    .ZN(\u_multiplier/_3717_ ));
 NOR4_X4 \u_multiplier/_4537_  (.A1(\u_multiplier/_3334_ ),
    .A2(\u_multiplier/_3715_ ),
    .A3(\u_multiplier/_3716_ ),
    .A4(\u_multiplier/_3717_ ),
    .ZN(product[13]));
 OR2_X2 \u_multiplier/_4538_  (.A1(\u_multiplier/_3712_ ),
    .A2(\u_multiplier/_3717_ ),
    .ZN(\u_multiplier/_3718_ ));
 NOR2_X1 \u_multiplier/_4539_  (.A1(\u_multiplier/_3716_ ),
    .A2(\u_multiplier/_3718_ ),
    .ZN(\u_multiplier/_3719_ ));
 AOI21_X1 \u_multiplier/_4540_  (.A(\u_multiplier/_3709_ ),
    .B1(\u_multiplier/_3710_ ),
    .B2(\u_multiplier/_3694_ ),
    .ZN(\u_multiplier/_3720_ ));
 MUX2_X1 \u_multiplier/_4541_  (.A(\u_multiplier/_3200_ ),
    .B(\u_multiplier/_3202_ ),
    .S(net17),
    .Z(\u_multiplier/_3721_ ));
 MUX2_X1 \u_multiplier/_4542_  (.A(\u_multiplier/_3685_ ),
    .B(\u_multiplier/_3721_ ),
    .S(\u_multiplier/_3113_ ),
    .Z(\u_multiplier/_3722_ ));
 MUX2_X1 \u_multiplier/_4543_  (.A(\u_multiplier/_3655_ ),
    .B(\u_multiplier/_3722_ ),
    .S(\u_multiplier/_3114_ ),
    .Z(\u_multiplier/_3723_ ));
 AND2_X1 \u_multiplier/_4544_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/_3598_ ),
    .ZN(\u_multiplier/_3724_ ));
 AOI21_X2 \u_multiplier/_4545_  (.A(\u_multiplier/_3724_ ),
    .B1(\u_multiplier/_3723_ ),
    .B2(\u_multiplier/_3112_ ),
    .ZN(\u_multiplier/_3725_ ));
 MUX2_X2 \u_multiplier/_4546_  (.A(\u_multiplier/_3478_ ),
    .B(\u_multiplier/_3725_ ),
    .S(\u_multiplier/_3115_ ),
    .Z(\u_multiplier/_3726_ ));
 OAI21_X1 \u_multiplier/_4547_  (.A(\u_multiplier/_3118_ ),
    .B1(\u_multiplier/_3726_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_3727_ ));
 MUX2_X1 \u_multiplier/_4548_  (.A(\u_multiplier/_3200_ ),
    .B(\u_multiplier/_3211_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_3728_ ));
 MUX2_X1 \u_multiplier/_4549_  (.A(\u_multiplier/_3728_ ),
    .B(\u_multiplier/_3662_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_3729_ ));
 OR2_X1 \u_multiplier/_4550_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_3729_ ),
    .ZN(\u_multiplier/_3730_ ));
 OAI21_X1 \u_multiplier/_4551_  (.A(\u_multiplier/_3730_ ),
    .B1(\u_multiplier/_3603_ ),
    .B2(\u_multiplier/_3110_ ),
    .ZN(\u_multiplier/_3731_ ));
 MUX2_X2 \u_multiplier/_4552_  (.A(\u_multiplier/_3485_ ),
    .B(\u_multiplier/_3731_ ),
    .S(\u_multiplier/_3111_ ),
    .Z(\u_multiplier/_3732_ ));
 NOR2_X2 \u_multiplier/_4553_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_3732_ ),
    .ZN(\u_multiplier/_3733_ ));
 MUX2_X1 \u_multiplier/_4554_  (.A(\u_multiplier/_3202_ ),
    .B(\u_multiplier/_3213_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_3734_ ));
 MUX2_X1 \u_multiplier/_4555_  (.A(\u_multiplier/_3734_ ),
    .B(\u_multiplier/_3669_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_3735_ ));
 OR2_X1 \u_multiplier/_4556_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_3735_ ),
    .ZN(\u_multiplier/_3736_ ));
 OAI21_X2 \u_multiplier/_4557_  (.A(\u_multiplier/_3736_ ),
    .B1(\u_multiplier/_3608_ ),
    .B2(\u_multiplier/_3106_ ),
    .ZN(\u_multiplier/_3737_ ));
 MUX2_X2 \u_multiplier/_4558_  (.A(\u_multiplier/_3492_ ),
    .B(\u_multiplier/_3737_ ),
    .S(\u_multiplier/_3107_ ),
    .Z(\u_multiplier/_3738_ ));
 NOR2_X2 \u_multiplier/_4559_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_3738_ ),
    .ZN(\u_multiplier/_3739_ ));
 XOR2_X2 \u_multiplier/_4560_  (.A(\u_multiplier/_3733_ ),
    .B(\u_multiplier/_3739_ ),
    .Z(\u_multiplier/_3740_ ));
 AND2_X1 \u_multiplier/_4561_  (.A1(\u_multiplier/_3727_ ),
    .A2(\u_multiplier/_3740_ ),
    .ZN(\u_multiplier/_3741_ ));
 XOR2_X1 \u_multiplier/_4562_  (.A(\u_multiplier/_3727_ ),
    .B(\u_multiplier/_3740_ ),
    .Z(\u_multiplier/_3742_ ));
 INV_X1 \u_multiplier/_4563_  (.A(\u_multiplier/_3742_ ),
    .ZN(\u_multiplier/_3743_ ));
 NOR2_X1 \u_multiplier/_4564_  (.A1(\u_multiplier/_3720_ ),
    .A2(\u_multiplier/_3743_ ),
    .ZN(\u_multiplier/_3744_ ));
 XNOR2_X1 \u_multiplier/_4565_  (.A(\u_multiplier/_3720_ ),
    .B(\u_multiplier/_3743_ ),
    .ZN(\u_multiplier/_3745_ ));
 INV_X1 \u_multiplier/_4566_  (.A(\u_multiplier/_3745_ ),
    .ZN(\u_multiplier/_3746_ ));
 NOR2_X1 \u_multiplier/_4567_  (.A1(\u_multiplier/_3719_ ),
    .A2(\u_multiplier/_3745_ ),
    .ZN(\u_multiplier/_3747_ ));
 NOR3_X1 \u_multiplier/_4568_  (.A1(\u_multiplier/_3716_ ),
    .A2(\u_multiplier/_3718_ ),
    .A3(\u_multiplier/_3746_ ),
    .ZN(\u_multiplier/_3748_ ));
 NOR3_X1 \u_multiplier/_4569_  (.A1(\u_multiplier/_3334_ ),
    .A2(\u_multiplier/_3747_ ),
    .A3(\u_multiplier/_3748_ ),
    .ZN(product[14]));
 AOI21_X2 \u_multiplier/_4570_  (.A(\u_multiplier/_3741_ ),
    .B1(\u_multiplier/_3739_ ),
    .B2(\u_multiplier/_3733_ ),
    .ZN(\u_multiplier/_3749_ ));
 INV_X1 \u_multiplier/_4571_  (.A(\u_multiplier/_3749_ ),
    .ZN(\u_multiplier/_3750_ ));
 MUX2_X1 \u_multiplier/_4572_  (.A(\u_multiplier/_3204_ ),
    .B(\u_multiplier/_3206_ ),
    .S(net17),
    .Z(\u_multiplier/_3751_ ));
 AND2_X1 \u_multiplier/_4573_  (.A1(\u_multiplier/_3113_ ),
    .A2(\u_multiplier/_3751_ ),
    .ZN(\u_multiplier/_2003_ ));
 AOI21_X1 \u_multiplier/_4574_  (.A(\u_multiplier/_2003_ ),
    .B1(\u_multiplier/_3721_ ),
    .B2(\u_multiplier/K [0]),
    .ZN(\u_multiplier/_2004_ ));
 NAND2_X1 \u_multiplier/_4575_  (.A1(\u_multiplier/K [1]),
    .A2(\u_multiplier/_3686_ ),
    .ZN(\u_multiplier/_2005_ ));
 OAI21_X1 \u_multiplier/_4576_  (.A(\u_multiplier/_2005_ ),
    .B1(\u_multiplier/_2004_ ),
    .B2(\u_multiplier/K [1]),
    .ZN(\u_multiplier/_2006_ ));
 MUX2_X1 \u_multiplier/_4577_  (.A(\u_multiplier/_3625_ ),
    .B(\u_multiplier/_2006_ ),
    .S(\u_multiplier/_3112_ ),
    .Z(\u_multiplier/_2007_ ));
 NAND2_X1 \u_multiplier/_4578_  (.A1(\u_multiplier/_3115_ ),
    .A2(\u_multiplier/_2007_ ),
    .ZN(\u_multiplier/_2008_ ));
 OAI21_X4 \u_multiplier/_4579_  (.A(\u_multiplier/_2008_ ),
    .B1(\u_multiplier/_3509_ ),
    .B2(\u_multiplier/_3115_ ),
    .ZN(\u_multiplier/_2009_ ));
 AOI21_X2 \u_multiplier/_4580_  (.A(\u_multiplier/dec_out [15]),
    .B1(\u_multiplier/_2009_ ),
    .B2(\u_multiplier/_3116_ ),
    .ZN(\u_multiplier/_2010_ ));
 MUX2_X1 \u_multiplier/_4581_  (.A(\u_multiplier/_3204_ ),
    .B(\u_multiplier/_3200_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_2011_ ));
 MUX2_X1 \u_multiplier/_4582_  (.A(\u_multiplier/_2011_ ),
    .B(\u_multiplier/_3695_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_2012_ ));
 MUX2_X1 \u_multiplier/_4583_  (.A(\u_multiplier/_3631_ ),
    .B(\u_multiplier/_2012_ ),
    .S(\u_multiplier/_3110_ ),
    .Z(\u_multiplier/_2013_ ));
 NAND2_X1 \u_multiplier/_4584_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_3515_ ),
    .ZN(\u_multiplier/_2014_ ));
 OAI21_X2 \u_multiplier/_4585_  (.A(\u_multiplier/_2014_ ),
    .B1(\u_multiplier/_2013_ ),
    .B2(\u_multiplier/code_x [3]),
    .ZN(\u_multiplier/_2015_ ));
 NOR2_X2 \u_multiplier/_4586_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2015_ ),
    .ZN(\u_multiplier/_2016_ ));
 MUX2_X1 \u_multiplier/_4587_  (.A(\u_multiplier/_3202_ ),
    .B(\u_multiplier/_3206_ ),
    .S(\u_multiplier/_3105_ ),
    .Z(\u_multiplier/_2017_ ));
 MUX2_X1 \u_multiplier/_4588_  (.A(\u_multiplier/_2017_ ),
    .B(\u_multiplier/_3702_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_2018_ ));
 OR2_X1 \u_multiplier/_4589_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_2018_ ),
    .ZN(\u_multiplier/_2019_ ));
 OAI21_X2 \u_multiplier/_4590_  (.A(\u_multiplier/_2019_ ),
    .B1(\u_multiplier/_3637_ ),
    .B2(\u_multiplier/_3106_ ),
    .ZN(\u_multiplier/_2020_ ));
 MUX2_X2 \u_multiplier/_4591_  (.A(\u_multiplier/_3520_ ),
    .B(\u_multiplier/_2020_ ),
    .S(\u_multiplier/_3107_ ),
    .Z(\u_multiplier/_2021_ ));
 NOR2_X2 \u_multiplier/_4592_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_2021_ ),
    .ZN(\u_multiplier/_2022_ ));
 XNOR2_X2 \u_multiplier/_4593_  (.A(\u_multiplier/_2016_ ),
    .B(\u_multiplier/_2022_ ),
    .ZN(\u_multiplier/_2023_ ));
 NOR2_X1 \u_multiplier/_4594_  (.A1(\u_multiplier/_2010_ ),
    .A2(\u_multiplier/_2023_ ),
    .ZN(\u_multiplier/_2024_ ));
 XOR2_X2 \u_multiplier/_4595_  (.A(\u_multiplier/_2010_ ),
    .B(\u_multiplier/_2023_ ),
    .Z(\u_multiplier/_2025_ ));
 NAND2_X1 \u_multiplier/_4596_  (.A1(\u_multiplier/_3750_ ),
    .A2(\u_multiplier/_2025_ ),
    .ZN(\u_multiplier/_2026_ ));
 XNOR2_X2 \u_multiplier/_4597_  (.A(\u_multiplier/_3749_ ),
    .B(\u_multiplier/_2025_ ),
    .ZN(\u_multiplier/_2027_ ));
 OR3_X1 \u_multiplier/_4598_  (.A1(\u_multiplier/_3744_ ),
    .A2(\u_multiplier/_3747_ ),
    .A3(\u_multiplier/_2027_ ),
    .ZN(\u_multiplier/_2028_ ));
 OAI211_X4 \u_multiplier/_4599_  (.A(\u_multiplier/_3746_ ),
    .B(\u_multiplier/_2027_ ),
    .C1(\u_multiplier/_3716_ ),
    .C2(\u_multiplier/_3718_ ),
    .ZN(\u_multiplier/_2029_ ));
 NAND2_X1 \u_multiplier/_4600_  (.A1(\u_multiplier/_3744_ ),
    .A2(\u_multiplier/_2027_ ),
    .ZN(\u_multiplier/_2030_ ));
 AND4_X2 \u_multiplier/_4601_  (.A1(net21),
    .A2(\u_multiplier/_2028_ ),
    .A3(\u_multiplier/_2029_ ),
    .A4(\u_multiplier/_2030_ ),
    .ZN(product[15]));
 AND2_X1 \u_multiplier/_4602_  (.A1(\u_multiplier/_2026_ ),
    .A2(\u_multiplier/_2030_ ),
    .ZN(\u_multiplier/_2031_ ));
 NAND2_X2 \u_multiplier/_4603_  (.A1(\u_multiplier/_2029_ ),
    .A2(\u_multiplier/_2031_ ),
    .ZN(\u_multiplier/_2032_ ));
 AOI21_X2 \u_multiplier/_4604_  (.A(\u_multiplier/_2024_ ),
    .B1(\u_multiplier/_2022_ ),
    .B2(\u_multiplier/_2016_ ),
    .ZN(\u_multiplier/_2033_ ));
 MUX2_X1 \u_multiplier/_4605_  (.A(\u_multiplier/_3262_ ),
    .B(\u_multiplier/_3261_ ),
    .S(net17),
    .Z(\u_multiplier/_2034_ ));
 MUX2_X1 \u_multiplier/_4606_  (.A(\u_multiplier/_3751_ ),
    .B(\u_multiplier/_2034_ ),
    .S(\u_multiplier/_3113_ ),
    .Z(\u_multiplier/_2035_ ));
 MUX2_X1 \u_multiplier/_4607_  (.A(\u_multiplier/_3722_ ),
    .B(\u_multiplier/_2035_ ),
    .S(\u_multiplier/_3114_ ),
    .Z(\u_multiplier/_2036_ ));
 MUX2_X1 \u_multiplier/_4608_  (.A(\u_multiplier/_3656_ ),
    .B(\u_multiplier/_2036_ ),
    .S(\u_multiplier/_3112_ ),
    .Z(\u_multiplier/_2037_ ));
 AND2_X1 \u_multiplier/_4609_  (.A1(\u_multiplier/_3115_ ),
    .A2(\u_multiplier/_2037_ ),
    .ZN(\u_multiplier/_2038_ ));
 AOI21_X2 \u_multiplier/_4610_  (.A(\u_multiplier/_2038_ ),
    .B1(\u_multiplier/_3537_ ),
    .B2(\u_multiplier/K [3]),
    .ZN(\u_multiplier/_2039_ ));
 OR2_X1 \u_multiplier/_4611_  (.A1(\u_multiplier/K [4]),
    .A2(\u_multiplier/_2039_ ),
    .ZN(\u_multiplier/_2040_ ));
 NAND3_X1 \u_multiplier/_4612_  (.A1(\u_multiplier/_3115_ ),
    .A2(\u_multiplier/K [4]),
    .A3(\u_multiplier/_3320_ ),
    .ZN(\u_multiplier/_2041_ ));
 AND3_X2 \u_multiplier/_4613_  (.A1(\u_multiplier/_3119_ ),
    .A2(\u_multiplier/_2040_ ),
    .A3(\u_multiplier/_2041_ ),
    .ZN(\u_multiplier/_2042_ ));
 MUX2_X1 \u_multiplier/_4614_  (.A(\u_multiplier/_3262_ ),
    .B(\u_multiplier/_3204_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_2043_ ));
 MUX2_X1 \u_multiplier/_4615_  (.A(\u_multiplier/_2043_ ),
    .B(\u_multiplier/_3728_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_2044_ ));
 MUX2_X1 \u_multiplier/_4616_  (.A(\u_multiplier/_3663_ ),
    .B(\u_multiplier/_2044_ ),
    .S(\u_multiplier/_3110_ ),
    .Z(\u_multiplier/_2045_ ));
 NAND2_X1 \u_multiplier/_4617_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_3543_ ),
    .ZN(\u_multiplier/_2046_ ));
 OAI21_X1 \u_multiplier/_4618_  (.A(\u_multiplier/_2046_ ),
    .B1(\u_multiplier/_2045_ ),
    .B2(\u_multiplier/code_x [3]),
    .ZN(\u_multiplier/_2047_ ));
 MUX2_X1 \u_multiplier/_4619_  (.A(\u_multiplier/_3326_ ),
    .B(\u_multiplier/_2047_ ),
    .S(\u_multiplier/_3109_ ),
    .Z(\u_multiplier/_2048_ ));
 MUX2_X1 \u_multiplier/_4620_  (.A(\u_multiplier/_3206_ ),
    .B(\u_multiplier/_3261_ ),
    .S(\u_multiplier/_3105_ ),
    .Z(\u_multiplier/_2049_ ));
 MUX2_X1 \u_multiplier/_4621_  (.A(\u_multiplier/_2049_ ),
    .B(\u_multiplier/_3734_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_2050_ ));
 MUX2_X1 \u_multiplier/_4622_  (.A(\u_multiplier/_3670_ ),
    .B(\u_multiplier/_2050_ ),
    .S(\u_multiplier/_3106_ ),
    .Z(\u_multiplier/_2051_ ));
 NAND2_X1 \u_multiplier/_4623_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_3550_ ),
    .ZN(\u_multiplier/_2052_ ));
 OAI21_X1 \u_multiplier/_4624_  (.A(\u_multiplier/_2052_ ),
    .B1(\u_multiplier/_2051_ ),
    .B2(\u_multiplier/code_y [3]),
    .ZN(\u_multiplier/_2053_ ));
 MUX2_X2 \u_multiplier/_4625_  (.A(\u_multiplier/_3329_ ),
    .B(\u_multiplier/_2053_ ),
    .S(\u_multiplier/_3108_ ),
    .Z(\u_multiplier/_2054_ ));
 NOR2_X1 \u_multiplier/_4626_  (.A1(\u_multiplier/_2048_ ),
    .A2(\u_multiplier/_2054_ ),
    .ZN(\u_multiplier/_2055_ ));
 XNOR2_X2 \u_multiplier/_4627_  (.A(\u_multiplier/_2048_ ),
    .B(\u_multiplier/_2054_ ),
    .ZN(\u_multiplier/_2056_ ));
 NOR2_X1 \u_multiplier/_4628_  (.A1(\u_multiplier/_2042_ ),
    .A2(\u_multiplier/_2056_ ),
    .ZN(\u_multiplier/_2057_ ));
 XNOR2_X2 \u_multiplier/_4629_  (.A(\u_multiplier/_2042_ ),
    .B(\u_multiplier/_2056_ ),
    .ZN(\u_multiplier/_2058_ ));
 OR2_X1 \u_multiplier/_4630_  (.A1(\u_multiplier/_2033_ ),
    .A2(\u_multiplier/_2058_ ),
    .ZN(\u_multiplier/_2059_ ));
 XOR2_X2 \u_multiplier/_4631_  (.A(\u_multiplier/_2033_ ),
    .B(\u_multiplier/_2058_ ),
    .Z(\u_multiplier/_2060_ ));
 INV_X1 \u_multiplier/_4632_  (.A(\u_multiplier/_2060_ ),
    .ZN(\u_multiplier/_2061_ ));
 NAND2_X1 \u_multiplier/_4633_  (.A1(\u_multiplier/_2032_ ),
    .A2(\u_multiplier/_2060_ ),
    .ZN(\u_multiplier/_2062_ ));
 OAI21_X2 \u_multiplier/_4634_  (.A(net21),
    .B1(\u_multiplier/_2032_ ),
    .B2(\u_multiplier/_2060_ ),
    .ZN(\u_multiplier/_2063_ ));
 AOI21_X4 \u_multiplier/_4635_  (.A(\u_multiplier/_2063_ ),
    .B1(\u_multiplier/_2060_ ),
    .B2(\u_multiplier/_2032_ ),
    .ZN(product[16]));
 NOR2_X1 \u_multiplier/_4636_  (.A1(\u_multiplier/_2055_ ),
    .A2(\u_multiplier/_2057_ ),
    .ZN(\u_multiplier/_2064_ ));
 MUX2_X1 \u_multiplier/_4637_  (.A(\u_multiplier/_3257_ ),
    .B(\u_multiplier/_3255_ ),
    .S(net17),
    .Z(\u_multiplier/_2065_ ));
 AND2_X1 \u_multiplier/_4638_  (.A1(\u_multiplier/_3113_ ),
    .A2(\u_multiplier/_2065_ ),
    .ZN(\u_multiplier/_2066_ ));
 AOI21_X1 \u_multiplier/_4639_  (.A(\u_multiplier/_2066_ ),
    .B1(\u_multiplier/_2034_ ),
    .B2(\u_multiplier/K [0]),
    .ZN(\u_multiplier/_2067_ ));
 MUX2_X1 \u_multiplier/_4640_  (.A(\u_multiplier/_2004_ ),
    .B(\u_multiplier/_2067_ ),
    .S(\u_multiplier/_3114_ ),
    .Z(\u_multiplier/_2068_ ));
 NOR2_X1 \u_multiplier/_4641_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/_2068_ ),
    .ZN(\u_multiplier/_2069_ ));
 AOI21_X2 \u_multiplier/_4642_  (.A(\u_multiplier/_2069_ ),
    .B1(\u_multiplier/_3687_ ),
    .B2(\u_multiplier/K [2]),
    .ZN(\u_multiplier/_2070_ ));
 MUX2_X1 \u_multiplier/_4643_  (.A(\u_multiplier/_3567_ ),
    .B(\u_multiplier/_2070_ ),
    .S(\u_multiplier/_3115_ ),
    .Z(\u_multiplier/_2071_ ));
 AOI21_X1 \u_multiplier/_4644_  (.A(\u_multiplier/dec_out [17]),
    .B1(\u_multiplier/_3341_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2072_ ));
 OAI21_X2 \u_multiplier/_4645_  (.A(\u_multiplier/_2072_ ),
    .B1(\u_multiplier/_2071_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2073_ ));
 MUX2_X1 \u_multiplier/_4646_  (.A(\u_multiplier/_3257_ ),
    .B(\u_multiplier/_3262_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_2074_ ));
 MUX2_X1 \u_multiplier/_4647_  (.A(\u_multiplier/_2074_ ),
    .B(\u_multiplier/_2011_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_2075_ ));
 MUX2_X1 \u_multiplier/_4648_  (.A(\u_multiplier/_3696_ ),
    .B(\u_multiplier/_2075_ ),
    .S(\u_multiplier/_3110_ ),
    .Z(\u_multiplier/_2076_ ));
 NOR2_X1 \u_multiplier/_4649_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_2076_ ),
    .ZN(\u_multiplier/_2077_ ));
 AOI21_X2 \u_multiplier/_4650_  (.A(\u_multiplier/_2077_ ),
    .B1(\u_multiplier/_3574_ ),
    .B2(\u_multiplier/code_x [3]),
    .ZN(\u_multiplier/_2078_ ));
 NOR2_X1 \u_multiplier/_4651_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2078_ ),
    .ZN(\u_multiplier/_2079_ ));
 AOI21_X1 \u_multiplier/_4652_  (.A(\u_multiplier/_3109_ ),
    .B1(\u_multiplier/_3111_ ),
    .B2(\u_multiplier/_3345_ ),
    .ZN(\u_multiplier/_2080_ ));
 NOR2_X1 \u_multiplier/_4653_  (.A1(\u_multiplier/_2079_ ),
    .A2(\u_multiplier/_2080_ ),
    .ZN(\u_multiplier/_2081_ ));
 MUX2_X1 \u_multiplier/_4654_  (.A(\u_multiplier/_3255_ ),
    .B(\u_multiplier/_3261_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_2082_ ));
 MUX2_X1 \u_multiplier/_4655_  (.A(\u_multiplier/_2082_ ),
    .B(\u_multiplier/_2017_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_2083_ ));
 MUX2_X1 \u_multiplier/_4656_  (.A(\u_multiplier/_3703_ ),
    .B(\u_multiplier/_2083_ ),
    .S(\u_multiplier/_3106_ ),
    .Z(\u_multiplier/_2084_ ));
 NAND2_X1 \u_multiplier/_4657_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_3581_ ),
    .ZN(\u_multiplier/_2085_ ));
 OAI21_X1 \u_multiplier/_4658_  (.A(\u_multiplier/_2085_ ),
    .B1(\u_multiplier/_2084_ ),
    .B2(\u_multiplier/code_y [3]),
    .ZN(\u_multiplier/_2086_ ));
 MUX2_X1 \u_multiplier/_4659_  (.A(\u_multiplier/_3350_ ),
    .B(\u_multiplier/_2086_ ),
    .S(\u_multiplier/_3108_ ),
    .Z(\u_multiplier/_2087_ ));
 OR3_X1 \u_multiplier/_4660_  (.A1(\u_multiplier/_2079_ ),
    .A2(\u_multiplier/_2080_ ),
    .A3(\u_multiplier/_2087_ ),
    .ZN(\u_multiplier/_2088_ ));
 XNOR2_X2 \u_multiplier/_4661_  (.A(\u_multiplier/_2081_ ),
    .B(\u_multiplier/_2087_ ),
    .ZN(\u_multiplier/_2089_ ));
 NAND2_X1 \u_multiplier/_4662_  (.A1(\u_multiplier/_2073_ ),
    .A2(\u_multiplier/_2089_ ),
    .ZN(\u_multiplier/_2090_ ));
 XNOR2_X2 \u_multiplier/_4663_  (.A(\u_multiplier/_2073_ ),
    .B(\u_multiplier/_2089_ ),
    .ZN(\u_multiplier/_2091_ ));
 OR2_X1 \u_multiplier/_4664_  (.A1(\u_multiplier/_2064_ ),
    .A2(\u_multiplier/_2091_ ),
    .ZN(\u_multiplier/_2092_ ));
 INV_X1 \u_multiplier/_4665_  (.A(\u_multiplier/_2092_ ),
    .ZN(\u_multiplier/_2093_ ));
 XOR2_X1 \u_multiplier/_4666_  (.A(\u_multiplier/_2064_ ),
    .B(\u_multiplier/_2091_ ),
    .Z(\u_multiplier/_2094_ ));
 INV_X1 \u_multiplier/_4667_  (.A(\u_multiplier/_2094_ ),
    .ZN(\u_multiplier/_2095_ ));
 NOR2_X1 \u_multiplier/_4668_  (.A1(\u_multiplier/_2059_ ),
    .A2(\u_multiplier/_2095_ ),
    .ZN(\u_multiplier/_2096_ ));
 AOI211_X2 \u_multiplier/_4669_  (.A(\u_multiplier/_2061_ ),
    .B(\u_multiplier/_2095_ ),
    .C1(\u_multiplier/_2029_ ),
    .C2(\u_multiplier/_2031_ ),
    .ZN(\u_multiplier/_2097_ ));
 NOR2_X1 \u_multiplier/_4670_  (.A1(\u_multiplier/_2096_ ),
    .A2(\u_multiplier/_2097_ ),
    .ZN(\u_multiplier/_2098_ ));
 NAND3_X1 \u_multiplier/_4671_  (.A1(\u_multiplier/_2059_ ),
    .A2(\u_multiplier/_2062_ ),
    .A3(\u_multiplier/_2095_ ),
    .ZN(\u_multiplier/_2099_ ));
 AND3_X2 \u_multiplier/_4672_  (.A1(net21),
    .A2(\u_multiplier/_2098_ ),
    .A3(\u_multiplier/_2099_ ),
    .ZN(product[17]));
 NAND2_X1 \u_multiplier/_4673_  (.A1(\u_multiplier/_2088_ ),
    .A2(\u_multiplier/_2090_ ),
    .ZN(\u_multiplier/_2100_ ));
 MUX2_X1 \u_multiplier/_4674_  (.A(\u_multiplier/_3250_ ),
    .B(\u_multiplier/_3252_ ),
    .S(net17),
    .Z(\u_multiplier/_2101_ ));
 MUX2_X1 \u_multiplier/_4675_  (.A(\u_multiplier/_2065_ ),
    .B(\u_multiplier/_2101_ ),
    .S(\u_multiplier/_3113_ ),
    .Z(\u_multiplier/_2102_ ));
 MUX2_X1 \u_multiplier/_4676_  (.A(\u_multiplier/_2035_ ),
    .B(\u_multiplier/_2102_ ),
    .S(\u_multiplier/_3114_ ),
    .Z(\u_multiplier/_2103_ ));
 MUX2_X1 \u_multiplier/_4677_  (.A(\u_multiplier/_3723_ ),
    .B(\u_multiplier/_2103_ ),
    .S(\u_multiplier/_3112_ ),
    .Z(\u_multiplier/_2104_ ));
 AND2_X1 \u_multiplier/_4678_  (.A1(\u_multiplier/K [3]),
    .A2(\u_multiplier/_3599_ ),
    .ZN(\u_multiplier/_2105_ ));
 AOI21_X1 \u_multiplier/_4679_  (.A(\u_multiplier/_2105_ ),
    .B1(\u_multiplier/_2104_ ),
    .B2(\u_multiplier/_3115_ ),
    .ZN(\u_multiplier/_2106_ ));
 NOR4_X2 \u_multiplier/_4680_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/K [3]),
    .A3(\u_multiplier/_3116_ ),
    .A4(\u_multiplier/_3360_ ),
    .ZN(\u_multiplier/_2107_ ));
 OAI21_X1 \u_multiplier/_4681_  (.A(\u_multiplier/_3120_ ),
    .B1(\u_multiplier/_2106_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2108_ ));
 NOR2_X1 \u_multiplier/_4682_  (.A1(\u_multiplier/_2107_ ),
    .A2(\u_multiplier/_2108_ ),
    .ZN(\u_multiplier/_2109_ ));
 MUX2_X1 \u_multiplier/_4683_  (.A(\u_multiplier/_3250_ ),
    .B(\u_multiplier/_3257_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_2110_ ));
 MUX2_X1 \u_multiplier/_4684_  (.A(\u_multiplier/_2110_ ),
    .B(\u_multiplier/_2043_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_2111_ ));
 OR2_X1 \u_multiplier/_4685_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_2111_ ),
    .ZN(\u_multiplier/_2112_ ));
 OAI21_X1 \u_multiplier/_4686_  (.A(\u_multiplier/_2112_ ),
    .B1(\u_multiplier/_3729_ ),
    .B2(\u_multiplier/_3110_ ),
    .ZN(\u_multiplier/_2113_ ));
 MUX2_X1 \u_multiplier/_4687_  (.A(\u_multiplier/_3605_ ),
    .B(\u_multiplier/_2113_ ),
    .S(\u_multiplier/_3111_ ),
    .Z(\u_multiplier/_2114_ ));
 AND2_X1 \u_multiplier/_4688_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_3366_ ),
    .ZN(\u_multiplier/_2115_ ));
 AOI21_X2 \u_multiplier/_4689_  (.A(\u_multiplier/_2115_ ),
    .B1(\u_multiplier/_2114_ ),
    .B2(\u_multiplier/_3109_ ),
    .ZN(\u_multiplier/_2116_ ));
 MUX2_X1 \u_multiplier/_4690_  (.A(\u_multiplier/_3252_ ),
    .B(\u_multiplier/_3255_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_2117_ ));
 MUX2_X1 \u_multiplier/_4691_  (.A(\u_multiplier/_2117_ ),
    .B(\u_multiplier/_2049_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_2118_ ));
 OR2_X1 \u_multiplier/_4692_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_2118_ ),
    .ZN(\u_multiplier/_2119_ ));
 OAI21_X1 \u_multiplier/_4693_  (.A(\u_multiplier/_2119_ ),
    .B1(\u_multiplier/_3735_ ),
    .B2(\u_multiplier/_3106_ ),
    .ZN(\u_multiplier/_2120_ ));
 MUX2_X1 \u_multiplier/_4694_  (.A(\u_multiplier/_3610_ ),
    .B(\u_multiplier/_2120_ ),
    .S(\u_multiplier/_3107_ ),
    .Z(\u_multiplier/_2121_ ));
 AND2_X1 \u_multiplier/_4695_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_3371_ ),
    .ZN(\u_multiplier/_2122_ ));
 AOI21_X2 \u_multiplier/_4696_  (.A(\u_multiplier/_2122_ ),
    .B1(\u_multiplier/_2121_ ),
    .B2(\u_multiplier/_3108_ ),
    .ZN(\u_multiplier/_2123_ ));
 NAND2_X1 \u_multiplier/_4697_  (.A1(\u_multiplier/_2116_ ),
    .A2(\u_multiplier/_2123_ ),
    .ZN(\u_multiplier/_2124_ ));
 XOR2_X2 \u_multiplier/_4698_  (.A(\u_multiplier/_2116_ ),
    .B(\u_multiplier/_2123_ ),
    .Z(\u_multiplier/_2125_ ));
 OAI21_X2 \u_multiplier/_4699_  (.A(\u_multiplier/_2125_ ),
    .B1(\u_multiplier/_2108_ ),
    .B2(\u_multiplier/_2107_ ),
    .ZN(\u_multiplier/_2126_ ));
 XOR2_X2 \u_multiplier/_4700_  (.A(\u_multiplier/_2109_ ),
    .B(\u_multiplier/_2125_ ),
    .Z(\u_multiplier/_2127_ ));
 AOI21_X2 \u_multiplier/_4701_  (.A(\u_multiplier/_2127_ ),
    .B1(\u_multiplier/_2090_ ),
    .B2(\u_multiplier/_2088_ ),
    .ZN(\u_multiplier/_2128_ ));
 XOR2_X2 \u_multiplier/_4702_  (.A(\u_multiplier/_2100_ ),
    .B(\u_multiplier/_2127_ ),
    .Z(\u_multiplier/_2129_ ));
 INV_X1 \u_multiplier/_4703_  (.A(\u_multiplier/_2129_ ),
    .ZN(\u_multiplier/_2130_ ));
 OR3_X2 \u_multiplier/_4704_  (.A1(\u_multiplier/_2093_ ),
    .A2(\u_multiplier/_2096_ ),
    .A3(\u_multiplier/_2097_ ),
    .ZN(\u_multiplier/_2131_ ));
 AND2_X1 \u_multiplier/_4705_  (.A1(\u_multiplier/_2130_ ),
    .A2(\u_multiplier/_2131_ ),
    .ZN(\u_multiplier/_2132_ ));
 OAI21_X1 \u_multiplier/_4706_  (.A(\u_multiplier/_3333_ ),
    .B1(\u_multiplier/_2130_ ),
    .B2(\u_multiplier/_2131_ ),
    .ZN(\u_multiplier/_2133_ ));
 NOR2_X1 \u_multiplier/_4707_  (.A1(\u_multiplier/_2132_ ),
    .A2(\u_multiplier/_2133_ ),
    .ZN(product[18]));
 NOR2_X1 \u_multiplier/_4708_  (.A1(\u_multiplier/_2128_ ),
    .A2(\u_multiplier/_2132_ ),
    .ZN(\u_multiplier/_2134_ ));
 MUX2_X1 \u_multiplier/_4709_  (.A(\u_multiplier/_3248_ ),
    .B(\u_multiplier/_3246_ ),
    .S(net17),
    .Z(\u_multiplier/_2135_ ));
 MUX2_X1 \u_multiplier/_4710_  (.A(\u_multiplier/_2101_ ),
    .B(\u_multiplier/_2135_ ),
    .S(\u_multiplier/_3113_ ),
    .Z(\u_multiplier/_2136_ ));
 NAND2_X1 \u_multiplier/_4711_  (.A1(\u_multiplier/K [1]),
    .A2(\u_multiplier/_2067_ ),
    .ZN(\u_multiplier/_2137_ ));
 OAI21_X1 \u_multiplier/_4712_  (.A(\u_multiplier/_2137_ ),
    .B1(\u_multiplier/_2136_ ),
    .B2(\u_multiplier/K [1]),
    .ZN(\u_multiplier/_2138_ ));
 NOR2_X1 \u_multiplier/_4713_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/_2138_ ),
    .ZN(\u_multiplier/_2139_ ));
 AOI21_X2 \u_multiplier/_4714_  (.A(\u_multiplier/_2139_ ),
    .B1(\u_multiplier/_2006_ ),
    .B2(\u_multiplier/K [2]),
    .ZN(\u_multiplier/_2140_ ));
 NOR2_X1 \u_multiplier/_4715_  (.A1(\u_multiplier/K [3]),
    .A2(\u_multiplier/_2140_ ),
    .ZN(\u_multiplier/_2141_ ));
 AOI21_X2 \u_multiplier/_4716_  (.A(\u_multiplier/_2141_ ),
    .B1(\u_multiplier/_3627_ ),
    .B2(\u_multiplier/K [3]),
    .ZN(\u_multiplier/_2142_ ));
 NOR2_X1 \u_multiplier/_4717_  (.A1(\u_multiplier/K [4]),
    .A2(\u_multiplier/_2142_ ),
    .ZN(\u_multiplier/_2143_ ));
 AOI211_X2 \u_multiplier/_4718_  (.A(\u_multiplier/dec_out [19]),
    .B(\u_multiplier/_2143_ ),
    .C1(\u_multiplier/_3391_ ),
    .C2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2144_ ));
 MUX2_X1 \u_multiplier/_4719_  (.A(\u_multiplier/_3248_ ),
    .B(\u_multiplier/_3250_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_2145_ ));
 MUX2_X1 \u_multiplier/_4720_  (.A(\u_multiplier/_2145_ ),
    .B(\u_multiplier/_2074_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_2146_ ));
 MUX2_X1 \u_multiplier/_4721_  (.A(\u_multiplier/_2012_ ),
    .B(\u_multiplier/_2146_ ),
    .S(\u_multiplier/_3110_ ),
    .Z(\u_multiplier/_2147_ ));
 MUX2_X1 \u_multiplier/_4722_  (.A(\u_multiplier/_3632_ ),
    .B(\u_multiplier/_2147_ ),
    .S(\u_multiplier/_3111_ ),
    .Z(\u_multiplier/_2148_ ));
 NOR2_X1 \u_multiplier/_4723_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2148_ ),
    .ZN(\u_multiplier/_2149_ ));
 AOI21_X2 \u_multiplier/_4724_  (.A(\u_multiplier/_2149_ ),
    .B1(\u_multiplier/_3396_ ),
    .B2(\u_multiplier/code_x [4]),
    .ZN(\u_multiplier/_2150_ ));
 MUX2_X1 \u_multiplier/_4725_  (.A(\u_multiplier/_3246_ ),
    .B(\u_multiplier/_3252_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_2151_ ));
 MUX2_X1 \u_multiplier/_4726_  (.A(\u_multiplier/_2151_ ),
    .B(\u_multiplier/_2082_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_2152_ ));
 MUX2_X1 \u_multiplier/_4727_  (.A(\u_multiplier/_2018_ ),
    .B(\u_multiplier/_2152_ ),
    .S(\u_multiplier/_3106_ ),
    .Z(\u_multiplier/_2153_ ));
 NOR2_X1 \u_multiplier/_4728_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_2153_ ),
    .ZN(\u_multiplier/_2154_ ));
 AOI21_X2 \u_multiplier/_4729_  (.A(\u_multiplier/_2154_ ),
    .B1(\u_multiplier/_3639_ ),
    .B2(\u_multiplier/code_y [3]),
    .ZN(\u_multiplier/_2155_ ));
 NAND2_X1 \u_multiplier/_4730_  (.A1(\u_multiplier/_3108_ ),
    .A2(\u_multiplier/_2155_ ),
    .ZN(\u_multiplier/_2156_ ));
 OAI21_X1 \u_multiplier/_4731_  (.A(\u_multiplier/_2156_ ),
    .B1(\u_multiplier/_3400_ ),
    .B2(\u_multiplier/_3108_ ),
    .ZN(\u_multiplier/_2157_ ));
 XOR2_X1 \u_multiplier/_4732_  (.A(\u_multiplier/_2150_ ),
    .B(\u_multiplier/_2157_ ),
    .Z(\u_multiplier/_2158_ ));
 INV_X1 \u_multiplier/_4733_  (.A(\u_multiplier/_2158_ ),
    .ZN(\u_multiplier/_2159_ ));
 NOR2_X1 \u_multiplier/_4734_  (.A1(\u_multiplier/_2144_ ),
    .A2(\u_multiplier/_2159_ ),
    .ZN(\u_multiplier/_2160_ ));
 XNOR2_X1 \u_multiplier/_4735_  (.A(\u_multiplier/_2144_ ),
    .B(\u_multiplier/_2159_ ),
    .ZN(\u_multiplier/_2161_ ));
 AOI21_X2 \u_multiplier/_4736_  (.A(\u_multiplier/_2161_ ),
    .B1(\u_multiplier/_2126_ ),
    .B2(\u_multiplier/_2124_ ),
    .ZN(\u_multiplier/_2162_ ));
 AND3_X2 \u_multiplier/_4737_  (.A1(\u_multiplier/_2124_ ),
    .A2(\u_multiplier/_2126_ ),
    .A3(\u_multiplier/_2161_ ),
    .ZN(\u_multiplier/_2163_ ));
 OR2_X1 \u_multiplier/_4738_  (.A1(\u_multiplier/_2162_ ),
    .A2(\u_multiplier/_2163_ ),
    .ZN(\u_multiplier/_2164_ ));
 OAI21_X1 \u_multiplier/_4739_  (.A(\u_multiplier/_3333_ ),
    .B1(\u_multiplier/_2134_ ),
    .B2(\u_multiplier/_2164_ ),
    .ZN(\u_multiplier/_2165_ ));
 AOI21_X1 \u_multiplier/_4740_  (.A(\u_multiplier/_2165_ ),
    .B1(\u_multiplier/_2164_ ),
    .B2(\u_multiplier/_2134_ ),
    .ZN(product[19]));
 AOI21_X2 \u_multiplier/_4741_  (.A(\u_multiplier/_2160_ ),
    .B1(\u_multiplier/_2157_ ),
    .B2(\u_multiplier/_2150_ ),
    .ZN(\u_multiplier/_2166_ ));
 MUX2_X1 \u_multiplier/_4742_  (.A(\u_multiplier/_3241_ ),
    .B(\u_multiplier/_3240_ ),
    .S(\u_multiplier/_3313_ ),
    .Z(\u_multiplier/_2167_ ));
 MUX2_X1 \u_multiplier/_4743_  (.A(\u_multiplier/_2135_ ),
    .B(\u_multiplier/_2167_ ),
    .S(\u_multiplier/_3113_ ),
    .Z(\u_multiplier/_2168_ ));
 MUX2_X1 \u_multiplier/_4744_  (.A(\u_multiplier/_2102_ ),
    .B(\u_multiplier/_2168_ ),
    .S(\u_multiplier/_3114_ ),
    .Z(\u_multiplier/_2169_ ));
 MUX2_X1 \u_multiplier/_4745_  (.A(\u_multiplier/_2036_ ),
    .B(\u_multiplier/_2169_ ),
    .S(\u_multiplier/_3112_ ),
    .Z(\u_multiplier/_2170_ ));
 AND2_X1 \u_multiplier/_4746_  (.A1(\u_multiplier/_3115_ ),
    .A2(\u_multiplier/_2170_ ),
    .ZN(\u_multiplier/_2171_ ));
 AOI21_X4 \u_multiplier/_4747_  (.A(\u_multiplier/_2171_ ),
    .B1(\u_multiplier/_3657_ ),
    .B2(\u_multiplier/K [3]),
    .ZN(\u_multiplier/_2172_ ));
 AOI21_X2 \u_multiplier/_4748_  (.A(\u_multiplier/dec_out [20]),
    .B1(\u_multiplier/_3416_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2173_ ));
 OAI21_X4 \u_multiplier/_4749_  (.A(\u_multiplier/_2173_ ),
    .B1(\u_multiplier/_2172_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2174_ ));
 MUX2_X1 \u_multiplier/_4750_  (.A(\u_multiplier/_3241_ ),
    .B(\u_multiplier/_3248_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_2175_ ));
 MUX2_X1 \u_multiplier/_4751_  (.A(\u_multiplier/_2175_ ),
    .B(\u_multiplier/_2110_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_2176_ ));
 OR2_X1 \u_multiplier/_4752_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_2176_ ),
    .ZN(\u_multiplier/_2177_ ));
 OAI21_X1 \u_multiplier/_4753_  (.A(\u_multiplier/_2177_ ),
    .B1(\u_multiplier/_2044_ ),
    .B2(\u_multiplier/_3110_ ),
    .ZN(\u_multiplier/_2178_ ));
 MUX2_X1 \u_multiplier/_4754_  (.A(\u_multiplier/_3665_ ),
    .B(\u_multiplier/_2178_ ),
    .S(\u_multiplier/_3111_ ),
    .Z(\u_multiplier/_2179_ ));
 MUX2_X1 \u_multiplier/_4755_  (.A(\u_multiplier/_3422_ ),
    .B(\u_multiplier/_2179_ ),
    .S(\u_multiplier/_3109_ ),
    .Z(\u_multiplier/_2180_ ));
 MUX2_X1 \u_multiplier/_4756_  (.A(\u_multiplier/_3240_ ),
    .B(\u_multiplier/_3246_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_2181_ ));
 MUX2_X1 \u_multiplier/_4757_  (.A(\u_multiplier/_2181_ ),
    .B(\u_multiplier/_2117_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_2182_ ));
 OR2_X1 \u_multiplier/_4758_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_2182_ ),
    .ZN(\u_multiplier/_2183_ ));
 OAI21_X2 \u_multiplier/_4759_  (.A(\u_multiplier/_2183_ ),
    .B1(\u_multiplier/_2050_ ),
    .B2(\u_multiplier/_3106_ ),
    .ZN(\u_multiplier/_2184_ ));
 MUX2_X1 \u_multiplier/_4760_  (.A(\u_multiplier/_3672_ ),
    .B(\u_multiplier/_2184_ ),
    .S(\u_multiplier/_3107_ ),
    .Z(\u_multiplier/_2185_ ));
 MUX2_X1 \u_multiplier/_4761_  (.A(\u_multiplier/_3429_ ),
    .B(\u_multiplier/_2185_ ),
    .S(\u_multiplier/_3108_ ),
    .Z(\u_multiplier/_2186_ ));
 NOR2_X1 \u_multiplier/_4762_  (.A1(\u_multiplier/_2180_ ),
    .A2(\u_multiplier/_2186_ ),
    .ZN(\u_multiplier/_2187_ ));
 XNOR2_X1 \u_multiplier/_4763_  (.A(\u_multiplier/_2180_ ),
    .B(\u_multiplier/_2186_ ),
    .ZN(\u_multiplier/_2188_ ));
 INV_X2 \u_multiplier/_4764_  (.A(\u_multiplier/_2188_ ),
    .ZN(\u_multiplier/_2189_ ));
 XNOR2_X2 \u_multiplier/_4765_  (.A(\u_multiplier/_2174_ ),
    .B(\u_multiplier/_2189_ ),
    .ZN(\u_multiplier/_2190_ ));
 NOR2_X1 \u_multiplier/_4766_  (.A1(\u_multiplier/_2166_ ),
    .A2(\u_multiplier/_2190_ ),
    .ZN(\u_multiplier/_2191_ ));
 XNOR2_X2 \u_multiplier/_4767_  (.A(\u_multiplier/_2166_ ),
    .B(\u_multiplier/_2190_ ),
    .ZN(\u_multiplier/_2192_ ));
 AOI211_X2 \u_multiplier/_4768_  (.A(\u_multiplier/_2128_ ),
    .B(\u_multiplier/_2162_ ),
    .C1(\u_multiplier/_2131_ ),
    .C2(\u_multiplier/_2130_ ),
    .ZN(\u_multiplier/_2193_ ));
 NOR3_X2 \u_multiplier/_4769_  (.A1(\u_multiplier/_2163_ ),
    .A2(\u_multiplier/_2192_ ),
    .A3(\u_multiplier/_2193_ ),
    .ZN(\u_multiplier/_2194_ ));
 OAI21_X1 \u_multiplier/_4770_  (.A(\u_multiplier/_2192_ ),
    .B1(\u_multiplier/_2193_ ),
    .B2(\u_multiplier/_2163_ ),
    .ZN(\u_multiplier/_2195_ ));
 NAND2_X1 \u_multiplier/_4771_  (.A1(\u_multiplier/_3333_ ),
    .A2(\u_multiplier/_2195_ ),
    .ZN(\u_multiplier/_2196_ ));
 NOR2_X2 \u_multiplier/_4772_  (.A1(\u_multiplier/_2194_ ),
    .A2(\u_multiplier/_2196_ ),
    .ZN(product[20]));
 AOI21_X4 \u_multiplier/_4773_  (.A(\u_multiplier/_2187_ ),
    .B1(\u_multiplier/_2189_ ),
    .B2(\u_multiplier/_2174_ ),
    .ZN(\u_multiplier/_2197_ ));
 MUX2_X1 \u_multiplier/_4774_  (.A(\u_multiplier/_3238_ ),
    .B(\u_multiplier/_3236_ ),
    .S(\u_multiplier/_3313_ ),
    .Z(\u_multiplier/_2198_ ));
 MUX2_X1 \u_multiplier/_4775_  (.A(\u_multiplier/_2167_ ),
    .B(\u_multiplier/_2198_ ),
    .S(\u_multiplier/_3113_ ),
    .Z(\u_multiplier/_2199_ ));
 MUX2_X1 \u_multiplier/_4776_  (.A(\u_multiplier/_2136_ ),
    .B(\u_multiplier/_2199_ ),
    .S(\u_multiplier/_3114_ ),
    .Z(\u_multiplier/_2200_ ));
 NAND2_X1 \u_multiplier/_4777_  (.A1(\u_multiplier/_3112_ ),
    .A2(\u_multiplier/_2200_ ),
    .ZN(\u_multiplier/_2201_ ));
 OAI21_X1 \u_multiplier/_4778_  (.A(\u_multiplier/_2201_ ),
    .B1(\u_multiplier/_2068_ ),
    .B2(\u_multiplier/_3112_ ),
    .ZN(\u_multiplier/_2202_ ));
 MUX2_X1 \u_multiplier/_4779_  (.A(\u_multiplier/_3689_ ),
    .B(\u_multiplier/_2202_ ),
    .S(\u_multiplier/_3115_ ),
    .Z(\u_multiplier/_2203_ ));
 AND2_X1 \u_multiplier/_4780_  (.A1(\u_multiplier/_3116_ ),
    .A2(\u_multiplier/_2203_ ),
    .ZN(\u_multiplier/_2204_ ));
 AOI211_X2 \u_multiplier/_4781_  (.A(\u_multiplier/dec_out [21]),
    .B(\u_multiplier/_2204_ ),
    .C1(\u_multiplier/_3447_ ),
    .C2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2205_ ));
 MUX2_X1 \u_multiplier/_4782_  (.A(\u_multiplier/_3238_ ),
    .B(\u_multiplier/_3241_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_2206_ ));
 MUX2_X1 \u_multiplier/_4783_  (.A(\u_multiplier/_2206_ ),
    .B(\u_multiplier/_2145_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_2207_ ));
 OR2_X1 \u_multiplier/_4784_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_2207_ ),
    .ZN(\u_multiplier/_2208_ ));
 OAI21_X1 \u_multiplier/_4785_  (.A(\u_multiplier/_2208_ ),
    .B1(\u_multiplier/_2075_ ),
    .B2(\u_multiplier/_3110_ ),
    .ZN(\u_multiplier/_2209_ ));
 MUX2_X1 \u_multiplier/_4786_  (.A(\u_multiplier/_3698_ ),
    .B(\u_multiplier/_2209_ ),
    .S(\u_multiplier/_3111_ ),
    .Z(\u_multiplier/_2210_ ));
 MUX2_X1 \u_multiplier/_4787_  (.A(\u_multiplier/_3454_ ),
    .B(\u_multiplier/_2210_ ),
    .S(\u_multiplier/_3109_ ),
    .Z(\u_multiplier/_2211_ ));
 MUX2_X1 \u_multiplier/_4788_  (.A(\u_multiplier/_3236_ ),
    .B(\u_multiplier/_3240_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_2212_ ));
 MUX2_X1 \u_multiplier/_4789_  (.A(\u_multiplier/_2212_ ),
    .B(\u_multiplier/_2151_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_2213_ ));
 MUX2_X1 \u_multiplier/_4790_  (.A(\u_multiplier/_2083_ ),
    .B(\u_multiplier/_2213_ ),
    .S(\u_multiplier/_3106_ ),
    .Z(\u_multiplier/_2214_ ));
 NAND2_X1 \u_multiplier/_4791_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_3705_ ),
    .ZN(\u_multiplier/_2215_ ));
 OAI21_X2 \u_multiplier/_4792_  (.A(\u_multiplier/_2215_ ),
    .B1(\u_multiplier/_2214_ ),
    .B2(\u_multiplier/code_y [3]),
    .ZN(\u_multiplier/_2216_ ));
 MUX2_X1 \u_multiplier/_4793_  (.A(\u_multiplier/_3462_ ),
    .B(\u_multiplier/_2216_ ),
    .S(\u_multiplier/_3108_ ),
    .Z(\u_multiplier/_2217_ ));
 NOR2_X1 \u_multiplier/_4794_  (.A1(\u_multiplier/_2211_ ),
    .A2(\u_multiplier/_2217_ ),
    .ZN(\u_multiplier/_2218_ ));
 XNOR2_X2 \u_multiplier/_4795_  (.A(\u_multiplier/_2211_ ),
    .B(\u_multiplier/_2217_ ),
    .ZN(\u_multiplier/_2219_ ));
 NOR2_X1 \u_multiplier/_4796_  (.A1(\u_multiplier/_2205_ ),
    .A2(\u_multiplier/_2219_ ),
    .ZN(\u_multiplier/_2220_ ));
 XNOR2_X2 \u_multiplier/_4797_  (.A(\u_multiplier/_2205_ ),
    .B(\u_multiplier/_2219_ ),
    .ZN(\u_multiplier/_2221_ ));
 XOR2_X2 \u_multiplier/_4798_  (.A(\u_multiplier/_2197_ ),
    .B(\u_multiplier/_2221_ ),
    .Z(\u_multiplier/_2222_ ));
 INV_X1 \u_multiplier/_4799_  (.A(\u_multiplier/_2222_ ),
    .ZN(\u_multiplier/_2223_ ));
 OAI21_X1 \u_multiplier/_4800_  (.A(\u_multiplier/_2223_ ),
    .B1(\u_multiplier/_2190_ ),
    .B2(\u_multiplier/_2166_ ),
    .ZN(\u_multiplier/_2224_ ));
 NOR4_X4 \u_multiplier/_4801_  (.A1(\u_multiplier/_2163_ ),
    .A2(\u_multiplier/_2192_ ),
    .A3(\u_multiplier/_2193_ ),
    .A4(\u_multiplier/_2223_ ),
    .ZN(\u_multiplier/_2225_ ));
 NAND2_X2 \u_multiplier/_4802_  (.A1(\u_multiplier/_2191_ ),
    .A2(\u_multiplier/_2222_ ),
    .ZN(\u_multiplier/_2226_ ));
 OAI21_X2 \u_multiplier/_4803_  (.A(\u_multiplier/_2226_ ),
    .B1(\u_multiplier/_2224_ ),
    .B2(\u_multiplier/_2194_ ),
    .ZN(\u_multiplier/_2227_ ));
 NOR3_X4 \u_multiplier/_4804_  (.A1(\u_multiplier/_3334_ ),
    .A2(\u_multiplier/_2225_ ),
    .A3(\u_multiplier/_2227_ ),
    .ZN(product[21]));
 OAI21_X4 \u_multiplier/_4805_  (.A(\u_multiplier/_2226_ ),
    .B1(\u_multiplier/_2221_ ),
    .B2(\u_multiplier/_2197_ ),
    .ZN(\u_multiplier/_2228_ ));
 OR2_X1 \u_multiplier/_4806_  (.A1(\u_multiplier/_2225_ ),
    .A2(\u_multiplier/_2228_ ),
    .ZN(\u_multiplier/_2229_ ));
 NOR2_X2 \u_multiplier/_4807_  (.A1(\u_multiplier/_2218_ ),
    .A2(\u_multiplier/_2220_ ),
    .ZN(\u_multiplier/_2230_ ));
 MUX2_X1 \u_multiplier/_4808_  (.A(\u_multiplier/_3226_ ),
    .B(\u_multiplier/_3227_ ),
    .S(\u_multiplier/_3313_ ),
    .Z(\u_multiplier/_2231_ ));
 MUX2_X1 \u_multiplier/_4809_  (.A(\u_multiplier/_2198_ ),
    .B(\u_multiplier/_2231_ ),
    .S(\u_multiplier/_3113_ ),
    .Z(\u_multiplier/_2232_ ));
 MUX2_X1 \u_multiplier/_4810_  (.A(\u_multiplier/_2168_ ),
    .B(\u_multiplier/_2232_ ),
    .S(\u_multiplier/_3114_ ),
    .Z(\u_multiplier/_2233_ ));
 MUX2_X2 \u_multiplier/_4811_  (.A(\u_multiplier/_2103_ ),
    .B(\u_multiplier/_2233_ ),
    .S(\u_multiplier/_3112_ ),
    .Z(\u_multiplier/_2234_ ));
 NOR2_X1 \u_multiplier/_4812_  (.A1(\u_multiplier/_3115_ ),
    .A2(\u_multiplier/_3725_ ),
    .ZN(\u_multiplier/_2235_ ));
 AOI21_X4 \u_multiplier/_4813_  (.A(\u_multiplier/_2235_ ),
    .B1(\u_multiplier/_2234_ ),
    .B2(\u_multiplier/_3115_ ),
    .ZN(\u_multiplier/_2236_ ));
 AOI21_X1 \u_multiplier/_4814_  (.A(\u_multiplier/dec_out [22]),
    .B1(\u_multiplier/_3479_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2237_ ));
 OAI21_X2 \u_multiplier/_4815_  (.A(\u_multiplier/_2237_ ),
    .B1(\u_multiplier/_2236_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2238_ ));
 MUX2_X1 \u_multiplier/_4816_  (.A(\u_multiplier/_3226_ ),
    .B(\u_multiplier/_3238_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_2239_ ));
 MUX2_X1 \u_multiplier/_4817_  (.A(\u_multiplier/_2239_ ),
    .B(\u_multiplier/_2175_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_2240_ ));
 MUX2_X1 \u_multiplier/_4818_  (.A(\u_multiplier/_2111_ ),
    .B(\u_multiplier/_2240_ ),
    .S(\u_multiplier/_3110_ ),
    .Z(\u_multiplier/_2241_ ));
 NAND2_X1 \u_multiplier/_4819_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_3731_ ),
    .ZN(\u_multiplier/_2242_ ));
 OAI21_X1 \u_multiplier/_4820_  (.A(\u_multiplier/_2242_ ),
    .B1(\u_multiplier/_2241_ ),
    .B2(\u_multiplier/code_x [3]),
    .ZN(\u_multiplier/_2243_ ));
 MUX2_X1 \u_multiplier/_4821_  (.A(\u_multiplier/_3486_ ),
    .B(\u_multiplier/_2243_ ),
    .S(\u_multiplier/_3109_ ),
    .Z(\u_multiplier/_2244_ ));
 MUX2_X1 \u_multiplier/_4822_  (.A(\u_multiplier/_3227_ ),
    .B(\u_multiplier/_3236_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_2245_ ));
 MUX2_X1 \u_multiplier/_4823_  (.A(\u_multiplier/_2245_ ),
    .B(\u_multiplier/_2181_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_2246_ ));
 MUX2_X2 \u_multiplier/_4824_  (.A(\u_multiplier/_2118_ ),
    .B(\u_multiplier/_2246_ ),
    .S(\u_multiplier/_3106_ ),
    .Z(\u_multiplier/_2247_ ));
 NAND2_X1 \u_multiplier/_4825_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_3737_ ),
    .ZN(\u_multiplier/_2248_ ));
 OAI21_X2 \u_multiplier/_4826_  (.A(\u_multiplier/_2248_ ),
    .B1(\u_multiplier/_2247_ ),
    .B2(\u_multiplier/code_y [3]),
    .ZN(\u_multiplier/_2249_ ));
 MUX2_X1 \u_multiplier/_4827_  (.A(\u_multiplier/_3493_ ),
    .B(\u_multiplier/_2249_ ),
    .S(\u_multiplier/_3108_ ),
    .Z(\u_multiplier/_2250_ ));
 NOR2_X1 \u_multiplier/_4828_  (.A1(\u_multiplier/_2244_ ),
    .A2(\u_multiplier/_2250_ ),
    .ZN(\u_multiplier/_2251_ ));
 XNOR2_X1 \u_multiplier/_4829_  (.A(\u_multiplier/_2244_ ),
    .B(\u_multiplier/_2250_ ),
    .ZN(\u_multiplier/_2252_ ));
 INV_X1 \u_multiplier/_4830_  (.A(\u_multiplier/_2252_ ),
    .ZN(\u_multiplier/_2253_ ));
 XNOR2_X2 \u_multiplier/_4831_  (.A(\u_multiplier/_2238_ ),
    .B(\u_multiplier/_2253_ ),
    .ZN(\u_multiplier/_2254_ ));
 OR2_X1 \u_multiplier/_4832_  (.A1(\u_multiplier/_2230_ ),
    .A2(\u_multiplier/_2254_ ),
    .ZN(\u_multiplier/_2255_ ));
 XOR2_X2 \u_multiplier/_4833_  (.A(\u_multiplier/_2230_ ),
    .B(\u_multiplier/_2254_ ),
    .Z(\u_multiplier/_2256_ ));
 NAND2_X1 \u_multiplier/_4834_  (.A1(\u_multiplier/_2229_ ),
    .A2(\u_multiplier/_2256_ ),
    .ZN(\u_multiplier/_2257_ ));
 OAI21_X1 \u_multiplier/_4835_  (.A(net21),
    .B1(\u_multiplier/_2229_ ),
    .B2(\u_multiplier/_2256_ ),
    .ZN(\u_multiplier/_2258_ ));
 AOI21_X1 \u_multiplier/_4836_  (.A(\u_multiplier/_2258_ ),
    .B1(\u_multiplier/_2256_ ),
    .B2(\u_multiplier/_2229_ ),
    .ZN(product[22]));
 AND2_X1 \u_multiplier/_4837_  (.A1(\u_multiplier/_2255_ ),
    .A2(\u_multiplier/_2257_ ),
    .ZN(\u_multiplier/_2259_ ));
 AOI21_X2 \u_multiplier/_4838_  (.A(\u_multiplier/_2251_ ),
    .B1(\u_multiplier/_2253_ ),
    .B2(\u_multiplier/_2238_ ),
    .ZN(\u_multiplier/_2260_ ));
 MUX2_X1 \u_multiplier/_4839_  (.A(\u_multiplier/_3231_ ),
    .B(\u_multiplier/_3229_ ),
    .S(\u_multiplier/_3313_ ),
    .Z(\u_multiplier/_2261_ ));
 MUX2_X1 \u_multiplier/_4840_  (.A(\u_multiplier/_2231_ ),
    .B(\u_multiplier/_2261_ ),
    .S(\u_multiplier/_3113_ ),
    .Z(\u_multiplier/_2262_ ));
 MUX2_X1 \u_multiplier/_4841_  (.A(\u_multiplier/_2199_ ),
    .B(\u_multiplier/_2262_ ),
    .S(\u_multiplier/_3114_ ),
    .Z(\u_multiplier/_2263_ ));
 NAND2_X1 \u_multiplier/_4842_  (.A1(\u_multiplier/_3112_ ),
    .A2(\u_multiplier/_2263_ ),
    .ZN(\u_multiplier/_2264_ ));
 OAI21_X2 \u_multiplier/_4843_  (.A(\u_multiplier/_2264_ ),
    .B1(\u_multiplier/_2138_ ),
    .B2(\u_multiplier/_3112_ ),
    .ZN(\u_multiplier/_2265_ ));
 AND2_X1 \u_multiplier/_4844_  (.A1(\u_multiplier/K [3]),
    .A2(\u_multiplier/_2007_ ),
    .ZN(\u_multiplier/_2266_ ));
 AOI21_X4 \u_multiplier/_4845_  (.A(\u_multiplier/_2266_ ),
    .B1(\u_multiplier/_2265_ ),
    .B2(\u_multiplier/_3115_ ),
    .ZN(\u_multiplier/_2267_ ));
 AOI21_X1 \u_multiplier/_4846_  (.A(\u_multiplier/dec_out [23]),
    .B1(\u_multiplier/_3510_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2268_ ));
 OAI21_X2 \u_multiplier/_4847_  (.A(\u_multiplier/_2268_ ),
    .B1(\u_multiplier/_2267_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2269_ ));
 MUX2_X1 \u_multiplier/_4848_  (.A(\u_multiplier/_3231_ ),
    .B(\u_multiplier/_3226_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_2270_ ));
 MUX2_X1 \u_multiplier/_4849_  (.A(\u_multiplier/_2270_ ),
    .B(\u_multiplier/_2206_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_2271_ ));
 MUX2_X1 \u_multiplier/_4850_  (.A(\u_multiplier/_2146_ ),
    .B(\u_multiplier/_2271_ ),
    .S(\u_multiplier/_3110_ ),
    .Z(\u_multiplier/_2272_ ));
 MUX2_X1 \u_multiplier/_4851_  (.A(\u_multiplier/_2013_ ),
    .B(\u_multiplier/_2272_ ),
    .S(\u_multiplier/_3111_ ),
    .Z(\u_multiplier/_2273_ ));
 NOR2_X1 \u_multiplier/_4852_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2273_ ),
    .ZN(\u_multiplier/_2274_ ));
 AOI21_X2 \u_multiplier/_4853_  (.A(\u_multiplier/_2274_ ),
    .B1(\u_multiplier/_3516_ ),
    .B2(\u_multiplier/code_x [4]),
    .ZN(\u_multiplier/_2275_ ));
 MUX2_X1 \u_multiplier/_4854_  (.A(\u_multiplier/_3227_ ),
    .B(\u_multiplier/_3229_ ),
    .S(\u_multiplier/_3105_ ),
    .Z(\u_multiplier/_2276_ ));
 MUX2_X1 \u_multiplier/_4855_  (.A(\u_multiplier/_2276_ ),
    .B(\u_multiplier/_2212_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_2277_ ));
 MUX2_X1 \u_multiplier/_4856_  (.A(\u_multiplier/_2152_ ),
    .B(\u_multiplier/_2277_ ),
    .S(\u_multiplier/_3106_ ),
    .Z(\u_multiplier/_2278_ ));
 NOR2_X1 \u_multiplier/_4857_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_2278_ ),
    .ZN(\u_multiplier/_2279_ ));
 AOI21_X2 \u_multiplier/_4858_  (.A(\u_multiplier/_2279_ ),
    .B1(\u_multiplier/_2020_ ),
    .B2(\u_multiplier/code_y [3]),
    .ZN(\u_multiplier/_2280_ ));
 NAND2_X1 \u_multiplier/_4859_  (.A1(\u_multiplier/_3108_ ),
    .A2(\u_multiplier/_2280_ ),
    .ZN(\u_multiplier/_2281_ ));
 OAI21_X2 \u_multiplier/_4860_  (.A(\u_multiplier/_2281_ ),
    .B1(\u_multiplier/_3521_ ),
    .B2(\u_multiplier/_3108_ ),
    .ZN(\u_multiplier/_2282_ ));
 NAND2_X1 \u_multiplier/_4861_  (.A1(\u_multiplier/_2275_ ),
    .A2(\u_multiplier/_2282_ ),
    .ZN(\u_multiplier/_2283_ ));
 XOR2_X2 \u_multiplier/_4862_  (.A(\u_multiplier/_2275_ ),
    .B(\u_multiplier/_2282_ ),
    .Z(\u_multiplier/_2284_ ));
 NAND2_X1 \u_multiplier/_4863_  (.A1(\u_multiplier/_2269_ ),
    .A2(\u_multiplier/_2284_ ),
    .ZN(\u_multiplier/_2285_ ));
 XNOR2_X2 \u_multiplier/_4864_  (.A(\u_multiplier/_2269_ ),
    .B(\u_multiplier/_2284_ ),
    .ZN(\u_multiplier/_2286_ ));
 OR2_X1 \u_multiplier/_4865_  (.A1(\u_multiplier/_2260_ ),
    .A2(\u_multiplier/_2286_ ),
    .ZN(\u_multiplier/_2287_ ));
 AND2_X1 \u_multiplier/_4866_  (.A1(\u_multiplier/_2260_ ),
    .A2(\u_multiplier/_2286_ ),
    .ZN(\u_multiplier/_2288_ ));
 XNOR2_X2 \u_multiplier/_4867_  (.A(\u_multiplier/_2260_ ),
    .B(\u_multiplier/_2286_ ),
    .ZN(\u_multiplier/_2289_ ));
 INV_X1 \u_multiplier/_4868_  (.A(\u_multiplier/_2289_ ),
    .ZN(\u_multiplier/_2290_ ));
 OAI21_X1 \u_multiplier/_4869_  (.A(net21),
    .B1(\u_multiplier/_2259_ ),
    .B2(\u_multiplier/_2289_ ),
    .ZN(\u_multiplier/_2291_ ));
 AOI21_X2 \u_multiplier/_4870_  (.A(\u_multiplier/_2291_ ),
    .B1(\u_multiplier/_2289_ ),
    .B2(\u_multiplier/_2259_ ),
    .ZN(product[23]));
 OAI211_X4 \u_multiplier/_4871_  (.A(\u_multiplier/_2256_ ),
    .B(\u_multiplier/_2290_ ),
    .C1(\u_multiplier/_2225_ ),
    .C2(\u_multiplier/_2228_ ),
    .ZN(\u_multiplier/_2292_ ));
 OAI21_X1 \u_multiplier/_4872_  (.A(\u_multiplier/_2287_ ),
    .B1(\u_multiplier/_2288_ ),
    .B2(\u_multiplier/_2255_ ),
    .ZN(\u_multiplier/_2293_ ));
 INV_X2 \u_multiplier/_4873_  (.A(\u_multiplier/_2293_ ),
    .ZN(\u_multiplier/_2294_ ));
 NAND2_X1 \u_multiplier/_4874_  (.A1(\u_multiplier/_2292_ ),
    .A2(\u_multiplier/_2294_ ),
    .ZN(\u_multiplier/_2295_ ));
 NAND2_X1 \u_multiplier/_4875_  (.A1(\u_multiplier/_2283_ ),
    .A2(\u_multiplier/_2285_ ),
    .ZN(\u_multiplier/_2296_ ));
 MUX2_X1 \u_multiplier/_4876_  (.A(\u_multiplier/_3292_ ),
    .B(\u_multiplier/_3291_ ),
    .S(\u_multiplier/_3313_ ),
    .Z(\u_multiplier/_2297_ ));
 MUX2_X1 \u_multiplier/_4877_  (.A(\u_multiplier/_2261_ ),
    .B(\u_multiplier/_2297_ ),
    .S(\u_multiplier/_3113_ ),
    .Z(\u_multiplier/_2298_ ));
 MUX2_X1 \u_multiplier/_4878_  (.A(\u_multiplier/_2232_ ),
    .B(\u_multiplier/_2298_ ),
    .S(\u_multiplier/_3114_ ),
    .Z(\u_multiplier/_2299_ ));
 MUX2_X1 \u_multiplier/_4879_  (.A(\u_multiplier/_2169_ ),
    .B(\u_multiplier/_2299_ ),
    .S(\u_multiplier/_3112_ ),
    .Z(\u_multiplier/_2300_ ));
 MUX2_X2 \u_multiplier/_4880_  (.A(\u_multiplier/_2037_ ),
    .B(\u_multiplier/_2300_ ),
    .S(\u_multiplier/_3115_ ),
    .Z(\u_multiplier/_2301_ ));
 MUX2_X1 \u_multiplier/_4881_  (.A(\u_multiplier/_3538_ ),
    .B(\u_multiplier/_2301_ ),
    .S(\u_multiplier/_3116_ ),
    .Z(\u_multiplier/_2302_ ));
 MUX2_X1 \u_multiplier/_4882_  (.A(\u_multiplier/_3292_ ),
    .B(\u_multiplier/_3231_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_2303_ ));
 MUX2_X1 \u_multiplier/_4883_  (.A(\u_multiplier/_2303_ ),
    .B(\u_multiplier/_2239_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_2304_ ));
 MUX2_X1 \u_multiplier/_4884_  (.A(\u_multiplier/_2176_ ),
    .B(\u_multiplier/_2304_ ),
    .S(\u_multiplier/_3110_ ),
    .Z(\u_multiplier/_2305_ ));
 MUX2_X1 \u_multiplier/_4885_  (.A(\u_multiplier/_2045_ ),
    .B(\u_multiplier/_2305_ ),
    .S(\u_multiplier/_3111_ ),
    .Z(\u_multiplier/_2306_ ));
 NOR2_X1 \u_multiplier/_4886_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2306_ ),
    .ZN(\u_multiplier/_2307_ ));
 AOI21_X1 \u_multiplier/_4887_  (.A(\u_multiplier/_2307_ ),
    .B1(\u_multiplier/_3545_ ),
    .B2(\u_multiplier/code_x [4]),
    .ZN(\u_multiplier/_2308_ ));
 MUX2_X1 \u_multiplier/_4888_  (.A(\u_multiplier/_3229_ ),
    .B(\u_multiplier/_3291_ ),
    .S(\u_multiplier/_3105_ ),
    .Z(\u_multiplier/_2309_ ));
 MUX2_X1 \u_multiplier/_4889_  (.A(\u_multiplier/_2309_ ),
    .B(\u_multiplier/_2245_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_2310_ ));
 MUX2_X1 \u_multiplier/_4890_  (.A(\u_multiplier/_2182_ ),
    .B(\u_multiplier/_2310_ ),
    .S(\u_multiplier/_3106_ ),
    .Z(\u_multiplier/_2311_ ));
 MUX2_X2 \u_multiplier/_4891_  (.A(\u_multiplier/_2051_ ),
    .B(\u_multiplier/_2311_ ),
    .S(\u_multiplier/_3107_ ),
    .Z(\u_multiplier/_2312_ ));
 NAND2_X1 \u_multiplier/_4892_  (.A1(\u_multiplier/_3108_ ),
    .A2(\u_multiplier/_2312_ ),
    .ZN(\u_multiplier/_2313_ ));
 OAI21_X1 \u_multiplier/_4893_  (.A(\u_multiplier/_2313_ ),
    .B1(\u_multiplier/_3552_ ),
    .B2(\u_multiplier/_3108_ ),
    .ZN(\u_multiplier/_2314_ ));
 NAND2_X1 \u_multiplier/_4894_  (.A1(\u_multiplier/_2308_ ),
    .A2(\u_multiplier/_2314_ ),
    .ZN(\u_multiplier/_2315_ ));
 XOR2_X1 \u_multiplier/_4895_  (.A(\u_multiplier/_2308_ ),
    .B(\u_multiplier/_2314_ ),
    .Z(\u_multiplier/_2316_ ));
 OAI21_X1 \u_multiplier/_4896_  (.A(\u_multiplier/_2316_ ),
    .B1(\u_multiplier/_2302_ ),
    .B2(\u_multiplier/dec_out [24]),
    .ZN(\u_multiplier/_2317_ ));
 OR3_X1 \u_multiplier/_4897_  (.A1(\u_multiplier/dec_out [24]),
    .A2(\u_multiplier/_2302_ ),
    .A3(\u_multiplier/_2316_ ),
    .ZN(\u_multiplier/_2318_ ));
 AND2_X1 \u_multiplier/_4898_  (.A1(\u_multiplier/_2317_ ),
    .A2(\u_multiplier/_2318_ ),
    .ZN(\u_multiplier/_2319_ ));
 NAND2_X1 \u_multiplier/_4899_  (.A1(\u_multiplier/_2296_ ),
    .A2(\u_multiplier/_2319_ ),
    .ZN(\u_multiplier/_2320_ ));
 XOR2_X2 \u_multiplier/_4900_  (.A(\u_multiplier/_2296_ ),
    .B(\u_multiplier/_2319_ ),
    .Z(\u_multiplier/_2321_ ));
 INV_X1 \u_multiplier/_4901_  (.A(\u_multiplier/_2321_ ),
    .ZN(\u_multiplier/_2322_ ));
 AOI21_X4 \u_multiplier/_4902_  (.A(\u_multiplier/_2322_ ),
    .B1(\u_multiplier/_2294_ ),
    .B2(\u_multiplier/_2292_ ),
    .ZN(\u_multiplier/_2323_ ));
 OAI21_X2 \u_multiplier/_4903_  (.A(net21),
    .B1(\u_multiplier/_2295_ ),
    .B2(\u_multiplier/_2321_ ),
    .ZN(\u_multiplier/_2324_ ));
 NOR2_X4 \u_multiplier/_4904_  (.A1(\u_multiplier/_2323_ ),
    .A2(\u_multiplier/_2324_ ),
    .ZN(product[24]));
 NAND2_X1 \u_multiplier/_4905_  (.A1(\u_multiplier/_2315_ ),
    .A2(\u_multiplier/_2317_ ),
    .ZN(\u_multiplier/_2325_ ));
 MUX2_X1 \u_multiplier/_4906_  (.A(\u_multiplier/_3289_ ),
    .B(\u_multiplier/_3287_ ),
    .S(\u_multiplier/_3313_ ),
    .Z(\u_multiplier/_2326_ ));
 MUX2_X1 \u_multiplier/_4907_  (.A(\u_multiplier/_2297_ ),
    .B(\u_multiplier/_2326_ ),
    .S(\u_multiplier/_3113_ ),
    .Z(\u_multiplier/_2327_ ));
 MUX2_X1 \u_multiplier/_4908_  (.A(\u_multiplier/_2262_ ),
    .B(\u_multiplier/_2327_ ),
    .S(\u_multiplier/_3114_ ),
    .Z(\u_multiplier/_2328_ ));
 MUX2_X1 \u_multiplier/_4909_  (.A(\u_multiplier/_2200_ ),
    .B(\u_multiplier/_2328_ ),
    .S(\u_multiplier/_3112_ ),
    .Z(\u_multiplier/_2329_ ));
 NAND2_X1 \u_multiplier/_4910_  (.A1(\u_multiplier/_3115_ ),
    .A2(\u_multiplier/_2329_ ),
    .ZN(\u_multiplier/_2330_ ));
 OAI21_X4 \u_multiplier/_4911_  (.A(\u_multiplier/_2330_ ),
    .B1(\u_multiplier/_2070_ ),
    .B2(\u_multiplier/_3115_ ),
    .ZN(\u_multiplier/_2331_ ));
 NOR2_X1 \u_multiplier/_4912_  (.A1(\u_multiplier/_3116_ ),
    .A2(\u_multiplier/_3569_ ),
    .ZN(\u_multiplier/_2332_ ));
 AOI211_X2 \u_multiplier/_4913_  (.A(\u_multiplier/dec_out [25]),
    .B(\u_multiplier/_2332_ ),
    .C1(\u_multiplier/_2331_ ),
    .C2(\u_multiplier/_3116_ ),
    .ZN(\u_multiplier/_2333_ ));
 MUX2_X1 \u_multiplier/_4914_  (.A(\u_multiplier/_3289_ ),
    .B(\u_multiplier/_3292_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_2334_ ));
 MUX2_X1 \u_multiplier/_4915_  (.A(\u_multiplier/_2334_ ),
    .B(\u_multiplier/_2270_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_2335_ ));
 MUX2_X1 \u_multiplier/_4916_  (.A(\u_multiplier/_2207_ ),
    .B(\u_multiplier/_2335_ ),
    .S(\u_multiplier/_3110_ ),
    .Z(\u_multiplier/_2336_ ));
 MUX2_X1 \u_multiplier/_4917_  (.A(\u_multiplier/_2076_ ),
    .B(\u_multiplier/_2336_ ),
    .S(\u_multiplier/_3111_ ),
    .Z(\u_multiplier/_2337_ ));
 NOR2_X1 \u_multiplier/_4918_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2337_ ),
    .ZN(\u_multiplier/_2338_ ));
 AOI21_X2 \u_multiplier/_4919_  (.A(\u_multiplier/_2338_ ),
    .B1(\u_multiplier/_3576_ ),
    .B2(\u_multiplier/code_x [4]),
    .ZN(\u_multiplier/_2339_ ));
 MUX2_X1 \u_multiplier/_4920_  (.A(\u_multiplier/_3287_ ),
    .B(\u_multiplier/_3291_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_2340_ ));
 MUX2_X1 \u_multiplier/_4921_  (.A(\u_multiplier/_2340_ ),
    .B(\u_multiplier/_2276_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_2341_ ));
 MUX2_X1 \u_multiplier/_4922_  (.A(\u_multiplier/_2213_ ),
    .B(\u_multiplier/_2341_ ),
    .S(\u_multiplier/_3106_ ),
    .Z(\u_multiplier/_2342_ ));
 MUX2_X2 \u_multiplier/_4923_  (.A(\u_multiplier/_2084_ ),
    .B(\u_multiplier/_2342_ ),
    .S(\u_multiplier/_3107_ ),
    .Z(\u_multiplier/_2343_ ));
 NAND2_X1 \u_multiplier/_4924_  (.A1(\u_multiplier/_3108_ ),
    .A2(\u_multiplier/_2343_ ),
    .ZN(\u_multiplier/_2344_ ));
 OAI21_X2 \u_multiplier/_4925_  (.A(\u_multiplier/_2344_ ),
    .B1(\u_multiplier/_3582_ ),
    .B2(\u_multiplier/_3108_ ),
    .ZN(\u_multiplier/_2345_ ));
 NAND2_X1 \u_multiplier/_4926_  (.A1(\u_multiplier/_2339_ ),
    .A2(\u_multiplier/_2345_ ),
    .ZN(\u_multiplier/_2346_ ));
 XOR2_X2 \u_multiplier/_4927_  (.A(\u_multiplier/_2339_ ),
    .B(\u_multiplier/_2345_ ),
    .Z(\u_multiplier/_2347_ ));
 INV_X1 \u_multiplier/_4928_  (.A(\u_multiplier/_2347_ ),
    .ZN(\u_multiplier/_2348_ ));
 XNOR2_X2 \u_multiplier/_4929_  (.A(\u_multiplier/_2333_ ),
    .B(\u_multiplier/_2347_ ),
    .ZN(\u_multiplier/_2349_ ));
 NAND2_X1 \u_multiplier/_4930_  (.A1(\u_multiplier/_2325_ ),
    .A2(\u_multiplier/_2349_ ),
    .ZN(\u_multiplier/_2350_ ));
 XNOR2_X2 \u_multiplier/_4931_  (.A(\u_multiplier/_2325_ ),
    .B(\u_multiplier/_2349_ ),
    .ZN(\u_multiplier/_2351_ ));
 NAND2_X1 \u_multiplier/_4932_  (.A1(\u_multiplier/_2320_ ),
    .A2(\u_multiplier/_2351_ ),
    .ZN(\u_multiplier/_2352_ ));
 AOI211_X2 \u_multiplier/_4933_  (.A(\u_multiplier/_2322_ ),
    .B(\u_multiplier/_2351_ ),
    .C1(\u_multiplier/_2292_ ),
    .C2(\u_multiplier/_2294_ ),
    .ZN(\u_multiplier/_2353_ ));
 OAI21_X1 \u_multiplier/_4934_  (.A(net21),
    .B1(\u_multiplier/_2320_ ),
    .B2(\u_multiplier/_2351_ ),
    .ZN(\u_multiplier/_2354_ ));
 NOR2_X1 \u_multiplier/_4935_  (.A1(\u_multiplier/_2353_ ),
    .A2(\u_multiplier/_2354_ ),
    .ZN(\u_multiplier/_2355_ ));
 OAI21_X2 \u_multiplier/_4936_  (.A(\u_multiplier/_2355_ ),
    .B1(\u_multiplier/_2352_ ),
    .B2(\u_multiplier/_2323_ ),
    .ZN(\u_multiplier/_2356_ ));
 INV_X1 \u_multiplier/_4937_  (.A(\u_multiplier/_2356_ ),
    .ZN(product[25]));
 OAI21_X2 \u_multiplier/_4938_  (.A(\u_multiplier/_2350_ ),
    .B1(\u_multiplier/_2351_ ),
    .B2(\u_multiplier/_2320_ ),
    .ZN(\u_multiplier/_2357_ ));
 NOR2_X1 \u_multiplier/_4939_  (.A1(\u_multiplier/_2353_ ),
    .A2(\u_multiplier/_2357_ ),
    .ZN(\u_multiplier/_2358_ ));
 OAI21_X2 \u_multiplier/_4940_  (.A(\u_multiplier/_2346_ ),
    .B1(\u_multiplier/_2348_ ),
    .B2(\u_multiplier/_2333_ ),
    .ZN(\u_multiplier/_2359_ ));
 MUX2_X1 \u_multiplier/_4941_  (.A(\u_multiplier/_3277_ ),
    .B(\u_multiplier/_3276_ ),
    .S(\u_multiplier/_3313_ ),
    .Z(\u_multiplier/_2360_ ));
 MUX2_X1 \u_multiplier/_4942_  (.A(\u_multiplier/_2326_ ),
    .B(\u_multiplier/_2360_ ),
    .S(\u_multiplier/_3113_ ),
    .Z(\u_multiplier/_2361_ ));
 MUX2_X1 \u_multiplier/_4943_  (.A(\u_multiplier/_2298_ ),
    .B(\u_multiplier/_2361_ ),
    .S(\u_multiplier/_3114_ ),
    .Z(\u_multiplier/_2362_ ));
 MUX2_X1 \u_multiplier/_4944_  (.A(\u_multiplier/_2233_ ),
    .B(\u_multiplier/_2362_ ),
    .S(\u_multiplier/_3112_ ),
    .Z(\u_multiplier/_2363_ ));
 MUX2_X2 \u_multiplier/_4945_  (.A(\u_multiplier/_2104_ ),
    .B(\u_multiplier/_2363_ ),
    .S(\u_multiplier/_3115_ ),
    .Z(\u_multiplier/_2364_ ));
 AND2_X1 \u_multiplier/_4946_  (.A1(\u_multiplier/_3116_ ),
    .A2(\u_multiplier/_2364_ ),
    .ZN(\u_multiplier/_2365_ ));
 AOI211_X2 \u_multiplier/_4947_  (.A(\u_multiplier/dec_out [26]),
    .B(\u_multiplier/_2365_ ),
    .C1(\u_multiplier/_3600_ ),
    .C2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2366_ ));
 MUX2_X1 \u_multiplier/_4948_  (.A(\u_multiplier/_3277_ ),
    .B(\u_multiplier/_3289_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_2367_ ));
 MUX2_X1 \u_multiplier/_4949_  (.A(\u_multiplier/_2367_ ),
    .B(\u_multiplier/_2303_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_2368_ ));
 MUX2_X1 \u_multiplier/_4950_  (.A(\u_multiplier/_2240_ ),
    .B(\u_multiplier/_2368_ ),
    .S(\u_multiplier/_3110_ ),
    .Z(\u_multiplier/_2369_ ));
 NAND2_X1 \u_multiplier/_4951_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_2113_ ),
    .ZN(\u_multiplier/_2370_ ));
 OAI21_X2 \u_multiplier/_4952_  (.A(\u_multiplier/_2370_ ),
    .B1(\u_multiplier/_2369_ ),
    .B2(\u_multiplier/code_x [3]),
    .ZN(\u_multiplier/_2371_ ));
 MUX2_X1 \u_multiplier/_4953_  (.A(\u_multiplier/_3606_ ),
    .B(\u_multiplier/_2371_ ),
    .S(\u_multiplier/_3109_ ),
    .Z(\u_multiplier/_2372_ ));
 MUX2_X1 \u_multiplier/_4954_  (.A(\u_multiplier/_3276_ ),
    .B(\u_multiplier/_3287_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_2373_ ));
 MUX2_X1 \u_multiplier/_4955_  (.A(\u_multiplier/_2373_ ),
    .B(\u_multiplier/_2309_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_2374_ ));
 MUX2_X1 \u_multiplier/_4956_  (.A(\u_multiplier/_2246_ ),
    .B(\u_multiplier/_2374_ ),
    .S(\u_multiplier/_3106_ ),
    .Z(\u_multiplier/_2375_ ));
 NAND2_X1 \u_multiplier/_4957_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_2120_ ),
    .ZN(\u_multiplier/_2376_ ));
 OAI21_X2 \u_multiplier/_4958_  (.A(\u_multiplier/_2376_ ),
    .B1(\u_multiplier/_2375_ ),
    .B2(\u_multiplier/code_y [3]),
    .ZN(\u_multiplier/_2377_ ));
 MUX2_X1 \u_multiplier/_4959_  (.A(\u_multiplier/_3611_ ),
    .B(\u_multiplier/_2377_ ),
    .S(\u_multiplier/_3108_ ),
    .Z(\u_multiplier/_2378_ ));
 OR2_X1 \u_multiplier/_4960_  (.A1(\u_multiplier/_2372_ ),
    .A2(\u_multiplier/_2378_ ),
    .ZN(\u_multiplier/_2379_ ));
 XNOR2_X2 \u_multiplier/_4961_  (.A(\u_multiplier/_2372_ ),
    .B(\u_multiplier/_2378_ ),
    .ZN(\u_multiplier/_2380_ ));
 XOR2_X2 \u_multiplier/_4962_  (.A(\u_multiplier/_2366_ ),
    .B(\u_multiplier/_2380_ ),
    .Z(\u_multiplier/_2381_ ));
 NAND2_X1 \u_multiplier/_4963_  (.A1(\u_multiplier/_2359_ ),
    .A2(\u_multiplier/_2381_ ),
    .ZN(\u_multiplier/_2382_ ));
 XNOR2_X2 \u_multiplier/_4964_  (.A(\u_multiplier/_2359_ ),
    .B(\u_multiplier/_2381_ ),
    .ZN(\u_multiplier/_2383_ ));
 INV_X1 \u_multiplier/_4965_  (.A(\u_multiplier/_2383_ ),
    .ZN(\u_multiplier/_2384_ ));
 NOR2_X1 \u_multiplier/_4966_  (.A1(\u_multiplier/_2358_ ),
    .A2(\u_multiplier/_2383_ ),
    .ZN(\u_multiplier/_2385_ ));
 NOR3_X1 \u_multiplier/_4967_  (.A1(\u_multiplier/_2353_ ),
    .A2(\u_multiplier/_2357_ ),
    .A3(\u_multiplier/_2384_ ),
    .ZN(\u_multiplier/_2386_ ));
 NOR3_X1 \u_multiplier/_4968_  (.A1(\u_multiplier/_3334_ ),
    .A2(\u_multiplier/_2385_ ),
    .A3(\u_multiplier/_2386_ ),
    .ZN(product[26]));
 OAI21_X1 \u_multiplier/_4969_  (.A(\u_multiplier/_2382_ ),
    .B1(\u_multiplier/_2383_ ),
    .B2(\u_multiplier/_2358_ ),
    .ZN(\u_multiplier/_2387_ ));
 OAI21_X2 \u_multiplier/_4970_  (.A(\u_multiplier/_2379_ ),
    .B1(\u_multiplier/_2380_ ),
    .B2(\u_multiplier/_2366_ ),
    .ZN(\u_multiplier/_2388_ ));
 MUX2_X1 \u_multiplier/_4971_  (.A(\u_multiplier/_3282_ ),
    .B(\u_multiplier/_3280_ ),
    .S(\u_multiplier/_3313_ ),
    .Z(\u_multiplier/_2389_ ));
 MUX2_X1 \u_multiplier/_4972_  (.A(\u_multiplier/_2360_ ),
    .B(\u_multiplier/_2389_ ),
    .S(\u_multiplier/_3113_ ),
    .Z(\u_multiplier/_2390_ ));
 MUX2_X1 \u_multiplier/_4973_  (.A(\u_multiplier/_2327_ ),
    .B(\u_multiplier/_2390_ ),
    .S(\u_multiplier/_3114_ ),
    .Z(\u_multiplier/_2391_ ));
 MUX2_X1 \u_multiplier/_4974_  (.A(\u_multiplier/_2263_ ),
    .B(\u_multiplier/_2391_ ),
    .S(\u_multiplier/_3112_ ),
    .Z(\u_multiplier/_2392_ ));
 NAND2_X1 \u_multiplier/_4975_  (.A1(\u_multiplier/_3115_ ),
    .A2(\u_multiplier/_2392_ ),
    .ZN(\u_multiplier/_2393_ ));
 OAI21_X4 \u_multiplier/_4976_  (.A(\u_multiplier/_2393_ ),
    .B1(\u_multiplier/_2140_ ),
    .B2(\u_multiplier/_3115_ ),
    .ZN(\u_multiplier/_2394_ ));
 AND2_X1 \u_multiplier/_4977_  (.A1(\u_multiplier/K [4]),
    .A2(\u_multiplier/_3628_ ),
    .ZN(\u_multiplier/_2395_ ));
 AOI211_X2 \u_multiplier/_4978_  (.A(\u_multiplier/dec_out [27]),
    .B(\u_multiplier/_2395_ ),
    .C1(\u_multiplier/_2394_ ),
    .C2(\u_multiplier/_3116_ ),
    .ZN(\u_multiplier/_2396_ ));
 MUX2_X1 \u_multiplier/_4979_  (.A(\u_multiplier/_3282_ ),
    .B(\u_multiplier/_3277_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_2397_ ));
 MUX2_X1 \u_multiplier/_4980_  (.A(\u_multiplier/_2397_ ),
    .B(\u_multiplier/_2334_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_2398_ ));
 MUX2_X1 \u_multiplier/_4981_  (.A(\u_multiplier/_2271_ ),
    .B(\u_multiplier/_2398_ ),
    .S(\u_multiplier/_3110_ ),
    .Z(\u_multiplier/_2399_ ));
 MUX2_X2 \u_multiplier/_4982_  (.A(\u_multiplier/_2147_ ),
    .B(\u_multiplier/_2399_ ),
    .S(\u_multiplier/_3111_ ),
    .Z(\u_multiplier/_2400_ ));
 NOR2_X1 \u_multiplier/_4983_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2400_ ),
    .ZN(\u_multiplier/_2401_ ));
 AOI21_X2 \u_multiplier/_4984_  (.A(\u_multiplier/_2401_ ),
    .B1(\u_multiplier/_3634_ ),
    .B2(\u_multiplier/code_x [4]),
    .ZN(\u_multiplier/_2402_ ));
 MUX2_X1 \u_multiplier/_4985_  (.A(\u_multiplier/_3276_ ),
    .B(\u_multiplier/_3280_ ),
    .S(\u_multiplier/_3105_ ),
    .Z(\u_multiplier/_2403_ ));
 MUX2_X1 \u_multiplier/_4986_  (.A(\u_multiplier/_2403_ ),
    .B(\u_multiplier/_2340_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_2404_ ));
 MUX2_X1 \u_multiplier/_4987_  (.A(\u_multiplier/_2277_ ),
    .B(\u_multiplier/_2404_ ),
    .S(\u_multiplier/_3106_ ),
    .Z(\u_multiplier/_2405_ ));
 MUX2_X2 \u_multiplier/_4988_  (.A(\u_multiplier/_2153_ ),
    .B(\u_multiplier/_2405_ ),
    .S(\u_multiplier/_3107_ ),
    .Z(\u_multiplier/_2406_ ));
 NAND2_X1 \u_multiplier/_4989_  (.A1(\u_multiplier/_3108_ ),
    .A2(\u_multiplier/_2406_ ),
    .ZN(\u_multiplier/_2407_ ));
 OAI21_X2 \u_multiplier/_4990_  (.A(\u_multiplier/_2407_ ),
    .B1(\u_multiplier/_3640_ ),
    .B2(\u_multiplier/_3108_ ),
    .ZN(\u_multiplier/_2408_ ));
 NAND2_X1 \u_multiplier/_4991_  (.A1(\u_multiplier/_2402_ ),
    .A2(\u_multiplier/_2408_ ),
    .ZN(\u_multiplier/_2409_ ));
 XOR2_X2 \u_multiplier/_4992_  (.A(\u_multiplier/_2402_ ),
    .B(\u_multiplier/_2408_ ),
    .Z(\u_multiplier/_2410_ ));
 INV_X1 \u_multiplier/_4993_  (.A(\u_multiplier/_2410_ ),
    .ZN(\u_multiplier/_2411_ ));
 XNOR2_X2 \u_multiplier/_4994_  (.A(\u_multiplier/_2396_ ),
    .B(\u_multiplier/_2410_ ),
    .ZN(\u_multiplier/_2412_ ));
 NAND2_X1 \u_multiplier/_4995_  (.A1(\u_multiplier/_2388_ ),
    .A2(\u_multiplier/_2412_ ),
    .ZN(\u_multiplier/_2413_ ));
 NOR2_X1 \u_multiplier/_4996_  (.A1(\u_multiplier/_2388_ ),
    .A2(\u_multiplier/_2412_ ),
    .ZN(\u_multiplier/_2414_ ));
 XOR2_X2 \u_multiplier/_4997_  (.A(\u_multiplier/_2388_ ),
    .B(\u_multiplier/_2412_ ),
    .Z(\u_multiplier/_2415_ ));
 OAI21_X1 \u_multiplier/_4998_  (.A(net21),
    .B1(\u_multiplier/_2387_ ),
    .B2(\u_multiplier/_2415_ ),
    .ZN(\u_multiplier/_2416_ ));
 AOI21_X1 \u_multiplier/_4999_  (.A(\u_multiplier/_2416_ ),
    .B1(\u_multiplier/_2415_ ),
    .B2(\u_multiplier/_2387_ ),
    .ZN(product[27]));
 OAI211_X2 \u_multiplier/_5000_  (.A(\u_multiplier/_2384_ ),
    .B(\u_multiplier/_2415_ ),
    .C1(\u_multiplier/_2353_ ),
    .C2(\u_multiplier/_2357_ ),
    .ZN(\u_multiplier/_2417_ ));
 OAI21_X1 \u_multiplier/_5001_  (.A(\u_multiplier/_2413_ ),
    .B1(\u_multiplier/_2414_ ),
    .B2(\u_multiplier/_2382_ ),
    .ZN(\u_multiplier/_2418_ ));
 INV_X1 \u_multiplier/_5002_  (.A(\u_multiplier/_2418_ ),
    .ZN(\u_multiplier/_2419_ ));
 AND2_X1 \u_multiplier/_5003_  (.A1(\u_multiplier/_2417_ ),
    .A2(\u_multiplier/_2419_ ),
    .ZN(\u_multiplier/_2420_ ));
 OAI21_X2 \u_multiplier/_5004_  (.A(\u_multiplier/_2409_ ),
    .B1(\u_multiplier/_2411_ ),
    .B2(\u_multiplier/_2396_ ),
    .ZN(\u_multiplier/_2421_ ));
 MUX2_X1 \u_multiplier/_5005_  (.A(\u_multiplier/_3307_ ),
    .B(\u_multiplier/_3306_ ),
    .S(\u_multiplier/_3313_ ),
    .Z(\u_multiplier/_2422_ ));
 MUX2_X1 \u_multiplier/_5006_  (.A(\u_multiplier/_2389_ ),
    .B(\u_multiplier/_2422_ ),
    .S(\u_multiplier/_3113_ ),
    .Z(\u_multiplier/_2423_ ));
 MUX2_X1 \u_multiplier/_5007_  (.A(\u_multiplier/_2361_ ),
    .B(\u_multiplier/_2423_ ),
    .S(\u_multiplier/_3114_ ),
    .Z(\u_multiplier/_2424_ ));
 MUX2_X1 \u_multiplier/_5008_  (.A(\u_multiplier/_2299_ ),
    .B(\u_multiplier/_2424_ ),
    .S(\u_multiplier/_3112_ ),
    .Z(\u_multiplier/_2425_ ));
 MUX2_X2 \u_multiplier/_5009_  (.A(\u_multiplier/_2170_ ),
    .B(\u_multiplier/_2425_ ),
    .S(\u_multiplier/_3115_ ),
    .Z(\u_multiplier/_2426_ ));
 NOR2_X1 \u_multiplier/_5010_  (.A1(\u_multiplier/K [4]),
    .A2(\u_multiplier/_2426_ ),
    .ZN(\u_multiplier/_2427_ ));
 AOI21_X1 \u_multiplier/_5011_  (.A(\u_multiplier/_2427_ ),
    .B1(\u_multiplier/_3659_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2428_ ));
 MUX2_X1 \u_multiplier/_5012_  (.A(\u_multiplier/_3307_ ),
    .B(\u_multiplier/_3282_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_2429_ ));
 MUX2_X1 \u_multiplier/_5013_  (.A(\u_multiplier/_2429_ ),
    .B(\u_multiplier/_2367_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_2430_ ));
 MUX2_X1 \u_multiplier/_5014_  (.A(\u_multiplier/_2304_ ),
    .B(\u_multiplier/_2430_ ),
    .S(\u_multiplier/_3110_ ),
    .Z(\u_multiplier/_2431_ ));
 NOR2_X1 \u_multiplier/_5015_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_2431_ ),
    .ZN(\u_multiplier/_2432_ ));
 AOI21_X2 \u_multiplier/_5016_  (.A(\u_multiplier/_2432_ ),
    .B1(\u_multiplier/_2178_ ),
    .B2(\u_multiplier/code_x [3]),
    .ZN(\u_multiplier/_2433_ ));
 NOR2_X1 \u_multiplier/_5017_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2433_ ),
    .ZN(\u_multiplier/_2434_ ));
 AOI21_X1 \u_multiplier/_5018_  (.A(\u_multiplier/_2434_ ),
    .B1(\u_multiplier/_3667_ ),
    .B2(\u_multiplier/code_x [4]),
    .ZN(\u_multiplier/_2435_ ));
 MUX2_X1 \u_multiplier/_5019_  (.A(\u_multiplier/_3280_ ),
    .B(\u_multiplier/_3306_ ),
    .S(\u_multiplier/_3105_ ),
    .Z(\u_multiplier/_2436_ ));
 MUX2_X1 \u_multiplier/_5020_  (.A(\u_multiplier/_2436_ ),
    .B(\u_multiplier/_2373_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_2437_ ));
 MUX2_X1 \u_multiplier/_5021_  (.A(\u_multiplier/_2310_ ),
    .B(\u_multiplier/_2437_ ),
    .S(\u_multiplier/_3106_ ),
    .Z(\u_multiplier/_2438_ ));
 NOR2_X1 \u_multiplier/_5022_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_2438_ ),
    .ZN(\u_multiplier/_2439_ ));
 AOI21_X4 \u_multiplier/_5023_  (.A(\u_multiplier/_2439_ ),
    .B1(\u_multiplier/_2184_ ),
    .B2(\u_multiplier/code_y [3]),
    .ZN(\u_multiplier/_2440_ ));
 NAND2_X1 \u_multiplier/_5024_  (.A1(\u_multiplier/_3108_ ),
    .A2(\u_multiplier/_2440_ ),
    .ZN(\u_multiplier/_2441_ ));
 OAI21_X1 \u_multiplier/_5025_  (.A(\u_multiplier/_2441_ ),
    .B1(\u_multiplier/_3674_ ),
    .B2(\u_multiplier/_3108_ ),
    .ZN(\u_multiplier/_2442_ ));
 NAND2_X1 \u_multiplier/_5026_  (.A1(\u_multiplier/_2435_ ),
    .A2(\u_multiplier/_2442_ ),
    .ZN(\u_multiplier/_2443_ ));
 XOR2_X1 \u_multiplier/_5027_  (.A(\u_multiplier/_2435_ ),
    .B(\u_multiplier/_2442_ ),
    .Z(\u_multiplier/_2444_ ));
 OAI21_X1 \u_multiplier/_5028_  (.A(\u_multiplier/_2444_ ),
    .B1(\u_multiplier/_2428_ ),
    .B2(\u_multiplier/dec_out [28]),
    .ZN(\u_multiplier/_2445_ ));
 OR3_X1 \u_multiplier/_5029_  (.A1(\u_multiplier/dec_out [28]),
    .A2(\u_multiplier/_2428_ ),
    .A3(\u_multiplier/_2444_ ),
    .ZN(\u_multiplier/_2446_ ));
 AND2_X1 \u_multiplier/_5030_  (.A1(\u_multiplier/_2445_ ),
    .A2(\u_multiplier/_2446_ ),
    .ZN(\u_multiplier/_2447_ ));
 NAND2_X1 \u_multiplier/_5031_  (.A1(\u_multiplier/_2421_ ),
    .A2(\u_multiplier/_2447_ ),
    .ZN(\u_multiplier/_2448_ ));
 XNOR2_X2 \u_multiplier/_5032_  (.A(\u_multiplier/_2421_ ),
    .B(\u_multiplier/_2447_ ),
    .ZN(\u_multiplier/_2449_ ));
 NOR2_X1 \u_multiplier/_5033_  (.A1(\u_multiplier/_2420_ ),
    .A2(\u_multiplier/_2449_ ),
    .ZN(\u_multiplier/_2450_ ));
 AND2_X1 \u_multiplier/_5034_  (.A1(\u_multiplier/_2420_ ),
    .A2(\u_multiplier/_2449_ ),
    .ZN(\u_multiplier/_2451_ ));
 NOR3_X1 \u_multiplier/_5035_  (.A1(\u_multiplier/_3334_ ),
    .A2(\u_multiplier/_2450_ ),
    .A3(\u_multiplier/_2451_ ),
    .ZN(product[28]));
 NAND2_X1 \u_multiplier/_5036_  (.A1(\u_multiplier/_2443_ ),
    .A2(\u_multiplier/_2445_ ),
    .ZN(\u_multiplier/_2452_ ));
 MUX2_X1 \u_multiplier/_5037_  (.A(\u_multiplier/_3303_ ),
    .B(\u_multiplier/_3301_ ),
    .S(\u_multiplier/_3313_ ),
    .Z(\u_multiplier/_2453_ ));
 MUX2_X1 \u_multiplier/_5038_  (.A(\u_multiplier/_2422_ ),
    .B(\u_multiplier/_2453_ ),
    .S(\u_multiplier/_3113_ ),
    .Z(\u_multiplier/_2454_ ));
 MUX2_X1 \u_multiplier/_5039_  (.A(\u_multiplier/_2390_ ),
    .B(\u_multiplier/_2454_ ),
    .S(\u_multiplier/_3114_ ),
    .Z(\u_multiplier/_2455_ ));
 MUX2_X1 \u_multiplier/_5040_  (.A(\u_multiplier/_2328_ ),
    .B(\u_multiplier/_2455_ ),
    .S(\u_multiplier/_3112_ ),
    .Z(\u_multiplier/_2456_ ));
 MUX2_X2 \u_multiplier/_5041_  (.A(\u_multiplier/_2202_ ),
    .B(\u_multiplier/_2456_ ),
    .S(\u_multiplier/_3115_ ),
    .Z(\u_multiplier/_2457_ ));
 NOR2_X1 \u_multiplier/_5042_  (.A1(\u_multiplier/_3116_ ),
    .A2(\u_multiplier/_3691_ ),
    .ZN(\u_multiplier/_2458_ ));
 AOI211_X2 \u_multiplier/_5043_  (.A(\u_multiplier/dec_out [29]),
    .B(\u_multiplier/_2458_ ),
    .C1(\u_multiplier/_2457_ ),
    .C2(\u_multiplier/_3116_ ),
    .ZN(\u_multiplier/_2459_ ));
 MUX2_X1 \u_multiplier/_5044_  (.A(\u_multiplier/_3303_ ),
    .B(\u_multiplier/_3307_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_2460_ ));
 MUX2_X1 \u_multiplier/_5045_  (.A(\u_multiplier/_2460_ ),
    .B(\u_multiplier/_2397_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_2461_ ));
 MUX2_X1 \u_multiplier/_5046_  (.A(\u_multiplier/_2335_ ),
    .B(\u_multiplier/_2461_ ),
    .S(\u_multiplier/_3110_ ),
    .Z(\u_multiplier/_2462_ ));
 NOR2_X1 \u_multiplier/_5047_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_2462_ ),
    .ZN(\u_multiplier/_2463_ ));
 AOI21_X2 \u_multiplier/_5048_  (.A(\u_multiplier/_2463_ ),
    .B1(\u_multiplier/_2209_ ),
    .B2(\u_multiplier/code_x [3]),
    .ZN(\u_multiplier/_2464_ ));
 NOR2_X1 \u_multiplier/_5049_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2464_ ),
    .ZN(\u_multiplier/_2465_ ));
 AOI21_X2 \u_multiplier/_5050_  (.A(\u_multiplier/_2465_ ),
    .B1(\u_multiplier/_3700_ ),
    .B2(\u_multiplier/code_x [4]),
    .ZN(\u_multiplier/_2466_ ));
 MUX2_X1 \u_multiplier/_5051_  (.A(\u_multiplier/_3301_ ),
    .B(\u_multiplier/_3306_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_2467_ ));
 MUX2_X2 \u_multiplier/_5052_  (.A(\u_multiplier/_2467_ ),
    .B(\u_multiplier/_2403_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_2468_ ));
 MUX2_X1 \u_multiplier/_5053_  (.A(\u_multiplier/_2341_ ),
    .B(\u_multiplier/_2468_ ),
    .S(\u_multiplier/_3106_ ),
    .Z(\u_multiplier/_2469_ ));
 MUX2_X2 \u_multiplier/_5054_  (.A(\u_multiplier/_2214_ ),
    .B(\u_multiplier/_2469_ ),
    .S(\u_multiplier/_3107_ ),
    .Z(\u_multiplier/_2470_ ));
 NOR2_X1 \u_multiplier/_5055_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_2470_ ),
    .ZN(\u_multiplier/_2471_ ));
 AOI21_X2 \u_multiplier/_5056_  (.A(\u_multiplier/_2471_ ),
    .B1(\u_multiplier/_3707_ ),
    .B2(\u_multiplier/code_y [4]),
    .ZN(\u_multiplier/_2472_ ));
 NAND2_X1 \u_multiplier/_5057_  (.A1(\u_multiplier/_2466_ ),
    .A2(\u_multiplier/_2472_ ),
    .ZN(\u_multiplier/_2473_ ));
 XNOR2_X2 \u_multiplier/_5058_  (.A(\u_multiplier/_2466_ ),
    .B(\u_multiplier/_2472_ ),
    .ZN(\u_multiplier/_2474_ ));
 XOR2_X2 \u_multiplier/_5059_  (.A(\u_multiplier/_2459_ ),
    .B(\u_multiplier/_2474_ ),
    .Z(\u_multiplier/_2475_ ));
 XNOR2_X2 \u_multiplier/_5060_  (.A(\u_multiplier/_2452_ ),
    .B(\u_multiplier/_2475_ ),
    .ZN(\u_multiplier/_2476_ ));
 NAND2_X1 \u_multiplier/_5061_  (.A1(\u_multiplier/_2448_ ),
    .A2(\u_multiplier/_2476_ ),
    .ZN(\u_multiplier/_2477_ ));
 AOI211_X2 \u_multiplier/_5062_  (.A(\u_multiplier/_2449_ ),
    .B(\u_multiplier/_2476_ ),
    .C1(\u_multiplier/_2417_ ),
    .C2(\u_multiplier/_2419_ ),
    .ZN(\u_multiplier/_2478_ ));
 NOR2_X1 \u_multiplier/_5063_  (.A1(\u_multiplier/_2448_ ),
    .A2(\u_multiplier/_2476_ ),
    .ZN(\u_multiplier/_2479_ ));
 NOR3_X1 \u_multiplier/_5064_  (.A1(\u_multiplier/_3334_ ),
    .A2(\u_multiplier/_2478_ ),
    .A3(\u_multiplier/_2479_ ),
    .ZN(\u_multiplier/_2480_ ));
 OAI21_X2 \u_multiplier/_5065_  (.A(\u_multiplier/_2480_ ),
    .B1(\u_multiplier/_2477_ ),
    .B2(\u_multiplier/_2450_ ),
    .ZN(\u_multiplier/_2481_ ));
 INV_X2 \u_multiplier/_5066_  (.A(\u_multiplier/_2481_ ),
    .ZN(product[29]));
 AOI21_X1 \u_multiplier/_5067_  (.A(\u_multiplier/_2479_ ),
    .B1(\u_multiplier/_2475_ ),
    .B2(\u_multiplier/_2452_ ),
    .ZN(\u_multiplier/_2482_ ));
 INV_X1 \u_multiplier/_5068_  (.A(\u_multiplier/_2482_ ),
    .ZN(\u_multiplier/_2483_ ));
 NOR2_X1 \u_multiplier/_5069_  (.A1(\u_multiplier/_2478_ ),
    .A2(\u_multiplier/_2483_ ),
    .ZN(\u_multiplier/_2484_ ));
 OAI21_X2 \u_multiplier/_5070_  (.A(\u_multiplier/_2473_ ),
    .B1(\u_multiplier/_2474_ ),
    .B2(\u_multiplier/_2459_ ),
    .ZN(\u_multiplier/_2485_ ));
 AND2_X1 \u_multiplier/_5071_  (.A1(\u_multiplier/_3129_ ),
    .A2(\u_multiplier/_3131_ ),
    .ZN(\u_multiplier/_2486_ ));
 MUX2_X1 \u_multiplier/_5072_  (.A(\u_multiplier/_2453_ ),
    .B(\u_multiplier/_2486_ ),
    .S(\u_multiplier/_3113_ ),
    .Z(\u_multiplier/_2487_ ));
 MUX2_X1 \u_multiplier/_5073_  (.A(\u_multiplier/_2423_ ),
    .B(\u_multiplier/_2487_ ),
    .S(\u_multiplier/_3114_ ),
    .Z(\u_multiplier/_2488_ ));
 MUX2_X1 \u_multiplier/_5074_  (.A(\u_multiplier/_2362_ ),
    .B(\u_multiplier/_2488_ ),
    .S(\u_multiplier/_3112_ ),
    .Z(\u_multiplier/_2489_ ));
 MUX2_X2 \u_multiplier/_5075_  (.A(\u_multiplier/_2234_ ),
    .B(\u_multiplier/_2489_ ),
    .S(\u_multiplier/_3115_ ),
    .Z(\u_multiplier/_2490_ ));
 NOR2_X1 \u_multiplier/_5076_  (.A1(\u_multiplier/_3116_ ),
    .A2(\u_multiplier/_3726_ ),
    .ZN(\u_multiplier/_2491_ ));
 AOI211_X2 \u_multiplier/_5077_  (.A(\u_multiplier/dec_out [30]),
    .B(\u_multiplier/_2491_ ),
    .C1(\u_multiplier/_2490_ ),
    .C2(\u_multiplier/_3116_ ),
    .ZN(\u_multiplier/_2492_ ));
 MUX2_X1 \u_multiplier/_5078_  (.A(\u_multiplier/_3131_ ),
    .B(\u_multiplier/_3303_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_2493_ ));
 MUX2_X1 \u_multiplier/_5079_  (.A(\u_multiplier/_2493_ ),
    .B(\u_multiplier/_2429_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_2494_ ));
 MUX2_X1 \u_multiplier/_5080_  (.A(\u_multiplier/_2368_ ),
    .B(\u_multiplier/_2494_ ),
    .S(\u_multiplier/_3110_ ),
    .Z(\u_multiplier/_2495_ ));
 MUX2_X2 \u_multiplier/_5081_  (.A(\u_multiplier/_2241_ ),
    .B(\u_multiplier/_2495_ ),
    .S(\u_multiplier/_3111_ ),
    .Z(\u_multiplier/_2496_ ));
 NOR2_X1 \u_multiplier/_5082_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2496_ ),
    .ZN(\u_multiplier/_2497_ ));
 AOI21_X2 \u_multiplier/_5083_  (.A(\u_multiplier/_2497_ ),
    .B1(\u_multiplier/_3732_ ),
    .B2(\u_multiplier/code_x [4]),
    .ZN(\u_multiplier/_2498_ ));
 MUX2_X1 \u_multiplier/_5084_  (.A(\u_multiplier/_3129_ ),
    .B(\u_multiplier/_3301_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_2499_ ));
 MUX2_X1 \u_multiplier/_5085_  (.A(\u_multiplier/_2499_ ),
    .B(\u_multiplier/_2436_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_2500_ ));
 MUX2_X1 \u_multiplier/_5086_  (.A(\u_multiplier/_2374_ ),
    .B(\u_multiplier/_2500_ ),
    .S(\u_multiplier/_3106_ ),
    .Z(\u_multiplier/_2501_ ));
 MUX2_X2 \u_multiplier/_5087_  (.A(\u_multiplier/_2247_ ),
    .B(\u_multiplier/_2501_ ),
    .S(\u_multiplier/_3107_ ),
    .Z(\u_multiplier/_2502_ ));
 NOR2_X1 \u_multiplier/_5088_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_2502_ ),
    .ZN(\u_multiplier/_2503_ ));
 AOI21_X2 \u_multiplier/_5089_  (.A(\u_multiplier/_2503_ ),
    .B1(\u_multiplier/_3738_ ),
    .B2(\u_multiplier/code_y [4]),
    .ZN(\u_multiplier/_2504_ ));
 NAND2_X1 \u_multiplier/_5090_  (.A1(\u_multiplier/_2498_ ),
    .A2(\u_multiplier/_2504_ ),
    .ZN(\u_multiplier/_2505_ ));
 XNOR2_X2 \u_multiplier/_5091_  (.A(\u_multiplier/_2498_ ),
    .B(\u_multiplier/_2504_ ),
    .ZN(\u_multiplier/_2506_ ));
 XOR2_X2 \u_multiplier/_5092_  (.A(\u_multiplier/_2492_ ),
    .B(\u_multiplier/_2506_ ),
    .Z(\u_multiplier/_2507_ ));
 NAND2_X1 \u_multiplier/_5093_  (.A1(\u_multiplier/_2485_ ),
    .A2(\u_multiplier/_2507_ ),
    .ZN(\u_multiplier/_2508_ ));
 XNOR2_X2 \u_multiplier/_5094_  (.A(\u_multiplier/_2485_ ),
    .B(\u_multiplier/_2507_ ),
    .ZN(\u_multiplier/_2509_ ));
 INV_X1 \u_multiplier/_5095_  (.A(\u_multiplier/_2509_ ),
    .ZN(\u_multiplier/_2510_ ));
 NOR2_X1 \u_multiplier/_5096_  (.A1(\u_multiplier/_2484_ ),
    .A2(\u_multiplier/_2509_ ),
    .ZN(\u_multiplier/_2511_ ));
 NOR3_X1 \u_multiplier/_5097_  (.A1(\u_multiplier/_2478_ ),
    .A2(\u_multiplier/_2483_ ),
    .A3(\u_multiplier/_2510_ ),
    .ZN(\u_multiplier/_2512_ ));
 NOR3_X1 \u_multiplier/_5098_  (.A1(\u_multiplier/_3334_ ),
    .A2(\u_multiplier/_2511_ ),
    .A3(\u_multiplier/_2512_ ),
    .ZN(product[30]));
 OAI21_X1 \u_multiplier/_5099_  (.A(\u_multiplier/_2508_ ),
    .B1(\u_multiplier/_2509_ ),
    .B2(\u_multiplier/_2484_ ),
    .ZN(\u_multiplier/_2513_ ));
 OAI21_X2 \u_multiplier/_5100_  (.A(\u_multiplier/_2505_ ),
    .B1(\u_multiplier/_2506_ ),
    .B2(\u_multiplier/_2492_ ),
    .ZN(\u_multiplier/_2514_ ));
 AND2_X1 \u_multiplier/_5101_  (.A1(\u_multiplier/K [0]),
    .A2(\u_multiplier/_2486_ ),
    .ZN(\u_multiplier/_2515_ ));
 MUX2_X1 \u_multiplier/_5102_  (.A(\u_multiplier/_2454_ ),
    .B(\u_multiplier/_2515_ ),
    .S(\u_multiplier/_3114_ ),
    .Z(\u_multiplier/_2516_ ));
 MUX2_X1 \u_multiplier/_5103_  (.A(\u_multiplier/_2391_ ),
    .B(\u_multiplier/_2516_ ),
    .S(\u_multiplier/_3112_ ),
    .Z(\u_multiplier/_2517_ ));
 MUX2_X2 \u_multiplier/_5104_  (.A(\u_multiplier/_2265_ ),
    .B(\u_multiplier/_2517_ ),
    .S(\u_multiplier/_3115_ ),
    .Z(\u_multiplier/_2518_ ));
 MUX2_X1 \u_multiplier/_5105_  (.A(\u_multiplier/_2009_ ),
    .B(\u_multiplier/_2518_ ),
    .S(\u_multiplier/_3116_ ),
    .Z(\u_multiplier/_2519_ ));
 NOR2_X1 \u_multiplier/_5106_  (.A1(\u_multiplier/dec_out [31]),
    .A2(\u_multiplier/_2519_ ),
    .ZN(\u_multiplier/_2520_ ));
 NAND2_X1 \u_multiplier/_5107_  (.A1(\u_multiplier/code_x [0]),
    .A2(\u_multiplier/_3131_ ),
    .ZN(\u_multiplier/_2521_ ));
 NOR2_X1 \u_multiplier/_5108_  (.A1(\u_multiplier/code_x [1]),
    .A2(\u_multiplier/_2521_ ),
    .ZN(\u_multiplier/_2522_ ));
 AOI21_X4 \u_multiplier/_5109_  (.A(\u_multiplier/_2522_ ),
    .B1(\u_multiplier/_2460_ ),
    .B2(\u_multiplier/code_x [1]),
    .ZN(\u_multiplier/_2523_ ));
 NOR2_X1 \u_multiplier/_5110_  (.A1(\u_multiplier/_3110_ ),
    .A2(\u_multiplier/_2398_ ),
    .ZN(\u_multiplier/_2524_ ));
 AOI21_X1 \u_multiplier/_5111_  (.A(\u_multiplier/_2524_ ),
    .B1(\u_multiplier/_2523_ ),
    .B2(\u_multiplier/_3110_ ),
    .ZN(\u_multiplier/_2525_ ));
 MUX2_X2 \u_multiplier/_5112_  (.A(\u_multiplier/_2272_ ),
    .B(\u_multiplier/_2525_ ),
    .S(\u_multiplier/_3111_ ),
    .Z(\u_multiplier/_2526_ ));
 NAND2_X1 \u_multiplier/_5113_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2015_ ),
    .ZN(\u_multiplier/_2527_ ));
 OAI21_X2 \u_multiplier/_5114_  (.A(\u_multiplier/_2527_ ),
    .B1(\u_multiplier/_2526_ ),
    .B2(\u_multiplier/code_x [4]),
    .ZN(\u_multiplier/_2528_ ));
 NOR3_X2 \u_multiplier/_5115_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_3105_ ),
    .A3(\u_multiplier/_3130_ ),
    .ZN(\u_multiplier/_2529_ ));
 AOI21_X4 \u_multiplier/_5116_  (.A(\u_multiplier/_2529_ ),
    .B1(\u_multiplier/_2467_ ),
    .B2(\u_multiplier/code_y [1]),
    .ZN(\u_multiplier/_2530_ ));
 NOR2_X1 \u_multiplier/_5117_  (.A1(\u_multiplier/_3106_ ),
    .A2(\u_multiplier/_2404_ ),
    .ZN(\u_multiplier/_2531_ ));
 AOI21_X2 \u_multiplier/_5118_  (.A(\u_multiplier/_2531_ ),
    .B1(\u_multiplier/_2530_ ),
    .B2(\u_multiplier/_3106_ ),
    .ZN(\u_multiplier/_2532_ ));
 MUX2_X2 \u_multiplier/_5119_  (.A(\u_multiplier/_2278_ ),
    .B(\u_multiplier/_2532_ ),
    .S(\u_multiplier/_3107_ ),
    .Z(\u_multiplier/_2533_ ));
 NAND2_X1 \u_multiplier/_5120_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_2021_ ),
    .ZN(\u_multiplier/_2534_ ));
 OAI21_X2 \u_multiplier/_5121_  (.A(\u_multiplier/_2534_ ),
    .B1(\u_multiplier/_2533_ ),
    .B2(\u_multiplier/code_y [4]),
    .ZN(\u_multiplier/_2535_ ));
 XOR2_X2 \u_multiplier/_5122_  (.A(\u_multiplier/_2528_ ),
    .B(\u_multiplier/_2535_ ),
    .Z(\u_multiplier/_2536_ ));
 OAI21_X1 \u_multiplier/_5123_  (.A(\u_multiplier/_2536_ ),
    .B1(\u_multiplier/_2519_ ),
    .B2(\u_multiplier/dec_out [31]),
    .ZN(\u_multiplier/_2537_ ));
 XNOR2_X2 \u_multiplier/_5124_  (.A(\u_multiplier/_2520_ ),
    .B(\u_multiplier/_2536_ ),
    .ZN(\u_multiplier/_2538_ ));
 NAND2_X1 \u_multiplier/_5125_  (.A1(\u_multiplier/_2514_ ),
    .A2(\u_multiplier/_2538_ ),
    .ZN(\u_multiplier/_2539_ ));
 NOR2_X1 \u_multiplier/_5126_  (.A1(\u_multiplier/_2514_ ),
    .A2(\u_multiplier/_2538_ ),
    .ZN(\u_multiplier/_2540_ ));
 XOR2_X2 \u_multiplier/_5127_  (.A(\u_multiplier/_2514_ ),
    .B(\u_multiplier/_2538_ ),
    .Z(\u_multiplier/_2541_ ));
 OAI21_X1 \u_multiplier/_5128_  (.A(net21),
    .B1(\u_multiplier/_2513_ ),
    .B2(\u_multiplier/_2541_ ),
    .ZN(\u_multiplier/_2542_ ));
 AOI21_X1 \u_multiplier/_5129_  (.A(\u_multiplier/_2542_ ),
    .B1(\u_multiplier/_2541_ ),
    .B2(\u_multiplier/_2513_ ),
    .ZN(product[31]));
 OAI211_X4 \u_multiplier/_5130_  (.A(\u_multiplier/_2510_ ),
    .B(\u_multiplier/_2541_ ),
    .C1(\u_multiplier/_2478_ ),
    .C2(\u_multiplier/_2483_ ),
    .ZN(\u_multiplier/_2543_ ));
 OAI21_X1 \u_multiplier/_5131_  (.A(\u_multiplier/_2539_ ),
    .B1(\u_multiplier/_2540_ ),
    .B2(\u_multiplier/_2508_ ),
    .ZN(\u_multiplier/_2544_ ));
 INV_X1 \u_multiplier/_5132_  (.A(\u_multiplier/_2544_ ),
    .ZN(\u_multiplier/_2545_ ));
 AND2_X1 \u_multiplier/_5133_  (.A1(\u_multiplier/_2543_ ),
    .A2(\u_multiplier/_2545_ ),
    .ZN(\u_multiplier/_2546_ ));
 OAI21_X2 \u_multiplier/_5134_  (.A(\u_multiplier/_2537_ ),
    .B1(\u_multiplier/_2535_ ),
    .B2(\u_multiplier/_2528_ ),
    .ZN(\u_multiplier/_2547_ ));
 AND2_X1 \u_multiplier/_5135_  (.A1(\u_multiplier/K [1]),
    .A2(\u_multiplier/_2487_ ),
    .ZN(\u_multiplier/_2548_ ));
 MUX2_X1 \u_multiplier/_5136_  (.A(\u_multiplier/_2424_ ),
    .B(\u_multiplier/_2548_ ),
    .S(\u_multiplier/_3112_ ),
    .Z(\u_multiplier/_2549_ ));
 MUX2_X2 \u_multiplier/_5137_  (.A(\u_multiplier/_2300_ ),
    .B(\u_multiplier/_2549_ ),
    .S(\u_multiplier/_3115_ ),
    .Z(\u_multiplier/_2550_ ));
 AOI21_X2 \u_multiplier/_5138_  (.A(\u_multiplier/dec_out [32]),
    .B1(\u_multiplier/_2550_ ),
    .B2(\u_multiplier/_3116_ ),
    .ZN(\u_multiplier/_2551_ ));
 OAI21_X4 \u_multiplier/_5139_  (.A(\u_multiplier/_2551_ ),
    .B1(\u_multiplier/_2039_ ),
    .B2(\u_multiplier/_3116_ ),
    .ZN(\u_multiplier/_2552_ ));
 AND2_X1 \u_multiplier/_5140_  (.A1(\u_multiplier/code_x [1]),
    .A2(\u_multiplier/_2493_ ),
    .ZN(\u_multiplier/_2553_ ));
 OR2_X1 \u_multiplier/_5141_  (.A1(\u_multiplier/_3110_ ),
    .A2(\u_multiplier/_2430_ ),
    .ZN(\u_multiplier/_2554_ ));
 OAI21_X2 \u_multiplier/_5142_  (.A(\u_multiplier/_2554_ ),
    .B1(\u_multiplier/_2553_ ),
    .B2(\u_multiplier/code_x [2]),
    .ZN(\u_multiplier/_2555_ ));
 NOR2_X1 \u_multiplier/_5143_  (.A1(\u_multiplier/_3111_ ),
    .A2(\u_multiplier/_2305_ ),
    .ZN(\u_multiplier/_2556_ ));
 AOI21_X2 \u_multiplier/_5144_  (.A(\u_multiplier/_2556_ ),
    .B1(\u_multiplier/_2555_ ),
    .B2(\u_multiplier/_3111_ ),
    .ZN(\u_multiplier/_2557_ ));
 NAND2_X1 \u_multiplier/_5145_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2047_ ),
    .ZN(\u_multiplier/_2558_ ));
 OAI21_X2 \u_multiplier/_5146_  (.A(\u_multiplier/_2558_ ),
    .B1(\u_multiplier/_2557_ ),
    .B2(\u_multiplier/code_x [4]),
    .ZN(\u_multiplier/_2559_ ));
 AND2_X2 \u_multiplier/_5147_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_2499_ ),
    .ZN(\u_multiplier/_2560_ ));
 OR2_X1 \u_multiplier/_5148_  (.A1(\u_multiplier/_3106_ ),
    .A2(\u_multiplier/_2437_ ),
    .ZN(\u_multiplier/_2561_ ));
 OAI21_X4 \u_multiplier/_5149_  (.A(\u_multiplier/_2561_ ),
    .B1(\u_multiplier/_2560_ ),
    .B2(\u_multiplier/code_y [2]),
    .ZN(\u_multiplier/_2562_ ));
 NOR2_X1 \u_multiplier/_5150_  (.A1(\u_multiplier/_3107_ ),
    .A2(\u_multiplier/_2311_ ),
    .ZN(\u_multiplier/_2563_ ));
 AOI21_X4 \u_multiplier/_5151_  (.A(\u_multiplier/_2563_ ),
    .B1(\u_multiplier/_2562_ ),
    .B2(\u_multiplier/_3107_ ),
    .ZN(\u_multiplier/_2564_ ));
 NAND2_X1 \u_multiplier/_5152_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_2053_ ),
    .ZN(\u_multiplier/_2565_ ));
 OAI21_X2 \u_multiplier/_5153_  (.A(\u_multiplier/_2565_ ),
    .B1(\u_multiplier/_2564_ ),
    .B2(\u_multiplier/code_y [4]),
    .ZN(\u_multiplier/_2566_ ));
 NOR2_X1 \u_multiplier/_5154_  (.A1(\u_multiplier/_2559_ ),
    .A2(\u_multiplier/_2566_ ),
    .ZN(\u_multiplier/_2567_ ));
 XOR2_X2 \u_multiplier/_5155_  (.A(\u_multiplier/_2559_ ),
    .B(\u_multiplier/_2566_ ),
    .Z(\u_multiplier/_2568_ ));
 XOR2_X2 \u_multiplier/_5156_  (.A(\u_multiplier/_2552_ ),
    .B(\u_multiplier/_2568_ ),
    .Z(\u_multiplier/_2569_ ));
 AND2_X1 \u_multiplier/_5157_  (.A1(\u_multiplier/_2547_ ),
    .A2(\u_multiplier/_2569_ ),
    .ZN(\u_multiplier/_2570_ ));
 XNOR2_X2 \u_multiplier/_5158_  (.A(\u_multiplier/_2547_ ),
    .B(\u_multiplier/_2569_ ),
    .ZN(\u_multiplier/_2571_ ));
 NOR2_X1 \u_multiplier/_5159_  (.A1(\u_multiplier/_2546_ ),
    .A2(\u_multiplier/_2571_ ),
    .ZN(\u_multiplier/_2572_ ));
 AND2_X1 \u_multiplier/_5160_  (.A1(\u_multiplier/_2546_ ),
    .A2(\u_multiplier/_2571_ ),
    .ZN(\u_multiplier/_2573_ ));
 NOR3_X1 \u_multiplier/_5161_  (.A1(\u_multiplier/_3334_ ),
    .A2(\u_multiplier/_2572_ ),
    .A3(\u_multiplier/_2573_ ),
    .ZN(product[32]));
 AOI21_X2 \u_multiplier/_5162_  (.A(\u_multiplier/_2567_ ),
    .B1(\u_multiplier/_2568_ ),
    .B2(\u_multiplier/_2552_ ),
    .ZN(\u_multiplier/_2574_ ));
 INV_X1 \u_multiplier/_5163_  (.A(\u_multiplier/_2574_ ),
    .ZN(\u_multiplier/_2575_ ));
 NAND2_X1 \u_multiplier/_5164_  (.A1(\u_multiplier/K [1]),
    .A2(\u_multiplier/_2515_ ),
    .ZN(\u_multiplier/_2576_ ));
 NAND2_X1 \u_multiplier/_5165_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/_2455_ ),
    .ZN(\u_multiplier/_2577_ ));
 OAI21_X2 \u_multiplier/_5166_  (.A(\u_multiplier/_2577_ ),
    .B1(\u_multiplier/_2576_ ),
    .B2(\u_multiplier/K [2]),
    .ZN(\u_multiplier/_2578_ ));
 MUX2_X2 \u_multiplier/_5167_  (.A(\u_multiplier/_2329_ ),
    .B(\u_multiplier/_2578_ ),
    .S(\u_multiplier/_3115_ ),
    .Z(\u_multiplier/_2579_ ));
 NOR2_X1 \u_multiplier/_5168_  (.A1(\u_multiplier/K [4]),
    .A2(\u_multiplier/_2579_ ),
    .ZN(\u_multiplier/_2580_ ));
 AOI21_X1 \u_multiplier/_5169_  (.A(\u_multiplier/_2580_ ),
    .B1(\u_multiplier/_2071_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2581_ ));
 NOR2_X1 \u_multiplier/_5170_  (.A1(\u_multiplier/dec_out [33]),
    .A2(\u_multiplier/_2581_ ),
    .ZN(\u_multiplier/_2582_ ));
 NAND3_X1 \u_multiplier/_5171_  (.A1(\u_multiplier/code_x [0]),
    .A2(\u_multiplier/code_x [1]),
    .A3(\u_multiplier/_3131_ ),
    .ZN(\u_multiplier/_2583_ ));
 NAND2_X1 \u_multiplier/_5172_  (.A1(\u_multiplier/_3110_ ),
    .A2(\u_multiplier/_2583_ ),
    .ZN(\u_multiplier/_2584_ ));
 OAI21_X2 \u_multiplier/_5173_  (.A(\u_multiplier/_2584_ ),
    .B1(\u_multiplier/_2461_ ),
    .B2(\u_multiplier/_3110_ ),
    .ZN(\u_multiplier/_2585_ ));
 NOR2_X1 \u_multiplier/_5174_  (.A1(\u_multiplier/_3111_ ),
    .A2(\u_multiplier/_2336_ ),
    .ZN(\u_multiplier/_2586_ ));
 AOI21_X2 \u_multiplier/_5175_  (.A(\u_multiplier/_2586_ ),
    .B1(\u_multiplier/_2585_ ),
    .B2(\u_multiplier/_3111_ ),
    .ZN(\u_multiplier/_2587_ ));
 OR2_X1 \u_multiplier/_5176_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2587_ ),
    .ZN(\u_multiplier/_2588_ ));
 OAI21_X2 \u_multiplier/_5177_  (.A(\u_multiplier/_2588_ ),
    .B1(\u_multiplier/_2078_ ),
    .B2(\u_multiplier/_3109_ ),
    .ZN(\u_multiplier/_2589_ ));
 NAND3_X1 \u_multiplier/_5178_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/code_y [0]),
    .A3(\u_multiplier/_3129_ ),
    .ZN(\u_multiplier/_2590_ ));
 NAND2_X1 \u_multiplier/_5179_  (.A1(\u_multiplier/_3106_ ),
    .A2(\u_multiplier/_2590_ ),
    .ZN(\u_multiplier/_2591_ ));
 OAI21_X4 \u_multiplier/_5180_  (.A(\u_multiplier/_2591_ ),
    .B1(\u_multiplier/_2468_ ),
    .B2(\u_multiplier/_3106_ ),
    .ZN(\u_multiplier/_2592_ ));
 NOR2_X1 \u_multiplier/_5181_  (.A1(\u_multiplier/_3107_ ),
    .A2(\u_multiplier/_2342_ ),
    .ZN(\u_multiplier/_2593_ ));
 AOI21_X4 \u_multiplier/_5182_  (.A(\u_multiplier/_2593_ ),
    .B1(\u_multiplier/_2592_ ),
    .B2(\u_multiplier/_3107_ ),
    .ZN(\u_multiplier/_2594_ ));
 NAND2_X1 \u_multiplier/_5183_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_2086_ ),
    .ZN(\u_multiplier/_2595_ ));
 OAI21_X2 \u_multiplier/_5184_  (.A(\u_multiplier/_2595_ ),
    .B1(\u_multiplier/_2594_ ),
    .B2(\u_multiplier/code_y [4]),
    .ZN(\u_multiplier/_2596_ ));
 XOR2_X2 \u_multiplier/_5185_  (.A(\u_multiplier/_2589_ ),
    .B(\u_multiplier/_2596_ ),
    .Z(\u_multiplier/_2597_ ));
 OAI21_X1 \u_multiplier/_5186_  (.A(\u_multiplier/_2597_ ),
    .B1(\u_multiplier/_2581_ ),
    .B2(\u_multiplier/dec_out [33]),
    .ZN(\u_multiplier/_2598_ ));
 XNOR2_X2 \u_multiplier/_5187_  (.A(\u_multiplier/_2582_ ),
    .B(\u_multiplier/_2597_ ),
    .ZN(\u_multiplier/_2599_ ));
 NAND2_X1 \u_multiplier/_5188_  (.A1(\u_multiplier/_2575_ ),
    .A2(\u_multiplier/_2599_ ),
    .ZN(\u_multiplier/_2600_ ));
 XNOR2_X2 \u_multiplier/_5189_  (.A(\u_multiplier/_2574_ ),
    .B(\u_multiplier/_2599_ ),
    .ZN(\u_multiplier/_2601_ ));
 INV_X1 \u_multiplier/_5190_  (.A(\u_multiplier/_2601_ ),
    .ZN(\u_multiplier/_2602_ ));
 AOI211_X2 \u_multiplier/_5191_  (.A(\u_multiplier/_2571_ ),
    .B(\u_multiplier/_2602_ ),
    .C1(\u_multiplier/_2543_ ),
    .C2(\u_multiplier/_2545_ ),
    .ZN(\u_multiplier/_2603_ ));
 NOR3_X2 \u_multiplier/_5192_  (.A1(\u_multiplier/_2570_ ),
    .A2(\u_multiplier/_2572_ ),
    .A3(\u_multiplier/_2601_ ),
    .ZN(\u_multiplier/_2604_ ));
 NAND2_X1 \u_multiplier/_5193_  (.A1(\u_multiplier/_2570_ ),
    .A2(\u_multiplier/_2601_ ),
    .ZN(\u_multiplier/_2605_ ));
 NAND2_X1 \u_multiplier/_5194_  (.A1(net21),
    .A2(\u_multiplier/_2605_ ),
    .ZN(\u_multiplier/_2606_ ));
 NOR3_X4 \u_multiplier/_5195_  (.A1(\u_multiplier/_2603_ ),
    .A2(\u_multiplier/_2604_ ),
    .A3(\u_multiplier/_2606_ ),
    .ZN(product[33]));
 NAND2_X1 \u_multiplier/_5196_  (.A1(\u_multiplier/_2600_ ),
    .A2(\u_multiplier/_2605_ ),
    .ZN(\u_multiplier/_2607_ ));
 OR2_X1 \u_multiplier/_5197_  (.A1(\u_multiplier/_2603_ ),
    .A2(\u_multiplier/_2607_ ),
    .ZN(\u_multiplier/_2608_ ));
 OAI21_X1 \u_multiplier/_5198_  (.A(\u_multiplier/_2598_ ),
    .B1(\u_multiplier/_2596_ ),
    .B2(\u_multiplier/_2589_ ),
    .ZN(\u_multiplier/_2609_ ));
 AND2_X1 \u_multiplier/_5199_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/_2488_ ),
    .ZN(\u_multiplier/_2610_ ));
 MUX2_X1 \u_multiplier/_5200_  (.A(\u_multiplier/_2363_ ),
    .B(\u_multiplier/_2610_ ),
    .S(\u_multiplier/_3115_ ),
    .Z(\u_multiplier/_2611_ ));
 NOR2_X1 \u_multiplier/_5201_  (.A1(\u_multiplier/K [4]),
    .A2(\u_multiplier/_2611_ ),
    .ZN(\u_multiplier/_2612_ ));
 AOI21_X1 \u_multiplier/_5202_  (.A(\u_multiplier/_2612_ ),
    .B1(\u_multiplier/_2106_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2613_ ));
 NOR2_X1 \u_multiplier/_5203_  (.A1(\u_multiplier/dec_out [34]),
    .A2(\u_multiplier/_2613_ ),
    .ZN(\u_multiplier/_2614_ ));
 AND2_X1 \u_multiplier/_5204_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_2494_ ),
    .ZN(\u_multiplier/_2615_ ));
 MUX2_X1 \u_multiplier/_5205_  (.A(\u_multiplier/_2369_ ),
    .B(\u_multiplier/_2615_ ),
    .S(\u_multiplier/_3111_ ),
    .Z(\u_multiplier/_2616_ ));
 NAND2_X1 \u_multiplier/_5206_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2114_ ),
    .ZN(\u_multiplier/_2617_ ));
 OAI21_X2 \u_multiplier/_5207_  (.A(\u_multiplier/_2617_ ),
    .B1(\u_multiplier/_2616_ ),
    .B2(\u_multiplier/code_x [4]),
    .ZN(\u_multiplier/_2618_ ));
 AND2_X1 \u_multiplier/_5208_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_2500_ ),
    .ZN(\u_multiplier/_2619_ ));
 MUX2_X2 \u_multiplier/_5209_  (.A(\u_multiplier/_2375_ ),
    .B(\u_multiplier/_2619_ ),
    .S(\u_multiplier/_3107_ ),
    .Z(\u_multiplier/_2620_ ));
 NAND2_X1 \u_multiplier/_5210_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_2121_ ),
    .ZN(\u_multiplier/_2621_ ));
 OAI21_X2 \u_multiplier/_5211_  (.A(\u_multiplier/_2621_ ),
    .B1(\u_multiplier/_2620_ ),
    .B2(\u_multiplier/code_y [4]),
    .ZN(\u_multiplier/_2622_ ));
 XOR2_X2 \u_multiplier/_5212_  (.A(\u_multiplier/_2618_ ),
    .B(\u_multiplier/_2622_ ),
    .Z(\u_multiplier/_2623_ ));
 OAI21_X1 \u_multiplier/_5213_  (.A(\u_multiplier/_2623_ ),
    .B1(\u_multiplier/_2613_ ),
    .B2(\u_multiplier/dec_out [34]),
    .ZN(\u_multiplier/_2624_ ));
 XNOR2_X2 \u_multiplier/_5214_  (.A(\u_multiplier/_2614_ ),
    .B(\u_multiplier/_2623_ ),
    .ZN(\u_multiplier/_2625_ ));
 AND2_X1 \u_multiplier/_5215_  (.A1(\u_multiplier/_2609_ ),
    .A2(\u_multiplier/_2625_ ),
    .ZN(\u_multiplier/_2626_ ));
 XOR2_X2 \u_multiplier/_5216_  (.A(\u_multiplier/_2609_ ),
    .B(\u_multiplier/_2625_ ),
    .Z(\u_multiplier/_2627_ ));
 AND2_X1 \u_multiplier/_5217_  (.A1(\u_multiplier/_2608_ ),
    .A2(\u_multiplier/_2627_ ),
    .ZN(\u_multiplier/_2628_ ));
 OAI21_X2 \u_multiplier/_5218_  (.A(net21),
    .B1(\u_multiplier/_2608_ ),
    .B2(\u_multiplier/_2627_ ),
    .ZN(\u_multiplier/_2629_ ));
 NOR2_X4 \u_multiplier/_5219_  (.A1(\u_multiplier/_2628_ ),
    .A2(\u_multiplier/_2629_ ),
    .ZN(product[34]));
 OR2_X2 \u_multiplier/_5220_  (.A1(\u_multiplier/_2626_ ),
    .A2(\u_multiplier/_2628_ ),
    .ZN(\u_multiplier/_2630_ ));
 OAI21_X2 \u_multiplier/_5221_  (.A(\u_multiplier/_2624_ ),
    .B1(\u_multiplier/_2622_ ),
    .B2(\u_multiplier/_2618_ ),
    .ZN(\u_multiplier/_2631_ ));
 AND2_X1 \u_multiplier/_5222_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/_2516_ ),
    .ZN(\u_multiplier/_2632_ ));
 MUX2_X2 \u_multiplier/_5223_  (.A(\u_multiplier/_2392_ ),
    .B(\u_multiplier/_2632_ ),
    .S(\u_multiplier/_3115_ ),
    .Z(\u_multiplier/_2633_ ));
 NOR2_X1 \u_multiplier/_5224_  (.A1(\u_multiplier/_3116_ ),
    .A2(\u_multiplier/_2142_ ),
    .ZN(\u_multiplier/_2634_ ));
 AOI211_X2 \u_multiplier/_5225_  (.A(\u_multiplier/dec_out [35]),
    .B(\u_multiplier/_2634_ ),
    .C1(\u_multiplier/_2633_ ),
    .C2(\u_multiplier/_3116_ ),
    .ZN(\u_multiplier/_2635_ ));
 NOR2_X1 \u_multiplier/_5226_  (.A1(\u_multiplier/_3110_ ),
    .A2(\u_multiplier/_2523_ ),
    .ZN(\u_multiplier/_2636_ ));
 MUX2_X1 \u_multiplier/_5227_  (.A(\u_multiplier/_2399_ ),
    .B(\u_multiplier/_2636_ ),
    .S(\u_multiplier/_3111_ ),
    .Z(\u_multiplier/_2637_ ));
 MUX2_X1 \u_multiplier/_5228_  (.A(\u_multiplier/_2148_ ),
    .B(\u_multiplier/_2637_ ),
    .S(\u_multiplier/_3109_ ),
    .Z(\u_multiplier/_2638_ ));
 NOR2_X1 \u_multiplier/_5229_  (.A1(\u_multiplier/_3106_ ),
    .A2(\u_multiplier/_2530_ ),
    .ZN(\u_multiplier/_2639_ ));
 MUX2_X1 \u_multiplier/_5230_  (.A(\u_multiplier/_2405_ ),
    .B(\u_multiplier/_2639_ ),
    .S(\u_multiplier/_3107_ ),
    .Z(\u_multiplier/_2640_ ));
 MUX2_X1 \u_multiplier/_5231_  (.A(\u_multiplier/_2155_ ),
    .B(\u_multiplier/_2640_ ),
    .S(\u_multiplier/_3108_ ),
    .Z(\u_multiplier/_2641_ ));
 NAND2_X1 \u_multiplier/_5232_  (.A1(\u_multiplier/_2638_ ),
    .A2(\u_multiplier/_2641_ ),
    .ZN(\u_multiplier/_2642_ ));
 XNOR2_X2 \u_multiplier/_5233_  (.A(\u_multiplier/_2638_ ),
    .B(\u_multiplier/_2641_ ),
    .ZN(\u_multiplier/_2643_ ));
 XOR2_X2 \u_multiplier/_5234_  (.A(\u_multiplier/_2635_ ),
    .B(\u_multiplier/_2643_ ),
    .Z(\u_multiplier/_2644_ ));
 NAND2_X1 \u_multiplier/_5235_  (.A1(\u_multiplier/_2631_ ),
    .A2(\u_multiplier/_2644_ ),
    .ZN(\u_multiplier/_2645_ ));
 XOR2_X2 \u_multiplier/_5236_  (.A(\u_multiplier/_2631_ ),
    .B(\u_multiplier/_2644_ ),
    .Z(\u_multiplier/_2646_ ));
 OAI21_X2 \u_multiplier/_5237_  (.A(net21),
    .B1(\u_multiplier/_2630_ ),
    .B2(\u_multiplier/_2646_ ),
    .ZN(\u_multiplier/_2647_ ));
 AOI21_X4 \u_multiplier/_5238_  (.A(\u_multiplier/_2647_ ),
    .B1(\u_multiplier/_2646_ ),
    .B2(\u_multiplier/_2630_ ),
    .ZN(product[35]));
 OAI211_X2 \u_multiplier/_5239_  (.A(\u_multiplier/_2627_ ),
    .B(\u_multiplier/_2646_ ),
    .C1(\u_multiplier/_2603_ ),
    .C2(\u_multiplier/_2607_ ),
    .ZN(\u_multiplier/_2648_ ));
 OAI21_X1 \u_multiplier/_5240_  (.A(\u_multiplier/_2626_ ),
    .B1(\u_multiplier/_2631_ ),
    .B2(\u_multiplier/_2644_ ),
    .ZN(\u_multiplier/_2649_ ));
 NAND2_X1 \u_multiplier/_5241_  (.A1(\u_multiplier/_2645_ ),
    .A2(\u_multiplier/_2649_ ),
    .ZN(\u_multiplier/_2650_ ));
 INV_X1 \u_multiplier/_5242_  (.A(\u_multiplier/_2650_ ),
    .ZN(\u_multiplier/_2651_ ));
 AND2_X1 \u_multiplier/_5243_  (.A1(\u_multiplier/_2648_ ),
    .A2(\u_multiplier/_2651_ ),
    .ZN(\u_multiplier/_2652_ ));
 OAI21_X2 \u_multiplier/_5244_  (.A(\u_multiplier/_2642_ ),
    .B1(\u_multiplier/_2643_ ),
    .B2(\u_multiplier/_2635_ ),
    .ZN(\u_multiplier/_2653_ ));
 AND2_X1 \u_multiplier/_5245_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/_2548_ ),
    .ZN(\u_multiplier/_2654_ ));
 MUX2_X2 \u_multiplier/_5246_  (.A(\u_multiplier/_2425_ ),
    .B(\u_multiplier/_2654_ ),
    .S(\u_multiplier/_3115_ ),
    .Z(\u_multiplier/_2655_ ));
 NOR2_X1 \u_multiplier/_5247_  (.A1(\u_multiplier/_3116_ ),
    .A2(\u_multiplier/_2172_ ),
    .ZN(\u_multiplier/_2656_ ));
 AOI211_X2 \u_multiplier/_5248_  (.A(\u_multiplier/dec_out [36]),
    .B(\u_multiplier/_2656_ ),
    .C1(\u_multiplier/_2655_ ),
    .C2(\u_multiplier/_3116_ ),
    .ZN(\u_multiplier/_2657_ ));
 INV_X1 \u_multiplier/_5249_  (.A(\u_multiplier/_2657_ ),
    .ZN(\u_multiplier/_2658_ ));
 NAND2_X1 \u_multiplier/_5250_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_2553_ ),
    .ZN(\u_multiplier/_2659_ ));
 NOR2_X1 \u_multiplier/_5251_  (.A1(\u_multiplier/_3111_ ),
    .A2(\u_multiplier/_2431_ ),
    .ZN(\u_multiplier/_2660_ ));
 AOI21_X2 \u_multiplier/_5252_  (.A(\u_multiplier/_2660_ ),
    .B1(\u_multiplier/_2659_ ),
    .B2(\u_multiplier/_3111_ ),
    .ZN(\u_multiplier/_2661_ ));
 NAND2_X1 \u_multiplier/_5253_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2179_ ),
    .ZN(\u_multiplier/_2662_ ));
 OAI21_X2 \u_multiplier/_5254_  (.A(\u_multiplier/_2662_ ),
    .B1(\u_multiplier/_2661_ ),
    .B2(\u_multiplier/code_x [4]),
    .ZN(\u_multiplier/_2663_ ));
 AOI21_X1 \u_multiplier/_5255_  (.A(\u_multiplier/code_y [3]),
    .B1(\u_multiplier/_2560_ ),
    .B2(\u_multiplier/code_y [2]),
    .ZN(\u_multiplier/_2664_ ));
 NOR2_X1 \u_multiplier/_5256_  (.A1(\u_multiplier/_3107_ ),
    .A2(\u_multiplier/_2438_ ),
    .ZN(\u_multiplier/_2665_ ));
 NOR2_X2 \u_multiplier/_5257_  (.A1(\u_multiplier/_2664_ ),
    .A2(\u_multiplier/_2665_ ),
    .ZN(\u_multiplier/_2666_ ));
 NAND2_X1 \u_multiplier/_5258_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_2185_ ),
    .ZN(\u_multiplier/_2667_ ));
 OAI21_X2 \u_multiplier/_5259_  (.A(\u_multiplier/_2667_ ),
    .B1(\u_multiplier/_2666_ ),
    .B2(\u_multiplier/code_y [4]),
    .ZN(\u_multiplier/_2668_ ));
 NOR2_X1 \u_multiplier/_5260_  (.A1(\u_multiplier/_2663_ ),
    .A2(\u_multiplier/_2668_ ),
    .ZN(\u_multiplier/_2669_ ));
 XOR2_X2 \u_multiplier/_5261_  (.A(\u_multiplier/_2663_ ),
    .B(\u_multiplier/_2668_ ),
    .Z(\u_multiplier/_2670_ ));
 XNOR2_X2 \u_multiplier/_5262_  (.A(\u_multiplier/_2657_ ),
    .B(\u_multiplier/_2670_ ),
    .ZN(\u_multiplier/_2671_ ));
 NAND2_X1 \u_multiplier/_5263_  (.A1(\u_multiplier/_2653_ ),
    .A2(\u_multiplier/_2671_ ),
    .ZN(\u_multiplier/_2672_ ));
 XNOR2_X2 \u_multiplier/_5264_  (.A(\u_multiplier/_2653_ ),
    .B(\u_multiplier/_2671_ ),
    .ZN(\u_multiplier/_2673_ ));
 NOR2_X1 \u_multiplier/_5265_  (.A1(\u_multiplier/_2652_ ),
    .A2(\u_multiplier/_2673_ ),
    .ZN(\u_multiplier/_2674_ ));
 AND2_X1 \u_multiplier/_5266_  (.A1(\u_multiplier/_2652_ ),
    .A2(\u_multiplier/_2673_ ),
    .ZN(\u_multiplier/_2675_ ));
 NOR3_X2 \u_multiplier/_5267_  (.A1(\u_multiplier/_3334_ ),
    .A2(\u_multiplier/_2674_ ),
    .A3(\u_multiplier/_2675_ ),
    .ZN(product[36]));
 AOI21_X2 \u_multiplier/_5268_  (.A(\u_multiplier/_2669_ ),
    .B1(\u_multiplier/_2670_ ),
    .B2(\u_multiplier/_2658_ ),
    .ZN(\u_multiplier/_2676_ ));
 INV_X1 \u_multiplier/_5269_  (.A(\u_multiplier/_2676_ ),
    .ZN(\u_multiplier/_2677_ ));
 NOR2_X2 \u_multiplier/_5270_  (.A1(\u_multiplier/_3112_ ),
    .A2(\u_multiplier/_2576_ ),
    .ZN(\u_multiplier/_2678_ ));
 MUX2_X1 \u_multiplier/_5271_  (.A(\u_multiplier/_2456_ ),
    .B(\u_multiplier/_2678_ ),
    .S(\u_multiplier/_3115_ ),
    .Z(\u_multiplier/_2679_ ));
 MUX2_X1 \u_multiplier/_5272_  (.A(\u_multiplier/_2203_ ),
    .B(\u_multiplier/_2679_ ),
    .S(\u_multiplier/_3116_ ),
    .Z(\u_multiplier/_2680_ ));
 NOR2_X1 \u_multiplier/_5273_  (.A1(\u_multiplier/dec_out [37]),
    .A2(\u_multiplier/_2680_ ),
    .ZN(\u_multiplier/_2681_ ));
 OR2_X1 \u_multiplier/_5274_  (.A1(\u_multiplier/_3110_ ),
    .A2(\u_multiplier/_2583_ ),
    .ZN(\u_multiplier/_2682_ ));
 NOR2_X1 \u_multiplier/_5275_  (.A1(\u_multiplier/_3111_ ),
    .A2(\u_multiplier/_2462_ ),
    .ZN(\u_multiplier/_2683_ ));
 AOI21_X2 \u_multiplier/_5276_  (.A(\u_multiplier/_2683_ ),
    .B1(\u_multiplier/_2682_ ),
    .B2(\u_multiplier/_3111_ ),
    .ZN(\u_multiplier/_2684_ ));
 NAND2_X1 \u_multiplier/_5277_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2210_ ),
    .ZN(\u_multiplier/_2685_ ));
 OAI21_X2 \u_multiplier/_5278_  (.A(\u_multiplier/_2685_ ),
    .B1(\u_multiplier/_2684_ ),
    .B2(\u_multiplier/code_x [4]),
    .ZN(\u_multiplier/_2686_ ));
 OR2_X1 \u_multiplier/_5279_  (.A1(\u_multiplier/_3106_ ),
    .A2(\u_multiplier/_2590_ ),
    .ZN(\u_multiplier/_2687_ ));
 NOR2_X1 \u_multiplier/_5280_  (.A1(\u_multiplier/_3107_ ),
    .A2(\u_multiplier/_2469_ ),
    .ZN(\u_multiplier/_2688_ ));
 AOI21_X2 \u_multiplier/_5281_  (.A(\u_multiplier/_2688_ ),
    .B1(\u_multiplier/_2687_ ),
    .B2(\u_multiplier/_3107_ ),
    .ZN(\u_multiplier/_2689_ ));
 NAND2_X1 \u_multiplier/_5282_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_2216_ ),
    .ZN(\u_multiplier/_2690_ ));
 OAI21_X2 \u_multiplier/_5283_  (.A(\u_multiplier/_2690_ ),
    .B1(\u_multiplier/_2689_ ),
    .B2(\u_multiplier/code_y [4]),
    .ZN(\u_multiplier/_2691_ ));
 XOR2_X2 \u_multiplier/_5284_  (.A(\u_multiplier/_2686_ ),
    .B(\u_multiplier/_2691_ ),
    .Z(\u_multiplier/_2692_ ));
 OAI21_X1 \u_multiplier/_5285_  (.A(\u_multiplier/_2692_ ),
    .B1(\u_multiplier/_2680_ ),
    .B2(\u_multiplier/dec_out [37]),
    .ZN(\u_multiplier/_2693_ ));
 XNOR2_X2 \u_multiplier/_5286_  (.A(\u_multiplier/_2681_ ),
    .B(\u_multiplier/_2692_ ),
    .ZN(\u_multiplier/_2694_ ));
 NAND2_X1 \u_multiplier/_5287_  (.A1(\u_multiplier/_2677_ ),
    .A2(\u_multiplier/_2694_ ),
    .ZN(\u_multiplier/_2695_ ));
 XOR2_X2 \u_multiplier/_5288_  (.A(\u_multiplier/_2676_ ),
    .B(\u_multiplier/_2694_ ),
    .Z(\u_multiplier/_2696_ ));
 NAND2_X1 \u_multiplier/_5289_  (.A1(\u_multiplier/_2672_ ),
    .A2(\u_multiplier/_2696_ ),
    .ZN(\u_multiplier/_2697_ ));
 AOI211_X2 \u_multiplier/_5290_  (.A(\u_multiplier/_2673_ ),
    .B(\u_multiplier/_2696_ ),
    .C1(\u_multiplier/_2648_ ),
    .C2(\u_multiplier/_2651_ ),
    .ZN(\u_multiplier/_2698_ ));
 OR2_X1 \u_multiplier/_5291_  (.A1(\u_multiplier/_2672_ ),
    .A2(\u_multiplier/_2696_ ),
    .ZN(\u_multiplier/_2699_ ));
 OAI21_X1 \u_multiplier/_5292_  (.A(\u_multiplier/_2699_ ),
    .B1(\u_multiplier/_2697_ ),
    .B2(\u_multiplier/_2674_ ),
    .ZN(\u_multiplier/_2700_ ));
 NOR3_X2 \u_multiplier/_5293_  (.A1(\u_multiplier/_3334_ ),
    .A2(\u_multiplier/_2698_ ),
    .A3(\u_multiplier/_2700_ ),
    .ZN(product[37]));
 NAND2_X2 \u_multiplier/_5294_  (.A1(\u_multiplier/_2695_ ),
    .A2(\u_multiplier/_2699_ ),
    .ZN(\u_multiplier/_2701_ ));
 OR2_X1 \u_multiplier/_5295_  (.A1(\u_multiplier/_2698_ ),
    .A2(\u_multiplier/_2701_ ),
    .ZN(\u_multiplier/_2702_ ));
 OAI21_X2 \u_multiplier/_5296_  (.A(\u_multiplier/_2693_ ),
    .B1(\u_multiplier/_2691_ ),
    .B2(\u_multiplier/_2686_ ),
    .ZN(\u_multiplier/_2703_ ));
 INV_X1 \u_multiplier/_5297_  (.A(\u_multiplier/_2703_ ),
    .ZN(\u_multiplier/_2704_ ));
 NAND2_X2 \u_multiplier/_5298_  (.A1(\u_multiplier/K [3]),
    .A2(\u_multiplier/_2489_ ),
    .ZN(\u_multiplier/_2705_ ));
 NOR2_X1 \u_multiplier/_5299_  (.A1(\u_multiplier/K [4]),
    .A2(\u_multiplier/_2705_ ),
    .ZN(\u_multiplier/_2706_ ));
 NOR2_X1 \u_multiplier/_5300_  (.A1(\u_multiplier/dec_out [38]),
    .A2(\u_multiplier/_2706_ ),
    .ZN(\u_multiplier/_2707_ ));
 OAI21_X2 \u_multiplier/_5301_  (.A(\u_multiplier/_2707_ ),
    .B1(\u_multiplier/_2236_ ),
    .B2(\u_multiplier/_3116_ ),
    .ZN(\u_multiplier/_2708_ ));
 AND2_X1 \u_multiplier/_5302_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_2495_ ),
    .ZN(\u_multiplier/_2709_ ));
 NAND2_X1 \u_multiplier/_5303_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2243_ ),
    .ZN(\u_multiplier/_2710_ ));
 OAI21_X2 \u_multiplier/_5304_  (.A(\u_multiplier/_2710_ ),
    .B1(\u_multiplier/_2709_ ),
    .B2(\u_multiplier/code_x [4]),
    .ZN(\u_multiplier/_2711_ ));
 AND2_X1 \u_multiplier/_5305_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_2501_ ),
    .ZN(\u_multiplier/_2712_ ));
 NAND2_X1 \u_multiplier/_5306_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_2249_ ),
    .ZN(\u_multiplier/_2713_ ));
 OAI21_X2 \u_multiplier/_5307_  (.A(\u_multiplier/_2713_ ),
    .B1(\u_multiplier/_2712_ ),
    .B2(\u_multiplier/code_y [4]),
    .ZN(\u_multiplier/_2714_ ));
 NOR2_X1 \u_multiplier/_5308_  (.A1(\u_multiplier/_2711_ ),
    .A2(\u_multiplier/_2714_ ),
    .ZN(\u_multiplier/_2715_ ));
 XOR2_X2 \u_multiplier/_5309_  (.A(\u_multiplier/_2711_ ),
    .B(\u_multiplier/_2714_ ),
    .Z(\u_multiplier/_2716_ ));
 XNOR2_X2 \u_multiplier/_5310_  (.A(\u_multiplier/_2708_ ),
    .B(\u_multiplier/_2716_ ),
    .ZN(\u_multiplier/_2717_ ));
 NOR2_X2 \u_multiplier/_5311_  (.A1(\u_multiplier/_2704_ ),
    .A2(\u_multiplier/_2717_ ),
    .ZN(\u_multiplier/_2718_ ));
 XNOR2_X2 \u_multiplier/_5312_  (.A(\u_multiplier/_2703_ ),
    .B(\u_multiplier/_2717_ ),
    .ZN(\u_multiplier/_2719_ ));
 AND2_X1 \u_multiplier/_5313_  (.A1(\u_multiplier/_2702_ ),
    .A2(\u_multiplier/_2719_ ),
    .ZN(\u_multiplier/_2720_ ));
 OAI21_X1 \u_multiplier/_5314_  (.A(net21),
    .B1(\u_multiplier/_2702_ ),
    .B2(\u_multiplier/_2719_ ),
    .ZN(\u_multiplier/_2721_ ));
 NOR2_X2 \u_multiplier/_5315_  (.A1(\u_multiplier/_2720_ ),
    .A2(\u_multiplier/_2721_ ),
    .ZN(product[38]));
 NOR2_X2 \u_multiplier/_5316_  (.A1(\u_multiplier/_2718_ ),
    .A2(\u_multiplier/_2720_ ),
    .ZN(\u_multiplier/_2722_ ));
 AOI21_X2 \u_multiplier/_5317_  (.A(\u_multiplier/_2715_ ),
    .B1(\u_multiplier/_2716_ ),
    .B2(\u_multiplier/_2708_ ),
    .ZN(\u_multiplier/_2723_ ));
 OR2_X1 \u_multiplier/_5318_  (.A1(\u_multiplier/_3116_ ),
    .A2(\u_multiplier/_2267_ ),
    .ZN(\u_multiplier/_2724_ ));
 NAND2_X2 \u_multiplier/_5319_  (.A1(\u_multiplier/K [3]),
    .A2(\u_multiplier/_2517_ ),
    .ZN(\u_multiplier/_2725_ ));
 NOR2_X1 \u_multiplier/_5320_  (.A1(\u_multiplier/K [4]),
    .A2(\u_multiplier/_2725_ ),
    .ZN(\u_multiplier/_2726_ ));
 NOR2_X1 \u_multiplier/_5321_  (.A1(\u_multiplier/dec_out [39]),
    .A2(\u_multiplier/_2726_ ),
    .ZN(\u_multiplier/_2727_ ));
 AND2_X1 \u_multiplier/_5322_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_2525_ ),
    .ZN(\u_multiplier/_2728_ ));
 MUX2_X1 \u_multiplier/_5323_  (.A(\u_multiplier/_2273_ ),
    .B(\u_multiplier/_2728_ ),
    .S(\u_multiplier/_3109_ ),
    .Z(\u_multiplier/_2729_ ));
 AND2_X1 \u_multiplier/_5324_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_2532_ ),
    .ZN(\u_multiplier/_2730_ ));
 MUX2_X1 \u_multiplier/_5325_  (.A(\u_multiplier/_2280_ ),
    .B(\u_multiplier/_2730_ ),
    .S(\u_multiplier/_3108_ ),
    .Z(\u_multiplier/_2731_ ));
 XNOR2_X1 \u_multiplier/_5326_  (.A(\u_multiplier/_2729_ ),
    .B(\u_multiplier/_2731_ ),
    .ZN(\u_multiplier/_2732_ ));
 AOI21_X2 \u_multiplier/_5327_  (.A(\u_multiplier/_2732_ ),
    .B1(\u_multiplier/_2727_ ),
    .B2(\u_multiplier/_2724_ ),
    .ZN(\u_multiplier/_2733_ ));
 AND3_X1 \u_multiplier/_5328_  (.A1(\u_multiplier/_2724_ ),
    .A2(\u_multiplier/_2727_ ),
    .A3(\u_multiplier/_2732_ ),
    .ZN(\u_multiplier/_2734_ ));
 OR2_X1 \u_multiplier/_5329_  (.A1(\u_multiplier/_2733_ ),
    .A2(\u_multiplier/_2734_ ),
    .ZN(\u_multiplier/_2735_ ));
 NOR2_X1 \u_multiplier/_5330_  (.A1(\u_multiplier/_2723_ ),
    .A2(\u_multiplier/_2735_ ),
    .ZN(\u_multiplier/_2736_ ));
 NAND2_X1 \u_multiplier/_5331_  (.A1(\u_multiplier/_2723_ ),
    .A2(\u_multiplier/_2735_ ),
    .ZN(\u_multiplier/_2737_ ));
 XNOR2_X2 \u_multiplier/_5332_  (.A(\u_multiplier/_2723_ ),
    .B(\u_multiplier/_2735_ ),
    .ZN(\u_multiplier/_2738_ ));
 INV_X1 \u_multiplier/_5333_  (.A(\u_multiplier/_2738_ ),
    .ZN(\u_multiplier/_2739_ ));
 OAI21_X2 \u_multiplier/_5334_  (.A(net21),
    .B1(\u_multiplier/_2722_ ),
    .B2(\u_multiplier/_2738_ ),
    .ZN(\u_multiplier/_2740_ ));
 AOI21_X4 \u_multiplier/_5335_  (.A(\u_multiplier/_2740_ ),
    .B1(\u_multiplier/_2738_ ),
    .B2(\u_multiplier/_2722_ ),
    .ZN(product[39]));
 OAI211_X4 \u_multiplier/_5336_  (.A(\u_multiplier/_2719_ ),
    .B(\u_multiplier/_2739_ ),
    .C1(\u_multiplier/_2698_ ),
    .C2(\u_multiplier/_2701_ ),
    .ZN(\u_multiplier/_2741_ ));
 AOI21_X4 \u_multiplier/_5337_  (.A(\u_multiplier/_2736_ ),
    .B1(\u_multiplier/_2737_ ),
    .B2(\u_multiplier/_2718_ ),
    .ZN(\u_multiplier/_2742_ ));
 NAND2_X1 \u_multiplier/_5338_  (.A1(\u_multiplier/_2741_ ),
    .A2(\u_multiplier/_2742_ ),
    .ZN(\u_multiplier/_2743_ ));
 AOI21_X2 \u_multiplier/_5339_  (.A(\u_multiplier/_2733_ ),
    .B1(\u_multiplier/_2731_ ),
    .B2(\u_multiplier/_2729_ ),
    .ZN(\u_multiplier/_2744_ ));
 NAND2_X2 \u_multiplier/_5340_  (.A1(\u_multiplier/K [3]),
    .A2(\u_multiplier/_2549_ ),
    .ZN(\u_multiplier/_2745_ ));
 AOI21_X1 \u_multiplier/_5341_  (.A(\u_multiplier/dec_out [40]),
    .B1(\u_multiplier/_2301_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2746_ ));
 OAI21_X2 \u_multiplier/_5342_  (.A(\u_multiplier/_2746_ ),
    .B1(\u_multiplier/_2745_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2747_ ));
 INV_X1 \u_multiplier/_5343_  (.A(\u_multiplier/_2747_ ),
    .ZN(\u_multiplier/_2748_ ));
 NOR2_X1 \u_multiplier/_5344_  (.A1(\u_multiplier/_3111_ ),
    .A2(\u_multiplier/_2555_ ),
    .ZN(\u_multiplier/_2749_ ));
 MUX2_X1 \u_multiplier/_5345_  (.A(\u_multiplier/_2306_ ),
    .B(\u_multiplier/_2749_ ),
    .S(\u_multiplier/_3109_ ),
    .Z(\u_multiplier/_2750_ ));
 NOR2_X2 \u_multiplier/_5346_  (.A1(\u_multiplier/_3107_ ),
    .A2(\u_multiplier/_2562_ ),
    .ZN(\u_multiplier/_2751_ ));
 MUX2_X1 \u_multiplier/_5347_  (.A(\u_multiplier/_2312_ ),
    .B(\u_multiplier/_2751_ ),
    .S(\u_multiplier/_3108_ ),
    .Z(\u_multiplier/_2752_ ));
 XNOR2_X2 \u_multiplier/_5348_  (.A(\u_multiplier/_2750_ ),
    .B(\u_multiplier/_2752_ ),
    .ZN(\u_multiplier/_2753_ ));
 NOR2_X1 \u_multiplier/_5349_  (.A1(\u_multiplier/_2748_ ),
    .A2(\u_multiplier/_2753_ ),
    .ZN(\u_multiplier/_2754_ ));
 XOR2_X2 \u_multiplier/_5350_  (.A(\u_multiplier/_2747_ ),
    .B(\u_multiplier/_2753_ ),
    .Z(\u_multiplier/_2755_ ));
 NOR2_X1 \u_multiplier/_5351_  (.A1(\u_multiplier/_2744_ ),
    .A2(\u_multiplier/_2755_ ),
    .ZN(\u_multiplier/_2756_ ));
 XOR2_X2 \u_multiplier/_5352_  (.A(\u_multiplier/_2744_ ),
    .B(\u_multiplier/_2755_ ),
    .Z(\u_multiplier/_2757_ ));
 INV_X1 \u_multiplier/_5353_  (.A(\u_multiplier/_2757_ ),
    .ZN(\u_multiplier/_2758_ ));
 AOI21_X4 \u_multiplier/_5354_  (.A(\u_multiplier/_2758_ ),
    .B1(\u_multiplier/_2742_ ),
    .B2(\u_multiplier/_2741_ ),
    .ZN(\u_multiplier/_2759_ ));
 OAI21_X2 \u_multiplier/_5355_  (.A(net21),
    .B1(\u_multiplier/_2743_ ),
    .B2(\u_multiplier/_2757_ ),
    .ZN(\u_multiplier/_2760_ ));
 NOR2_X4 \u_multiplier/_5356_  (.A1(\u_multiplier/_2759_ ),
    .A2(\u_multiplier/_2760_ ),
    .ZN(product[40]));
 AOI21_X2 \u_multiplier/_5357_  (.A(\u_multiplier/_2754_ ),
    .B1(\u_multiplier/_2752_ ),
    .B2(\u_multiplier/_2750_ ),
    .ZN(\u_multiplier/_2761_ ));
 NAND2_X2 \u_multiplier/_5358_  (.A1(\u_multiplier/K [3]),
    .A2(\u_multiplier/_2578_ ),
    .ZN(\u_multiplier/_2762_ ));
 AOI21_X1 \u_multiplier/_5359_  (.A(\u_multiplier/dec_out [41]),
    .B1(\u_multiplier/_2331_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2763_ ));
 OAI21_X2 \u_multiplier/_5360_  (.A(\u_multiplier/_2763_ ),
    .B1(\u_multiplier/_2762_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2764_ ));
 INV_X1 \u_multiplier/_5361_  (.A(\u_multiplier/_2764_ ),
    .ZN(\u_multiplier/_2765_ ));
 NOR2_X1 \u_multiplier/_5362_  (.A1(\u_multiplier/_3111_ ),
    .A2(\u_multiplier/_2585_ ),
    .ZN(\u_multiplier/_2766_ ));
 MUX2_X1 \u_multiplier/_5363_  (.A(\u_multiplier/_2337_ ),
    .B(\u_multiplier/_2766_ ),
    .S(\u_multiplier/_3109_ ),
    .Z(\u_multiplier/_2767_ ));
 NOR2_X2 \u_multiplier/_5364_  (.A1(\u_multiplier/_3107_ ),
    .A2(\u_multiplier/_2592_ ),
    .ZN(\u_multiplier/_2768_ ));
 MUX2_X1 \u_multiplier/_5365_  (.A(\u_multiplier/_2343_ ),
    .B(\u_multiplier/_2768_ ),
    .S(\u_multiplier/_3108_ ),
    .Z(\u_multiplier/_2769_ ));
 XNOR2_X2 \u_multiplier/_5366_  (.A(\u_multiplier/_2767_ ),
    .B(\u_multiplier/_2769_ ),
    .ZN(\u_multiplier/_2770_ ));
 NOR2_X1 \u_multiplier/_5367_  (.A1(\u_multiplier/_2765_ ),
    .A2(\u_multiplier/_2770_ ),
    .ZN(\u_multiplier/_2771_ ));
 XOR2_X2 \u_multiplier/_5368_  (.A(\u_multiplier/_2764_ ),
    .B(\u_multiplier/_2770_ ),
    .Z(\u_multiplier/_2772_ ));
 NOR2_X1 \u_multiplier/_5369_  (.A1(\u_multiplier/_2761_ ),
    .A2(\u_multiplier/_2772_ ),
    .ZN(\u_multiplier/_2773_ ));
 XOR2_X2 \u_multiplier/_5370_  (.A(\u_multiplier/_2761_ ),
    .B(\u_multiplier/_2772_ ),
    .Z(\u_multiplier/_2774_ ));
 INV_X1 \u_multiplier/_5371_  (.A(\u_multiplier/_2774_ ),
    .ZN(\u_multiplier/_2775_ ));
 NOR3_X2 \u_multiplier/_5372_  (.A1(\u_multiplier/_2756_ ),
    .A2(\u_multiplier/_2759_ ),
    .A3(\u_multiplier/_2774_ ),
    .ZN(\u_multiplier/_2776_ ));
 AOI211_X2 \u_multiplier/_5373_  (.A(\u_multiplier/_2758_ ),
    .B(\u_multiplier/_2775_ ),
    .C1(\u_multiplier/_2741_ ),
    .C2(\u_multiplier/_2742_ ),
    .ZN(\u_multiplier/_2777_ ));
 AND2_X1 \u_multiplier/_5374_  (.A1(\u_multiplier/_2756_ ),
    .A2(\u_multiplier/_2774_ ),
    .ZN(\u_multiplier/_2778_ ));
 NOR4_X4 \u_multiplier/_5375_  (.A1(\u_multiplier/_3334_ ),
    .A2(\u_multiplier/_2776_ ),
    .A3(\u_multiplier/_2777_ ),
    .A4(\u_multiplier/_2778_ ),
    .ZN(product[41]));
 OR2_X2 \u_multiplier/_5376_  (.A1(\u_multiplier/_2773_ ),
    .A2(\u_multiplier/_2778_ ),
    .ZN(\u_multiplier/_2779_ ));
 NOR2_X2 \u_multiplier/_5377_  (.A1(\u_multiplier/_2777_ ),
    .A2(\u_multiplier/_2779_ ),
    .ZN(\u_multiplier/_2780_ ));
 AOI21_X2 \u_multiplier/_5378_  (.A(\u_multiplier/_2771_ ),
    .B1(\u_multiplier/_2769_ ),
    .B2(\u_multiplier/_2767_ ),
    .ZN(\u_multiplier/_2781_ ));
 INV_X1 \u_multiplier/_5379_  (.A(\u_multiplier/_2781_ ),
    .ZN(\u_multiplier/_2782_ ));
 AND2_X1 \u_multiplier/_5380_  (.A1(\u_multiplier/K [4]),
    .A2(\u_multiplier/_2364_ ),
    .ZN(\u_multiplier/_2783_ ));
 AND2_X2 \u_multiplier/_5381_  (.A1(\u_multiplier/K [3]),
    .A2(\u_multiplier/_2610_ ),
    .ZN(\u_multiplier/_2784_ ));
 AOI211_X2 \u_multiplier/_5382_  (.A(\u_multiplier/dec_out [42]),
    .B(\u_multiplier/_2783_ ),
    .C1(\u_multiplier/_2784_ ),
    .C2(\u_multiplier/_3116_ ),
    .ZN(\u_multiplier/_2785_ ));
 INV_X1 \u_multiplier/_5383_  (.A(\u_multiplier/_2785_ ),
    .ZN(\u_multiplier/_2786_ ));
 AND2_X1 \u_multiplier/_5384_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_2615_ ),
    .ZN(\u_multiplier/_2787_ ));
 NAND2_X1 \u_multiplier/_5385_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2371_ ),
    .ZN(\u_multiplier/_2788_ ));
 OAI21_X2 \u_multiplier/_5386_  (.A(\u_multiplier/_2788_ ),
    .B1(\u_multiplier/_2787_ ),
    .B2(\u_multiplier/code_x [4]),
    .ZN(\u_multiplier/_2789_ ));
 AND2_X2 \u_multiplier/_5387_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_2619_ ),
    .ZN(\u_multiplier/_2790_ ));
 NAND2_X1 \u_multiplier/_5388_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_2377_ ),
    .ZN(\u_multiplier/_2791_ ));
 OAI21_X2 \u_multiplier/_5389_  (.A(\u_multiplier/_2791_ ),
    .B1(\u_multiplier/_2790_ ),
    .B2(\u_multiplier/code_y [4]),
    .ZN(\u_multiplier/_2792_ ));
 NOR2_X1 \u_multiplier/_5390_  (.A1(\u_multiplier/_2789_ ),
    .A2(\u_multiplier/_2792_ ),
    .ZN(\u_multiplier/_2793_ ));
 XOR2_X2 \u_multiplier/_5391_  (.A(\u_multiplier/_2789_ ),
    .B(\u_multiplier/_2792_ ),
    .Z(\u_multiplier/_2794_ ));
 XNOR2_X2 \u_multiplier/_5392_  (.A(\u_multiplier/_2785_ ),
    .B(\u_multiplier/_2794_ ),
    .ZN(\u_multiplier/_2795_ ));
 NAND2_X1 \u_multiplier/_5393_  (.A1(\u_multiplier/_2782_ ),
    .A2(\u_multiplier/_2795_ ),
    .ZN(\u_multiplier/_2796_ ));
 XOR2_X2 \u_multiplier/_5394_  (.A(\u_multiplier/_2781_ ),
    .B(\u_multiplier/_2795_ ),
    .Z(\u_multiplier/_2797_ ));
 INV_X1 \u_multiplier/_5395_  (.A(\u_multiplier/_2797_ ),
    .ZN(\u_multiplier/_2798_ ));
 OAI21_X1 \u_multiplier/_5396_  (.A(\u_multiplier/_2798_ ),
    .B1(\u_multiplier/_2779_ ),
    .B2(\u_multiplier/_2777_ ),
    .ZN(\u_multiplier/_2799_ ));
 NAND2_X1 \u_multiplier/_5397_  (.A1(net21),
    .A2(\u_multiplier/_2799_ ),
    .ZN(\u_multiplier/_2800_ ));
 AOI21_X4 \u_multiplier/_5398_  (.A(\u_multiplier/_2800_ ),
    .B1(\u_multiplier/_2797_ ),
    .B2(\u_multiplier/_2780_ ),
    .ZN(product[42]));
 NAND2_X1 \u_multiplier/_5399_  (.A1(\u_multiplier/_2796_ ),
    .A2(\u_multiplier/_2799_ ),
    .ZN(\u_multiplier/_2801_ ));
 AOI21_X2 \u_multiplier/_5400_  (.A(\u_multiplier/_2793_ ),
    .B1(\u_multiplier/_2794_ ),
    .B2(\u_multiplier/_2786_ ),
    .ZN(\u_multiplier/_2802_ ));
 AND2_X1 \u_multiplier/_5401_  (.A1(\u_multiplier/K [4]),
    .A2(\u_multiplier/_2394_ ),
    .ZN(\u_multiplier/_2803_ ));
 AND2_X2 \u_multiplier/_5402_  (.A1(\u_multiplier/K [3]),
    .A2(\u_multiplier/_2632_ ),
    .ZN(\u_multiplier/_2804_ ));
 AOI211_X2 \u_multiplier/_5403_  (.A(\u_multiplier/dec_out [43]),
    .B(\u_multiplier/_2803_ ),
    .C1(\u_multiplier/_2804_ ),
    .C2(\u_multiplier/_3116_ ),
    .ZN(\u_multiplier/_2805_ ));
 INV_X1 \u_multiplier/_5404_  (.A(\u_multiplier/_2805_ ),
    .ZN(\u_multiplier/_2806_ ));
 NOR3_X4 \u_multiplier/_5405_  (.A1(\u_multiplier/_3110_ ),
    .A2(\u_multiplier/_3111_ ),
    .A3(\u_multiplier/_2523_ ),
    .ZN(\u_multiplier/_2807_ ));
 OR2_X1 \u_multiplier/_5406_  (.A1(\u_multiplier/_3109_ ),
    .A2(\u_multiplier/_2400_ ),
    .ZN(\u_multiplier/_2808_ ));
 OAI21_X2 \u_multiplier/_5407_  (.A(\u_multiplier/_2808_ ),
    .B1(\u_multiplier/_2807_ ),
    .B2(\u_multiplier/code_x [4]),
    .ZN(\u_multiplier/_2809_ ));
 NOR3_X4 \u_multiplier/_5408_  (.A1(\u_multiplier/_3106_ ),
    .A2(\u_multiplier/_3107_ ),
    .A3(\u_multiplier/_2530_ ),
    .ZN(\u_multiplier/_2810_ ));
 OR2_X1 \u_multiplier/_5409_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_2810_ ),
    .ZN(\u_multiplier/_2811_ ));
 OAI21_X2 \u_multiplier/_5410_  (.A(\u_multiplier/_2811_ ),
    .B1(\u_multiplier/_2406_ ),
    .B2(\u_multiplier/_3108_ ),
    .ZN(\u_multiplier/_2812_ ));
 NOR2_X1 \u_multiplier/_5411_  (.A1(\u_multiplier/_2809_ ),
    .A2(\u_multiplier/_2812_ ),
    .ZN(\u_multiplier/_2813_ ));
 XOR2_X2 \u_multiplier/_5412_  (.A(\u_multiplier/_2809_ ),
    .B(\u_multiplier/_2812_ ),
    .Z(\u_multiplier/_2814_ ));
 XOR2_X2 \u_multiplier/_5413_  (.A(\u_multiplier/_2805_ ),
    .B(\u_multiplier/_2814_ ),
    .Z(\u_multiplier/_2815_ ));
 NOR2_X1 \u_multiplier/_5414_  (.A1(\u_multiplier/_2802_ ),
    .A2(\u_multiplier/_2815_ ),
    .ZN(\u_multiplier/_2816_ ));
 XOR2_X2 \u_multiplier/_5415_  (.A(\u_multiplier/_2802_ ),
    .B(\u_multiplier/_2815_ ),
    .Z(\u_multiplier/_2817_ ));
 OAI21_X1 \u_multiplier/_5416_  (.A(net21),
    .B1(\u_multiplier/_2801_ ),
    .B2(\u_multiplier/_2817_ ),
    .ZN(\u_multiplier/_2818_ ));
 AOI21_X1 \u_multiplier/_5417_  (.A(\u_multiplier/_2818_ ),
    .B1(\u_multiplier/_2817_ ),
    .B2(\u_multiplier/_2801_ ),
    .ZN(product[43]));
 OAI211_X2 \u_multiplier/_5418_  (.A(\u_multiplier/_2798_ ),
    .B(\u_multiplier/_2817_ ),
    .C1(\u_multiplier/_2777_ ),
    .C2(\u_multiplier/_2779_ ),
    .ZN(\u_multiplier/_2819_ ));
 AOI21_X1 \u_multiplier/_5419_  (.A(\u_multiplier/_2796_ ),
    .B1(\u_multiplier/_2802_ ),
    .B2(\u_multiplier/_2815_ ),
    .ZN(\u_multiplier/_2820_ ));
 NOR2_X2 \u_multiplier/_5420_  (.A1(\u_multiplier/_2816_ ),
    .A2(\u_multiplier/_2820_ ),
    .ZN(\u_multiplier/_2821_ ));
 NAND2_X1 \u_multiplier/_5421_  (.A1(\u_multiplier/_2819_ ),
    .A2(\u_multiplier/_2821_ ),
    .ZN(\u_multiplier/_2822_ ));
 AOI21_X2 \u_multiplier/_5422_  (.A(\u_multiplier/_2813_ ),
    .B1(\u_multiplier/_2814_ ),
    .B2(\u_multiplier/_2806_ ),
    .ZN(\u_multiplier/_2823_ ));
 NAND2_X2 \u_multiplier/_5423_  (.A1(\u_multiplier/K [3]),
    .A2(\u_multiplier/_2654_ ),
    .ZN(\u_multiplier/_2824_ ));
 INV_X1 \u_multiplier/_5424_  (.A(\u_multiplier/_2824_ ),
    .ZN(\u_multiplier/_2825_ ));
 AOI21_X1 \u_multiplier/_5425_  (.A(\u_multiplier/dec_out [44]),
    .B1(\u_multiplier/_2426_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2826_ ));
 OAI21_X2 \u_multiplier/_5426_  (.A(\u_multiplier/_2826_ ),
    .B1(\u_multiplier/_2824_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2827_ ));
 OAI21_X2 \u_multiplier/_5427_  (.A(\u_multiplier/_3109_ ),
    .B1(\u_multiplier/_3111_ ),
    .B2(\u_multiplier/_2659_ ),
    .ZN(\u_multiplier/_2828_ ));
 OAI21_X2 \u_multiplier/_5428_  (.A(\u_multiplier/_2828_ ),
    .B1(\u_multiplier/_2433_ ),
    .B2(\u_multiplier/_3109_ ),
    .ZN(\u_multiplier/_2829_ ));
 NAND3_X4 \u_multiplier/_5429_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/code_y [3]),
    .A3(\u_multiplier/_2560_ ),
    .ZN(\u_multiplier/_2830_ ));
 NAND2_X1 \u_multiplier/_5430_  (.A1(\u_multiplier/_3108_ ),
    .A2(\u_multiplier/_2830_ ),
    .ZN(\u_multiplier/_2831_ ));
 OAI21_X2 \u_multiplier/_5431_  (.A(\u_multiplier/_2831_ ),
    .B1(\u_multiplier/_2440_ ),
    .B2(\u_multiplier/_3108_ ),
    .ZN(\u_multiplier/_2832_ ));
 NOR2_X1 \u_multiplier/_5432_  (.A1(\u_multiplier/_2829_ ),
    .A2(\u_multiplier/_2832_ ),
    .ZN(\u_multiplier/_2833_ ));
 XOR2_X2 \u_multiplier/_5433_  (.A(\u_multiplier/_2829_ ),
    .B(\u_multiplier/_2832_ ),
    .Z(\u_multiplier/_2834_ ));
 XNOR2_X2 \u_multiplier/_5434_  (.A(\u_multiplier/_2827_ ),
    .B(\u_multiplier/_2834_ ),
    .ZN(\u_multiplier/_2835_ ));
 XOR2_X2 \u_multiplier/_5435_  (.A(\u_multiplier/_2823_ ),
    .B(\u_multiplier/_2835_ ),
    .Z(\u_multiplier/_2836_ ));
 INV_X1 \u_multiplier/_5436_  (.A(\u_multiplier/_2836_ ),
    .ZN(\u_multiplier/_2837_ ));
 AOI21_X1 \u_multiplier/_5437_  (.A(\u_multiplier/_2837_ ),
    .B1(\u_multiplier/_2821_ ),
    .B2(\u_multiplier/_2819_ ),
    .ZN(\u_multiplier/_2838_ ));
 OAI21_X1 \u_multiplier/_5438_  (.A(net21),
    .B1(\u_multiplier/_2822_ ),
    .B2(\u_multiplier/_2836_ ),
    .ZN(\u_multiplier/_2839_ ));
 NOR2_X1 \u_multiplier/_5439_  (.A1(\u_multiplier/_2838_ ),
    .A2(\u_multiplier/_2839_ ),
    .ZN(product[44]));
 AOI21_X2 \u_multiplier/_5440_  (.A(\u_multiplier/_2833_ ),
    .B1(\u_multiplier/_2834_ ),
    .B2(\u_multiplier/_2827_ ),
    .ZN(\u_multiplier/_2840_ ));
 NAND2_X2 \u_multiplier/_5441_  (.A1(\u_multiplier/K [3]),
    .A2(\u_multiplier/_2678_ ),
    .ZN(\u_multiplier/_2841_ ));
 AOI21_X1 \u_multiplier/_5442_  (.A(\u_multiplier/dec_out [45]),
    .B1(\u_multiplier/_2457_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2842_ ));
 OAI21_X2 \u_multiplier/_5443_  (.A(\u_multiplier/_2842_ ),
    .B1(\u_multiplier/_2841_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2843_ ));
 NOR2_X2 \u_multiplier/_5444_  (.A1(\u_multiplier/_3111_ ),
    .A2(\u_multiplier/_2682_ ),
    .ZN(\u_multiplier/_2844_ ));
 MUX2_X1 \u_multiplier/_5445_  (.A(\u_multiplier/_2464_ ),
    .B(\u_multiplier/_2844_ ),
    .S(\u_multiplier/_3109_ ),
    .Z(\u_multiplier/_2845_ ));
 NOR2_X2 \u_multiplier/_5446_  (.A1(\u_multiplier/_3107_ ),
    .A2(\u_multiplier/_2687_ ),
    .ZN(\u_multiplier/_2846_ ));
 MUX2_X1 \u_multiplier/_5447_  (.A(\u_multiplier/_2470_ ),
    .B(\u_multiplier/_2846_ ),
    .S(\u_multiplier/_3108_ ),
    .Z(\u_multiplier/_2847_ ));
 AND2_X1 \u_multiplier/_5448_  (.A1(\u_multiplier/_2845_ ),
    .A2(\u_multiplier/_2847_ ),
    .ZN(\u_multiplier/_2848_ ));
 XOR2_X2 \u_multiplier/_5449_  (.A(\u_multiplier/_2845_ ),
    .B(\u_multiplier/_2847_ ),
    .Z(\u_multiplier/_2849_ ));
 XNOR2_X2 \u_multiplier/_5450_  (.A(\u_multiplier/_2843_ ),
    .B(\u_multiplier/_2849_ ),
    .ZN(\u_multiplier/_2850_ ));
 NOR2_X1 \u_multiplier/_5451_  (.A1(\u_multiplier/_2840_ ),
    .A2(\u_multiplier/_2850_ ),
    .ZN(\u_multiplier/_2851_ ));
 XOR2_X1 \u_multiplier/_5452_  (.A(\u_multiplier/_2840_ ),
    .B(\u_multiplier/_2850_ ),
    .Z(\u_multiplier/_2852_ ));
 INV_X1 \u_multiplier/_5453_  (.A(\u_multiplier/_2852_ ),
    .ZN(\u_multiplier/_2853_ ));
 AOI211_X2 \u_multiplier/_5454_  (.A(\u_multiplier/_2837_ ),
    .B(\u_multiplier/_2853_ ),
    .C1(\u_multiplier/_2819_ ),
    .C2(\u_multiplier/_2821_ ),
    .ZN(\u_multiplier/_2854_ ));
 OAI21_X1 \u_multiplier/_5455_  (.A(\u_multiplier/_2853_ ),
    .B1(\u_multiplier/_2835_ ),
    .B2(\u_multiplier/_2823_ ),
    .ZN(\u_multiplier/_2855_ ));
 NOR2_X1 \u_multiplier/_5456_  (.A1(\u_multiplier/_2838_ ),
    .A2(\u_multiplier/_2855_ ),
    .ZN(\u_multiplier/_2856_ ));
 NOR3_X1 \u_multiplier/_5457_  (.A1(\u_multiplier/_2823_ ),
    .A2(\u_multiplier/_2835_ ),
    .A3(\u_multiplier/_2853_ ),
    .ZN(\u_multiplier/_2857_ ));
 NOR4_X1 \u_multiplier/_5458_  (.A1(\u_multiplier/_3334_ ),
    .A2(\u_multiplier/_2854_ ),
    .A3(\u_multiplier/_2856_ ),
    .A4(\u_multiplier/_2857_ ),
    .ZN(product[45]));
 NOR2_X1 \u_multiplier/_5459_  (.A1(\u_multiplier/_2851_ ),
    .A2(\u_multiplier/_2857_ ),
    .ZN(\u_multiplier/_2858_ ));
 INV_X1 \u_multiplier/_5460_  (.A(\u_multiplier/_2858_ ),
    .ZN(\u_multiplier/_2859_ ));
 NOR2_X1 \u_multiplier/_5461_  (.A1(\u_multiplier/_2854_ ),
    .A2(\u_multiplier/_2859_ ),
    .ZN(\u_multiplier/_2860_ ));
 AOI21_X1 \u_multiplier/_5462_  (.A(\u_multiplier/_2848_ ),
    .B1(\u_multiplier/_2849_ ),
    .B2(\u_multiplier/_2843_ ),
    .ZN(\u_multiplier/_2861_ ));
 AND2_X1 \u_multiplier/_5463_  (.A1(\u_multiplier/K [4]),
    .A2(\u_multiplier/_2490_ ),
    .ZN(\u_multiplier/_2862_ ));
 NOR2_X1 \u_multiplier/_5464_  (.A1(\u_multiplier/dec_out [46]),
    .A2(\u_multiplier/_2862_ ),
    .ZN(\u_multiplier/_2863_ ));
 NAND2_X2 \u_multiplier/_5465_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2496_ ),
    .ZN(\u_multiplier/_2864_ ));
 NAND2_X1 \u_multiplier/_5466_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_2502_ ),
    .ZN(\u_multiplier/_2865_ ));
 XOR2_X2 \u_multiplier/_5467_  (.A(\u_multiplier/_2864_ ),
    .B(\u_multiplier/_2865_ ),
    .Z(\u_multiplier/_2866_ ));
 OAI21_X1 \u_multiplier/_5468_  (.A(\u_multiplier/_2866_ ),
    .B1(\u_multiplier/_2862_ ),
    .B2(\u_multiplier/dec_out [46]),
    .ZN(\u_multiplier/_2867_ ));
 XOR2_X2 \u_multiplier/_5469_  (.A(\u_multiplier/_2863_ ),
    .B(\u_multiplier/_2866_ ),
    .Z(\u_multiplier/_2868_ ));
 OR2_X1 \u_multiplier/_5470_  (.A1(\u_multiplier/_2861_ ),
    .A2(\u_multiplier/_2868_ ),
    .ZN(\u_multiplier/_2869_ ));
 XNOR2_X1 \u_multiplier/_5471_  (.A(\u_multiplier/_2861_ ),
    .B(\u_multiplier/_2868_ ),
    .ZN(\u_multiplier/_2870_ ));
 INV_X1 \u_multiplier/_5472_  (.A(\u_multiplier/_2870_ ),
    .ZN(\u_multiplier/_2871_ ));
 OAI21_X1 \u_multiplier/_5473_  (.A(\u_multiplier/_2871_ ),
    .B1(\u_multiplier/_2859_ ),
    .B2(\u_multiplier/_2854_ ),
    .ZN(\u_multiplier/_2872_ ));
 NAND2_X1 \u_multiplier/_5474_  (.A1(net21),
    .A2(\u_multiplier/_2872_ ),
    .ZN(\u_multiplier/_2873_ ));
 AOI21_X1 \u_multiplier/_5475_  (.A(\u_multiplier/_2873_ ),
    .B1(\u_multiplier/_2870_ ),
    .B2(\u_multiplier/_2860_ ),
    .ZN(product[46]));
 NAND2_X1 \u_multiplier/_5476_  (.A1(\u_multiplier/_2869_ ),
    .A2(\u_multiplier/_2872_ ),
    .ZN(\u_multiplier/_2874_ ));
 OAI21_X2 \u_multiplier/_5477_  (.A(\u_multiplier/_2867_ ),
    .B1(\u_multiplier/_2865_ ),
    .B2(\u_multiplier/_2864_ ),
    .ZN(\u_multiplier/_2875_ ));
 AND2_X1 \u_multiplier/_5478_  (.A1(\u_multiplier/K [4]),
    .A2(\u_multiplier/_2518_ ),
    .ZN(\u_multiplier/_2876_ ));
 OR2_X1 \u_multiplier/_5479_  (.A1(\u_multiplier/dec_out [47]),
    .A2(\u_multiplier/_2876_ ),
    .ZN(\u_multiplier/_2877_ ));
 INV_X1 \u_multiplier/_5480_  (.A(\u_multiplier/_2877_ ),
    .ZN(\u_multiplier/_2878_ ));
 NAND2_X1 \u_multiplier/_5481_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2526_ ),
    .ZN(\u_multiplier/_2879_ ));
 NAND2_X1 \u_multiplier/_5482_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_2533_ ),
    .ZN(\u_multiplier/_2880_ ));
 OR2_X1 \u_multiplier/_5483_  (.A1(\u_multiplier/_2879_ ),
    .A2(\u_multiplier/_2880_ ),
    .ZN(\u_multiplier/_2881_ ));
 XNOR2_X2 \u_multiplier/_5484_  (.A(\u_multiplier/_2879_ ),
    .B(\u_multiplier/_2880_ ),
    .ZN(\u_multiplier/_2882_ ));
 XNOR2_X2 \u_multiplier/_5485_  (.A(\u_multiplier/_2877_ ),
    .B(\u_multiplier/_2882_ ),
    .ZN(\u_multiplier/_2883_ ));
 NAND2_X1 \u_multiplier/_5486_  (.A1(\u_multiplier/_2875_ ),
    .A2(\u_multiplier/_2883_ ),
    .ZN(\u_multiplier/_2884_ ));
 NOR2_X1 \u_multiplier/_5487_  (.A1(\u_multiplier/_2875_ ),
    .A2(\u_multiplier/_2883_ ),
    .ZN(\u_multiplier/_2885_ ));
 XOR2_X2 \u_multiplier/_5488_  (.A(\u_multiplier/_2875_ ),
    .B(\u_multiplier/_2883_ ),
    .Z(\u_multiplier/_2886_ ));
 OAI21_X1 \u_multiplier/_5489_  (.A(net21),
    .B1(\u_multiplier/_2874_ ),
    .B2(\u_multiplier/_2886_ ),
    .ZN(\u_multiplier/_2887_ ));
 AOI21_X1 \u_multiplier/_5490_  (.A(\u_multiplier/_2887_ ),
    .B1(\u_multiplier/_2886_ ),
    .B2(\u_multiplier/_2874_ ),
    .ZN(product[47]));
 OAI211_X4 \u_multiplier/_5491_  (.A(\u_multiplier/_2871_ ),
    .B(\u_multiplier/_2886_ ),
    .C1(\u_multiplier/_2854_ ),
    .C2(\u_multiplier/_2859_ ),
    .ZN(\u_multiplier/_2888_ ));
 OAI21_X1 \u_multiplier/_5492_  (.A(\u_multiplier/_2884_ ),
    .B1(\u_multiplier/_2885_ ),
    .B2(\u_multiplier/_2869_ ),
    .ZN(\u_multiplier/_2889_ ));
 INV_X1 \u_multiplier/_5493_  (.A(\u_multiplier/_2889_ ),
    .ZN(\u_multiplier/_2890_ ));
 NAND2_X1 \u_multiplier/_5494_  (.A1(\u_multiplier/_2888_ ),
    .A2(\u_multiplier/_2890_ ),
    .ZN(\u_multiplier/_2891_ ));
 OAI21_X1 \u_multiplier/_5495_  (.A(\u_multiplier/_2881_ ),
    .B1(\u_multiplier/_2882_ ),
    .B2(\u_multiplier/_2878_ ),
    .ZN(\u_multiplier/_2892_ ));
 INV_X1 \u_multiplier/_5496_  (.A(\u_multiplier/_2892_ ),
    .ZN(\u_multiplier/_2893_ ));
 AOI21_X4 \u_multiplier/_5497_  (.A(\u_multiplier/dec_out [48]),
    .B1(\u_multiplier/_2550_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2894_ ));
 NAND2_X1 \u_multiplier/_5498_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2557_ ),
    .ZN(\u_multiplier/_2895_ ));
 NAND2_X1 \u_multiplier/_5499_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_2564_ ),
    .ZN(\u_multiplier/_2896_ ));
 XNOR2_X2 \u_multiplier/_5500_  (.A(\u_multiplier/_2895_ ),
    .B(\u_multiplier/_2896_ ),
    .ZN(\u_multiplier/_2897_ ));
 OR2_X1 \u_multiplier/_5501_  (.A1(\u_multiplier/_2894_ ),
    .A2(\u_multiplier/_2897_ ),
    .ZN(\u_multiplier/_2898_ ));
 XNOR2_X2 \u_multiplier/_5502_  (.A(\u_multiplier/_2894_ ),
    .B(\u_multiplier/_2897_ ),
    .ZN(\u_multiplier/_2899_ ));
 XNOR2_X1 \u_multiplier/_5503_  (.A(\u_multiplier/_2892_ ),
    .B(\u_multiplier/_2899_ ),
    .ZN(\u_multiplier/_2900_ ));
 INV_X1 \u_multiplier/_5504_  (.A(\u_multiplier/_2900_ ),
    .ZN(\u_multiplier/_2901_ ));
 AOI21_X2 \u_multiplier/_5505_  (.A(\u_multiplier/_2901_ ),
    .B1(\u_multiplier/_2890_ ),
    .B2(\u_multiplier/_2888_ ),
    .ZN(\u_multiplier/_2902_ ));
 OAI21_X1 \u_multiplier/_5506_  (.A(net21),
    .B1(\u_multiplier/_2891_ ),
    .B2(\u_multiplier/_2900_ ),
    .ZN(\u_multiplier/_2903_ ));
 NOR2_X1 \u_multiplier/_5507_  (.A1(\u_multiplier/_2902_ ),
    .A2(\u_multiplier/_2903_ ),
    .ZN(product[48]));
 OAI21_X2 \u_multiplier/_5508_  (.A(\u_multiplier/_2898_ ),
    .B1(\u_multiplier/_2896_ ),
    .B2(\u_multiplier/_2895_ ),
    .ZN(\u_multiplier/_2904_ ));
 AOI21_X4 \u_multiplier/_5509_  (.A(\u_multiplier/dec_out [49]),
    .B1(\u_multiplier/_2579_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2905_ ));
 AND2_X1 \u_multiplier/_5510_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2587_ ),
    .ZN(\u_multiplier/_2906_ ));
 NAND2_X1 \u_multiplier/_5511_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_2594_ ),
    .ZN(\u_multiplier/_2907_ ));
 NAND3_X1 \u_multiplier/_5512_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_2594_ ),
    .A3(\u_multiplier/_2906_ ),
    .ZN(\u_multiplier/_2908_ ));
 XOR2_X2 \u_multiplier/_5513_  (.A(\u_multiplier/_2906_ ),
    .B(\u_multiplier/_2907_ ),
    .Z(\u_multiplier/_2909_ ));
 XOR2_X2 \u_multiplier/_5514_  (.A(\u_multiplier/_2905_ ),
    .B(\u_multiplier/_2909_ ),
    .Z(\u_multiplier/_2910_ ));
 XOR2_X2 \u_multiplier/_5515_  (.A(\u_multiplier/_2904_ ),
    .B(\u_multiplier/_2910_ ),
    .Z(\u_multiplier/_2911_ ));
 INV_X1 \u_multiplier/_5516_  (.A(\u_multiplier/_2911_ ),
    .ZN(\u_multiplier/_2912_ ));
 AOI211_X2 \u_multiplier/_5517_  (.A(\u_multiplier/_2901_ ),
    .B(\u_multiplier/_2912_ ),
    .C1(\u_multiplier/_2888_ ),
    .C2(\u_multiplier/_2890_ ),
    .ZN(\u_multiplier/_2913_ ));
 NAND2_X1 \u_multiplier/_5518_  (.A1(\u_multiplier/_2902_ ),
    .A2(\u_multiplier/_2911_ ),
    .ZN(\u_multiplier/_2914_ ));
 NOR3_X1 \u_multiplier/_5519_  (.A1(\u_multiplier/_2893_ ),
    .A2(\u_multiplier/_2899_ ),
    .A3(\u_multiplier/_2912_ ),
    .ZN(\u_multiplier/_2915_ ));
 OAI21_X1 \u_multiplier/_5520_  (.A(\u_multiplier/_2912_ ),
    .B1(\u_multiplier/_2899_ ),
    .B2(\u_multiplier/_2893_ ),
    .ZN(\u_multiplier/_2916_ ));
 OAI21_X1 \u_multiplier/_5521_  (.A(\u_multiplier/_2914_ ),
    .B1(\u_multiplier/_2916_ ),
    .B2(\u_multiplier/_2902_ ),
    .ZN(\u_multiplier/_2917_ ));
 NOR3_X1 \u_multiplier/_5522_  (.A1(\u_multiplier/_3334_ ),
    .A2(\u_multiplier/_2915_ ),
    .A3(\u_multiplier/_2917_ ),
    .ZN(product[49]));
 AOI21_X1 \u_multiplier/_5523_  (.A(\u_multiplier/_2915_ ),
    .B1(\u_multiplier/_2910_ ),
    .B2(\u_multiplier/_2904_ ),
    .ZN(\u_multiplier/_2918_ ));
 INV_X1 \u_multiplier/_5524_  (.A(\u_multiplier/_2918_ ),
    .ZN(\u_multiplier/_2919_ ));
 OAI21_X1 \u_multiplier/_5525_  (.A(\u_multiplier/_2908_ ),
    .B1(\u_multiplier/_2909_ ),
    .B2(\u_multiplier/_2905_ ),
    .ZN(\u_multiplier/_2920_ ));
 AOI21_X2 \u_multiplier/_5526_  (.A(\u_multiplier/dec_out [50]),
    .B1(\u_multiplier/_2611_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2921_ ));
 NAND2_X1 \u_multiplier/_5527_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2616_ ),
    .ZN(\u_multiplier/_2922_ ));
 NAND2_X2 \u_multiplier/_5528_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_2620_ ),
    .ZN(\u_multiplier/_2923_ ));
 XNOR2_X2 \u_multiplier/_5529_  (.A(\u_multiplier/_2922_ ),
    .B(\u_multiplier/_2923_ ),
    .ZN(\u_multiplier/_2924_ ));
 OR2_X1 \u_multiplier/_5530_  (.A1(\u_multiplier/_2921_ ),
    .A2(\u_multiplier/_2924_ ),
    .ZN(\u_multiplier/_2925_ ));
 XNOR2_X2 \u_multiplier/_5531_  (.A(\u_multiplier/_2921_ ),
    .B(\u_multiplier/_2924_ ),
    .ZN(\u_multiplier/_2926_ ));
 INV_X1 \u_multiplier/_5532_  (.A(\u_multiplier/_2926_ ),
    .ZN(\u_multiplier/_2927_ ));
 NAND2_X1 \u_multiplier/_5533_  (.A1(\u_multiplier/_2920_ ),
    .A2(\u_multiplier/_2927_ ),
    .ZN(\u_multiplier/_2928_ ));
 XNOR2_X1 \u_multiplier/_5534_  (.A(\u_multiplier/_2920_ ),
    .B(\u_multiplier/_2927_ ),
    .ZN(\u_multiplier/_2929_ ));
 INV_X1 \u_multiplier/_5535_  (.A(\u_multiplier/_2929_ ),
    .ZN(\u_multiplier/_2930_ ));
 OAI21_X1 \u_multiplier/_5536_  (.A(\u_multiplier/_2930_ ),
    .B1(\u_multiplier/_2919_ ),
    .B2(\u_multiplier/_2913_ ),
    .ZN(\u_multiplier/_2931_ ));
 NAND3_X1 \u_multiplier/_5537_  (.A1(\u_multiplier/_2914_ ),
    .A2(\u_multiplier/_2918_ ),
    .A3(\u_multiplier/_2929_ ),
    .ZN(\u_multiplier/_2932_ ));
 AND3_X1 \u_multiplier/_5538_  (.A1(net21),
    .A2(\u_multiplier/_2931_ ),
    .A3(\u_multiplier/_2932_ ),
    .ZN(product[50]));
 OAI21_X2 \u_multiplier/_5539_  (.A(\u_multiplier/_2925_ ),
    .B1(\u_multiplier/_2923_ ),
    .B2(\u_multiplier/_2922_ ),
    .ZN(\u_multiplier/_2933_ ));
 AOI21_X2 \u_multiplier/_5540_  (.A(\u_multiplier/dec_out [51]),
    .B1(\u_multiplier/_2633_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2934_ ));
 NAND2_X1 \u_multiplier/_5541_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2637_ ),
    .ZN(\u_multiplier/_2935_ ));
 NAND2_X1 \u_multiplier/_5542_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_2640_ ),
    .ZN(\u_multiplier/_2936_ ));
 XNOR2_X1 \u_multiplier/_5543_  (.A(\u_multiplier/_2935_ ),
    .B(\u_multiplier/_2936_ ),
    .ZN(\u_multiplier/_2937_ ));
 OR2_X1 \u_multiplier/_5544_  (.A1(\u_multiplier/_2934_ ),
    .A2(\u_multiplier/_2937_ ),
    .ZN(\u_multiplier/_2938_ ));
 XNOR2_X1 \u_multiplier/_5545_  (.A(\u_multiplier/_2934_ ),
    .B(\u_multiplier/_2937_ ),
    .ZN(\u_multiplier/_2939_ ));
 INV_X1 \u_multiplier/_5546_  (.A(\u_multiplier/_2939_ ),
    .ZN(\u_multiplier/_2940_ ));
 NAND2_X1 \u_multiplier/_5547_  (.A1(\u_multiplier/_2933_ ),
    .A2(\u_multiplier/_2940_ ),
    .ZN(\u_multiplier/_2941_ ));
 XNOR2_X2 \u_multiplier/_5548_  (.A(\u_multiplier/_2933_ ),
    .B(\u_multiplier/_2940_ ),
    .ZN(\u_multiplier/_2942_ ));
 INV_X1 \u_multiplier/_5549_  (.A(\u_multiplier/_2942_ ),
    .ZN(\u_multiplier/_2943_ ));
 NAND3_X1 \u_multiplier/_5550_  (.A1(\u_multiplier/_2928_ ),
    .A2(\u_multiplier/_2931_ ),
    .A3(\u_multiplier/_2942_ ),
    .ZN(\u_multiplier/_2944_ ));
 OAI211_X4 \u_multiplier/_5551_  (.A(\u_multiplier/_2930_ ),
    .B(\u_multiplier/_2943_ ),
    .C1(\u_multiplier/_2913_ ),
    .C2(\u_multiplier/_2919_ ),
    .ZN(\u_multiplier/_2945_ ));
 OR2_X1 \u_multiplier/_5552_  (.A1(\u_multiplier/_2928_ ),
    .A2(\u_multiplier/_2942_ ),
    .ZN(\u_multiplier/_2946_ ));
 AND4_X1 \u_multiplier/_5553_  (.A1(net21),
    .A2(\u_multiplier/_2944_ ),
    .A3(\u_multiplier/_2945_ ),
    .A4(\u_multiplier/_2946_ ),
    .ZN(product[51]));
 AND2_X1 \u_multiplier/_5554_  (.A1(\u_multiplier/_2941_ ),
    .A2(\u_multiplier/_2946_ ),
    .ZN(\u_multiplier/_2947_ ));
 AND2_X1 \u_multiplier/_5555_  (.A1(\u_multiplier/_2945_ ),
    .A2(\u_multiplier/_2947_ ),
    .ZN(\u_multiplier/_2948_ ));
 OAI21_X1 \u_multiplier/_5556_  (.A(\u_multiplier/_2938_ ),
    .B1(\u_multiplier/_2936_ ),
    .B2(\u_multiplier/_2935_ ),
    .ZN(\u_multiplier/_2949_ ));
 INV_X1 \u_multiplier/_5557_  (.A(\u_multiplier/_2949_ ),
    .ZN(\u_multiplier/_2950_ ));
 AOI21_X2 \u_multiplier/_5558_  (.A(\u_multiplier/dec_out [52]),
    .B1(\u_multiplier/_2655_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2951_ ));
 AND4_X1 \u_multiplier/_5559_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/code_x [4]),
    .A3(\u_multiplier/_2661_ ),
    .A4(\u_multiplier/_2666_ ),
    .ZN(\u_multiplier/_2952_ ));
 AOI22_X1 \u_multiplier/_5560_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2661_ ),
    .B1(\u_multiplier/_2666_ ),
    .B2(\u_multiplier/code_y [4]),
    .ZN(\u_multiplier/_2953_ ));
 OR2_X1 \u_multiplier/_5561_  (.A1(\u_multiplier/_2952_ ),
    .A2(\u_multiplier/_2953_ ),
    .ZN(\u_multiplier/_2954_ ));
 NOR2_X1 \u_multiplier/_5562_  (.A1(\u_multiplier/_2951_ ),
    .A2(\u_multiplier/_2954_ ),
    .ZN(\u_multiplier/_2955_ ));
 XNOR2_X1 \u_multiplier/_5563_  (.A(\u_multiplier/_2951_ ),
    .B(\u_multiplier/_2954_ ),
    .ZN(\u_multiplier/_2956_ ));
 NOR2_X1 \u_multiplier/_5564_  (.A1(\u_multiplier/_2950_ ),
    .A2(\u_multiplier/_2956_ ),
    .ZN(\u_multiplier/_2957_ ));
 XNOR2_X1 \u_multiplier/_5565_  (.A(\u_multiplier/_2949_ ),
    .B(\u_multiplier/_2956_ ),
    .ZN(\u_multiplier/_2958_ ));
 INV_X1 \u_multiplier/_5566_  (.A(\u_multiplier/_2958_ ),
    .ZN(\u_multiplier/_2959_ ));
 NOR2_X1 \u_multiplier/_5567_  (.A1(\u_multiplier/_2948_ ),
    .A2(\u_multiplier/_2959_ ),
    .ZN(\u_multiplier/_2960_ ));
 OAI21_X1 \u_multiplier/_5568_  (.A(net21),
    .B1(\u_multiplier/_2948_ ),
    .B2(\u_multiplier/_2959_ ),
    .ZN(\u_multiplier/_2961_ ));
 AOI21_X2 \u_multiplier/_5569_  (.A(\u_multiplier/_2961_ ),
    .B1(\u_multiplier/_2959_ ),
    .B2(\u_multiplier/_2948_ ),
    .ZN(product[52]));
 NOR2_X1 \u_multiplier/_5570_  (.A1(\u_multiplier/_2952_ ),
    .A2(\u_multiplier/_2955_ ),
    .ZN(\u_multiplier/_2962_ ));
 AOI21_X2 \u_multiplier/_5571_  (.A(\u_multiplier/dec_out [53]),
    .B1(\u_multiplier/_2679_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_2963_ ));
 NAND2_X1 \u_multiplier/_5572_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2684_ ),
    .ZN(\u_multiplier/_2964_ ));
 NAND2_X1 \u_multiplier/_5573_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_2689_ ),
    .ZN(\u_multiplier/_2965_ ));
 XOR2_X2 \u_multiplier/_5574_  (.A(\u_multiplier/_2964_ ),
    .B(\u_multiplier/_2965_ ),
    .Z(\u_multiplier/_2966_ ));
 INV_X1 \u_multiplier/_5575_  (.A(\u_multiplier/_2966_ ),
    .ZN(\u_multiplier/_2967_ ));
 OR2_X1 \u_multiplier/_5576_  (.A1(\u_multiplier/_2963_ ),
    .A2(\u_multiplier/_2967_ ),
    .ZN(\u_multiplier/_2968_ ));
 XNOR2_X2 \u_multiplier/_5577_  (.A(\u_multiplier/_2963_ ),
    .B(\u_multiplier/_2966_ ),
    .ZN(\u_multiplier/_2969_ ));
 INV_X1 \u_multiplier/_5578_  (.A(\u_multiplier/_2969_ ),
    .ZN(\u_multiplier/_2970_ ));
 NOR2_X1 \u_multiplier/_5579_  (.A1(\u_multiplier/_2962_ ),
    .A2(\u_multiplier/_2970_ ),
    .ZN(\u_multiplier/_2971_ ));
 XNOR2_X2 \u_multiplier/_5580_  (.A(\u_multiplier/_2962_ ),
    .B(\u_multiplier/_2969_ ),
    .ZN(\u_multiplier/_2972_ ));
 INV_X1 \u_multiplier/_5581_  (.A(\u_multiplier/_2972_ ),
    .ZN(\u_multiplier/_2973_ ));
 NOR3_X2 \u_multiplier/_5582_  (.A1(\u_multiplier/_2957_ ),
    .A2(\u_multiplier/_2960_ ),
    .A3(\u_multiplier/_2972_ ),
    .ZN(\u_multiplier/_2974_ ));
 AOI211_X2 \u_multiplier/_5583_  (.A(\u_multiplier/_2959_ ),
    .B(\u_multiplier/_2973_ ),
    .C1(\u_multiplier/_2945_ ),
    .C2(\u_multiplier/_2947_ ),
    .ZN(\u_multiplier/_2975_ ));
 AND2_X1 \u_multiplier/_5584_  (.A1(\u_multiplier/_2957_ ),
    .A2(\u_multiplier/_2972_ ),
    .ZN(\u_multiplier/_2976_ ));
 NOR4_X4 \u_multiplier/_5585_  (.A1(\u_multiplier/_3334_ ),
    .A2(\u_multiplier/_2974_ ),
    .A3(\u_multiplier/_2975_ ),
    .A4(\u_multiplier/_2976_ ),
    .ZN(product[53]));
 NOR2_X1 \u_multiplier/_5586_  (.A1(\u_multiplier/_2971_ ),
    .A2(\u_multiplier/_2976_ ),
    .ZN(\u_multiplier/_2977_ ));
 INV_X2 \u_multiplier/_5587_  (.A(\u_multiplier/_2977_ ),
    .ZN(\u_multiplier/_2978_ ));
 NOR2_X1 \u_multiplier/_5588_  (.A1(\u_multiplier/_2975_ ),
    .A2(\u_multiplier/_2978_ ),
    .ZN(\u_multiplier/_2979_ ));
 OAI21_X2 \u_multiplier/_5589_  (.A(\u_multiplier/_2968_ ),
    .B1(\u_multiplier/_2965_ ),
    .B2(\u_multiplier/_2964_ ),
    .ZN(\u_multiplier/_2980_ ));
 INV_X1 \u_multiplier/_5590_  (.A(\u_multiplier/_2980_ ),
    .ZN(\u_multiplier/_2981_ ));
 OAI21_X2 \u_multiplier/_5591_  (.A(\u_multiplier/_3121_ ),
    .B1(\u_multiplier/_2705_ ),
    .B2(\u_multiplier/_3116_ ),
    .ZN(\u_multiplier/_2982_ ));
 AND4_X1 \u_multiplier/_5592_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/code_x [4]),
    .A3(\u_multiplier/_2709_ ),
    .A4(\u_multiplier/_2712_ ),
    .ZN(\u_multiplier/_2983_ ));
 AOI22_X2 \u_multiplier/_5593_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2709_ ),
    .B1(\u_multiplier/_2712_ ),
    .B2(\u_multiplier/code_y [4]),
    .ZN(\u_multiplier/_2984_ ));
 NOR2_X2 \u_multiplier/_5594_  (.A1(\u_multiplier/_2983_ ),
    .A2(\u_multiplier/_2984_ ),
    .ZN(\u_multiplier/_2985_ ));
 XNOR2_X2 \u_multiplier/_5595_  (.A(\u_multiplier/_2982_ ),
    .B(\u_multiplier/_2985_ ),
    .ZN(\u_multiplier/_2986_ ));
 NOR2_X2 \u_multiplier/_5596_  (.A1(\u_multiplier/_2981_ ),
    .A2(\u_multiplier/_2986_ ),
    .ZN(\u_multiplier/_2987_ ));
 XOR2_X2 \u_multiplier/_5597_  (.A(\u_multiplier/_2980_ ),
    .B(\u_multiplier/_2986_ ),
    .Z(\u_multiplier/_2988_ ));
 INV_X1 \u_multiplier/_5598_  (.A(\u_multiplier/_2988_ ),
    .ZN(\u_multiplier/_2989_ ));
 NOR2_X2 \u_multiplier/_5599_  (.A1(\u_multiplier/_2979_ ),
    .A2(\u_multiplier/_2988_ ),
    .ZN(\u_multiplier/_2990_ ));
 NOR3_X2 \u_multiplier/_5600_  (.A1(\u_multiplier/_2975_ ),
    .A2(\u_multiplier/_2978_ ),
    .A3(\u_multiplier/_2989_ ),
    .ZN(\u_multiplier/_2991_ ));
 NOR3_X4 \u_multiplier/_5601_  (.A1(\u_multiplier/_3334_ ),
    .A2(\u_multiplier/_2990_ ),
    .A3(\u_multiplier/_2991_ ),
    .ZN(product[54]));
 AOI21_X2 \u_multiplier/_5602_  (.A(\u_multiplier/_2983_ ),
    .B1(\u_multiplier/_2985_ ),
    .B2(\u_multiplier/_2982_ ),
    .ZN(\u_multiplier/_2992_ ));
 OAI21_X2 \u_multiplier/_5603_  (.A(\u_multiplier/_3122_ ),
    .B1(\u_multiplier/_2725_ ),
    .B2(\u_multiplier/_3116_ ),
    .ZN(\u_multiplier/_2993_ ));
 NAND2_X1 \u_multiplier/_5604_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2728_ ),
    .ZN(\u_multiplier/_2994_ ));
 NAND2_X1 \u_multiplier/_5605_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_2730_ ),
    .ZN(\u_multiplier/_2995_ ));
 OR2_X1 \u_multiplier/_5606_  (.A1(\u_multiplier/_2994_ ),
    .A2(\u_multiplier/_2995_ ),
    .ZN(\u_multiplier/_2996_ ));
 XOR2_X2 \u_multiplier/_5607_  (.A(\u_multiplier/_2994_ ),
    .B(\u_multiplier/_2995_ ),
    .Z(\u_multiplier/_2997_ ));
 NAND2_X1 \u_multiplier/_5608_  (.A1(\u_multiplier/_2993_ ),
    .A2(\u_multiplier/_2997_ ),
    .ZN(\u_multiplier/_2998_ ));
 XNOR2_X2 \u_multiplier/_5609_  (.A(\u_multiplier/_2993_ ),
    .B(\u_multiplier/_2997_ ),
    .ZN(\u_multiplier/_2999_ ));
 NOR2_X1 \u_multiplier/_5610_  (.A1(\u_multiplier/_2992_ ),
    .A2(\u_multiplier/_2999_ ),
    .ZN(\u_multiplier/_3000_ ));
 XOR2_X2 \u_multiplier/_5611_  (.A(\u_multiplier/_2992_ ),
    .B(\u_multiplier/_2999_ ),
    .Z(\u_multiplier/_3001_ ));
 NOR3_X1 \u_multiplier/_5612_  (.A1(\u_multiplier/_2987_ ),
    .A2(\u_multiplier/_2990_ ),
    .A3(\u_multiplier/_3001_ ),
    .ZN(\u_multiplier/_3002_ ));
 OAI211_X4 \u_multiplier/_5613_  (.A(\u_multiplier/_2989_ ),
    .B(\u_multiplier/_3001_ ),
    .C1(\u_multiplier/_2975_ ),
    .C2(\u_multiplier/_2978_ ),
    .ZN(\u_multiplier/_3003_ ));
 AOI21_X1 \u_multiplier/_5614_  (.A(\u_multiplier/_3334_ ),
    .B1(\u_multiplier/_2987_ ),
    .B2(\u_multiplier/_3001_ ),
    .ZN(\u_multiplier/_3004_ ));
 NAND2_X1 \u_multiplier/_5615_  (.A1(\u_multiplier/_3003_ ),
    .A2(\u_multiplier/_3004_ ),
    .ZN(\u_multiplier/_3005_ ));
 NOR2_X1 \u_multiplier/_5616_  (.A1(\u_multiplier/_3002_ ),
    .A2(\u_multiplier/_3005_ ),
    .ZN(product[55]));
 AOI21_X2 \u_multiplier/_5617_  (.A(\u_multiplier/_3000_ ),
    .B1(\u_multiplier/_3001_ ),
    .B2(\u_multiplier/_2987_ ),
    .ZN(\u_multiplier/_3006_ ));
 NAND2_X1 \u_multiplier/_5618_  (.A1(\u_multiplier/_2996_ ),
    .A2(\u_multiplier/_2998_ ),
    .ZN(\u_multiplier/_3007_ ));
 OAI21_X2 \u_multiplier/_5619_  (.A(\u_multiplier/_3123_ ),
    .B1(\u_multiplier/_2745_ ),
    .B2(\u_multiplier/_3116_ ),
    .ZN(\u_multiplier/_3008_ ));
 NAND2_X1 \u_multiplier/_5620_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2749_ ),
    .ZN(\u_multiplier/_3009_ ));
 NAND2_X1 \u_multiplier/_5621_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_2751_ ),
    .ZN(\u_multiplier/_3010_ ));
 OR2_X1 \u_multiplier/_5622_  (.A1(\u_multiplier/_3009_ ),
    .A2(\u_multiplier/_3010_ ),
    .ZN(\u_multiplier/_3011_ ));
 XOR2_X2 \u_multiplier/_5623_  (.A(\u_multiplier/_3009_ ),
    .B(\u_multiplier/_3010_ ),
    .Z(\u_multiplier/_3012_ ));
 NAND2_X1 \u_multiplier/_5624_  (.A1(\u_multiplier/_3008_ ),
    .A2(\u_multiplier/_3012_ ),
    .ZN(\u_multiplier/_3013_ ));
 XNOR2_X2 \u_multiplier/_5625_  (.A(\u_multiplier/_3008_ ),
    .B(\u_multiplier/_3012_ ),
    .ZN(\u_multiplier/_3014_ ));
 AOI21_X1 \u_multiplier/_5626_  (.A(\u_multiplier/_3014_ ),
    .B1(\u_multiplier/_2998_ ),
    .B2(\u_multiplier/_2996_ ),
    .ZN(\u_multiplier/_3015_ ));
 XOR2_X2 \u_multiplier/_5627_  (.A(\u_multiplier/_3007_ ),
    .B(\u_multiplier/_3014_ ),
    .Z(\u_multiplier/_3016_ ));
 AOI21_X4 \u_multiplier/_5628_  (.A(\u_multiplier/_3016_ ),
    .B1(\u_multiplier/_3006_ ),
    .B2(\u_multiplier/_3003_ ),
    .ZN(\u_multiplier/_3017_ ));
 AND3_X1 \u_multiplier/_5629_  (.A1(\u_multiplier/_3003_ ),
    .A2(\u_multiplier/_3006_ ),
    .A3(\u_multiplier/_3016_ ),
    .ZN(\u_multiplier/_3018_ ));
 NOR3_X4 \u_multiplier/_5630_  (.A1(\u_multiplier/_3334_ ),
    .A2(\u_multiplier/_3017_ ),
    .A3(\u_multiplier/_3018_ ),
    .ZN(product[56]));
 NAND2_X1 \u_multiplier/_5631_  (.A1(\u_multiplier/_3011_ ),
    .A2(\u_multiplier/_3013_ ),
    .ZN(\u_multiplier/_3019_ ));
 OAI21_X1 \u_multiplier/_5632_  (.A(\u_multiplier/_3124_ ),
    .B1(\u_multiplier/_2762_ ),
    .B2(\u_multiplier/_3116_ ),
    .ZN(\u_multiplier/_3020_ ));
 NAND2_X1 \u_multiplier/_5633_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2766_ ),
    .ZN(\u_multiplier/_3021_ ));
 NAND2_X1 \u_multiplier/_5634_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_2768_ ),
    .ZN(\u_multiplier/_3022_ ));
 XOR2_X2 \u_multiplier/_5635_  (.A(\u_multiplier/_3021_ ),
    .B(\u_multiplier/_3022_ ),
    .Z(\u_multiplier/_3023_ ));
 NAND2_X1 \u_multiplier/_5636_  (.A1(\u_multiplier/_3020_ ),
    .A2(\u_multiplier/_3023_ ),
    .ZN(\u_multiplier/_3024_ ));
 XNOR2_X1 \u_multiplier/_5637_  (.A(\u_multiplier/_3020_ ),
    .B(\u_multiplier/_3023_ ),
    .ZN(\u_multiplier/_3025_ ));
 AOI21_X1 \u_multiplier/_5638_  (.A(\u_multiplier/_3025_ ),
    .B1(\u_multiplier/_3013_ ),
    .B2(\u_multiplier/_3011_ ),
    .ZN(\u_multiplier/_3026_ ));
 INV_X1 \u_multiplier/_5639_  (.A(\u_multiplier/_3026_ ),
    .ZN(\u_multiplier/_3027_ ));
 XOR2_X1 \u_multiplier/_5640_  (.A(\u_multiplier/_3019_ ),
    .B(\u_multiplier/_3025_ ),
    .Z(\u_multiplier/_3028_ ));
 INV_X1 \u_multiplier/_5641_  (.A(\u_multiplier/_3028_ ),
    .ZN(\u_multiplier/_3029_ ));
 OAI21_X2 \u_multiplier/_5642_  (.A(\u_multiplier/_3029_ ),
    .B1(\u_multiplier/_3017_ ),
    .B2(\u_multiplier/_3015_ ),
    .ZN(\u_multiplier/_3030_ ));
 OR3_X1 \u_multiplier/_5643_  (.A1(\u_multiplier/_3015_ ),
    .A2(\u_multiplier/_3017_ ),
    .A3(\u_multiplier/_3029_ ),
    .ZN(\u_multiplier/_3031_ ));
 AND3_X2 \u_multiplier/_5644_  (.A1(net21),
    .A2(\u_multiplier/_3030_ ),
    .A3(\u_multiplier/_3031_ ),
    .ZN(product[57]));
 OAI21_X1 \u_multiplier/_5645_  (.A(\u_multiplier/_3024_ ),
    .B1(\u_multiplier/_3022_ ),
    .B2(\u_multiplier/_3021_ ),
    .ZN(\u_multiplier/_3032_ ));
 AOI21_X2 \u_multiplier/_5646_  (.A(\u_multiplier/dec_out [58]),
    .B1(\u_multiplier/_2784_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_3033_ ));
 INV_X1 \u_multiplier/_5647_  (.A(\u_multiplier/_3033_ ),
    .ZN(\u_multiplier/_3034_ ));
 AND4_X1 \u_multiplier/_5648_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/code_x [4]),
    .A3(\u_multiplier/_2787_ ),
    .A4(\u_multiplier/_2790_ ),
    .ZN(\u_multiplier/_3035_ ));
 AOI22_X1 \u_multiplier/_5649_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2787_ ),
    .B1(\u_multiplier/_2790_ ),
    .B2(\u_multiplier/code_y [4]),
    .ZN(\u_multiplier/_3036_ ));
 NOR2_X1 \u_multiplier/_5650_  (.A1(\u_multiplier/_3035_ ),
    .A2(\u_multiplier/_3036_ ),
    .ZN(\u_multiplier/_3037_ ));
 XNOR2_X2 \u_multiplier/_5651_  (.A(\u_multiplier/_3033_ ),
    .B(\u_multiplier/_3037_ ),
    .ZN(\u_multiplier/_3038_ ));
 AND2_X1 \u_multiplier/_5652_  (.A1(\u_multiplier/_3032_ ),
    .A2(\u_multiplier/_3038_ ),
    .ZN(\u_multiplier/_3039_ ));
 XNOR2_X2 \u_multiplier/_5653_  (.A(\u_multiplier/_3032_ ),
    .B(\u_multiplier/_3038_ ),
    .ZN(\u_multiplier/_3040_ ));
 AOI21_X4 \u_multiplier/_5654_  (.A(\u_multiplier/_3040_ ),
    .B1(\u_multiplier/_3030_ ),
    .B2(\u_multiplier/_3027_ ),
    .ZN(\u_multiplier/_3041_ ));
 AND3_X1 \u_multiplier/_5655_  (.A1(\u_multiplier/_3027_ ),
    .A2(\u_multiplier/_3030_ ),
    .A3(\u_multiplier/_3040_ ),
    .ZN(\u_multiplier/_3042_ ));
 NOR3_X4 \u_multiplier/_5656_  (.A1(\u_multiplier/_3334_ ),
    .A2(\u_multiplier/_3041_ ),
    .A3(\u_multiplier/_3042_ ),
    .ZN(product[58]));
 AOI21_X1 \u_multiplier/_5657_  (.A(\u_multiplier/_3035_ ),
    .B1(\u_multiplier/_3037_ ),
    .B2(\u_multiplier/_3034_ ),
    .ZN(\u_multiplier/_3043_ ));
 INV_X1 \u_multiplier/_5658_  (.A(\u_multiplier/_3043_ ),
    .ZN(\u_multiplier/_3044_ ));
 AOI21_X2 \u_multiplier/_5659_  (.A(\u_multiplier/dec_out [59]),
    .B1(\u_multiplier/_2804_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_3045_ ));
 INV_X1 \u_multiplier/_5660_  (.A(\u_multiplier/_3045_ ),
    .ZN(\u_multiplier/_3046_ ));
 AND4_X1 \u_multiplier/_5661_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/code_x [4]),
    .A3(\u_multiplier/_2807_ ),
    .A4(\u_multiplier/_2810_ ),
    .ZN(\u_multiplier/_3047_ ));
 AOI22_X1 \u_multiplier/_5662_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2807_ ),
    .B1(\u_multiplier/_2810_ ),
    .B2(\u_multiplier/code_y [4]),
    .ZN(\u_multiplier/_3048_ ));
 NOR2_X1 \u_multiplier/_5663_  (.A1(\u_multiplier/_3047_ ),
    .A2(\u_multiplier/_3048_ ),
    .ZN(\u_multiplier/_3049_ ));
 XNOR2_X1 \u_multiplier/_5664_  (.A(\u_multiplier/_3045_ ),
    .B(\u_multiplier/_3049_ ),
    .ZN(\u_multiplier/_3050_ ));
 NAND2_X1 \u_multiplier/_5665_  (.A1(\u_multiplier/_3044_ ),
    .A2(\u_multiplier/_3050_ ),
    .ZN(\u_multiplier/_3051_ ));
 XOR2_X1 \u_multiplier/_5666_  (.A(\u_multiplier/_3043_ ),
    .B(\u_multiplier/_3050_ ),
    .Z(\u_multiplier/_3052_ ));
 INV_X1 \u_multiplier/_5667_  (.A(\u_multiplier/_3052_ ),
    .ZN(\u_multiplier/_3053_ ));
 OAI21_X2 \u_multiplier/_5668_  (.A(\u_multiplier/_3053_ ),
    .B1(\u_multiplier/_3041_ ),
    .B2(\u_multiplier/_3039_ ),
    .ZN(\u_multiplier/_3054_ ));
 OR3_X1 \u_multiplier/_5669_  (.A1(\u_multiplier/_3039_ ),
    .A2(\u_multiplier/_3041_ ),
    .A3(\u_multiplier/_3053_ ),
    .ZN(\u_multiplier/_3055_ ));
 AND3_X4 \u_multiplier/_5670_  (.A1(net21),
    .A2(\u_multiplier/_3054_ ),
    .A3(\u_multiplier/_3055_ ),
    .ZN(product[59]));
 AOI21_X1 \u_multiplier/_5671_  (.A(\u_multiplier/_3047_ ),
    .B1(\u_multiplier/_3049_ ),
    .B2(\u_multiplier/_3046_ ),
    .ZN(\u_multiplier/_3056_ ));
 AOI21_X1 \u_multiplier/_5672_  (.A(\u_multiplier/dec_out [60]),
    .B1(\u_multiplier/_2825_ ),
    .B2(\u_multiplier/K [4]),
    .ZN(\u_multiplier/_3057_ ));
 NAND4_X4 \u_multiplier/_5673_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/code_x [2]),
    .A3(\u_multiplier/code_x [3]),
    .A4(\u_multiplier/_2553_ ),
    .ZN(\u_multiplier/_3058_ ));
 NOR2_X1 \u_multiplier/_5674_  (.A1(\u_multiplier/_3108_ ),
    .A2(\u_multiplier/_2830_ ),
    .ZN(\u_multiplier/_3059_ ));
 NOR3_X1 \u_multiplier/_5675_  (.A1(\u_multiplier/_3108_ ),
    .A2(\u_multiplier/_2830_ ),
    .A3(\u_multiplier/_3058_ ),
    .ZN(\u_multiplier/_3060_ ));
 XOR2_X2 \u_multiplier/_5676_  (.A(\u_multiplier/_3058_ ),
    .B(\u_multiplier/_3059_ ),
    .Z(\u_multiplier/_3061_ ));
 NOR2_X1 \u_multiplier/_5677_  (.A1(\u_multiplier/_3057_ ),
    .A2(\u_multiplier/_3061_ ),
    .ZN(\u_multiplier/_3062_ ));
 XNOR2_X1 \u_multiplier/_5678_  (.A(\u_multiplier/_3057_ ),
    .B(\u_multiplier/_3061_ ),
    .ZN(\u_multiplier/_3063_ ));
 NOR2_X1 \u_multiplier/_5679_  (.A1(\u_multiplier/_3056_ ),
    .A2(\u_multiplier/_3063_ ),
    .ZN(\u_multiplier/_3064_ ));
 XOR2_X1 \u_multiplier/_5680_  (.A(\u_multiplier/_3056_ ),
    .B(\u_multiplier/_3063_ ),
    .Z(\u_multiplier/_3065_ ));
 INV_X1 \u_multiplier/_5681_  (.A(\u_multiplier/_3065_ ),
    .ZN(\u_multiplier/_3066_ ));
 AOI21_X2 \u_multiplier/_5682_  (.A(\u_multiplier/_3066_ ),
    .B1(\u_multiplier/_3054_ ),
    .B2(\u_multiplier/_3051_ ),
    .ZN(\u_multiplier/_3067_ ));
 NAND3_X1 \u_multiplier/_5683_  (.A1(\u_multiplier/_3051_ ),
    .A2(\u_multiplier/_3054_ ),
    .A3(\u_multiplier/_3066_ ),
    .ZN(\u_multiplier/_3068_ ));
 NAND2_X1 \u_multiplier/_5684_  (.A1(net21),
    .A2(\u_multiplier/_3068_ ),
    .ZN(\u_multiplier/_3069_ ));
 NOR2_X1 \u_multiplier/_5685_  (.A1(\u_multiplier/_3067_ ),
    .A2(\u_multiplier/_3069_ ),
    .ZN(product[60]));
 NOR2_X1 \u_multiplier/_5686_  (.A1(\u_multiplier/_3060_ ),
    .A2(\u_multiplier/_3062_ ),
    .ZN(\u_multiplier/_3070_ ));
 OAI21_X2 \u_multiplier/_5687_  (.A(\u_multiplier/_3125_ ),
    .B1(\u_multiplier/_2841_ ),
    .B2(\u_multiplier/_3116_ ),
    .ZN(\u_multiplier/_3071_ ));
 NAND2_X1 \u_multiplier/_5688_  (.A1(\u_multiplier/code_x [4]),
    .A2(\u_multiplier/_2844_ ),
    .ZN(\u_multiplier/_3072_ ));
 NAND2_X1 \u_multiplier/_5689_  (.A1(\u_multiplier/code_y [4]),
    .A2(\u_multiplier/_2846_ ),
    .ZN(\u_multiplier/_3073_ ));
 NOR2_X1 \u_multiplier/_5690_  (.A1(\u_multiplier/_3072_ ),
    .A2(\u_multiplier/_3073_ ),
    .ZN(\u_multiplier/_3074_ ));
 XOR2_X2 \u_multiplier/_5691_  (.A(\u_multiplier/_3072_ ),
    .B(\u_multiplier/_3073_ ),
    .Z(\u_multiplier/_3075_ ));
 XNOR2_X2 \u_multiplier/_5692_  (.A(\u_multiplier/_3071_ ),
    .B(\u_multiplier/_3075_ ),
    .ZN(\u_multiplier/_3076_ ));
 OR2_X1 \u_multiplier/_5693_  (.A1(\u_multiplier/_3070_ ),
    .A2(\u_multiplier/_3076_ ),
    .ZN(\u_multiplier/_3077_ ));
 XOR2_X2 \u_multiplier/_5694_  (.A(\u_multiplier/_3070_ ),
    .B(\u_multiplier/_3076_ ),
    .Z(\u_multiplier/_3078_ ));
 OAI21_X2 \u_multiplier/_5695_  (.A(\u_multiplier/_3078_ ),
    .B1(\u_multiplier/_3067_ ),
    .B2(\u_multiplier/_3064_ ),
    .ZN(\u_multiplier/_3079_ ));
 OR3_X1 \u_multiplier/_5696_  (.A1(\u_multiplier/_3064_ ),
    .A2(\u_multiplier/_3067_ ),
    .A3(\u_multiplier/_3078_ ),
    .ZN(\u_multiplier/_3080_ ));
 AND3_X1 \u_multiplier/_5697_  (.A1(net21),
    .A2(\u_multiplier/_3079_ ),
    .A3(\u_multiplier/_3080_ ),
    .ZN(product[61]));
 AOI21_X2 \u_multiplier/_5698_  (.A(\u_multiplier/_3074_ ),
    .B1(\u_multiplier/_3075_ ),
    .B2(\u_multiplier/_3071_ ),
    .ZN(\u_multiplier/_3081_ ));
 NOR2_X1 \u_multiplier/_5699_  (.A1(\u_multiplier/_3126_ ),
    .A2(\u_multiplier/_3081_ ),
    .ZN(\u_multiplier/_3082_ ));
 XNOR2_X1 \u_multiplier/_5700_  (.A(\u_multiplier/dec_out [62]),
    .B(\u_multiplier/_3081_ ),
    .ZN(\u_multiplier/_3083_ ));
 INV_X1 \u_multiplier/_5701_  (.A(\u_multiplier/_3083_ ),
    .ZN(\u_multiplier/_3084_ ));
 AOI21_X4 \u_multiplier/_5702_  (.A(\u_multiplier/_3084_ ),
    .B1(\u_multiplier/_3079_ ),
    .B2(\u_multiplier/_3077_ ),
    .ZN(\u_multiplier/_3085_ ));
 AND3_X1 \u_multiplier/_5703_  (.A1(\u_multiplier/_3077_ ),
    .A2(\u_multiplier/_3079_ ),
    .A3(\u_multiplier/_3084_ ),
    .ZN(\u_multiplier/_3086_ ));
 NOR3_X4 \u_multiplier/_5704_  (.A1(\u_multiplier/_3334_ ),
    .A2(\u_multiplier/_3085_ ),
    .A3(\u_multiplier/_3086_ ),
    .ZN(product[62]));
 OAI21_X1 \u_multiplier/_5705_  (.A(\u_multiplier/dec_out [63]),
    .B1(\u_multiplier/_3082_ ),
    .B2(\u_multiplier/_3085_ ),
    .ZN(\u_multiplier/_3087_ ));
 OR3_X1 \u_multiplier/_5706_  (.A1(\u_multiplier/dec_out [63]),
    .A2(\u_multiplier/_3082_ ),
    .A3(\u_multiplier/_3085_ ),
    .ZN(\u_multiplier/_3088_ ));
 AND3_X1 \u_multiplier/_5707_  (.A1(net21),
    .A2(\u_multiplier/_3087_ ),
    .A3(\u_multiplier/_3088_ ),
    .ZN(product[63]));
 NAND2_X1 \u_multiplier/_5708_  (.A1(\u_multiplier/code_y [0]),
    .A2(\u_multiplier/code_x [0]),
    .ZN(\u_multiplier/_3089_ ));
 NOR2_X1 \u_multiplier/_5709_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/code_x [1]),
    .ZN(\u_multiplier/_3090_ ));
 NAND2_X1 \u_multiplier/_5710_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/code_x [1]),
    .ZN(\u_multiplier/_3091_ ));
 XOR2_X2 \u_multiplier/_5711_  (.A(\u_multiplier/code_y [1]),
    .B(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_3092_ ));
 XNOR2_X2 \u_multiplier/_5712_  (.A(\u_multiplier/_3089_ ),
    .B(\u_multiplier/_3092_ ),
    .ZN(\u_multiplier/_1862_ ));
 OAI21_X2 \u_multiplier/_5713_  (.A(\u_multiplier/_3091_ ),
    .B1(\u_multiplier/_3090_ ),
    .B2(\u_multiplier/_3089_ ),
    .ZN(\u_multiplier/_3093_ ));
 NAND2_X1 \u_multiplier/_5714_  (.A1(\u_multiplier/_3106_ ),
    .A2(\u_multiplier/_3110_ ),
    .ZN(\u_multiplier/_3094_ ));
 NOR2_X1 \u_multiplier/_5715_  (.A1(\u_multiplier/_3106_ ),
    .A2(\u_multiplier/_3110_ ),
    .ZN(\u_multiplier/_3095_ ));
 XNOR2_X1 \u_multiplier/_5716_  (.A(\u_multiplier/code_y [2]),
    .B(\u_multiplier/code_x [2]),
    .ZN(\u_multiplier/_3096_ ));
 XNOR2_X2 \u_multiplier/_5717_  (.A(\u_multiplier/_3093_ ),
    .B(\u_multiplier/_3096_ ),
    .ZN(\u_multiplier/_1863_ ));
 AOI21_X4 \u_multiplier/_5718_  (.A(\u_multiplier/_3095_ ),
    .B1(\u_multiplier/_3094_ ),
    .B2(\u_multiplier/_3093_ ),
    .ZN(\u_multiplier/_3097_ ));
 NOR2_X1 \u_multiplier/_5719_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/code_x [3]),
    .ZN(\u_multiplier/_3098_ ));
 NAND2_X1 \u_multiplier/_5720_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/code_x [3]),
    .ZN(\u_multiplier/_3099_ ));
 XOR2_X2 \u_multiplier/_5721_  (.A(\u_multiplier/code_y [3]),
    .B(\u_multiplier/code_x [3]),
    .Z(\u_multiplier/_3100_ ));
 XNOR2_X2 \u_multiplier/_5722_  (.A(\u_multiplier/_3097_ ),
    .B(\u_multiplier/_3100_ ),
    .ZN(\u_multiplier/_1864_ ));
 XNOR2_X2 \u_multiplier/_5723_  (.A(\u_multiplier/code_y [4]),
    .B(\u_multiplier/code_x [4]),
    .ZN(\u_multiplier/_3101_ ));
 AOI21_X2 \u_multiplier/_5724_  (.A(\u_multiplier/_3098_ ),
    .B1(\u_multiplier/_3099_ ),
    .B2(\u_multiplier/_3097_ ),
    .ZN(\u_multiplier/_3102_ ));
 AOI211_X2 \u_multiplier/_5725_  (.A(\u_multiplier/_3098_ ),
    .B(\u_multiplier/_3101_ ),
    .C1(\u_multiplier/_3099_ ),
    .C2(\u_multiplier/_3097_ ),
    .ZN(\u_multiplier/_3103_ ));
 XNOR2_X2 \u_multiplier/_5726_  (.A(\u_multiplier/_3101_ ),
    .B(\u_multiplier/_3102_ ),
    .ZN(\u_multiplier/_1865_ ));
 XOR2_X2 \u_multiplier/_5727_  (.A(\u_multiplier/code_y [0]),
    .B(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_1861_ ));
 AOI21_X4 \u_multiplier/_5728_  (.A(\u_multiplier/_3103_ ),
    .B1(\u_multiplier/code_x [4]),
    .B2(\u_multiplier/code_y [4]),
    .ZN(\u_multiplier/_3104_ ));
 INV_X16 \u_multiplier/_5729_  (.A(\u_multiplier/_3104_ ),
    .ZN(\u_multiplier/_1866_ ));
 INV_X8 \u_multiplier/dec/_163_  (.A(\u_multiplier/_1866_ ),
    .ZN(\u_multiplier/dec/_143_ ));
 INV_X2 \u_multiplier/dec/_164_  (.A(\u_multiplier/_1862_ ),
    .ZN(\u_multiplier/dec/_144_ ));
 INV_X2 \u_multiplier/dec/_165_  (.A(\u_multiplier/_1861_ ),
    .ZN(\u_multiplier/dec/_145_ ));
 INV_X2 \u_multiplier/dec/_166_  (.A(\u_multiplier/_1863_ ),
    .ZN(\u_multiplier/dec/_146_ ));
 INV_X4 \u_multiplier/dec/_167_  (.A(net20),
    .ZN(\u_multiplier/dec/_147_ ));
 INV_X8 \u_multiplier/dec/_168_  (.A(net18),
    .ZN(\u_multiplier/dec/_148_ ));
 NOR2_X2 \u_multiplier/dec/_169_  (.A1(\u_multiplier/_1862_ ),
    .A2(\u_multiplier/_1861_ ),
    .ZN(\u_multiplier/dec/_149_ ));
 NOR3_X1 \u_multiplier/dec/_170_  (.A1(\u_multiplier/_1862_ ),
    .A2(\u_multiplier/_1861_ ),
    .A3(\u_multiplier/_1863_ ),
    .ZN(\u_multiplier/dec/_150_ ));
 OR4_X2 \u_multiplier/dec/_171_  (.A1(\u_multiplier/_1862_ ),
    .A2(\u_multiplier/_1861_ ),
    .A3(\u_multiplier/_1863_ ),
    .A4(\u_multiplier/_1864_ ),
    .ZN(\u_multiplier/dec/_151_ ));
 NOR3_X2 \u_multiplier/dec/_172_  (.A1(\u_multiplier/_1866_ ),
    .A2(\u_multiplier/_1865_ ),
    .A3(\u_multiplier/dec/_151_ ),
    .ZN(\u_multiplier/dec_out [0]));
 NAND4_X4 \u_multiplier/dec/_173_  (.A1(\u_multiplier/dec/_144_ ),
    .A2(\u_multiplier/_1861_ ),
    .A3(\u_multiplier/dec/_146_ ),
    .A4(\u_multiplier/dec/_147_ ),
    .ZN(\u_multiplier/dec/_152_ ));
 NOR3_X2 \u_multiplier/dec/_174_  (.A1(\u_multiplier/_1866_ ),
    .A2(\u_multiplier/_1865_ ),
    .A3(\u_multiplier/dec/_152_ ),
    .ZN(\u_multiplier/dec_out [1]));
 NAND4_X4 \u_multiplier/dec/_175_  (.A1(\u_multiplier/_1862_ ),
    .A2(\u_multiplier/dec/_145_ ),
    .A3(\u_multiplier/dec/_146_ ),
    .A4(\u_multiplier/dec/_147_ ),
    .ZN(\u_multiplier/dec/_153_ ));
 NOR3_X2 \u_multiplier/dec/_176_  (.A1(\u_multiplier/_1866_ ),
    .A2(\u_multiplier/_1865_ ),
    .A3(\u_multiplier/dec/_153_ ),
    .ZN(\u_multiplier/dec_out [2]));
 NAND2_X1 \u_multiplier/dec/_177_  (.A1(\u_multiplier/_1862_ ),
    .A2(\u_multiplier/_1861_ ),
    .ZN(\u_multiplier/dec/_154_ ));
 NOR2_X1 \u_multiplier/dec/_178_  (.A1(\u_multiplier/_1863_ ),
    .A2(\u_multiplier/dec/_154_ ),
    .ZN(\u_multiplier/dec/_155_ ));
 OR3_X4 \u_multiplier/dec/_179_  (.A1(\u_multiplier/_1863_ ),
    .A2(net20),
    .A3(\u_multiplier/dec/_154_ ),
    .ZN(\u_multiplier/dec/_156_ ));
 NOR3_X2 \u_multiplier/dec/_180_  (.A1(\u_multiplier/_1866_ ),
    .A2(\u_multiplier/_1865_ ),
    .A3(\u_multiplier/dec/_156_ ),
    .ZN(\u_multiplier/dec_out [3]));
 NAND2_X4 \u_multiplier/dec/_181_  (.A1(\u_multiplier/_1863_ ),
    .A2(\u_multiplier/dec/_149_ ),
    .ZN(\u_multiplier/dec/_157_ ));
 NOR4_X2 \u_multiplier/dec/_182_  (.A1(\u_multiplier/_1866_ ),
    .A2(\u_multiplier/_1864_ ),
    .A3(\u_multiplier/_1865_ ),
    .A4(\u_multiplier/dec/_157_ ),
    .ZN(\u_multiplier/dec_out [4]));
 NAND4_X4 \u_multiplier/dec/_183_  (.A1(\u_multiplier/dec/_144_ ),
    .A2(\u_multiplier/_1861_ ),
    .A3(\u_multiplier/_1863_ ),
    .A4(\u_multiplier/dec/_147_ ),
    .ZN(\u_multiplier/dec/_158_ ));
 NOR3_X1 \u_multiplier/dec/_184_  (.A1(\u_multiplier/_1866_ ),
    .A2(net19),
    .A3(\u_multiplier/dec/_158_ ),
    .ZN(\u_multiplier/dec_out [5]));
 NAND4_X2 \u_multiplier/dec/_185_  (.A1(\u_multiplier/_1862_ ),
    .A2(\u_multiplier/dec/_145_ ),
    .A3(\u_multiplier/_1863_ ),
    .A4(\u_multiplier/dec/_147_ ),
    .ZN(\u_multiplier/dec/_159_ ));
 NOR3_X1 \u_multiplier/dec/_186_  (.A1(\u_multiplier/_1866_ ),
    .A2(net19),
    .A3(\u_multiplier/dec/_159_ ),
    .ZN(\u_multiplier/dec_out [6]));
 NAND3_X2 \u_multiplier/dec/_187_  (.A1(\u_multiplier/_1862_ ),
    .A2(\u_multiplier/_1861_ ),
    .A3(\u_multiplier/_1863_ ),
    .ZN(\u_multiplier/dec/_160_ ));
 NOR4_X2 \u_multiplier/dec/_188_  (.A1(\u_multiplier/_1866_ ),
    .A2(net20),
    .A3(net19),
    .A4(\u_multiplier/dec/_160_ ),
    .ZN(\u_multiplier/dec_out [7]));
 NAND2_X1 \u_multiplier/dec/_189_  (.A1(net20),
    .A2(\u_multiplier/dec/_150_ ),
    .ZN(\u_multiplier/dec/_161_ ));
 NOR3_X2 \u_multiplier/dec/_190_  (.A1(\u_multiplier/_1866_ ),
    .A2(net19),
    .A3(\u_multiplier/dec/_161_ ),
    .ZN(\u_multiplier/dec_out [8]));
 NAND4_X2 \u_multiplier/dec/_191_  (.A1(\u_multiplier/dec/_144_ ),
    .A2(\u_multiplier/_1861_ ),
    .A3(\u_multiplier/dec/_146_ ),
    .A4(net20),
    .ZN(\u_multiplier/dec/_162_ ));
 NOR3_X1 \u_multiplier/dec/_192_  (.A1(\u_multiplier/_1866_ ),
    .A2(net18),
    .A3(\u_multiplier/dec/_162_ ),
    .ZN(\u_multiplier/dec_out [9]));
 NAND4_X4 \u_multiplier/dec/_193_  (.A1(\u_multiplier/_1862_ ),
    .A2(\u_multiplier/dec/_145_ ),
    .A3(\u_multiplier/dec/_146_ ),
    .A4(net20),
    .ZN(\u_multiplier/dec/_134_ ));
 NOR3_X2 \u_multiplier/dec/_194_  (.A1(\u_multiplier/_1866_ ),
    .A2(net19),
    .A3(\u_multiplier/dec/_134_ ),
    .ZN(\u_multiplier/dec_out [10]));
 OR4_X1 \u_multiplier/dec/_195_  (.A1(\u_multiplier/_1863_ ),
    .A2(\u_multiplier/dec/_147_ ),
    .A3(net18),
    .A4(\u_multiplier/dec/_154_ ),
    .ZN(\u_multiplier/dec/_135_ ));
 NOR2_X1 \u_multiplier/dec/_196_  (.A1(\u_multiplier/_1866_ ),
    .A2(\u_multiplier/dec/_135_ ),
    .ZN(\u_multiplier/dec_out [11]));
 NAND3_X1 \u_multiplier/dec/_197_  (.A1(\u_multiplier/_1863_ ),
    .A2(net20),
    .A3(\u_multiplier/dec/_149_ ),
    .ZN(\u_multiplier/dec/_136_ ));
 NOR3_X2 \u_multiplier/dec/_198_  (.A1(\u_multiplier/_1866_ ),
    .A2(net19),
    .A3(\u_multiplier/dec/_136_ ),
    .ZN(\u_multiplier/dec_out [12]));
 NAND4_X2 \u_multiplier/dec/_199_  (.A1(\u_multiplier/dec/_144_ ),
    .A2(\u_multiplier/_1861_ ),
    .A3(\u_multiplier/_1863_ ),
    .A4(net20),
    .ZN(\u_multiplier/dec/_137_ ));
 NOR3_X1 \u_multiplier/dec/_200_  (.A1(\u_multiplier/_1866_ ),
    .A2(net18),
    .A3(\u_multiplier/dec/_137_ ),
    .ZN(\u_multiplier/dec_out [13]));
 NAND4_X2 \u_multiplier/dec/_201_  (.A1(\u_multiplier/_1862_ ),
    .A2(\u_multiplier/dec/_145_ ),
    .A3(\u_multiplier/_1863_ ),
    .A4(net20),
    .ZN(\u_multiplier/dec/_138_ ));
 NOR3_X1 \u_multiplier/dec/_202_  (.A1(\u_multiplier/_1866_ ),
    .A2(net18),
    .A3(\u_multiplier/dec/_138_ ),
    .ZN(\u_multiplier/dec_out [14]));
 OR2_X1 \u_multiplier/dec/_203_  (.A1(\u_multiplier/dec/_147_ ),
    .A2(\u_multiplier/dec/_160_ ),
    .ZN(\u_multiplier/dec/_139_ ));
 NOR3_X1 \u_multiplier/dec/_204_  (.A1(\u_multiplier/_1866_ ),
    .A2(net18),
    .A3(\u_multiplier/dec/_139_ ),
    .ZN(\u_multiplier/dec_out [15]));
 OR2_X1 \u_multiplier/dec/_205_  (.A1(\u_multiplier/dec/_148_ ),
    .A2(\u_multiplier/dec/_151_ ),
    .ZN(\u_multiplier/dec/_140_ ));
 NOR2_X1 \u_multiplier/dec/_206_  (.A1(\u_multiplier/_1866_ ),
    .A2(\u_multiplier/dec/_140_ ),
    .ZN(\u_multiplier/dec_out [16]));
 NOR3_X1 \u_multiplier/dec/_207_  (.A1(\u_multiplier/_1866_ ),
    .A2(\u_multiplier/dec/_148_ ),
    .A3(\u_multiplier/dec/_152_ ),
    .ZN(\u_multiplier/dec_out [17]));
 NOR3_X1 \u_multiplier/dec/_208_  (.A1(\u_multiplier/_1866_ ),
    .A2(\u_multiplier/dec/_148_ ),
    .A3(\u_multiplier/dec/_153_ ),
    .ZN(\u_multiplier/dec_out [18]));
 NOR3_X1 \u_multiplier/dec/_209_  (.A1(\u_multiplier/_1866_ ),
    .A2(\u_multiplier/dec/_148_ ),
    .A3(\u_multiplier/dec/_156_ ),
    .ZN(\u_multiplier/dec_out [19]));
 NOR4_X2 \u_multiplier/dec/_210_  (.A1(\u_multiplier/_1866_ ),
    .A2(\u_multiplier/_1864_ ),
    .A3(\u_multiplier/dec/_148_ ),
    .A4(\u_multiplier/dec/_157_ ),
    .ZN(\u_multiplier/dec_out [20]));
 NOR3_X1 \u_multiplier/dec/_211_  (.A1(\u_multiplier/_1866_ ),
    .A2(\u_multiplier/dec/_148_ ),
    .A3(\u_multiplier/dec/_158_ ),
    .ZN(\u_multiplier/dec_out [21]));
 NOR3_X1 \u_multiplier/dec/_212_  (.A1(\u_multiplier/_1866_ ),
    .A2(\u_multiplier/dec/_148_ ),
    .A3(\u_multiplier/dec/_159_ ),
    .ZN(\u_multiplier/dec_out [22]));
 NOR4_X1 \u_multiplier/dec/_213_  (.A1(\u_multiplier/_1866_ ),
    .A2(net20),
    .A3(\u_multiplier/dec/_148_ ),
    .A4(\u_multiplier/dec/_160_ ),
    .ZN(\u_multiplier/dec_out [23]));
 NAND3_X1 \u_multiplier/dec/_214_  (.A1(net20),
    .A2(net19),
    .A3(\u_multiplier/dec/_150_ ),
    .ZN(\u_multiplier/dec/_141_ ));
 NOR2_X1 \u_multiplier/dec/_215_  (.A1(\u_multiplier/_1866_ ),
    .A2(\u_multiplier/dec/_141_ ),
    .ZN(\u_multiplier/dec_out [24]));
 NOR3_X1 \u_multiplier/dec/_216_  (.A1(\u_multiplier/_1866_ ),
    .A2(\u_multiplier/dec/_148_ ),
    .A3(\u_multiplier/dec/_162_ ),
    .ZN(\u_multiplier/dec_out [25]));
 NOR3_X1 \u_multiplier/dec/_217_  (.A1(\u_multiplier/_1866_ ),
    .A2(\u_multiplier/dec/_148_ ),
    .A3(\u_multiplier/dec/_134_ ),
    .ZN(\u_multiplier/dec_out [26]));
 AND4_X1 \u_multiplier/dec/_218_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(net20),
    .A3(net18),
    .A4(\u_multiplier/dec/_155_ ),
    .ZN(\u_multiplier/dec_out [27]));
 NAND4_X1 \u_multiplier/dec/_219_  (.A1(\u_multiplier/_1863_ ),
    .A2(net20),
    .A3(net19),
    .A4(\u_multiplier/dec/_149_ ),
    .ZN(\u_multiplier/dec/_142_ ));
 NOR2_X1 \u_multiplier/dec/_220_  (.A1(\u_multiplier/_1866_ ),
    .A2(\u_multiplier/dec/_142_ ),
    .ZN(\u_multiplier/dec_out [28]));
 NOR3_X1 \u_multiplier/dec/_221_  (.A1(\u_multiplier/_1866_ ),
    .A2(\u_multiplier/dec/_148_ ),
    .A3(\u_multiplier/dec/_137_ ),
    .ZN(\u_multiplier/dec_out [29]));
 NOR3_X1 \u_multiplier/dec/_222_  (.A1(\u_multiplier/_1866_ ),
    .A2(\u_multiplier/dec/_148_ ),
    .A3(\u_multiplier/dec/_138_ ),
    .ZN(\u_multiplier/dec_out [30]));
 NOR3_X1 \u_multiplier/dec/_223_  (.A1(\u_multiplier/_1866_ ),
    .A2(\u_multiplier/dec/_148_ ),
    .A3(\u_multiplier/dec/_139_ ),
    .ZN(\u_multiplier/dec_out [31]));
 NOR3_X1 \u_multiplier/dec/_224_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(\u_multiplier/_1865_ ),
    .A3(\u_multiplier/dec/_151_ ),
    .ZN(\u_multiplier/dec_out [32]));
 NOR3_X1 \u_multiplier/dec/_225_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(\u_multiplier/_1865_ ),
    .A3(\u_multiplier/dec/_152_ ),
    .ZN(\u_multiplier/dec_out [33]));
 NOR3_X1 \u_multiplier/dec/_226_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(\u_multiplier/_1865_ ),
    .A3(\u_multiplier/dec/_153_ ),
    .ZN(\u_multiplier/dec_out [34]));
 NOR3_X1 \u_multiplier/dec/_227_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(\u_multiplier/_1865_ ),
    .A3(\u_multiplier/dec/_156_ ),
    .ZN(\u_multiplier/dec_out [35]));
 NOR4_X1 \u_multiplier/dec/_228_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(\u_multiplier/_1864_ ),
    .A3(net19),
    .A4(\u_multiplier/dec/_157_ ),
    .ZN(\u_multiplier/dec_out [36]));
 NOR3_X1 \u_multiplier/dec/_229_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(net19),
    .A3(\u_multiplier/dec/_158_ ),
    .ZN(\u_multiplier/dec_out [37]));
 NOR3_X1 \u_multiplier/dec/_230_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(net19),
    .A3(\u_multiplier/dec/_159_ ),
    .ZN(\u_multiplier/dec_out [38]));
 NOR4_X1 \u_multiplier/dec/_231_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(net20),
    .A3(net19),
    .A4(\u_multiplier/dec/_160_ ),
    .ZN(\u_multiplier/dec_out [39]));
 NOR3_X1 \u_multiplier/dec/_232_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(net19),
    .A3(\u_multiplier/dec/_161_ ),
    .ZN(\u_multiplier/dec_out [40]));
 NOR3_X1 \u_multiplier/dec/_233_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(net19),
    .A3(\u_multiplier/dec/_162_ ),
    .ZN(\u_multiplier/dec_out [41]));
 NOR3_X1 \u_multiplier/dec/_234_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(net19),
    .A3(\u_multiplier/dec/_134_ ),
    .ZN(\u_multiplier/dec_out [42]));
 NOR2_X1 \u_multiplier/dec/_235_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(\u_multiplier/dec/_135_ ),
    .ZN(\u_multiplier/dec_out [43]));
 NOR3_X1 \u_multiplier/dec/_236_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(net19),
    .A3(\u_multiplier/dec/_136_ ),
    .ZN(\u_multiplier/dec_out [44]));
 NOR3_X1 \u_multiplier/dec/_237_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(net18),
    .A3(\u_multiplier/dec/_137_ ),
    .ZN(\u_multiplier/dec_out [45]));
 NOR3_X1 \u_multiplier/dec/_238_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(net18),
    .A3(\u_multiplier/dec/_138_ ),
    .ZN(\u_multiplier/dec_out [46]));
 NOR3_X1 \u_multiplier/dec/_239_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(net18),
    .A3(\u_multiplier/dec/_139_ ),
    .ZN(\u_multiplier/dec_out [47]));
 NOR2_X1 \u_multiplier/dec/_240_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(\u_multiplier/dec/_140_ ),
    .ZN(\u_multiplier/dec_out [48]));
 NOR3_X2 \u_multiplier/dec/_241_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(\u_multiplier/dec/_148_ ),
    .A3(\u_multiplier/dec/_152_ ),
    .ZN(\u_multiplier/dec_out [49]));
 NOR3_X1 \u_multiplier/dec/_242_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(\u_multiplier/dec/_148_ ),
    .A3(\u_multiplier/dec/_153_ ),
    .ZN(\u_multiplier/dec_out [50]));
 NOR3_X1 \u_multiplier/dec/_243_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(\u_multiplier/dec/_148_ ),
    .A3(\u_multiplier/dec/_156_ ),
    .ZN(\u_multiplier/dec_out [51]));
 NOR4_X2 \u_multiplier/dec/_244_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(\u_multiplier/_1864_ ),
    .A3(\u_multiplier/dec/_148_ ),
    .A4(\u_multiplier/dec/_157_ ),
    .ZN(\u_multiplier/dec_out [52]));
 NOR3_X1 \u_multiplier/dec/_245_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(\u_multiplier/dec/_148_ ),
    .A3(\u_multiplier/dec/_158_ ),
    .ZN(\u_multiplier/dec_out [53]));
 NOR3_X1 \u_multiplier/dec/_246_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(\u_multiplier/dec/_148_ ),
    .A3(\u_multiplier/dec/_159_ ),
    .ZN(\u_multiplier/dec_out [54]));
 NOR4_X1 \u_multiplier/dec/_247_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(net20),
    .A3(\u_multiplier/dec/_148_ ),
    .A4(\u_multiplier/dec/_160_ ),
    .ZN(\u_multiplier/dec_out [55]));
 NOR2_X1 \u_multiplier/dec/_248_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(\u_multiplier/dec/_141_ ),
    .ZN(\u_multiplier/dec_out [56]));
 NOR3_X1 \u_multiplier/dec/_249_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(\u_multiplier/dec/_148_ ),
    .A3(\u_multiplier/dec/_162_ ),
    .ZN(\u_multiplier/dec_out [57]));
 NOR3_X1 \u_multiplier/dec/_250_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(\u_multiplier/dec/_148_ ),
    .A3(\u_multiplier/dec/_134_ ),
    .ZN(\u_multiplier/dec_out [58]));
 AND4_X1 \u_multiplier/dec/_251_  (.A1(\u_multiplier/_1866_ ),
    .A2(net20),
    .A3(net18),
    .A4(\u_multiplier/dec/_155_ ),
    .ZN(\u_multiplier/dec_out [59]));
 NOR2_X1 \u_multiplier/dec/_252_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(\u_multiplier/dec/_142_ ),
    .ZN(\u_multiplier/dec_out [60]));
 NOR3_X1 \u_multiplier/dec/_253_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(\u_multiplier/dec/_148_ ),
    .A3(\u_multiplier/dec/_137_ ),
    .ZN(\u_multiplier/dec_out [61]));
 NOR3_X1 \u_multiplier/dec/_254_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(\u_multiplier/dec/_148_ ),
    .A3(\u_multiplier/dec/_138_ ),
    .ZN(\u_multiplier/dec_out [62]));
 NOR3_X1 \u_multiplier/dec/_255_  (.A1(\u_multiplier/dec/_143_ ),
    .A2(\u_multiplier/dec/_148_ ),
    .A3(\u_multiplier/dec/_139_ ),
    .ZN(\u_multiplier/dec_out [63]));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_219_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_220_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_221_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_222_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_223_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_224_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_225_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_226_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_227_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_228_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_229_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_2_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_2_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_2_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_2_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_2_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_2_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_2_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_2_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_2_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_2_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_2_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_2_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_2_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_2_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_2_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_2_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_2_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_2_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_2_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_2_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_2_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_2_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_2_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_2_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_2_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_2_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_2_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_2_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_2_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_2_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_2_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_2_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_2_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_2_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_2_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_2_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_2_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_2_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_2_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_2_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_2_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_2_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_2_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_2_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_2_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_2_Right_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_2_Right_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_2_Right_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_2_Right_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_2_Right_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_2_Right_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_2_Right_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_2_Right_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_2_Right_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_2_Right_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_2_Right_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_2_Right_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_2_Right_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_2_Right_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_2_Right_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_2_Right_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_2_Right_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_2_Right_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_2_Right_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_2_Right_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_2_Right_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_2_Right_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_2_Right_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_2_Right_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_2_Right_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_2_Right_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_2_Right_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_2_Right_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_2_Right_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_2_Right_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_2_Right_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_2_Right_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_2_Right_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_2_Right_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_2_Right_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_2_Right_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_2_Right_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_2_Right_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_2_Right_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_2_Right_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_2_Right_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_2_Right_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_2_Right_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_2_Right_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_2_Right_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_2_Right_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_2_Right_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_2_Right_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_2_Right_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_2_Right_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_2_Right_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_2_Right_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_2_Right_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_2_Right_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_2_Right_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_2_Right_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_2_Right_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_2_Right_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_2_Right_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_2_Right_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_2_Right_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_2_Right_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_2_Right_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_2_Right_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_2_Right_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_2_Right_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_2_Right_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_2_Right_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_2_Right_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_2_Right_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_2_Right_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_2_Right_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_2_Right_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_2_Right_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_2_Right_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_2_Right_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_2_Right_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_2_Right_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_2_Right_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_2_Right_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_2_Right_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_2_Right_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_2_Right_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_2_Right_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_2_Right_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_2_Right_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_2_Right_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_2_Right_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_2_Right_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_2_Right_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_2_Right_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_2_Right_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_2_Right_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_2_Right_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_2_Right_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_2_Right_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_2_Right_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_2_Right_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_2_Right_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_2_Right_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_2_Right_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_2_Right_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_2_Right_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_2_Right_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_2_Right_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_2_Right_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_2_Right_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_2_Right_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_2_Right_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_2_Right_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_2_Right_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_2_Right_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_2_Right_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_2_Right_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_2_Right_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_2_Right_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_2_Right_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_2_Right_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_2_Right_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_2_Right_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_2_Right_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_2_Right_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_2_Right_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_265 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_266 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_267 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_268 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_269 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_1_Left_270 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_1_Left_271 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_1_Left_272 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_1_Left_273 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_1_Left_274 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_1_Left_275 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_1_Left_276 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_1_Left_277 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_1_Left_278 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_1_Left_279 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_1_Left_280 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_1_Left_281 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_1_Left_282 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_1_Left_283 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_1_Left_284 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_1_Left_285 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_1_Left_286 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_1_Left_287 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_1_Left_288 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_1_Left_289 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_1_Left_290 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_1_Left_291 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_1_Left_292 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_1_Left_293 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_1_Left_294 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_1_Left_295 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_1_Left_296 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_1_Left_297 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_1_Left_298 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_1_Left_299 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_1_Left_300 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_1_Left_301 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_1_Left_302 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_1_Left_303 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_1_Left_304 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_1_Left_305 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_1_Left_306 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_1_Left_307 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_1_Left_308 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_1_Left_309 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_1_Left_310 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_1_Left_311 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_1_Left_312 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_1_Left_313 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_1_Left_314 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_1_Left_315 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_1_Left_316 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_1_Left_317 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_1_Left_318 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_1_Left_319 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_1_Left_320 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_1_Left_321 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_1_Left_322 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_1_Left_323 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_1_Left_324 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_1_Left_325 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_1_Left_326 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_1_Left_327 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_1_Left_328 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_1_Left_329 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_1_Left_330 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_1_Left_331 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_1_Left_332 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_1_Left_333 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_1_Left_334 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_1_Left_335 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_1_Left_336 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_1_Left_337 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_1_Left_338 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_1_Left_339 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_1_Left_340 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_1_Left_341 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_1_Left_342 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_1_Left_343 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_1_Left_344 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_1_Left_345 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_1_Left_346 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_1_Left_347 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_1_Left_348 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_1_Left_349 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_1_Left_350 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_1_Left_351 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_1_Left_352 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_1_Left_353 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_1_Left_354 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_1_Left_355 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_1_Left_356 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_1_Left_357 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_1_Left_358 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_1_Left_359 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_1_Left_360 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_1_Left_361 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_1_Left_362 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_1_Left_363 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_1_Left_364 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_1_Left_365 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_1_Left_366 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_1_Left_367 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_1_Left_368 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_1_Left_369 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_1_Left_370 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_1_Left_371 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_1_Left_372 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_1_Left_373 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_1_Left_374 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_1_Left_375 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_1_Left_376 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_1_Left_377 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_1_Left_378 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_1_Left_379 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_1_Left_380 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_1_Left_381 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_1_Left_382 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_1_Left_383 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_1_Left_384 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_1_Left_385 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_1_Left_386 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_1_Left_387 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_1_Left_388 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_1_Left_389 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_1_Left_390 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_1_Left_391 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_1_Left_392 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_1_Left_393 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_1_Left_394 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_1_Left_395 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_1_Left_396 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_1_Left_397 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_1_Left_398 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_1_Left_399 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_1_Left_400 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_1_Left_401 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_1_Left_402 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_1_Left_403 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_1_Left_404 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_1_Left_405 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_1_Left_406 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_1_Left_407 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_1_Left_408 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_1_Left_409 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_1_Left_410 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_1_Left_411 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_1_Left_412 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_1_Left_413 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_1_Left_414 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_1_Left_415 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_1_Left_416 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_1_Left_417 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_1_Left_418 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_1_Left_419 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_1_Left_420 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_1_Left_421 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_1_Left_422 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_1_Left_423 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_1_Left_424 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_1_Left_425 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_1_Left_426 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_1_Left_427 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_1_Left_428 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_1_Left_429 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_1_Left_430 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_1_Left_431 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_1_Left_432 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_1_Left_433 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_1_Left_434 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_1_Left_435 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_1_Left_436 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Left_437 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Left_438 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Left_439 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Left_440 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Left_441 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Left_442 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Left_443 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Left_444 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Left_445 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Left_446 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Left_447 ();
 TAPCELL_X1 PHY_EDGE_ROW_219_Left_448 ();
 TAPCELL_X1 PHY_EDGE_ROW_220_Left_449 ();
 TAPCELL_X1 PHY_EDGE_ROW_221_Left_450 ();
 TAPCELL_X1 PHY_EDGE_ROW_222_Left_451 ();
 TAPCELL_X1 PHY_EDGE_ROW_223_Left_452 ();
 TAPCELL_X1 PHY_EDGE_ROW_224_Left_453 ();
 TAPCELL_X1 PHY_EDGE_ROW_225_Left_454 ();
 TAPCELL_X1 PHY_EDGE_ROW_226_Left_455 ();
 TAPCELL_X1 PHY_EDGE_ROW_227_Left_456 ();
 TAPCELL_X1 PHY_EDGE_ROW_228_Left_457 ();
 TAPCELL_X1 PHY_EDGE_ROW_229_Left_458 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_1_Left_459 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_2_Left_460 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_2_Left_461 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_2_Left_462 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_2_Left_463 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_2_Left_464 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_2_Left_465 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_2_Left_466 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_2_Left_467 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_2_Left_468 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_2_Left_469 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_2_Left_470 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_2_Left_471 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_2_Left_472 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_2_Left_473 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_2_Left_474 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_2_Left_475 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_2_Left_476 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_2_Left_477 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_2_Left_478 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_2_Left_479 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_2_Left_480 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_2_Left_481 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_2_Left_482 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_2_Left_483 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_2_Left_484 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_2_Left_485 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_2_Left_486 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_2_Left_487 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_2_Left_488 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_2_Left_489 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_2_Left_490 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_2_Left_491 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_2_Left_492 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_2_Left_493 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_2_Left_494 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_2_Left_495 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_2_Left_496 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_2_Left_497 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_2_Left_498 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_2_Left_499 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_2_Left_500 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_2_Left_501 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_2_Left_502 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_2_Left_503 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_2_Left_504 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_2_Left_505 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_2_Left_506 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_2_Left_507 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_2_Left_508 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_2_Left_509 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_2_Left_510 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_2_Left_511 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_2_Left_512 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_2_Left_513 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_2_Left_514 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_2_Left_515 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_2_Left_516 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_2_Left_517 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_2_Left_518 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_2_Left_519 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_2_Left_520 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_2_Left_521 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_2_Left_522 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_2_Left_523 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_2_Left_524 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_2_Left_525 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_2_Left_526 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_2_Left_527 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_2_Left_528 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_2_Left_529 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_2_Left_530 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_2_Left_531 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_2_Left_532 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_2_Left_533 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_2_Left_534 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_2_Left_535 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_2_Left_536 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_2_Left_537 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_2_Left_538 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_2_Left_539 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_2_Left_540 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_2_Left_541 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_2_Left_542 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_2_Left_543 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_2_Left_544 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_2_Left_545 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_2_Left_546 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_2_Left_547 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_2_Left_548 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_2_Left_549 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_2_Left_550 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_2_Left_551 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_2_Left_552 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_2_Left_553 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_2_Left_554 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_2_Left_555 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_2_Left_556 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_2_Left_557 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_2_Left_558 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_2_Left_559 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_2_Left_560 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_2_Left_561 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_2_Left_562 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_2_Left_563 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_2_Left_564 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_2_Left_565 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_2_Left_566 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_2_Left_567 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_2_Left_568 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_2_Left_569 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_2_Left_570 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_2_Left_571 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_2_Left_572 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_2_Left_573 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_2_Left_574 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_2_Left_575 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_2_Left_576 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_2_Left_577 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_2_Left_578 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_2_Left_579 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_2_Left_580 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_2_Left_581 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_2_Left_582 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_2_Left_583 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_2_Left_584 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_2_Left_585 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_2_Left_586 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_2_Left_587 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_2_Left_588 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_2_Left_589 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_2_Left_590 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_2_Left_591 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_2_Left_592 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_2_Left_593 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_2_Left_594 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_2_Left_595 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_2_Left_596 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_2_Left_597 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_2_Left_598 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_2_Left_599 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_2_Left_600 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_2_Left_601 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_2_Left_602 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_2_Left_603 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_2_Left_604 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_2_Left_605 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_2_Left_606 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_2_Left_607 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_2_Left_608 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_2_Left_609 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_2_Left_610 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_2_Left_611 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_2_Left_612 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_2_Left_613 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_2_Left_614 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_2_Left_615 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_2_Left_616 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_2_Left_617 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_2_Left_618 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_2_Left_619 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_2_Left_620 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_2_Left_621 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_2_Left_622 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_2_Left_623 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_2_Left_624 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_2_Left_625 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_2_Left_626 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_2_Left_627 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_1_Right_628 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_1_Right_629 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_1_Right_630 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_1_Right_631 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_1_Right_632 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_1_Right_633 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_1_Right_634 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_1_Right_635 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_1_Right_636 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_1_Right_637 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_1_Right_638 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_1_Right_639 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_1_Right_640 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_1_Right_641 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_1_Right_642 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_1_Right_643 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_1_Right_644 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_1_Right_645 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_1_Right_646 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_1_Right_647 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_1_Right_648 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_1_Right_649 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_1_Right_650 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_1_Right_651 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_1_Right_652 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_1_Right_653 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_1_Right_654 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_1_Right_655 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_1_Right_656 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_1_Right_657 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_1_Right_658 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_1_Right_659 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_1_Right_660 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_1_Right_661 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_1_Right_662 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_1_Right_663 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_1_Right_664 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_1_Right_665 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_1_Right_666 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_1_Right_667 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_1_Right_668 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_1_Right_669 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_1_Right_670 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_1_Right_671 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_1_Right_672 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_1_Right_673 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_1_Right_674 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_1_Right_675 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_1_Right_676 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_1_Right_677 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_1_Right_678 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_1_Right_679 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_1_Right_680 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_1_Right_681 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_1_Right_682 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_1_Right_683 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_1_Right_684 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_1_Right_685 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_1_Right_686 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_1_Right_687 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_1_Right_688 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_1_Right_689 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_1_Right_690 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_1_Right_691 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_1_Right_692 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_1_Right_693 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_1_Right_694 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_1_Right_695 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_1_Right_696 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_1_Right_697 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_1_Right_698 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_1_Right_699 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_1_Right_700 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_1_Right_701 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_1_Right_702 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_1_Right_703 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_1_Right_704 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_1_Right_705 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_1_Right_706 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_1_Right_707 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_1_Right_708 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_1_Right_709 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_1_Right_710 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_1_Right_711 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_1_Right_712 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_1_Right_713 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_1_Right_714 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_1_Right_715 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_1_Right_716 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_1_Right_717 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_1_Right_718 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_1_Right_719 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_1_Right_720 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_1_Right_721 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_1_Right_722 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_1_Right_723 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_1_Right_724 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_1_Right_725 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_1_Right_726 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_1_Right_727 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_1_Right_728 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_1_Right_729 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_1_Right_730 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_1_Right_731 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_1_Right_732 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_1_Right_733 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_1_Right_734 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_1_Right_735 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_1_Right_736 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_1_Right_737 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_1_Right_738 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_1_Right_739 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_1_Right_740 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_1_Right_741 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_1_Right_742 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_1_Right_743 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_1_Right_744 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_1_Right_745 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_1_Right_746 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_1_Right_747 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_1_Right_748 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_1_Right_749 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_1_Right_750 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_1_Right_751 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_1_Right_752 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_1_Right_753 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_1_Right_754 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_1_Right_755 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_1_Right_756 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_1_Right_757 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_1_Right_758 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_1_Right_759 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_1_Right_760 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_1_Right_761 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_1_Right_762 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_1_Right_763 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_1_Right_764 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_1_Right_765 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_1_Right_766 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_1_Right_767 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_1_Right_768 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_1_Right_769 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_1_Right_770 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_1_Right_771 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_1_Right_772 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_1_Right_773 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_1_Right_774 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_1_Right_775 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_1_Right_776 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_1_Right_777 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_1_Right_778 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_1_Right_779 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_1_Right_780 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_1_Right_781 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_1_Right_782 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_1_Right_783 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_1_Right_784 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_1_Right_785 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_1_Right_786 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_1_Right_787 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_1_Right_788 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_1_Right_789 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_1_Right_790 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_1_Right_791 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_1_Right_792 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_1_Right_793 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_1_Right_794 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_1_Right_795 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_796 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_797 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_798 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_799 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_800 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_801 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_802 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_803 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_804 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_805 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_806 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_807 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_808 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_809 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_810 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_811 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_812 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_813 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_814 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_815 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_816 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_817 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_818 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_819 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_820 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_821 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_822 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_823 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_824 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_825 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_826 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_827 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_828 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_829 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_830 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_831 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_832 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_833 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_834 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_835 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_836 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_837 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_208_838 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_208_839 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_209_840 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_210_841 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_211_842 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_212_843 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_213_844 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_214_845 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_215_846 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_216_847 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_217_848 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_218_849 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_219_850 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_220_851 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_221_852 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_222_853 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_223_854 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_224_855 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_225_856 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_226_857 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_227_858 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_228_859 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_229_860 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_229_861 ();
 LOGIC1_X1 \u_multiplier/NOD/nod_cels[29].Nod_bits/_07__125  (.Z(net125));
 CLKBUF_X1 hold126 (.A(net202),
    .Z(net126));
 BUF_X16 max_cap17 (.A(\u_multiplier/_3313_ ),
    .Z(net17));
 BUF_X8 max_cap18 (.A(net19),
    .Z(net18));
 BUF_X8 wire19 (.A(\u_multiplier/_1865_ ),
    .Z(net19));
 BUF_X8 max_cap20 (.A(\u_multiplier/_1864_ ),
    .Z(net20));
 BUF_X16 max_cap21 (.A(\u_multiplier/_3333_ ),
    .Z(net21));
 BUF_X16 max_length22 (.A(_0304_),
    .Z(net22));
 BUF_X16 max_length23 (.A(_0304_),
    .Z(net23));
 BUF_X4 input24 (.A(data_in[0]),
    .Z(net24));
 BUF_X4 input25 (.A(data_in[10]),
    .Z(net25));
 BUF_X2 input26 (.A(data_in[11]),
    .Z(net26));
 BUF_X1 input27 (.A(data_in[12]),
    .Z(net27));
 CLKBUF_X3 input28 (.A(data_in[13]),
    .Z(net28));
 BUF_X4 input29 (.A(data_in[14]),
    .Z(net29));
 BUF_X1 input30 (.A(data_in[15]),
    .Z(net30));
 BUF_X2 input31 (.A(data_in[16]),
    .Z(net31));
 CLKBUF_X3 input32 (.A(data_in[17]),
    .Z(net32));
 BUF_X1 input33 (.A(data_in[18]),
    .Z(net33));
 BUF_X4 input34 (.A(data_in[19]),
    .Z(net34));
 CLKBUF_X2 input35 (.A(data_in[1]),
    .Z(net35));
 CLKBUF_X3 input36 (.A(data_in[20]),
    .Z(net36));
 CLKBUF_X3 input37 (.A(data_in[21]),
    .Z(net37));
 CLKBUF_X3 input38 (.A(data_in[22]),
    .Z(net38));
 BUF_X4 input39 (.A(data_in[23]),
    .Z(net39));
 BUF_X1 input40 (.A(data_in[24]),
    .Z(net40));
 CLKBUF_X3 input41 (.A(data_in[25]),
    .Z(net41));
 BUF_X4 input42 (.A(data_in[26]),
    .Z(net42));
 BUF_X4 input43 (.A(data_in[27]),
    .Z(net43));
 BUF_X1 input44 (.A(data_in[28]),
    .Z(net44));
 CLKBUF_X2 input45 (.A(data_in[29]),
    .Z(net45));
 CLKBUF_X2 input46 (.A(data_in[2]),
    .Z(net46));
 BUF_X2 input47 (.A(data_in[30]),
    .Z(net47));
 BUF_X2 input48 (.A(data_in[31]),
    .Z(net48));
 BUF_X4 input49 (.A(data_in[3]),
    .Z(net49));
 BUF_X4 input50 (.A(data_in[4]),
    .Z(net50));
 CLKBUF_X3 input51 (.A(data_in[5]),
    .Z(net51));
 BUF_X1 input52 (.A(data_in[6]),
    .Z(net52));
 BUF_X2 input53 (.A(data_in[7]),
    .Z(net53));
 CLKBUF_X3 input54 (.A(data_in[8]),
    .Z(net54));
 BUF_X4 input55 (.A(data_in[9]),
    .Z(net55));
 BUF_X4 input56 (.A(init_enable),
    .Z(net56));
 BUF_X4 input57 (.A(pe_ce),
    .Z(net57));
 BUF_X32 input58 (.A(rst_n),
    .Z(net58));
 BUF_X1 output59 (.A(net59),
    .Z(curr_state[1]));
 BUF_X1 output60 (.A(net60),
    .Z(data_out[0]));
 BUF_X1 output61 (.A(net61),
    .Z(data_out[10]));
 BUF_X1 output62 (.A(net62),
    .Z(data_out[11]));
 BUF_X1 output63 (.A(net63),
    .Z(data_out[12]));
 BUF_X1 output64 (.A(net64),
    .Z(data_out[13]));
 BUF_X1 output65 (.A(net65),
    .Z(data_out[14]));
 BUF_X1 output66 (.A(net66),
    .Z(data_out[15]));
 BUF_X1 output67 (.A(net67),
    .Z(data_out[16]));
 BUF_X1 output68 (.A(net68),
    .Z(data_out[17]));
 BUF_X1 output69 (.A(net69),
    .Z(data_out[18]));
 BUF_X1 output70 (.A(net70),
    .Z(data_out[19]));
 BUF_X1 output71 (.A(net71),
    .Z(data_out[1]));
 BUF_X1 output72 (.A(net72),
    .Z(data_out[20]));
 BUF_X1 output73 (.A(net73),
    .Z(data_out[21]));
 BUF_X1 output74 (.A(net74),
    .Z(data_out[22]));
 BUF_X1 output75 (.A(net75),
    .Z(data_out[23]));
 BUF_X1 output76 (.A(net76),
    .Z(data_out[24]));
 BUF_X1 output77 (.A(net77),
    .Z(data_out[25]));
 BUF_X1 output78 (.A(net78),
    .Z(data_out[26]));
 BUF_X1 output79 (.A(net79),
    .Z(data_out[27]));
 BUF_X1 output80 (.A(net80),
    .Z(data_out[28]));
 BUF_X1 output81 (.A(net81),
    .Z(data_out[29]));
 BUF_X1 output82 (.A(net82),
    .Z(data_out[2]));
 BUF_X1 output83 (.A(net83),
    .Z(data_out[30]));
 BUF_X1 output84 (.A(net84),
    .Z(data_out[31]));
 BUF_X1 output85 (.A(net85),
    .Z(data_out[32]));
 BUF_X1 output86 (.A(net86),
    .Z(data_out[33]));
 BUF_X1 output87 (.A(net87),
    .Z(data_out[34]));
 BUF_X1 output88 (.A(net88),
    .Z(data_out[35]));
 BUF_X1 output89 (.A(net89),
    .Z(data_out[36]));
 BUF_X1 output90 (.A(net90),
    .Z(data_out[37]));
 BUF_X1 output91 (.A(net91),
    .Z(data_out[38]));
 BUF_X1 output92 (.A(net92),
    .Z(data_out[39]));
 BUF_X1 output93 (.A(net93),
    .Z(data_out[3]));
 BUF_X1 output94 (.A(net94),
    .Z(data_out[40]));
 BUF_X1 output95 (.A(net95),
    .Z(data_out[41]));
 BUF_X1 output96 (.A(net96),
    .Z(data_out[42]));
 BUF_X1 output97 (.A(net97),
    .Z(data_out[43]));
 BUF_X1 output98 (.A(net98),
    .Z(data_out[44]));
 BUF_X1 output99 (.A(net99),
    .Z(data_out[45]));
 BUF_X1 output100 (.A(net100),
    .Z(data_out[46]));
 BUF_X1 output101 (.A(net101),
    .Z(data_out[47]));
 BUF_X1 output102 (.A(net102),
    .Z(data_out[48]));
 BUF_X1 output103 (.A(net103),
    .Z(data_out[49]));
 BUF_X1 output104 (.A(net104),
    .Z(data_out[4]));
 BUF_X1 output105 (.A(net105),
    .Z(data_out[50]));
 BUF_X1 output106 (.A(net106),
    .Z(data_out[51]));
 BUF_X1 output107 (.A(net107),
    .Z(data_out[52]));
 BUF_X1 output108 (.A(net108),
    .Z(data_out[53]));
 BUF_X1 output109 (.A(net109),
    .Z(data_out[54]));
 BUF_X1 output110 (.A(net110),
    .Z(data_out[55]));
 BUF_X1 output111 (.A(net111),
    .Z(data_out[56]));
 BUF_X1 output112 (.A(net112),
    .Z(data_out[57]));
 BUF_X1 output113 (.A(net113),
    .Z(data_out[58]));
 BUF_X1 output114 (.A(net114),
    .Z(data_out[59]));
 BUF_X1 output115 (.A(net115),
    .Z(data_out[5]));
 BUF_X1 output116 (.A(net116),
    .Z(data_out[60]));
 BUF_X1 output117 (.A(net117),
    .Z(data_out[61]));
 BUF_X1 output118 (.A(net118),
    .Z(data_out[62]));
 BUF_X1 output119 (.A(net119),
    .Z(data_out[63]));
 BUF_X1 output120 (.A(net120),
    .Z(data_out[6]));
 BUF_X1 output121 (.A(net121),
    .Z(data_out[7]));
 BUF_X1 output122 (.A(net122),
    .Z(data_out[8]));
 BUF_X1 output123 (.A(net123),
    .Z(data_out[9]));
 BUF_X1 output124 (.A(net124),
    .Z(valid_reg_out));
 CLKBUF_X1 hold127 (.A(_0165_),
    .Z(net127));
 CLKBUF_X1 hold128 (.A(net9),
    .Z(net128));
 CLKBUF_X1 hold129 (.A(net184),
    .Z(net129));
 CLKBUF_X1 hold130 (.A(net189),
    .Z(net130));
 CLKBUF_X1 hold131 (.A(net160),
    .Z(net131));
 CLKBUF_X1 hold132 (.A(net167),
    .Z(net132));
 CLKBUF_X1 hold133 (.A(net194),
    .Z(net133));
 CLKBUF_X1 hold134 (.A(net196),
    .Z(net134));
 CLKBUF_X1 hold135 (.A(net157),
    .Z(net135));
 CLKBUF_X1 hold136 (.A(net173),
    .Z(net136));
 CLKBUF_X1 hold137 (.A(net176),
    .Z(net137));
 CLKBUF_X1 hold138 (.A(net179),
    .Z(net138));
 CLKBUF_X1 hold139 (.A(net201),
    .Z(net139));
 CLKBUF_X1 hold140 (.A(net192),
    .Z(net140));
 CLKBUF_X1 hold141 (.A(net207),
    .Z(net141));
 CLKBUF_X1 hold142 (.A(net212),
    .Z(net142));
 CLKBUF_X1 hold143 (.A(net198),
    .Z(net143));
 CLKBUF_X1 hold144 (.A(net203),
    .Z(net144));
 CLKBUF_X1 hold145 (.A(net210),
    .Z(net145));
 CLKBUF_X1 hold146 (.A(net209),
    .Z(net146));
 CLKBUF_X1 hold147 (.A(net204),
    .Z(net147));
 CLKBUF_X1 hold148 (.A(net200),
    .Z(net148));
 CLKBUF_X1 hold149 (.A(net213),
    .Z(net149));
 CLKBUF_X1 hold150 (.A(net211),
    .Z(net150));
 CLKBUF_X1 hold151 (.A(net208),
    .Z(net151));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_1_0_0_clk));
 CLKBUF_X3 clkbuf_1_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_1_1_0_clk));
 CLKBUF_X3 clkbuf_2_0_0_clk (.A(clknet_1_0_0_clk),
    .Z(clknet_2_0_0_clk));
 CLKBUF_X3 clkbuf_2_1_0_clk (.A(clknet_1_0_0_clk),
    .Z(clknet_2_1_0_clk));
 CLKBUF_X3 clkbuf_2_2_0_clk (.A(clknet_1_1_0_clk),
    .Z(clknet_2_2_0_clk));
 CLKBUF_X3 clkbuf_2_3_0_clk (.A(clknet_1_1_0_clk),
    .Z(clknet_2_3_0_clk));
 CLKBUF_X3 clkbuf_4_0__f_clk (.A(clknet_2_0_0_clk),
    .Z(clknet_4_0__leaf_clk));
 CLKBUF_X3 clkbuf_4_1__f_clk (.A(clknet_2_0_0_clk),
    .Z(clknet_4_1__leaf_clk));
 CLKBUF_X3 clkbuf_4_2__f_clk (.A(clknet_2_0_0_clk),
    .Z(clknet_4_2__leaf_clk));
 CLKBUF_X3 clkbuf_4_3__f_clk (.A(clknet_2_0_0_clk),
    .Z(clknet_4_3__leaf_clk));
 CLKBUF_X3 clkbuf_4_4__f_clk (.A(clknet_2_1_0_clk),
    .Z(clknet_4_4__leaf_clk));
 CLKBUF_X3 clkbuf_4_5__f_clk (.A(clknet_2_1_0_clk),
    .Z(clknet_4_5__leaf_clk));
 CLKBUF_X3 clkbuf_4_6__f_clk (.A(clknet_2_1_0_clk),
    .Z(clknet_4_6__leaf_clk));
 CLKBUF_X3 clkbuf_4_7__f_clk (.A(clknet_2_1_0_clk),
    .Z(clknet_4_7__leaf_clk));
 CLKBUF_X3 clkbuf_4_8__f_clk (.A(clknet_2_2_0_clk),
    .Z(clknet_4_8__leaf_clk));
 CLKBUF_X3 clkbuf_4_9__f_clk (.A(clknet_2_2_0_clk),
    .Z(clknet_4_9__leaf_clk));
 CLKBUF_X3 clkbuf_4_10__f_clk (.A(clknet_2_2_0_clk),
    .Z(clknet_4_10__leaf_clk));
 CLKBUF_X3 clkbuf_4_11__f_clk (.A(clknet_2_2_0_clk),
    .Z(clknet_4_11__leaf_clk));
 CLKBUF_X3 clkbuf_4_12__f_clk (.A(clknet_2_3_0_clk),
    .Z(clknet_4_12__leaf_clk));
 CLKBUF_X3 clkbuf_4_13__f_clk (.A(clknet_2_3_0_clk),
    .Z(clknet_4_13__leaf_clk));
 CLKBUF_X3 clkbuf_4_14__f_clk (.A(clknet_2_3_0_clk),
    .Z(clknet_4_14__leaf_clk));
 CLKBUF_X3 clkbuf_4_15__f_clk (.A(clknet_2_3_0_clk),
    .Z(clknet_4_15__leaf_clk));
 INV_X2 clkload0 (.A(clknet_4_0__leaf_clk));
 INV_X2 clkload1 (.A(clknet_4_1__leaf_clk));
 INV_X2 clkload2 (.A(clknet_4_2__leaf_clk));
 INV_X2 clkload3 (.A(clknet_4_4__leaf_clk));
 INV_X2 clkload4 (.A(clknet_4_6__leaf_clk));
 INV_X4 clkload5 (.A(clknet_4_7__leaf_clk));
 INV_X4 clkload6 (.A(clknet_4_8__leaf_clk));
 INV_X2 clkload7 (.A(clknet_4_9__leaf_clk));
 INV_X2 clkload8 (.A(clknet_4_11__leaf_clk));
 CLKBUF_X1 clkload9 (.A(clknet_4_12__leaf_clk));
 INV_X2 clkload10 (.A(clknet_4_14__leaf_clk));
 INV_X1 clkload11 (.A(clknet_4_15__leaf_clk));
 CLKBUF_X1 hold1 (.A(net214),
    .Z(net1));
 CLKBUF_X1 hold2 (.A(net215),
    .Z(net2));
 CLKBUF_X1 hold3 (.A(net219),
    .Z(net3));
 CLKBUF_X1 hold4 (.A(net217),
    .Z(net4));
 CLKBUF_X1 hold5 (.A(net222),
    .Z(net5));
 CLKBUF_X1 hold6 (.A(net223),
    .Z(net6));
 CLKBUF_X1 hold7 (.A(net216),
    .Z(net7));
 CLKBUF_X1 hold8 (.A(data_in_reg[5]),
    .Z(net8));
 CLKBUF_X1 hold9 (.A(_0668_),
    .Z(net9));
 CLKBUF_X1 hold10 (.A(net128),
    .Z(net10));
 CLKBUF_X1 hold11 (.A(_0270_),
    .Z(net11));
 CLKBUF_X1 hold12 (.A(curr_state[0]),
    .Z(net12));
 CLKBUF_X1 hold13 (.A(_0372_),
    .Z(net13));
 CLKBUF_X1 hold14 (.A(_0663_),
    .Z(net14));
 CLKBUF_X1 hold15 (.A(_0427_),
    .Z(net15));
 CLKBUF_X1 hold16 (.A(net218),
    .Z(net16));
 CLKBUF_X1 hold17 (.A(net220),
    .Z(net152));
 CLKBUF_X1 hold18 (.A(_0662_),
    .Z(net153));
 CLKBUF_X1 hold19 (.A(_0425_),
    .Z(net154));
 CLKBUF_X1 hold20 (.A(data_in_reg[0]),
    .Z(net155));
 CLKBUF_X1 hold21 (.A(net225),
    .Z(net156));
 CLKBUF_X1 hold22 (.A(_0669_),
    .Z(net157));
 CLKBUF_X1 hold23 (.A(net135),
    .Z(net158));
 CLKBUF_X1 hold24 (.A(_0271_),
    .Z(net159));
 CLKBUF_X1 hold25 (.A(_0658_),
    .Z(net160));
 CLKBUF_X1 hold26 (.A(net131),
    .Z(net161));
 CLKBUF_X1 hold27 (.A(_0164_),
    .Z(net162));
 CLKBUF_X1 hold28 (.A(_0592_),
    .Z(net163));
 CLKBUF_X1 hold29 (.A(_0386_),
    .Z(net164));
 CLKBUF_X1 hold30 (.A(_0307_),
    .Z(net165));
 CLKBUF_X1 hold31 (.A(data_in_reg[18]),
    .Z(net166));
 CLKBUF_X1 hold32 (.A(_0664_),
    .Z(net167));
 CLKBUF_X1 hold33 (.A(net132),
    .Z(net168));
 CLKBUF_X1 hold34 (.A(_0266_),
    .Z(net169));
 CLKBUF_X1 hold35 (.A(data_in_reg[13]),
    .Z(net170));
 CLKBUF_X1 hold36 (.A(_0683_[29]),
    .Z(net171));
 CLKBUF_X1 hold37 (.A(net221),
    .Z(net172));
 CLKBUF_X1 hold38 (.A(_0667_),
    .Z(net173));
 CLKBUF_X1 hold39 (.A(net136),
    .Z(net174));
 CLKBUF_X1 hold40 (.A(_0269_),
    .Z(net175));
 CLKBUF_X1 hold41 (.A(_0666_),
    .Z(net176));
 CLKBUF_X1 hold42 (.A(net137),
    .Z(net177));
 CLKBUF_X1 hold43 (.A(_0268_),
    .Z(net178));
 CLKBUF_X1 hold44 (.A(_0665_),
    .Z(net179));
 CLKBUF_X1 hold45 (.A(net138),
    .Z(net180));
 CLKBUF_X1 hold46 (.A(_0267_),
    .Z(net181));
 CLKBUF_X1 hold47 (.A(data_in_reg[6]),
    .Z(net182));
 CLKBUF_X1 hold48 (.A(\u_multiplier/LODx/z [11]),
    .Z(net183));
 CLKBUF_X1 hold49 (.A(addr_ptr[4]),
    .Z(net184));
 CLKBUF_X1 hold50 (.A(net129),
    .Z(net185));
 CLKBUF_X1 hold51 (.A(\u_multiplier/LODx/z [3]),
    .Z(net186));
 CLKBUF_X1 hold52 (.A(data_in_reg[10]),
    .Z(net187));
 CLKBUF_X1 hold53 (.A(\u_multiplier/LODx/z [15]),
    .Z(net188));
 CLKBUF_X1 hold54 (.A(addr_ptr[5]),
    .Z(net189));
 CLKBUF_X1 hold55 (.A(net130),
    .Z(net190));
 CLKBUF_X1 hold56 (.A(data_in_reg[16]),
    .Z(net191));
 CLKBUF_X1 hold57 (.A(_0660_),
    .Z(net192));
 CLKBUF_X1 hold58 (.A(net140),
    .Z(net193));
 CLKBUF_X1 hold59 (.A(addr_ptr[2]),
    .Z(net194));
 CLKBUF_X1 hold60 (.A(net133),
    .Z(net195));
 CLKBUF_X1 hold61 (.A(addr_ptr[3]),
    .Z(net196));
 CLKBUF_X1 hold62 (.A(net134),
    .Z(net197));
 CLKBUF_X1 hold63 (.A(data_in_reg[24]),
    .Z(net198));
 CLKBUF_X1 hold64 (.A(net143),
    .Z(net199));
 CLKBUF_X1 hold65 (.A(_0683_[26]),
    .Z(net200));
 CLKBUF_X1 hold66 (.A(addr_ptr[1]),
    .Z(net201));
 CLKBUF_X1 hold67 (.A(_0659_),
    .Z(net202));
 CLKBUF_X1 hold68 (.A(\u_multiplier/LODx/z [31]),
    .Z(net203));
 CLKBUF_X1 hold69 (.A(_0661_),
    .Z(net204));
 CLKBUF_X1 hold70 (.A(curr_state[2]),
    .Z(net205));
 CLKBUF_X1 hold71 (.A(_0683_[30]),
    .Z(net206));
 CLKBUF_X1 hold72 (.A(addr_ptr[0]),
    .Z(net207));
 CLKBUF_X1 hold73 (.A(data_in_reg[12]),
    .Z(net208));
 CLKBUF_X1 hold74 (.A(data_in_reg[21]),
    .Z(net209));
 CLKBUF_X1 hold75 (.A(_0683_[25]),
    .Z(net210));
 CLKBUF_X1 hold76 (.A(\u_multiplier/LODx/z [23]),
    .Z(net211));
 CLKBUF_X1 hold77 (.A(data_in_reg[20]),
    .Z(net212));
 CLKBUF_X1 hold78 (.A(_0683_[28]),
    .Z(net213));
 CLKBUF_X1 hold79 (.A(\u_multiplier/LODx/z [27]),
    .Z(net214));
 CLKBUF_X1 hold80 (.A(data_in_reg[4]),
    .Z(net215));
 CLKBUF_X1 hold81 (.A(data_in_reg[1]),
    .Z(net216));
 CLKBUF_X1 hold82 (.A(data_in_reg[22]),
    .Z(net217));
 CLKBUF_X1 hold83 (.A(\u_multiplier/LODx/z [19]),
    .Z(net218));
 CLKBUF_X1 hold84 (.A(data_in_reg[14]),
    .Z(net219));
 CLKBUF_X1 hold85 (.A(data_in_reg[9]),
    .Z(net220));
 CLKBUF_X1 hold86 (.A(data_in_reg[17]),
    .Z(net221));
 CLKBUF_X1 hold87 (.A(data_in_reg[8]),
    .Z(net222));
 CLKBUF_X1 hold88 (.A(data_in_reg[2]),
    .Z(net223));
 CLKBUF_X1 hold89 (.A(init_count[5]),
    .Z(net224));
 CLKBUF_X1 hold90 (.A(\u_multiplier/LODx/z [7]),
    .Z(net225));
 FILLCELL_X4 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_8 ();
 FILLCELL_X4 FILLER_0_40 ();
 FILLCELL_X32 FILLER_0_47 ();
 FILLCELL_X32 FILLER_0_79 ();
 FILLCELL_X4 FILLER_0_111 ();
 FILLCELL_X32 FILLER_0_118 ();
 FILLCELL_X16 FILLER_0_150 ();
 FILLCELL_X8 FILLER_0_166 ();
 FILLCELL_X4 FILLER_0_174 ();
 FILLCELL_X2 FILLER_0_178 ();
 FILLCELL_X32 FILLER_0_184 ();
 FILLCELL_X32 FILLER_0_216 ();
 FILLCELL_X2 FILLER_0_248 ();
 FILLCELL_X1 FILLER_0_250 ();
 FILLCELL_X32 FILLER_0_254 ();
 FILLCELL_X32 FILLER_0_286 ();
 FILLCELL_X2 FILLER_0_318 ();
 FILLCELL_X1 FILLER_0_320 ();
 FILLCELL_X32 FILLER_0_324 ();
 FILLCELL_X16 FILLER_0_356 ();
 FILLCELL_X8 FILLER_0_372 ();
 FILLCELL_X4 FILLER_0_380 ();
 FILLCELL_X2 FILLER_0_384 ();
 FILLCELL_X16 FILLER_0_389 ();
 FILLCELL_X8 FILLER_0_405 ();
 FILLCELL_X2 FILLER_0_413 ();
 FILLCELL_X16 FILLER_0_419 ();
 FILLCELL_X2 FILLER_0_435 ();
 FILLCELL_X1 FILLER_0_437 ();
 FILLCELL_X8 FILLER_0_442 ();
 FILLCELL_X4 FILLER_0_450 ();
 FILLCELL_X2 FILLER_0_454 ();
 FILLCELL_X1 FILLER_0_456 ();
 FILLCELL_X4 FILLER_0_460 ();
 FILLCELL_X1 FILLER_0_464 ();
 FILLCELL_X8 FILLER_0_469 ();
 FILLCELL_X2 FILLER_0_477 ();
 FILLCELL_X1 FILLER_0_479 ();
 FILLCELL_X32 FILLER_0_489 ();
 FILLCELL_X1 FILLER_0_521 ();
 FILLCELL_X8 FILLER_0_525 ();
 FILLCELL_X2 FILLER_0_533 ();
 FILLCELL_X1 FILLER_0_535 ();
 FILLCELL_X8 FILLER_0_541 ();
 FILLCELL_X2 FILLER_0_549 ();
 FILLCELL_X1 FILLER_0_551 ();
 FILLCELL_X8 FILLER_0_556 ();
 FILLCELL_X4 FILLER_0_568 ();
 FILLCELL_X16 FILLER_0_575 ();
 FILLCELL_X1 FILLER_0_591 ();
 FILLCELL_X8 FILLER_0_595 ();
 FILLCELL_X4 FILLER_0_603 ();
 FILLCELL_X4 FILLER_0_611 ();
 FILLCELL_X8 FILLER_0_618 ();
 FILLCELL_X4 FILLER_0_626 ();
 FILLCELL_X1 FILLER_0_630 ();
 FILLCELL_X4 FILLER_0_632 ();
 FILLCELL_X1 FILLER_0_636 ();
 FILLCELL_X4 FILLER_0_639 ();
 FILLCELL_X16 FILLER_0_647 ();
 FILLCELL_X16 FILLER_0_667 ();
 FILLCELL_X2 FILLER_0_683 ();
 FILLCELL_X4 FILLER_0_688 ();
 FILLCELL_X4 FILLER_0_695 ();
 FILLCELL_X8 FILLER_0_701 ();
 FILLCELL_X4 FILLER_0_713 ();
 FILLCELL_X1 FILLER_0_717 ();
 FILLCELL_X4 FILLER_0_721 ();
 FILLCELL_X8 FILLER_0_729 ();
 FILLCELL_X4 FILLER_0_741 ();
 FILLCELL_X8 FILLER_0_752 ();
 FILLCELL_X1 FILLER_0_760 ();
 FILLCELL_X4 FILLER_0_764 ();
 FILLCELL_X8 FILLER_0_770 ();
 FILLCELL_X1 FILLER_0_778 ();
 FILLCELL_X16 FILLER_0_783 ();
 FILLCELL_X16 FILLER_0_802 ();
 FILLCELL_X8 FILLER_0_818 ();
 FILLCELL_X2 FILLER_0_826 ();
 FILLCELL_X1 FILLER_0_828 ();
 FILLCELL_X4 FILLER_0_831 ();
 FILLCELL_X8 FILLER_0_838 ();
 FILLCELL_X2 FILLER_0_846 ();
 FILLCELL_X8 FILLER_0_852 ();
 FILLCELL_X2 FILLER_0_860 ();
 FILLCELL_X8 FILLER_0_871 ();
 FILLCELL_X1 FILLER_0_879 ();
 FILLCELL_X4 FILLER_0_887 ();
 FILLCELL_X4 FILLER_0_894 ();
 FILLCELL_X16 FILLER_0_905 ();
 FILLCELL_X4 FILLER_0_924 ();
 FILLCELL_X4 FILLER_0_931 ();
 FILLCELL_X2 FILLER_0_935 ();
 FILLCELL_X1 FILLER_0_937 ();
 FILLCELL_X4 FILLER_0_942 ();
 FILLCELL_X8 FILLER_0_950 ();
 FILLCELL_X4 FILLER_0_958 ();
 FILLCELL_X1 FILLER_0_962 ();
 FILLCELL_X4 FILLER_0_966 ();
 FILLCELL_X2 FILLER_0_970 ();
 FILLCELL_X1 FILLER_0_972 ();
 FILLCELL_X16 FILLER_0_976 ();
 FILLCELL_X8 FILLER_0_992 ();
 FILLCELL_X4 FILLER_0_1000 ();
 FILLCELL_X1 FILLER_0_1004 ();
 FILLCELL_X4 FILLER_0_1008 ();
 FILLCELL_X2 FILLER_0_1012 ();
 FILLCELL_X16 FILLER_0_1023 ();
 FILLCELL_X1 FILLER_0_1039 ();
 FILLCELL_X8 FILLER_0_1049 ();
 FILLCELL_X2 FILLER_0_1057 ();
 FILLCELL_X4 FILLER_0_1066 ();
 FILLCELL_X4 FILLER_0_1073 ();
 FILLCELL_X4 FILLER_0_1080 ();
 FILLCELL_X8 FILLER_0_1087 ();
 FILLCELL_X4 FILLER_0_1095 ();
 FILLCELL_X1 FILLER_0_1099 ();
 FILLCELL_X32 FILLER_0_1103 ();
 FILLCELL_X4 FILLER_0_1135 ();
 FILLCELL_X1 FILLER_0_1139 ();
 FILLCELL_X4 FILLER_0_1143 ();
 FILLCELL_X4 FILLER_0_1151 ();
 FILLCELL_X4 FILLER_0_1162 ();
 FILLCELL_X16 FILLER_0_1173 ();
 FILLCELL_X4 FILLER_0_1189 ();
 FILLCELL_X2 FILLER_0_1193 ();
 FILLCELL_X1 FILLER_0_1195 ();
 FILLCELL_X4 FILLER_0_1200 ();
 FILLCELL_X2 FILLER_0_1204 ();
 FILLCELL_X4 FILLER_0_1213 ();
 FILLCELL_X32 FILLER_0_1221 ();
 FILLCELL_X8 FILLER_0_1253 ();
 FILLCELL_X1 FILLER_0_1261 ();
 FILLCELL_X8 FILLER_0_1263 ();
 FILLCELL_X4 FILLER_0_1271 ();
 FILLCELL_X1 FILLER_0_1275 ();
 FILLCELL_X32 FILLER_0_1279 ();
 FILLCELL_X32 FILLER_0_1311 ();
 FILLCELL_X4 FILLER_0_1343 ();
 FILLCELL_X32 FILLER_0_1350 ();
 FILLCELL_X16 FILLER_0_1382 ();
 FILLCELL_X8 FILLER_0_1398 ();
 FILLCELL_X4 FILLER_0_1406 ();
 FILLCELL_X2 FILLER_0_1410 ();
 FILLCELL_X32 FILLER_0_1415 ();
 FILLCELL_X32 FILLER_0_1447 ();
 FILLCELL_X4 FILLER_0_1479 ();
 FILLCELL_X32 FILLER_0_1486 ();
 FILLCELL_X16 FILLER_0_1518 ();
 FILLCELL_X8 FILLER_0_1534 ();
 FILLCELL_X4 FILLER_0_1542 ();
 FILLCELL_X1 FILLER_0_1546 ();
 FILLCELL_X32 FILLER_0_1550 ();
 FILLCELL_X32 FILLER_0_1582 ();
 FILLCELL_X4 FILLER_0_1614 ();
 FILLCELL_X32 FILLER_0_1621 ();
 FILLCELL_X32 FILLER_0_1653 ();
 FILLCELL_X4 FILLER_0_1685 ();
 FILLCELL_X8 FILLER_0_1692 ();
 FILLCELL_X1 FILLER_0_1700 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X32 FILLER_1_257 ();
 FILLCELL_X32 FILLER_1_289 ();
 FILLCELL_X32 FILLER_1_321 ();
 FILLCELL_X16 FILLER_1_353 ();
 FILLCELL_X8 FILLER_1_369 ();
 FILLCELL_X4 FILLER_1_377 ();
 FILLCELL_X1 FILLER_1_381 ();
 FILLCELL_X8 FILLER_1_401 ();
 FILLCELL_X8 FILLER_1_426 ();
 FILLCELL_X1 FILLER_1_434 ();
 FILLCELL_X4 FILLER_1_452 ();
 FILLCELL_X4 FILLER_1_473 ();
 FILLCELL_X4 FILLER_1_486 ();
 FILLCELL_X8 FILLER_1_507 ();
 FILLCELL_X4 FILLER_1_515 ();
 FILLCELL_X1 FILLER_1_519 ();
 FILLCELL_X4 FILLER_1_533 ();
 FILLCELL_X4 FILLER_1_541 ();
 FILLCELL_X8 FILLER_1_550 ();
 FILLCELL_X1 FILLER_1_558 ();
 FILLCELL_X4 FILLER_1_563 ();
 FILLCELL_X4 FILLER_1_571 ();
 FILLCELL_X4 FILLER_1_582 ();
 FILLCELL_X8 FILLER_1_593 ();
 FILLCELL_X4 FILLER_1_605 ();
 FILLCELL_X4 FILLER_1_613 ();
 FILLCELL_X4 FILLER_1_626 ();
 FILLCELL_X8 FILLER_1_640 ();
 FILLCELL_X2 FILLER_1_648 ();
 FILLCELL_X4 FILLER_1_657 ();
 FILLCELL_X2 FILLER_1_661 ();
 FILLCELL_X1 FILLER_1_663 ();
 FILLCELL_X4 FILLER_1_678 ();
 FILLCELL_X8 FILLER_1_692 ();
 FILLCELL_X1 FILLER_1_700 ();
 FILLCELL_X4 FILLER_1_718 ();
 FILLCELL_X8 FILLER_1_741 ();
 FILLCELL_X1 FILLER_1_749 ();
 FILLCELL_X8 FILLER_1_759 ();
 FILLCELL_X4 FILLER_1_774 ();
 FILLCELL_X4 FILLER_1_796 ();
 FILLCELL_X4 FILLER_1_817 ();
 FILLCELL_X4 FILLER_1_823 ();
 FILLCELL_X4 FILLER_1_833 ();
 FILLCELL_X2 FILLER_1_837 ();
 FILLCELL_X4 FILLER_1_845 ();
 FILLCELL_X8 FILLER_1_855 ();
 FILLCELL_X2 FILLER_1_863 ();
 FILLCELL_X8 FILLER_1_878 ();
 FILLCELL_X2 FILLER_1_886 ();
 FILLCELL_X4 FILLER_1_897 ();
 FILLCELL_X4 FILLER_1_914 ();
 FILLCELL_X4 FILLER_1_928 ();
 FILLCELL_X4 FILLER_1_939 ();
 FILLCELL_X4 FILLER_1_952 ();
 FILLCELL_X1 FILLER_1_956 ();
 FILLCELL_X8 FILLER_1_961 ();
 FILLCELL_X2 FILLER_1_969 ();
 FILLCELL_X8 FILLER_1_988 ();
 FILLCELL_X2 FILLER_1_996 ();
 FILLCELL_X4 FILLER_1_1015 ();
 FILLCELL_X4 FILLER_1_1033 ();
 FILLCELL_X4 FILLER_1_1050 ();
 FILLCELL_X4 FILLER_1_1063 ();
 FILLCELL_X4 FILLER_1_1076 ();
 FILLCELL_X4 FILLER_1_1084 ();
 FILLCELL_X1 FILLER_1_1088 ();
 FILLCELL_X4 FILLER_1_1102 ();
 FILLCELL_X4 FILLER_1_1115 ();
 FILLCELL_X4 FILLER_1_1136 ();
 FILLCELL_X4 FILLER_1_1157 ();
 FILLCELL_X8 FILLER_1_1168 ();
 FILLCELL_X1 FILLER_1_1176 ();
 FILLCELL_X4 FILLER_1_1186 ();
 FILLCELL_X4 FILLER_1_1209 ();
 FILLCELL_X1 FILLER_1_1213 ();
 FILLCELL_X32 FILLER_1_1231 ();
 FILLCELL_X32 FILLER_1_1264 ();
 FILLCELL_X32 FILLER_1_1296 ();
 FILLCELL_X32 FILLER_1_1328 ();
 FILLCELL_X32 FILLER_1_1360 ();
 FILLCELL_X32 FILLER_1_1392 ();
 FILLCELL_X16 FILLER_1_1424 ();
 FILLCELL_X8 FILLER_1_1440 ();
 FILLCELL_X4 FILLER_1_1448 ();
 FILLCELL_X1 FILLER_1_1452 ();
 FILLCELL_X8 FILLER_1_1457 ();
 FILLCELL_X1 FILLER_1_1465 ();
 FILLCELL_X16 FILLER_1_1483 ();
 FILLCELL_X8 FILLER_1_1499 ();
 FILLCELL_X4 FILLER_1_1507 ();
 FILLCELL_X2 FILLER_1_1511 ();
 FILLCELL_X1 FILLER_1_1513 ();
 FILLCELL_X32 FILLER_1_1518 ();
 FILLCELL_X32 FILLER_1_1550 ();
 FILLCELL_X32 FILLER_1_1582 ();
 FILLCELL_X32 FILLER_1_1614 ();
 FILLCELL_X32 FILLER_1_1646 ();
 FILLCELL_X8 FILLER_1_1678 ();
 FILLCELL_X4 FILLER_1_1686 ();
 FILLCELL_X2 FILLER_1_1690 ();
 FILLCELL_X1 FILLER_1_1692 ();
 FILLCELL_X4 FILLER_1_1697 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X32 FILLER_2_289 ();
 FILLCELL_X32 FILLER_2_321 ();
 FILLCELL_X32 FILLER_2_353 ();
 FILLCELL_X4 FILLER_2_385 ();
 FILLCELL_X4 FILLER_2_393 ();
 FILLCELL_X8 FILLER_2_401 ();
 FILLCELL_X4 FILLER_2_409 ();
 FILLCELL_X1 FILLER_2_413 ();
 FILLCELL_X4 FILLER_2_418 ();
 FILLCELL_X1 FILLER_2_422 ();
 FILLCELL_X4 FILLER_2_425 ();
 FILLCELL_X4 FILLER_2_433 ();
 FILLCELL_X4 FILLER_2_443 ();
 FILLCELL_X4 FILLER_2_451 ();
 FILLCELL_X16 FILLER_2_458 ();
 FILLCELL_X4 FILLER_2_477 ();
 FILLCELL_X8 FILLER_2_485 ();
 FILLCELL_X2 FILLER_2_493 ();
 FILLCELL_X1 FILLER_2_495 ();
 FILLCELL_X4 FILLER_2_500 ();
 FILLCELL_X2 FILLER_2_504 ();
 FILLCELL_X1 FILLER_2_506 ();
 FILLCELL_X4 FILLER_2_514 ();
 FILLCELL_X2 FILLER_2_518 ();
 FILLCELL_X8 FILLER_2_529 ();
 FILLCELL_X2 FILLER_2_537 ();
 FILLCELL_X4 FILLER_2_543 ();
 FILLCELL_X4 FILLER_2_551 ();
 FILLCELL_X8 FILLER_2_561 ();
 FILLCELL_X1 FILLER_2_569 ();
 FILLCELL_X4 FILLER_2_574 ();
 FILLCELL_X8 FILLER_2_589 ();
 FILLCELL_X4 FILLER_2_597 ();
 FILLCELL_X1 FILLER_2_601 ();
 FILLCELL_X8 FILLER_2_620 ();
 FILLCELL_X2 FILLER_2_628 ();
 FILLCELL_X1 FILLER_2_630 ();
 FILLCELL_X4 FILLER_2_632 ();
 FILLCELL_X4 FILLER_2_645 ();
 FILLCELL_X1 FILLER_2_649 ();
 FILLCELL_X4 FILLER_2_655 ();
 FILLCELL_X4 FILLER_2_662 ();
 FILLCELL_X4 FILLER_2_669 ();
 FILLCELL_X2 FILLER_2_673 ();
 FILLCELL_X4 FILLER_2_684 ();
 FILLCELL_X4 FILLER_2_695 ();
 FILLCELL_X32 FILLER_2_703 ();
 FILLCELL_X8 FILLER_2_735 ();
 FILLCELL_X4 FILLER_2_747 ();
 FILLCELL_X8 FILLER_2_755 ();
 FILLCELL_X2 FILLER_2_763 ();
 FILLCELL_X4 FILLER_2_775 ();
 FILLCELL_X4 FILLER_2_782 ();
 FILLCELL_X16 FILLER_2_788 ();
 FILLCELL_X4 FILLER_2_804 ();
 FILLCELL_X2 FILLER_2_808 ();
 FILLCELL_X8 FILLER_2_814 ();
 FILLCELL_X16 FILLER_2_826 ();
 FILLCELL_X4 FILLER_2_842 ();
 FILLCELL_X2 FILLER_2_846 ();
 FILLCELL_X1 FILLER_2_848 ();
 FILLCELL_X4 FILLER_2_853 ();
 FILLCELL_X2 FILLER_2_857 ();
 FILLCELL_X16 FILLER_2_863 ();
 FILLCELL_X2 FILLER_2_879 ();
 FILLCELL_X1 FILLER_2_881 ();
 FILLCELL_X8 FILLER_2_886 ();
 FILLCELL_X4 FILLER_2_899 ();
 FILLCELL_X4 FILLER_2_912 ();
 FILLCELL_X4 FILLER_2_920 ();
 FILLCELL_X4 FILLER_2_928 ();
 FILLCELL_X4 FILLER_2_936 ();
 FILLCELL_X4 FILLER_2_943 ();
 FILLCELL_X4 FILLER_2_951 ();
 FILLCELL_X4 FILLER_2_962 ();
 FILLCELL_X16 FILLER_2_979 ();
 FILLCELL_X2 FILLER_2_995 ();
 FILLCELL_X4 FILLER_2_1002 ();
 FILLCELL_X4 FILLER_2_1009 ();
 FILLCELL_X1 FILLER_2_1013 ();
 FILLCELL_X16 FILLER_2_1021 ();
 FILLCELL_X1 FILLER_2_1037 ();
 FILLCELL_X4 FILLER_2_1041 ();
 FILLCELL_X2 FILLER_2_1045 ();
 FILLCELL_X8 FILLER_2_1052 ();
 FILLCELL_X1 FILLER_2_1060 ();
 FILLCELL_X4 FILLER_2_1065 ();
 FILLCELL_X4 FILLER_2_1082 ();
 FILLCELL_X4 FILLER_2_1089 ();
 FILLCELL_X2 FILLER_2_1093 ();
 FILLCELL_X1 FILLER_2_1095 ();
 FILLCELL_X4 FILLER_2_1103 ();
 FILLCELL_X8 FILLER_2_1112 ();
 FILLCELL_X1 FILLER_2_1120 ();
 FILLCELL_X4 FILLER_2_1128 ();
 FILLCELL_X4 FILLER_2_1136 ();
 FILLCELL_X16 FILLER_2_1143 ();
 FILLCELL_X2 FILLER_2_1159 ();
 FILLCELL_X1 FILLER_2_1161 ();
 FILLCELL_X4 FILLER_2_1165 ();
 FILLCELL_X2 FILLER_2_1169 ();
 FILLCELL_X4 FILLER_2_1176 ();
 FILLCELL_X2 FILLER_2_1180 ();
 FILLCELL_X8 FILLER_2_1189 ();
 FILLCELL_X4 FILLER_2_1197 ();
 FILLCELL_X2 FILLER_2_1201 ();
 FILLCELL_X1 FILLER_2_1203 ();
 FILLCELL_X4 FILLER_2_1211 ();
 FILLCELL_X2 FILLER_2_1215 ();
 FILLCELL_X32 FILLER_2_1224 ();
 FILLCELL_X32 FILLER_2_1256 ();
 FILLCELL_X32 FILLER_2_1288 ();
 FILLCELL_X8 FILLER_2_1320 ();
 FILLCELL_X4 FILLER_2_1328 ();
 FILLCELL_X8 FILLER_2_1336 ();
 FILLCELL_X32 FILLER_2_1363 ();
 FILLCELL_X32 FILLER_2_1395 ();
 FILLCELL_X32 FILLER_2_1427 ();
 FILLCELL_X32 FILLER_2_1459 ();
 FILLCELL_X32 FILLER_2_1491 ();
 FILLCELL_X32 FILLER_2_1523 ();
 FILLCELL_X32 FILLER_2_1555 ();
 FILLCELL_X32 FILLER_2_1587 ();
 FILLCELL_X32 FILLER_2_1619 ();
 FILLCELL_X32 FILLER_2_1651 ();
 FILLCELL_X16 FILLER_2_1683 ();
 FILLCELL_X2 FILLER_2_1699 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X32 FILLER_3_289 ();
 FILLCELL_X32 FILLER_3_321 ();
 FILLCELL_X32 FILLER_3_353 ();
 FILLCELL_X16 FILLER_3_385 ();
 FILLCELL_X4 FILLER_3_401 ();
 FILLCELL_X1 FILLER_3_405 ();
 FILLCELL_X8 FILLER_3_411 ();
 FILLCELL_X1 FILLER_3_419 ();
 FILLCELL_X16 FILLER_3_437 ();
 FILLCELL_X8 FILLER_3_453 ();
 FILLCELL_X4 FILLER_3_461 ();
 FILLCELL_X1 FILLER_3_465 ();
 FILLCELL_X4 FILLER_3_469 ();
 FILLCELL_X4 FILLER_3_482 ();
 FILLCELL_X4 FILLER_3_490 ();
 FILLCELL_X8 FILLER_3_496 ();
 FILLCELL_X4 FILLER_3_504 ();
 FILLCELL_X4 FILLER_3_510 ();
 FILLCELL_X2 FILLER_3_514 ();
 FILLCELL_X4 FILLER_3_520 ();
 FILLCELL_X2 FILLER_3_524 ();
 FILLCELL_X4 FILLER_3_535 ();
 FILLCELL_X8 FILLER_3_545 ();
 FILLCELL_X2 FILLER_3_553 ();
 FILLCELL_X4 FILLER_3_559 ();
 FILLCELL_X4 FILLER_3_568 ();
 FILLCELL_X2 FILLER_3_572 ();
 FILLCELL_X1 FILLER_3_574 ();
 FILLCELL_X4 FILLER_3_578 ();
 FILLCELL_X4 FILLER_3_591 ();
 FILLCELL_X4 FILLER_3_602 ();
 FILLCELL_X2 FILLER_3_606 ();
 FILLCELL_X1 FILLER_3_608 ();
 FILLCELL_X8 FILLER_3_627 ();
 FILLCELL_X8 FILLER_3_648 ();
 FILLCELL_X2 FILLER_3_656 ();
 FILLCELL_X4 FILLER_3_663 ();
 FILLCELL_X8 FILLER_3_670 ();
 FILLCELL_X16 FILLER_3_680 ();
 FILLCELL_X4 FILLER_3_696 ();
 FILLCELL_X8 FILLER_3_707 ();
 FILLCELL_X1 FILLER_3_715 ();
 FILLCELL_X4 FILLER_3_719 ();
 FILLCELL_X16 FILLER_3_726 ();
 FILLCELL_X4 FILLER_3_742 ();
 FILLCELL_X1 FILLER_3_746 ();
 FILLCELL_X8 FILLER_3_752 ();
 FILLCELL_X4 FILLER_3_760 ();
 FILLCELL_X1 FILLER_3_764 ();
 FILLCELL_X4 FILLER_3_768 ();
 FILLCELL_X4 FILLER_3_775 ();
 FILLCELL_X4 FILLER_3_782 ();
 FILLCELL_X4 FILLER_3_796 ();
 FILLCELL_X2 FILLER_3_800 ();
 FILLCELL_X4 FILLER_3_809 ();
 FILLCELL_X4 FILLER_3_822 ();
 FILLCELL_X4 FILLER_3_833 ();
 FILLCELL_X8 FILLER_3_843 ();
 FILLCELL_X4 FILLER_3_855 ();
 FILLCELL_X4 FILLER_3_862 ();
 FILLCELL_X1 FILLER_3_866 ();
 FILLCELL_X8 FILLER_3_869 ();
 FILLCELL_X4 FILLER_3_877 ();
 FILLCELL_X4 FILLER_3_884 ();
 FILLCELL_X4 FILLER_3_897 ();
 FILLCELL_X8 FILLER_3_905 ();
 FILLCELL_X2 FILLER_3_913 ();
 FILLCELL_X1 FILLER_3_915 ();
 FILLCELL_X4 FILLER_3_925 ();
 FILLCELL_X2 FILLER_3_929 ();
 FILLCELL_X1 FILLER_3_931 ();
 FILLCELL_X4 FILLER_3_939 ();
 FILLCELL_X8 FILLER_3_947 ();
 FILLCELL_X1 FILLER_3_955 ();
 FILLCELL_X4 FILLER_3_960 ();
 FILLCELL_X2 FILLER_3_964 ();
 FILLCELL_X4 FILLER_3_975 ();
 FILLCELL_X2 FILLER_3_979 ();
 FILLCELL_X1 FILLER_3_981 ();
 FILLCELL_X4 FILLER_3_995 ();
 FILLCELL_X1 FILLER_3_999 ();
 FILLCELL_X4 FILLER_3_1013 ();
 FILLCELL_X2 FILLER_3_1017 ();
 FILLCELL_X4 FILLER_3_1028 ();
 FILLCELL_X2 FILLER_3_1032 ();
 FILLCELL_X8 FILLER_3_1052 ();
 FILLCELL_X4 FILLER_3_1060 ();
 FILLCELL_X1 FILLER_3_1064 ();
 FILLCELL_X32 FILLER_3_1069 ();
 FILLCELL_X1 FILLER_3_1101 ();
 FILLCELL_X4 FILLER_3_1111 ();
 FILLCELL_X4 FILLER_3_1118 ();
 FILLCELL_X8 FILLER_3_1125 ();
 FILLCELL_X2 FILLER_3_1133 ();
 FILLCELL_X1 FILLER_3_1135 ();
 FILLCELL_X4 FILLER_3_1139 ();
 FILLCELL_X2 FILLER_3_1143 ();
 FILLCELL_X1 FILLER_3_1145 ();
 FILLCELL_X8 FILLER_3_1150 ();
 FILLCELL_X2 FILLER_3_1158 ();
 FILLCELL_X1 FILLER_3_1160 ();
 FILLCELL_X4 FILLER_3_1164 ();
 FILLCELL_X2 FILLER_3_1168 ();
 FILLCELL_X4 FILLER_3_1177 ();
 FILLCELL_X4 FILLER_3_1188 ();
 FILLCELL_X4 FILLER_3_1199 ();
 FILLCELL_X2 FILLER_3_1203 ();
 FILLCELL_X4 FILLER_3_1212 ();
 FILLCELL_X4 FILLER_3_1223 ();
 FILLCELL_X2 FILLER_3_1227 ();
 FILLCELL_X8 FILLER_3_1238 ();
 FILLCELL_X2 FILLER_3_1246 ();
 FILLCELL_X1 FILLER_3_1248 ();
 FILLCELL_X8 FILLER_3_1253 ();
 FILLCELL_X2 FILLER_3_1261 ();
 FILLCELL_X4 FILLER_3_1264 ();
 FILLCELL_X32 FILLER_3_1272 ();
 FILLCELL_X32 FILLER_3_1304 ();
 FILLCELL_X32 FILLER_3_1336 ();
 FILLCELL_X32 FILLER_3_1368 ();
 FILLCELL_X32 FILLER_3_1400 ();
 FILLCELL_X32 FILLER_3_1432 ();
 FILLCELL_X32 FILLER_3_1464 ();
 FILLCELL_X32 FILLER_3_1496 ();
 FILLCELL_X32 FILLER_3_1528 ();
 FILLCELL_X32 FILLER_3_1560 ();
 FILLCELL_X32 FILLER_3_1592 ();
 FILLCELL_X32 FILLER_3_1624 ();
 FILLCELL_X32 FILLER_3_1656 ();
 FILLCELL_X8 FILLER_3_1688 ();
 FILLCELL_X4 FILLER_3_1696 ();
 FILLCELL_X1 FILLER_3_1700 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X32 FILLER_4_289 ();
 FILLCELL_X32 FILLER_4_321 ();
 FILLCELL_X2 FILLER_4_353 ();
 FILLCELL_X8 FILLER_4_374 ();
 FILLCELL_X4 FILLER_4_382 ();
 FILLCELL_X1 FILLER_4_386 ();
 FILLCELL_X4 FILLER_4_391 ();
 FILLCELL_X4 FILLER_4_399 ();
 FILLCELL_X4 FILLER_4_407 ();
 FILLCELL_X8 FILLER_4_414 ();
 FILLCELL_X1 FILLER_4_422 ();
 FILLCELL_X4 FILLER_4_425 ();
 FILLCELL_X8 FILLER_4_431 ();
 FILLCELL_X1 FILLER_4_439 ();
 FILLCELL_X4 FILLER_4_446 ();
 FILLCELL_X4 FILLER_4_453 ();
 FILLCELL_X4 FILLER_4_459 ();
 FILLCELL_X4 FILLER_4_468 ();
 FILLCELL_X1 FILLER_4_472 ();
 FILLCELL_X4 FILLER_4_477 ();
 FILLCELL_X2 FILLER_4_481 ();
 FILLCELL_X1 FILLER_4_483 ();
 FILLCELL_X4 FILLER_4_488 ();
 FILLCELL_X1 FILLER_4_492 ();
 FILLCELL_X4 FILLER_4_497 ();
 FILLCELL_X4 FILLER_4_505 ();
 FILLCELL_X2 FILLER_4_509 ();
 FILLCELL_X1 FILLER_4_511 ();
 FILLCELL_X8 FILLER_4_515 ();
 FILLCELL_X4 FILLER_4_523 ();
 FILLCELL_X2 FILLER_4_527 ();
 FILLCELL_X4 FILLER_4_532 ();
 FILLCELL_X4 FILLER_4_539 ();
 FILLCELL_X4 FILLER_4_550 ();
 FILLCELL_X4 FILLER_4_560 ();
 FILLCELL_X2 FILLER_4_564 ();
 FILLCELL_X8 FILLER_4_570 ();
 FILLCELL_X4 FILLER_4_578 ();
 FILLCELL_X1 FILLER_4_582 ();
 FILLCELL_X4 FILLER_4_586 ();
 FILLCELL_X4 FILLER_4_599 ();
 FILLCELL_X1 FILLER_4_603 ();
 FILLCELL_X4 FILLER_4_607 ();
 FILLCELL_X4 FILLER_4_614 ();
 FILLCELL_X4 FILLER_4_627 ();
 FILLCELL_X4 FILLER_4_632 ();
 FILLCELL_X4 FILLER_4_643 ();
 FILLCELL_X4 FILLER_4_651 ();
 FILLCELL_X2 FILLER_4_655 ();
 FILLCELL_X1 FILLER_4_657 ();
 FILLCELL_X4 FILLER_4_663 ();
 FILLCELL_X4 FILLER_4_671 ();
 FILLCELL_X4 FILLER_4_678 ();
 FILLCELL_X1 FILLER_4_682 ();
 FILLCELL_X4 FILLER_4_692 ();
 FILLCELL_X8 FILLER_4_699 ();
 FILLCELL_X1 FILLER_4_707 ();
 FILLCELL_X8 FILLER_4_711 ();
 FILLCELL_X4 FILLER_4_723 ();
 FILLCELL_X4 FILLER_4_731 ();
 FILLCELL_X4 FILLER_4_737 ();
 FILLCELL_X4 FILLER_4_758 ();
 FILLCELL_X16 FILLER_4_769 ();
 FILLCELL_X1 FILLER_4_785 ();
 FILLCELL_X4 FILLER_4_788 ();
 FILLCELL_X4 FILLER_4_802 ();
 FILLCELL_X2 FILLER_4_806 ();
 FILLCELL_X8 FILLER_4_812 ();
 FILLCELL_X4 FILLER_4_820 ();
 FILLCELL_X4 FILLER_4_827 ();
 FILLCELL_X4 FILLER_4_834 ();
 FILLCELL_X4 FILLER_4_842 ();
 FILLCELL_X8 FILLER_4_855 ();
 FILLCELL_X2 FILLER_4_863 ();
 FILLCELL_X4 FILLER_4_878 ();
 FILLCELL_X1 FILLER_4_882 ();
 FILLCELL_X4 FILLER_4_886 ();
 FILLCELL_X4 FILLER_4_899 ();
 FILLCELL_X2 FILLER_4_903 ();
 FILLCELL_X16 FILLER_4_909 ();
 FILLCELL_X4 FILLER_4_925 ();
 FILLCELL_X1 FILLER_4_929 ();
 FILLCELL_X4 FILLER_4_943 ();
 FILLCELL_X8 FILLER_4_954 ();
 FILLCELL_X8 FILLER_4_969 ();
 FILLCELL_X8 FILLER_4_990 ();
 FILLCELL_X4 FILLER_4_998 ();
 FILLCELL_X1 FILLER_4_1002 ();
 FILLCELL_X4 FILLER_4_1008 ();
 FILLCELL_X2 FILLER_4_1012 ();
 FILLCELL_X1 FILLER_4_1014 ();
 FILLCELL_X16 FILLER_4_1022 ();
 FILLCELL_X4 FILLER_4_1038 ();
 FILLCELL_X2 FILLER_4_1042 ();
 FILLCELL_X4 FILLER_4_1053 ();
 FILLCELL_X8 FILLER_4_1064 ();
 FILLCELL_X2 FILLER_4_1072 ();
 FILLCELL_X4 FILLER_4_1081 ();
 FILLCELL_X1 FILLER_4_1085 ();
 FILLCELL_X4 FILLER_4_1093 ();
 FILLCELL_X1 FILLER_4_1097 ();
 FILLCELL_X8 FILLER_4_1111 ();
 FILLCELL_X2 FILLER_4_1119 ();
 FILLCELL_X4 FILLER_4_1128 ();
 FILLCELL_X2 FILLER_4_1132 ();
 FILLCELL_X1 FILLER_4_1134 ();
 FILLCELL_X8 FILLER_4_1139 ();
 FILLCELL_X1 FILLER_4_1147 ();
 FILLCELL_X4 FILLER_4_1155 ();
 FILLCELL_X4 FILLER_4_1163 ();
 FILLCELL_X4 FILLER_4_1170 ();
 FILLCELL_X8 FILLER_4_1181 ();
 FILLCELL_X4 FILLER_4_1189 ();
 FILLCELL_X2 FILLER_4_1193 ();
 FILLCELL_X4 FILLER_4_1198 ();
 FILLCELL_X32 FILLER_4_1205 ();
 FILLCELL_X4 FILLER_4_1244 ();
 FILLCELL_X4 FILLER_4_1267 ();
 FILLCELL_X4 FILLER_4_1290 ();
 FILLCELL_X2 FILLER_4_1294 ();
 FILLCELL_X4 FILLER_4_1300 ();
 FILLCELL_X4 FILLER_4_1307 ();
 FILLCELL_X4 FILLER_4_1313 ();
 FILLCELL_X32 FILLER_4_1319 ();
 FILLCELL_X32 FILLER_4_1351 ();
 FILLCELL_X32 FILLER_4_1383 ();
 FILLCELL_X32 FILLER_4_1415 ();
 FILLCELL_X32 FILLER_4_1447 ();
 FILLCELL_X32 FILLER_4_1479 ();
 FILLCELL_X32 FILLER_4_1511 ();
 FILLCELL_X32 FILLER_4_1543 ();
 FILLCELL_X32 FILLER_4_1575 ();
 FILLCELL_X32 FILLER_4_1607 ();
 FILLCELL_X32 FILLER_4_1639 ();
 FILLCELL_X16 FILLER_4_1671 ();
 FILLCELL_X8 FILLER_4_1687 ();
 FILLCELL_X4 FILLER_4_1695 ();
 FILLCELL_X2 FILLER_4_1699 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X32 FILLER_5_257 ();
 FILLCELL_X32 FILLER_5_289 ();
 FILLCELL_X32 FILLER_5_321 ();
 FILLCELL_X16 FILLER_5_353 ();
 FILLCELL_X4 FILLER_5_369 ();
 FILLCELL_X1 FILLER_5_373 ();
 FILLCELL_X4 FILLER_5_377 ();
 FILLCELL_X2 FILLER_5_381 ();
 FILLCELL_X4 FILLER_5_385 ();
 FILLCELL_X8 FILLER_5_392 ();
 FILLCELL_X1 FILLER_5_400 ();
 FILLCELL_X4 FILLER_5_410 ();
 FILLCELL_X4 FILLER_5_418 ();
 FILLCELL_X2 FILLER_5_422 ();
 FILLCELL_X4 FILLER_5_428 ();
 FILLCELL_X16 FILLER_5_434 ();
 FILLCELL_X2 FILLER_5_450 ();
 FILLCELL_X4 FILLER_5_456 ();
 FILLCELL_X2 FILLER_5_460 ();
 FILLCELL_X8 FILLER_5_465 ();
 FILLCELL_X2 FILLER_5_473 ();
 FILLCELL_X4 FILLER_5_479 ();
 FILLCELL_X1 FILLER_5_483 ();
 FILLCELL_X4 FILLER_5_491 ();
 FILLCELL_X1 FILLER_5_495 ();
 FILLCELL_X4 FILLER_5_503 ();
 FILLCELL_X4 FILLER_5_513 ();
 FILLCELL_X8 FILLER_5_519 ();
 FILLCELL_X2 FILLER_5_527 ();
 FILLCELL_X8 FILLER_5_543 ();
 FILLCELL_X8 FILLER_5_553 ();
 FILLCELL_X2 FILLER_5_561 ();
 FILLCELL_X1 FILLER_5_563 ();
 FILLCELL_X16 FILLER_5_567 ();
 FILLCELL_X8 FILLER_5_583 ();
 FILLCELL_X4 FILLER_5_591 ();
 FILLCELL_X2 FILLER_5_595 ();
 FILLCELL_X1 FILLER_5_597 ();
 FILLCELL_X4 FILLER_5_602 ();
 FILLCELL_X4 FILLER_5_610 ();
 FILLCELL_X2 FILLER_5_614 ();
 FILLCELL_X1 FILLER_5_616 ();
 FILLCELL_X8 FILLER_5_635 ();
 FILLCELL_X16 FILLER_5_647 ();
 FILLCELL_X8 FILLER_5_663 ();
 FILLCELL_X4 FILLER_5_671 ();
 FILLCELL_X2 FILLER_5_675 ();
 FILLCELL_X4 FILLER_5_684 ();
 FILLCELL_X2 FILLER_5_688 ();
 FILLCELL_X1 FILLER_5_690 ();
 FILLCELL_X4 FILLER_5_695 ();
 FILLCELL_X4 FILLER_5_703 ();
 FILLCELL_X4 FILLER_5_709 ();
 FILLCELL_X8 FILLER_5_722 ();
 FILLCELL_X2 FILLER_5_730 ();
 FILLCELL_X4 FILLER_5_737 ();
 FILLCELL_X4 FILLER_5_750 ();
 FILLCELL_X4 FILLER_5_757 ();
 FILLCELL_X1 FILLER_5_761 ();
 FILLCELL_X4 FILLER_5_776 ();
 FILLCELL_X4 FILLER_5_790 ();
 FILLCELL_X2 FILLER_5_794 ();
 FILLCELL_X8 FILLER_5_800 ();
 FILLCELL_X4 FILLER_5_812 ();
 FILLCELL_X1 FILLER_5_816 ();
 FILLCELL_X8 FILLER_5_820 ();
 FILLCELL_X4 FILLER_5_828 ();
 FILLCELL_X2 FILLER_5_832 ();
 FILLCELL_X1 FILLER_5_834 ();
 FILLCELL_X4 FILLER_5_842 ();
 FILLCELL_X2 FILLER_5_846 ();
 FILLCELL_X4 FILLER_5_851 ();
 FILLCELL_X2 FILLER_5_855 ();
 FILLCELL_X1 FILLER_5_857 ();
 FILLCELL_X4 FILLER_5_868 ();
 FILLCELL_X8 FILLER_5_879 ();
 FILLCELL_X1 FILLER_5_887 ();
 FILLCELL_X16 FILLER_5_895 ();
 FILLCELL_X2 FILLER_5_911 ();
 FILLCELL_X16 FILLER_5_923 ();
 FILLCELL_X8 FILLER_5_939 ();
 FILLCELL_X4 FILLER_5_947 ();
 FILLCELL_X16 FILLER_5_954 ();
 FILLCELL_X4 FILLER_5_970 ();
 FILLCELL_X2 FILLER_5_974 ();
 FILLCELL_X1 FILLER_5_976 ();
 FILLCELL_X8 FILLER_5_984 ();
 FILLCELL_X4 FILLER_5_992 ();
 FILLCELL_X1 FILLER_5_996 ();
 FILLCELL_X4 FILLER_5_1002 ();
 FILLCELL_X16 FILLER_5_1011 ();
 FILLCELL_X8 FILLER_5_1030 ();
 FILLCELL_X4 FILLER_5_1038 ();
 FILLCELL_X1 FILLER_5_1042 ();
 FILLCELL_X4 FILLER_5_1047 ();
 FILLCELL_X4 FILLER_5_1064 ();
 FILLCELL_X2 FILLER_5_1068 ();
 FILLCELL_X1 FILLER_5_1070 ();
 FILLCELL_X8 FILLER_5_1078 ();
 FILLCELL_X8 FILLER_5_1091 ();
 FILLCELL_X2 FILLER_5_1099 ();
 FILLCELL_X1 FILLER_5_1101 ();
 FILLCELL_X8 FILLER_5_1106 ();
 FILLCELL_X2 FILLER_5_1114 ();
 FILLCELL_X1 FILLER_5_1116 ();
 FILLCELL_X4 FILLER_5_1120 ();
 FILLCELL_X8 FILLER_5_1131 ();
 FILLCELL_X2 FILLER_5_1139 ();
 FILLCELL_X8 FILLER_5_1144 ();
 FILLCELL_X4 FILLER_5_1152 ();
 FILLCELL_X1 FILLER_5_1156 ();
 FILLCELL_X16 FILLER_5_1161 ();
 FILLCELL_X4 FILLER_5_1177 ();
 FILLCELL_X16 FILLER_5_1185 ();
 FILLCELL_X1 FILLER_5_1201 ();
 FILLCELL_X8 FILLER_5_1209 ();
 FILLCELL_X4 FILLER_5_1217 ();
 FILLCELL_X2 FILLER_5_1221 ();
 FILLCELL_X4 FILLER_5_1230 ();
 FILLCELL_X4 FILLER_5_1241 ();
 FILLCELL_X8 FILLER_5_1252 ();
 FILLCELL_X2 FILLER_5_1260 ();
 FILLCELL_X1 FILLER_5_1262 ();
 FILLCELL_X16 FILLER_5_1264 ();
 FILLCELL_X2 FILLER_5_1280 ();
 FILLCELL_X1 FILLER_5_1282 ();
 FILLCELL_X4 FILLER_5_1287 ();
 FILLCELL_X4 FILLER_5_1295 ();
 FILLCELL_X2 FILLER_5_1299 ();
 FILLCELL_X1 FILLER_5_1301 ();
 FILLCELL_X4 FILLER_5_1309 ();
 FILLCELL_X1 FILLER_5_1313 ();
 FILLCELL_X8 FILLER_5_1317 ();
 FILLCELL_X2 FILLER_5_1325 ();
 FILLCELL_X32 FILLER_5_1329 ();
 FILLCELL_X32 FILLER_5_1361 ();
 FILLCELL_X32 FILLER_5_1393 ();
 FILLCELL_X32 FILLER_5_1425 ();
 FILLCELL_X32 FILLER_5_1457 ();
 FILLCELL_X32 FILLER_5_1489 ();
 FILLCELL_X4 FILLER_5_1521 ();
 FILLCELL_X2 FILLER_5_1525 ();
 FILLCELL_X4 FILLER_5_1531 ();
 FILLCELL_X32 FILLER_5_1554 ();
 FILLCELL_X32 FILLER_5_1586 ();
 FILLCELL_X32 FILLER_5_1618 ();
 FILLCELL_X32 FILLER_5_1650 ();
 FILLCELL_X16 FILLER_5_1682 ();
 FILLCELL_X2 FILLER_5_1698 ();
 FILLCELL_X1 FILLER_5_1700 ();
 FILLCELL_X4 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_9 ();
 FILLCELL_X32 FILLER_6_41 ();
 FILLCELL_X32 FILLER_6_73 ();
 FILLCELL_X32 FILLER_6_105 ();
 FILLCELL_X32 FILLER_6_137 ();
 FILLCELL_X32 FILLER_6_169 ();
 FILLCELL_X32 FILLER_6_201 ();
 FILLCELL_X32 FILLER_6_233 ();
 FILLCELL_X32 FILLER_6_265 ();
 FILLCELL_X32 FILLER_6_297 ();
 FILLCELL_X16 FILLER_6_329 ();
 FILLCELL_X8 FILLER_6_345 ();
 FILLCELL_X4 FILLER_6_353 ();
 FILLCELL_X2 FILLER_6_357 ();
 FILLCELL_X1 FILLER_6_359 ();
 FILLCELL_X4 FILLER_6_364 ();
 FILLCELL_X4 FILLER_6_372 ();
 FILLCELL_X2 FILLER_6_376 ();
 FILLCELL_X1 FILLER_6_378 ();
 FILLCELL_X4 FILLER_6_396 ();
 FILLCELL_X4 FILLER_6_402 ();
 FILLCELL_X2 FILLER_6_406 ();
 FILLCELL_X4 FILLER_6_411 ();
 FILLCELL_X1 FILLER_6_415 ();
 FILLCELL_X4 FILLER_6_422 ();
 FILLCELL_X4 FILLER_6_436 ();
 FILLCELL_X1 FILLER_6_440 ();
 FILLCELL_X4 FILLER_6_450 ();
 FILLCELL_X2 FILLER_6_454 ();
 FILLCELL_X8 FILLER_6_460 ();
 FILLCELL_X1 FILLER_6_468 ();
 FILLCELL_X4 FILLER_6_473 ();
 FILLCELL_X2 FILLER_6_477 ();
 FILLCELL_X1 FILLER_6_479 ();
 FILLCELL_X16 FILLER_6_484 ();
 FILLCELL_X4 FILLER_6_500 ();
 FILLCELL_X2 FILLER_6_504 ();
 FILLCELL_X4 FILLER_6_511 ();
 FILLCELL_X16 FILLER_6_528 ();
 FILLCELL_X4 FILLER_6_544 ();
 FILLCELL_X1 FILLER_6_548 ();
 FILLCELL_X4 FILLER_6_553 ();
 FILLCELL_X4 FILLER_6_561 ();
 FILLCELL_X4 FILLER_6_574 ();
 FILLCELL_X8 FILLER_6_596 ();
 FILLCELL_X16 FILLER_6_608 ();
 FILLCELL_X4 FILLER_6_624 ();
 FILLCELL_X2 FILLER_6_628 ();
 FILLCELL_X1 FILLER_6_630 ();
 FILLCELL_X4 FILLER_6_632 ();
 FILLCELL_X4 FILLER_6_643 ();
 FILLCELL_X2 FILLER_6_647 ();
 FILLCELL_X8 FILLER_6_653 ();
 FILLCELL_X2 FILLER_6_661 ();
 FILLCELL_X1 FILLER_6_663 ();
 FILLCELL_X4 FILLER_6_671 ();
 FILLCELL_X4 FILLER_6_680 ();
 FILLCELL_X4 FILLER_6_688 ();
 FILLCELL_X2 FILLER_6_692 ();
 FILLCELL_X4 FILLER_6_697 ();
 FILLCELL_X4 FILLER_6_708 ();
 FILLCELL_X2 FILLER_6_712 ();
 FILLCELL_X1 FILLER_6_714 ();
 FILLCELL_X4 FILLER_6_722 ();
 FILLCELL_X4 FILLER_6_736 ();
 FILLCELL_X2 FILLER_6_740 ();
 FILLCELL_X32 FILLER_6_744 ();
 FILLCELL_X8 FILLER_6_783 ();
 FILLCELL_X1 FILLER_6_791 ();
 FILLCELL_X4 FILLER_6_799 ();
 FILLCELL_X4 FILLER_6_807 ();
 FILLCELL_X4 FILLER_6_815 ();
 FILLCELL_X1 FILLER_6_819 ();
 FILLCELL_X4 FILLER_6_824 ();
 FILLCELL_X8 FILLER_6_833 ();
 FILLCELL_X1 FILLER_6_841 ();
 FILLCELL_X4 FILLER_6_846 ();
 FILLCELL_X4 FILLER_6_854 ();
 FILLCELL_X8 FILLER_6_861 ();
 FILLCELL_X2 FILLER_6_869 ();
 FILLCELL_X4 FILLER_6_880 ();
 FILLCELL_X1 FILLER_6_884 ();
 FILLCELL_X4 FILLER_6_888 ();
 FILLCELL_X8 FILLER_6_902 ();
 FILLCELL_X4 FILLER_6_917 ();
 FILLCELL_X4 FILLER_6_925 ();
 FILLCELL_X4 FILLER_6_932 ();
 FILLCELL_X4 FILLER_6_943 ();
 FILLCELL_X4 FILLER_6_951 ();
 FILLCELL_X1 FILLER_6_955 ();
 FILLCELL_X4 FILLER_6_960 ();
 FILLCELL_X4 FILLER_6_968 ();
 FILLCELL_X4 FILLER_6_975 ();
 FILLCELL_X4 FILLER_6_982 ();
 FILLCELL_X4 FILLER_6_988 ();
 FILLCELL_X2 FILLER_6_992 ();
 FILLCELL_X4 FILLER_6_1001 ();
 FILLCELL_X1 FILLER_6_1005 ();
 FILLCELL_X4 FILLER_6_1015 ();
 FILLCELL_X4 FILLER_6_1032 ();
 FILLCELL_X8 FILLER_6_1040 ();
 FILLCELL_X2 FILLER_6_1048 ();
 FILLCELL_X8 FILLER_6_1053 ();
 FILLCELL_X4 FILLER_6_1064 ();
 FILLCELL_X2 FILLER_6_1068 ();
 FILLCELL_X4 FILLER_6_1074 ();
 FILLCELL_X4 FILLER_6_1081 ();
 FILLCELL_X2 FILLER_6_1085 ();
 FILLCELL_X1 FILLER_6_1087 ();
 FILLCELL_X8 FILLER_6_1095 ();
 FILLCELL_X4 FILLER_6_1103 ();
 FILLCELL_X2 FILLER_6_1107 ();
 FILLCELL_X1 FILLER_6_1109 ();
 FILLCELL_X4 FILLER_6_1119 ();
 FILLCELL_X2 FILLER_6_1123 ();
 FILLCELL_X1 FILLER_6_1125 ();
 FILLCELL_X4 FILLER_6_1130 ();
 FILLCELL_X1 FILLER_6_1134 ();
 FILLCELL_X4 FILLER_6_1142 ();
 FILLCELL_X8 FILLER_6_1153 ();
 FILLCELL_X2 FILLER_6_1161 ();
 FILLCELL_X4 FILLER_6_1170 ();
 FILLCELL_X4 FILLER_6_1181 ();
 FILLCELL_X2 FILLER_6_1185 ();
 FILLCELL_X4 FILLER_6_1194 ();
 FILLCELL_X4 FILLER_6_1205 ();
 FILLCELL_X4 FILLER_6_1216 ();
 FILLCELL_X4 FILLER_6_1227 ();
 FILLCELL_X4 FILLER_6_1238 ();
 FILLCELL_X4 FILLER_6_1249 ();
 FILLCELL_X2 FILLER_6_1253 ();
 FILLCELL_X1 FILLER_6_1255 ();
 FILLCELL_X8 FILLER_6_1265 ();
 FILLCELL_X4 FILLER_6_1273 ();
 FILLCELL_X1 FILLER_6_1277 ();
 FILLCELL_X4 FILLER_6_1282 ();
 FILLCELL_X4 FILLER_6_1290 ();
 FILLCELL_X4 FILLER_6_1297 ();
 FILLCELL_X8 FILLER_6_1305 ();
 FILLCELL_X1 FILLER_6_1313 ();
 FILLCELL_X4 FILLER_6_1321 ();
 FILLCELL_X4 FILLER_6_1327 ();
 FILLCELL_X32 FILLER_6_1333 ();
 FILLCELL_X32 FILLER_6_1365 ();
 FILLCELL_X32 FILLER_6_1397 ();
 FILLCELL_X32 FILLER_6_1429 ();
 FILLCELL_X32 FILLER_6_1461 ();
 FILLCELL_X32 FILLER_6_1493 ();
 FILLCELL_X32 FILLER_6_1525 ();
 FILLCELL_X32 FILLER_6_1557 ();
 FILLCELL_X32 FILLER_6_1589 ();
 FILLCELL_X32 FILLER_6_1621 ();
 FILLCELL_X32 FILLER_6_1653 ();
 FILLCELL_X16 FILLER_6_1685 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X32 FILLER_7_257 ();
 FILLCELL_X32 FILLER_7_289 ();
 FILLCELL_X16 FILLER_7_321 ();
 FILLCELL_X8 FILLER_7_337 ();
 FILLCELL_X4 FILLER_7_345 ();
 FILLCELL_X8 FILLER_7_366 ();
 FILLCELL_X1 FILLER_7_374 ();
 FILLCELL_X4 FILLER_7_379 ();
 FILLCELL_X4 FILLER_7_387 ();
 FILLCELL_X4 FILLER_7_393 ();
 FILLCELL_X4 FILLER_7_406 ();
 FILLCELL_X4 FILLER_7_413 ();
 FILLCELL_X16 FILLER_7_419 ();
 FILLCELL_X4 FILLER_7_442 ();
 FILLCELL_X4 FILLER_7_455 ();
 FILLCELL_X2 FILLER_7_459 ();
 FILLCELL_X4 FILLER_7_465 ();
 FILLCELL_X2 FILLER_7_469 ();
 FILLCELL_X4 FILLER_7_473 ();
 FILLCELL_X4 FILLER_7_486 ();
 FILLCELL_X4 FILLER_7_494 ();
 FILLCELL_X2 FILLER_7_498 ();
 FILLCELL_X8 FILLER_7_507 ();
 FILLCELL_X4 FILLER_7_515 ();
 FILLCELL_X4 FILLER_7_523 ();
 FILLCELL_X8 FILLER_7_531 ();
 FILLCELL_X1 FILLER_7_539 ();
 FILLCELL_X8 FILLER_7_545 ();
 FILLCELL_X4 FILLER_7_560 ();
 FILLCELL_X8 FILLER_7_573 ();
 FILLCELL_X4 FILLER_7_581 ();
 FILLCELL_X8 FILLER_7_590 ();
 FILLCELL_X8 FILLER_7_601 ();
 FILLCELL_X2 FILLER_7_609 ();
 FILLCELL_X8 FILLER_7_613 ();
 FILLCELL_X2 FILLER_7_621 ();
 FILLCELL_X4 FILLER_7_632 ();
 FILLCELL_X4 FILLER_7_640 ();
 FILLCELL_X8 FILLER_7_651 ();
 FILLCELL_X4 FILLER_7_659 ();
 FILLCELL_X2 FILLER_7_663 ();
 FILLCELL_X8 FILLER_7_674 ();
 FILLCELL_X1 FILLER_7_682 ();
 FILLCELL_X4 FILLER_7_693 ();
 FILLCELL_X4 FILLER_7_707 ();
 FILLCELL_X4 FILLER_7_718 ();
 FILLCELL_X1 FILLER_7_722 ();
 FILLCELL_X4 FILLER_7_730 ();
 FILLCELL_X8 FILLER_7_739 ();
 FILLCELL_X2 FILLER_7_747 ();
 FILLCELL_X8 FILLER_7_751 ();
 FILLCELL_X4 FILLER_7_759 ();
 FILLCELL_X1 FILLER_7_763 ();
 FILLCELL_X8 FILLER_7_768 ();
 FILLCELL_X1 FILLER_7_776 ();
 FILLCELL_X4 FILLER_7_787 ();
 FILLCELL_X2 FILLER_7_791 ();
 FILLCELL_X4 FILLER_7_802 ();
 FILLCELL_X8 FILLER_7_808 ();
 FILLCELL_X8 FILLER_7_826 ();
 FILLCELL_X4 FILLER_7_834 ();
 FILLCELL_X8 FILLER_7_847 ();
 FILLCELL_X2 FILLER_7_855 ();
 FILLCELL_X1 FILLER_7_857 ();
 FILLCELL_X4 FILLER_7_868 ();
 FILLCELL_X2 FILLER_7_872 ();
 FILLCELL_X1 FILLER_7_874 ();
 FILLCELL_X16 FILLER_7_884 ();
 FILLCELL_X2 FILLER_7_900 ();
 FILLCELL_X4 FILLER_7_909 ();
 FILLCELL_X4 FILLER_7_922 ();
 FILLCELL_X8 FILLER_7_930 ();
 FILLCELL_X2 FILLER_7_938 ();
 FILLCELL_X1 FILLER_7_940 ();
 FILLCELL_X8 FILLER_7_945 ();
 FILLCELL_X2 FILLER_7_953 ();
 FILLCELL_X1 FILLER_7_955 ();
 FILLCELL_X4 FILLER_7_960 ();
 FILLCELL_X8 FILLER_7_977 ();
 FILLCELL_X4 FILLER_7_989 ();
 FILLCELL_X2 FILLER_7_993 ();
 FILLCELL_X8 FILLER_7_1004 ();
 FILLCELL_X4 FILLER_7_1012 ();
 FILLCELL_X2 FILLER_7_1016 ();
 FILLCELL_X1 FILLER_7_1018 ();
 FILLCELL_X4 FILLER_7_1028 ();
 FILLCELL_X2 FILLER_7_1032 ();
 FILLCELL_X1 FILLER_7_1034 ();
 FILLCELL_X8 FILLER_7_1044 ();
 FILLCELL_X2 FILLER_7_1052 ();
 FILLCELL_X1 FILLER_7_1054 ();
 FILLCELL_X8 FILLER_7_1059 ();
 FILLCELL_X4 FILLER_7_1067 ();
 FILLCELL_X8 FILLER_7_1074 ();
 FILLCELL_X4 FILLER_7_1085 ();
 FILLCELL_X2 FILLER_7_1089 ();
 FILLCELL_X8 FILLER_7_1095 ();
 FILLCELL_X2 FILLER_7_1103 ();
 FILLCELL_X4 FILLER_7_1114 ();
 FILLCELL_X16 FILLER_7_1123 ();
 FILLCELL_X2 FILLER_7_1139 ();
 FILLCELL_X4 FILLER_7_1148 ();
 FILLCELL_X8 FILLER_7_1161 ();
 FILLCELL_X4 FILLER_7_1169 ();
 FILLCELL_X2 FILLER_7_1173 ();
 FILLCELL_X16 FILLER_7_1182 ();
 FILLCELL_X8 FILLER_7_1198 ();
 FILLCELL_X2 FILLER_7_1206 ();
 FILLCELL_X4 FILLER_7_1212 ();
 FILLCELL_X4 FILLER_7_1223 ();
 FILLCELL_X4 FILLER_7_1234 ();
 FILLCELL_X1 FILLER_7_1238 ();
 FILLCELL_X4 FILLER_7_1246 ();
 FILLCELL_X4 FILLER_7_1259 ();
 FILLCELL_X8 FILLER_7_1264 ();
 FILLCELL_X8 FILLER_7_1276 ();
 FILLCELL_X4 FILLER_7_1286 ();
 FILLCELL_X2 FILLER_7_1290 ();
 FILLCELL_X4 FILLER_7_1299 ();
 FILLCELL_X4 FILLER_7_1305 ();
 FILLCELL_X1 FILLER_7_1309 ();
 FILLCELL_X8 FILLER_7_1314 ();
 FILLCELL_X2 FILLER_7_1322 ();
 FILLCELL_X4 FILLER_7_1331 ();
 FILLCELL_X32 FILLER_7_1338 ();
 FILLCELL_X32 FILLER_7_1370 ();
 FILLCELL_X32 FILLER_7_1402 ();
 FILLCELL_X32 FILLER_7_1434 ();
 FILLCELL_X32 FILLER_7_1466 ();
 FILLCELL_X4 FILLER_7_1498 ();
 FILLCELL_X2 FILLER_7_1502 ();
 FILLCELL_X1 FILLER_7_1504 ();
 FILLCELL_X4 FILLER_7_1509 ();
 FILLCELL_X1 FILLER_7_1513 ();
 FILLCELL_X32 FILLER_7_1531 ();
 FILLCELL_X32 FILLER_7_1563 ();
 FILLCELL_X32 FILLER_7_1595 ();
 FILLCELL_X32 FILLER_7_1627 ();
 FILLCELL_X32 FILLER_7_1659 ();
 FILLCELL_X8 FILLER_7_1691 ();
 FILLCELL_X2 FILLER_7_1699 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X32 FILLER_8_225 ();
 FILLCELL_X32 FILLER_8_257 ();
 FILLCELL_X32 FILLER_8_289 ();
 FILLCELL_X32 FILLER_8_321 ();
 FILLCELL_X16 FILLER_8_353 ();
 FILLCELL_X4 FILLER_8_369 ();
 FILLCELL_X1 FILLER_8_373 ();
 FILLCELL_X8 FILLER_8_377 ();
 FILLCELL_X4 FILLER_8_388 ();
 FILLCELL_X4 FILLER_8_399 ();
 FILLCELL_X1 FILLER_8_403 ();
 FILLCELL_X4 FILLER_8_408 ();
 FILLCELL_X4 FILLER_8_416 ();
 FILLCELL_X16 FILLER_8_429 ();
 FILLCELL_X4 FILLER_8_454 ();
 FILLCELL_X2 FILLER_8_458 ();
 FILLCELL_X1 FILLER_8_460 ();
 FILLCELL_X4 FILLER_8_470 ();
 FILLCELL_X2 FILLER_8_474 ();
 FILLCELL_X4 FILLER_8_480 ();
 FILLCELL_X8 FILLER_8_487 ();
 FILLCELL_X4 FILLER_8_495 ();
 FILLCELL_X8 FILLER_8_509 ();
 FILLCELL_X8 FILLER_8_524 ();
 FILLCELL_X1 FILLER_8_532 ();
 FILLCELL_X4 FILLER_8_537 ();
 FILLCELL_X2 FILLER_8_541 ();
 FILLCELL_X1 FILLER_8_543 ();
 FILLCELL_X4 FILLER_8_548 ();
 FILLCELL_X4 FILLER_8_556 ();
 FILLCELL_X16 FILLER_8_564 ();
 FILLCELL_X4 FILLER_8_580 ();
 FILLCELL_X4 FILLER_8_588 ();
 FILLCELL_X4 FILLER_8_596 ();
 FILLCELL_X2 FILLER_8_600 ();
 FILLCELL_X4 FILLER_8_606 ();
 FILLCELL_X4 FILLER_8_617 ();
 FILLCELL_X4 FILLER_8_625 ();
 FILLCELL_X2 FILLER_8_629 ();
 FILLCELL_X4 FILLER_8_632 ();
 FILLCELL_X16 FILLER_8_638 ();
 FILLCELL_X2 FILLER_8_654 ();
 FILLCELL_X1 FILLER_8_656 ();
 FILLCELL_X4 FILLER_8_670 ();
 FILLCELL_X1 FILLER_8_674 ();
 FILLCELL_X4 FILLER_8_678 ();
 FILLCELL_X8 FILLER_8_695 ();
 FILLCELL_X4 FILLER_8_703 ();
 FILLCELL_X2 FILLER_8_707 ();
 FILLCELL_X4 FILLER_8_719 ();
 FILLCELL_X4 FILLER_8_726 ();
 FILLCELL_X1 FILLER_8_730 ();
 FILLCELL_X4 FILLER_8_736 ();
 FILLCELL_X4 FILLER_8_750 ();
 FILLCELL_X4 FILLER_8_771 ();
 FILLCELL_X8 FILLER_8_780 ();
 FILLCELL_X4 FILLER_8_788 ();
 FILLCELL_X2 FILLER_8_792 ();
 FILLCELL_X4 FILLER_8_801 ();
 FILLCELL_X4 FILLER_8_814 ();
 FILLCELL_X2 FILLER_8_818 ();
 FILLCELL_X1 FILLER_8_820 ();
 FILLCELL_X4 FILLER_8_828 ();
 FILLCELL_X1 FILLER_8_832 ();
 FILLCELL_X4 FILLER_8_836 ();
 FILLCELL_X8 FILLER_8_842 ();
 FILLCELL_X2 FILLER_8_850 ();
 FILLCELL_X4 FILLER_8_859 ();
 FILLCELL_X4 FILLER_8_865 ();
 FILLCELL_X2 FILLER_8_869 ();
 FILLCELL_X1 FILLER_8_871 ();
 FILLCELL_X4 FILLER_8_877 ();
 FILLCELL_X2 FILLER_8_881 ();
 FILLCELL_X4 FILLER_8_892 ();
 FILLCELL_X8 FILLER_8_899 ();
 FILLCELL_X4 FILLER_8_907 ();
 FILLCELL_X2 FILLER_8_911 ();
 FILLCELL_X1 FILLER_8_913 ();
 FILLCELL_X8 FILLER_8_927 ();
 FILLCELL_X4 FILLER_8_935 ();
 FILLCELL_X2 FILLER_8_939 ();
 FILLCELL_X4 FILLER_8_958 ();
 FILLCELL_X4 FILLER_8_964 ();
 FILLCELL_X1 FILLER_8_968 ();
 FILLCELL_X4 FILLER_8_976 ();
 FILLCELL_X4 FILLER_8_986 ();
 FILLCELL_X4 FILLER_8_995 ();
 FILLCELL_X4 FILLER_8_1003 ();
 FILLCELL_X8 FILLER_8_1011 ();
 FILLCELL_X1 FILLER_8_1019 ();
 FILLCELL_X4 FILLER_8_1027 ();
 FILLCELL_X4 FILLER_8_1034 ();
 FILLCELL_X4 FILLER_8_1047 ();
 FILLCELL_X2 FILLER_8_1051 ();
 FILLCELL_X4 FILLER_8_1060 ();
 FILLCELL_X1 FILLER_8_1064 ();
 FILLCELL_X4 FILLER_8_1072 ();
 FILLCELL_X4 FILLER_8_1089 ();
 FILLCELL_X2 FILLER_8_1093 ();
 FILLCELL_X1 FILLER_8_1095 ();
 FILLCELL_X4 FILLER_8_1100 ();
 FILLCELL_X4 FILLER_8_1111 ();
 FILLCELL_X8 FILLER_8_1122 ();
 FILLCELL_X1 FILLER_8_1130 ();
 FILLCELL_X4 FILLER_8_1138 ();
 FILLCELL_X8 FILLER_8_1149 ();
 FILLCELL_X4 FILLER_8_1157 ();
 FILLCELL_X2 FILLER_8_1161 ();
 FILLCELL_X1 FILLER_8_1163 ();
 FILLCELL_X16 FILLER_8_1171 ();
 FILLCELL_X4 FILLER_8_1194 ();
 FILLCELL_X4 FILLER_8_1205 ();
 FILLCELL_X4 FILLER_8_1216 ();
 FILLCELL_X8 FILLER_8_1227 ();
 FILLCELL_X4 FILLER_8_1235 ();
 FILLCELL_X2 FILLER_8_1239 ();
 FILLCELL_X4 FILLER_8_1250 ();
 FILLCELL_X8 FILLER_8_1263 ();
 FILLCELL_X1 FILLER_8_1271 ();
 FILLCELL_X4 FILLER_8_1276 ();
 FILLCELL_X4 FILLER_8_1282 ();
 FILLCELL_X1 FILLER_8_1286 ();
 FILLCELL_X4 FILLER_8_1290 ();
 FILLCELL_X4 FILLER_8_1296 ();
 FILLCELL_X8 FILLER_8_1302 ();
 FILLCELL_X4 FILLER_8_1310 ();
 FILLCELL_X2 FILLER_8_1314 ();
 FILLCELL_X4 FILLER_8_1320 ();
 FILLCELL_X2 FILLER_8_1324 ();
 FILLCELL_X1 FILLER_8_1326 ();
 FILLCELL_X4 FILLER_8_1331 ();
 FILLCELL_X4 FILLER_8_1337 ();
 FILLCELL_X4 FILLER_8_1343 ();
 FILLCELL_X32 FILLER_8_1349 ();
 FILLCELL_X32 FILLER_8_1381 ();
 FILLCELL_X32 FILLER_8_1413 ();
 FILLCELL_X32 FILLER_8_1445 ();
 FILLCELL_X4 FILLER_8_1481 ();
 FILLCELL_X2 FILLER_8_1485 ();
 FILLCELL_X1 FILLER_8_1487 ();
 FILLCELL_X16 FILLER_8_1507 ();
 FILLCELL_X8 FILLER_8_1523 ();
 FILLCELL_X2 FILLER_8_1531 ();
 FILLCELL_X1 FILLER_8_1533 ();
 FILLCELL_X32 FILLER_8_1553 ();
 FILLCELL_X32 FILLER_8_1585 ();
 FILLCELL_X32 FILLER_8_1617 ();
 FILLCELL_X32 FILLER_8_1649 ();
 FILLCELL_X16 FILLER_8_1681 ();
 FILLCELL_X4 FILLER_8_1697 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X32 FILLER_9_257 ();
 FILLCELL_X32 FILLER_9_289 ();
 FILLCELL_X32 FILLER_9_321 ();
 FILLCELL_X4 FILLER_9_353 ();
 FILLCELL_X2 FILLER_9_357 ();
 FILLCELL_X8 FILLER_9_363 ();
 FILLCELL_X2 FILLER_9_371 ();
 FILLCELL_X1 FILLER_9_373 ();
 FILLCELL_X8 FILLER_9_376 ();
 FILLCELL_X2 FILLER_9_384 ();
 FILLCELL_X4 FILLER_9_390 ();
 FILLCELL_X4 FILLER_9_398 ();
 FILLCELL_X4 FILLER_9_408 ();
 FILLCELL_X4 FILLER_9_416 ();
 FILLCELL_X8 FILLER_9_422 ();
 FILLCELL_X16 FILLER_9_434 ();
 FILLCELL_X4 FILLER_9_469 ();
 FILLCELL_X16 FILLER_9_477 ();
 FILLCELL_X4 FILLER_9_493 ();
 FILLCELL_X8 FILLER_9_500 ();
 FILLCELL_X2 FILLER_9_508 ();
 FILLCELL_X8 FILLER_9_514 ();
 FILLCELL_X2 FILLER_9_522 ();
 FILLCELL_X4 FILLER_9_531 ();
 FILLCELL_X2 FILLER_9_535 ();
 FILLCELL_X1 FILLER_9_537 ();
 FILLCELL_X4 FILLER_9_542 ();
 FILLCELL_X8 FILLER_9_553 ();
 FILLCELL_X2 FILLER_9_561 ();
 FILLCELL_X1 FILLER_9_563 ();
 FILLCELL_X4 FILLER_9_568 ();
 FILLCELL_X8 FILLER_9_576 ();
 FILLCELL_X2 FILLER_9_584 ();
 FILLCELL_X1 FILLER_9_586 ();
 FILLCELL_X8 FILLER_9_594 ();
 FILLCELL_X4 FILLER_9_602 ();
 FILLCELL_X1 FILLER_9_606 ();
 FILLCELL_X4 FILLER_9_610 ();
 FILLCELL_X4 FILLER_9_618 ();
 FILLCELL_X1 FILLER_9_622 ();
 FILLCELL_X8 FILLER_9_630 ();
 FILLCELL_X4 FILLER_9_645 ();
 FILLCELL_X4 FILLER_9_658 ();
 FILLCELL_X4 FILLER_9_669 ();
 FILLCELL_X4 FILLER_9_676 ();
 FILLCELL_X4 FILLER_9_683 ();
 FILLCELL_X8 FILLER_9_690 ();
 FILLCELL_X4 FILLER_9_698 ();
 FILLCELL_X16 FILLER_9_709 ();
 FILLCELL_X1 FILLER_9_725 ();
 FILLCELL_X4 FILLER_9_735 ();
 FILLCELL_X4 FILLER_9_746 ();
 FILLCELL_X4 FILLER_9_755 ();
 FILLCELL_X4 FILLER_9_763 ();
 FILLCELL_X4 FILLER_9_771 ();
 FILLCELL_X8 FILLER_9_778 ();
 FILLCELL_X2 FILLER_9_786 ();
 FILLCELL_X4 FILLER_9_791 ();
 FILLCELL_X4 FILLER_9_802 ();
 FILLCELL_X16 FILLER_9_809 ();
 FILLCELL_X2 FILLER_9_825 ();
 FILLCELL_X8 FILLER_9_833 ();
 FILLCELL_X4 FILLER_9_841 ();
 FILLCELL_X4 FILLER_9_848 ();
 FILLCELL_X16 FILLER_9_861 ();
 FILLCELL_X4 FILLER_9_886 ();
 FILLCELL_X4 FILLER_9_897 ();
 FILLCELL_X32 FILLER_9_910 ();
 FILLCELL_X2 FILLER_9_942 ();
 FILLCELL_X8 FILLER_9_957 ();
 FILLCELL_X16 FILLER_9_972 ();
 FILLCELL_X1 FILLER_9_988 ();
 FILLCELL_X4 FILLER_9_992 ();
 FILLCELL_X8 FILLER_9_1000 ();
 FILLCELL_X4 FILLER_9_1017 ();
 FILLCELL_X4 FILLER_9_1026 ();
 FILLCELL_X4 FILLER_9_1035 ();
 FILLCELL_X2 FILLER_9_1039 ();
 FILLCELL_X4 FILLER_9_1048 ();
 FILLCELL_X8 FILLER_9_1055 ();
 FILLCELL_X4 FILLER_9_1063 ();
 FILLCELL_X8 FILLER_9_1071 ();
 FILLCELL_X4 FILLER_9_1079 ();
 FILLCELL_X1 FILLER_9_1083 ();
 FILLCELL_X4 FILLER_9_1093 ();
 FILLCELL_X1 FILLER_9_1097 ();
 FILLCELL_X8 FILLER_9_1105 ();
 FILLCELL_X2 FILLER_9_1113 ();
 FILLCELL_X8 FILLER_9_1122 ();
 FILLCELL_X2 FILLER_9_1130 ();
 FILLCELL_X4 FILLER_9_1139 ();
 FILLCELL_X2 FILLER_9_1143 ();
 FILLCELL_X4 FILLER_9_1152 ();
 FILLCELL_X1 FILLER_9_1156 ();
 FILLCELL_X8 FILLER_9_1164 ();
 FILLCELL_X4 FILLER_9_1172 ();
 FILLCELL_X1 FILLER_9_1176 ();
 FILLCELL_X4 FILLER_9_1184 ();
 FILLCELL_X32 FILLER_9_1195 ();
 FILLCELL_X4 FILLER_9_1227 ();
 FILLCELL_X1 FILLER_9_1231 ();
 FILLCELL_X16 FILLER_9_1239 ();
 FILLCELL_X8 FILLER_9_1255 ();
 FILLCELL_X4 FILLER_9_1264 ();
 FILLCELL_X1 FILLER_9_1268 ();
 FILLCELL_X4 FILLER_9_1273 ();
 FILLCELL_X1 FILLER_9_1277 ();
 FILLCELL_X4 FILLER_9_1281 ();
 FILLCELL_X2 FILLER_9_1285 ();
 FILLCELL_X1 FILLER_9_1287 ();
 FILLCELL_X4 FILLER_9_1295 ();
 FILLCELL_X2 FILLER_9_1299 ();
 FILLCELL_X16 FILLER_9_1312 ();
 FILLCELL_X4 FILLER_9_1332 ();
 FILLCELL_X4 FILLER_9_1339 ();
 FILLCELL_X2 FILLER_9_1343 ();
 FILLCELL_X1 FILLER_9_1345 ();
 FILLCELL_X4 FILLER_9_1350 ();
 FILLCELL_X32 FILLER_9_1371 ();
 FILLCELL_X32 FILLER_9_1403 ();
 FILLCELL_X32 FILLER_9_1435 ();
 FILLCELL_X32 FILLER_9_1467 ();
 FILLCELL_X16 FILLER_9_1499 ();
 FILLCELL_X4 FILLER_9_1515 ();
 FILLCELL_X1 FILLER_9_1519 ();
 FILLCELL_X32 FILLER_9_1524 ();
 FILLCELL_X32 FILLER_9_1556 ();
 FILLCELL_X32 FILLER_9_1588 ();
 FILLCELL_X32 FILLER_9_1620 ();
 FILLCELL_X32 FILLER_9_1652 ();
 FILLCELL_X16 FILLER_9_1684 ();
 FILLCELL_X1 FILLER_9_1700 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X32 FILLER_10_257 ();
 FILLCELL_X32 FILLER_10_289 ();
 FILLCELL_X16 FILLER_10_321 ();
 FILLCELL_X8 FILLER_10_337 ();
 FILLCELL_X2 FILLER_10_345 ();
 FILLCELL_X16 FILLER_10_366 ();
 FILLCELL_X1 FILLER_10_382 ();
 FILLCELL_X8 FILLER_10_386 ();
 FILLCELL_X2 FILLER_10_394 ();
 FILLCELL_X1 FILLER_10_396 ();
 FILLCELL_X16 FILLER_10_401 ();
 FILLCELL_X8 FILLER_10_417 ();
 FILLCELL_X4 FILLER_10_435 ();
 FILLCELL_X1 FILLER_10_439 ();
 FILLCELL_X16 FILLER_10_444 ();
 FILLCELL_X4 FILLER_10_460 ();
 FILLCELL_X1 FILLER_10_464 ();
 FILLCELL_X4 FILLER_10_468 ();
 FILLCELL_X16 FILLER_10_476 ();
 FILLCELL_X2 FILLER_10_492 ();
 FILLCELL_X4 FILLER_10_503 ();
 FILLCELL_X4 FILLER_10_510 ();
 FILLCELL_X2 FILLER_10_514 ();
 FILLCELL_X4 FILLER_10_519 ();
 FILLCELL_X4 FILLER_10_526 ();
 FILLCELL_X8 FILLER_10_532 ();
 FILLCELL_X4 FILLER_10_540 ();
 FILLCELL_X1 FILLER_10_544 ();
 FILLCELL_X4 FILLER_10_554 ();
 FILLCELL_X1 FILLER_10_558 ();
 FILLCELL_X4 FILLER_10_568 ();
 FILLCELL_X4 FILLER_10_579 ();
 FILLCELL_X1 FILLER_10_583 ();
 FILLCELL_X4 FILLER_10_597 ();
 FILLCELL_X4 FILLER_10_608 ();
 FILLCELL_X2 FILLER_10_612 ();
 FILLCELL_X4 FILLER_10_616 ();
 FILLCELL_X4 FILLER_10_627 ();
 FILLCELL_X4 FILLER_10_632 ();
 FILLCELL_X2 FILLER_10_636 ();
 FILLCELL_X4 FILLER_10_656 ();
 FILLCELL_X1 FILLER_10_660 ();
 FILLCELL_X4 FILLER_10_667 ();
 FILLCELL_X16 FILLER_10_673 ();
 FILLCELL_X8 FILLER_10_689 ();
 FILLCELL_X4 FILLER_10_700 ();
 FILLCELL_X4 FILLER_10_713 ();
 FILLCELL_X2 FILLER_10_717 ();
 FILLCELL_X4 FILLER_10_725 ();
 FILLCELL_X8 FILLER_10_742 ();
 FILLCELL_X2 FILLER_10_750 ();
 FILLCELL_X1 FILLER_10_752 ();
 FILLCELL_X16 FILLER_10_755 ();
 FILLCELL_X4 FILLER_10_771 ();
 FILLCELL_X1 FILLER_10_775 ();
 FILLCELL_X4 FILLER_10_783 ();
 FILLCELL_X8 FILLER_10_792 ();
 FILLCELL_X2 FILLER_10_800 ();
 FILLCELL_X1 FILLER_10_802 ();
 FILLCELL_X4 FILLER_10_810 ();
 FILLCELL_X4 FILLER_10_821 ();
 FILLCELL_X2 FILLER_10_825 ();
 FILLCELL_X1 FILLER_10_827 ();
 FILLCELL_X8 FILLER_10_833 ();
 FILLCELL_X4 FILLER_10_841 ();
 FILLCELL_X1 FILLER_10_845 ();
 FILLCELL_X4 FILLER_10_853 ();
 FILLCELL_X4 FILLER_10_860 ();
 FILLCELL_X8 FILLER_10_867 ();
 FILLCELL_X2 FILLER_10_875 ();
 FILLCELL_X1 FILLER_10_877 ();
 FILLCELL_X8 FILLER_10_891 ();
 FILLCELL_X2 FILLER_10_899 ();
 FILLCELL_X1 FILLER_10_901 ();
 FILLCELL_X8 FILLER_10_912 ();
 FILLCELL_X2 FILLER_10_920 ();
 FILLCELL_X1 FILLER_10_922 ();
 FILLCELL_X4 FILLER_10_933 ();
 FILLCELL_X8 FILLER_10_944 ();
 FILLCELL_X4 FILLER_10_959 ();
 FILLCELL_X16 FILLER_10_967 ();
 FILLCELL_X2 FILLER_10_983 ();
 FILLCELL_X1 FILLER_10_985 ();
 FILLCELL_X4 FILLER_10_999 ();
 FILLCELL_X4 FILLER_10_1012 ();
 FILLCELL_X4 FILLER_10_1023 ();
 FILLCELL_X4 FILLER_10_1040 ();
 FILLCELL_X8 FILLER_10_1047 ();
 FILLCELL_X8 FILLER_10_1062 ();
 FILLCELL_X4 FILLER_10_1070 ();
 FILLCELL_X2 FILLER_10_1074 ();
 FILLCELL_X4 FILLER_10_1079 ();
 FILLCELL_X4 FILLER_10_1090 ();
 FILLCELL_X8 FILLER_10_1098 ();
 FILLCELL_X2 FILLER_10_1106 ();
 FILLCELL_X4 FILLER_10_1112 ();
 FILLCELL_X32 FILLER_10_1120 ();
 FILLCELL_X2 FILLER_10_1152 ();
 FILLCELL_X4 FILLER_10_1158 ();
 FILLCELL_X4 FILLER_10_1166 ();
 FILLCELL_X16 FILLER_10_1174 ();
 FILLCELL_X2 FILLER_10_1190 ();
 FILLCELL_X4 FILLER_10_1199 ();
 FILLCELL_X16 FILLER_10_1210 ();
 FILLCELL_X4 FILLER_10_1226 ();
 FILLCELL_X1 FILLER_10_1230 ();
 FILLCELL_X4 FILLER_10_1240 ();
 FILLCELL_X4 FILLER_10_1253 ();
 FILLCELL_X4 FILLER_10_1266 ();
 FILLCELL_X8 FILLER_10_1274 ();
 FILLCELL_X1 FILLER_10_1282 ();
 FILLCELL_X8 FILLER_10_1290 ();
 FILLCELL_X1 FILLER_10_1298 ();
 FILLCELL_X8 FILLER_10_1310 ();
 FILLCELL_X1 FILLER_10_1318 ();
 FILLCELL_X4 FILLER_10_1326 ();
 FILLCELL_X4 FILLER_10_1334 ();
 FILLCELL_X32 FILLER_10_1341 ();
 FILLCELL_X32 FILLER_10_1373 ();
 FILLCELL_X32 FILLER_10_1405 ();
 FILLCELL_X32 FILLER_10_1437 ();
 FILLCELL_X32 FILLER_10_1469 ();
 FILLCELL_X32 FILLER_10_1501 ();
 FILLCELL_X32 FILLER_10_1533 ();
 FILLCELL_X32 FILLER_10_1565 ();
 FILLCELL_X32 FILLER_10_1597 ();
 FILLCELL_X32 FILLER_10_1629 ();
 FILLCELL_X32 FILLER_10_1661 ();
 FILLCELL_X1 FILLER_10_1693 ();
 FILLCELL_X4 FILLER_10_1697 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_11_193 ();
 FILLCELL_X32 FILLER_11_225 ();
 FILLCELL_X32 FILLER_11_257 ();
 FILLCELL_X32 FILLER_11_289 ();
 FILLCELL_X32 FILLER_11_321 ();
 FILLCELL_X8 FILLER_11_353 ();
 FILLCELL_X4 FILLER_11_361 ();
 FILLCELL_X2 FILLER_11_365 ();
 FILLCELL_X4 FILLER_11_370 ();
 FILLCELL_X4 FILLER_11_379 ();
 FILLCELL_X32 FILLER_11_386 ();
 FILLCELL_X1 FILLER_11_418 ();
 FILLCELL_X4 FILLER_11_423 ();
 FILLCELL_X4 FILLER_11_434 ();
 FILLCELL_X16 FILLER_11_448 ();
 FILLCELL_X4 FILLER_11_464 ();
 FILLCELL_X1 FILLER_11_468 ();
 FILLCELL_X4 FILLER_11_479 ();
 FILLCELL_X4 FILLER_11_487 ();
 FILLCELL_X4 FILLER_11_494 ();
 FILLCELL_X4 FILLER_11_502 ();
 FILLCELL_X4 FILLER_11_515 ();
 FILLCELL_X2 FILLER_11_519 ();
 FILLCELL_X4 FILLER_11_524 ();
 FILLCELL_X1 FILLER_11_528 ();
 FILLCELL_X8 FILLER_11_532 ();
 FILLCELL_X2 FILLER_11_540 ();
 FILLCELL_X32 FILLER_11_555 ();
 FILLCELL_X8 FILLER_11_587 ();
 FILLCELL_X8 FILLER_11_598 ();
 FILLCELL_X4 FILLER_11_606 ();
 FILLCELL_X2 FILLER_11_610 ();
 FILLCELL_X1 FILLER_11_612 ();
 FILLCELL_X8 FILLER_11_618 ();
 FILLCELL_X4 FILLER_11_628 ();
 FILLCELL_X4 FILLER_11_636 ();
 FILLCELL_X1 FILLER_11_640 ();
 FILLCELL_X4 FILLER_11_644 ();
 FILLCELL_X4 FILLER_11_657 ();
 FILLCELL_X4 FILLER_11_668 ();
 FILLCELL_X2 FILLER_11_672 ();
 FILLCELL_X1 FILLER_11_674 ();
 FILLCELL_X4 FILLER_11_684 ();
 FILLCELL_X8 FILLER_11_691 ();
 FILLCELL_X2 FILLER_11_699 ();
 FILLCELL_X4 FILLER_11_708 ();
 FILLCELL_X32 FILLER_11_719 ();
 FILLCELL_X2 FILLER_11_751 ();
 FILLCELL_X16 FILLER_11_757 ();
 FILLCELL_X2 FILLER_11_773 ();
 FILLCELL_X1 FILLER_11_775 ();
 FILLCELL_X4 FILLER_11_779 ();
 FILLCELL_X4 FILLER_11_786 ();
 FILLCELL_X1 FILLER_11_790 ();
 FILLCELL_X4 FILLER_11_798 ();
 FILLCELL_X4 FILLER_11_805 ();
 FILLCELL_X4 FILLER_11_812 ();
 FILLCELL_X2 FILLER_11_816 ();
 FILLCELL_X1 FILLER_11_818 ();
 FILLCELL_X4 FILLER_11_822 ();
 FILLCELL_X4 FILLER_11_833 ();
 FILLCELL_X4 FILLER_11_840 ();
 FILLCELL_X2 FILLER_11_844 ();
 FILLCELL_X8 FILLER_11_853 ();
 FILLCELL_X1 FILLER_11_861 ();
 FILLCELL_X8 FILLER_11_869 ();
 FILLCELL_X4 FILLER_11_877 ();
 FILLCELL_X8 FILLER_11_888 ();
 FILLCELL_X2 FILLER_11_896 ();
 FILLCELL_X4 FILLER_11_907 ();
 FILLCELL_X4 FILLER_11_921 ();
 FILLCELL_X8 FILLER_11_934 ();
 FILLCELL_X2 FILLER_11_942 ();
 FILLCELL_X1 FILLER_11_944 ();
 FILLCELL_X4 FILLER_11_954 ();
 FILLCELL_X4 FILLER_11_968 ();
 FILLCELL_X4 FILLER_11_982 ();
 FILLCELL_X1 FILLER_11_986 ();
 FILLCELL_X4 FILLER_11_996 ();
 FILLCELL_X4 FILLER_11_1009 ();
 FILLCELL_X8 FILLER_11_1016 ();
 FILLCELL_X4 FILLER_11_1024 ();
 FILLCELL_X4 FILLER_11_1031 ();
 FILLCELL_X4 FILLER_11_1042 ();
 FILLCELL_X8 FILLER_11_1055 ();
 FILLCELL_X4 FILLER_11_1063 ();
 FILLCELL_X2 FILLER_11_1067 ();
 FILLCELL_X1 FILLER_11_1069 ();
 FILLCELL_X4 FILLER_11_1074 ();
 FILLCELL_X2 FILLER_11_1078 ();
 FILLCELL_X8 FILLER_11_1087 ();
 FILLCELL_X1 FILLER_11_1095 ();
 FILLCELL_X8 FILLER_11_1103 ();
 FILLCELL_X2 FILLER_11_1111 ();
 FILLCELL_X1 FILLER_11_1113 ();
 FILLCELL_X4 FILLER_11_1121 ();
 FILLCELL_X4 FILLER_11_1132 ();
 FILLCELL_X4 FILLER_11_1143 ();
 FILLCELL_X4 FILLER_11_1154 ();
 FILLCELL_X4 FILLER_11_1165 ();
 FILLCELL_X4 FILLER_11_1176 ();
 FILLCELL_X4 FILLER_11_1187 ();
 FILLCELL_X4 FILLER_11_1195 ();
 FILLCELL_X2 FILLER_11_1199 ();
 FILLCELL_X4 FILLER_11_1210 ();
 FILLCELL_X1 FILLER_11_1214 ();
 FILLCELL_X4 FILLER_11_1219 ();
 FILLCELL_X8 FILLER_11_1230 ();
 FILLCELL_X1 FILLER_11_1238 ();
 FILLCELL_X4 FILLER_11_1246 ();
 FILLCELL_X4 FILLER_11_1259 ();
 FILLCELL_X8 FILLER_11_1264 ();
 FILLCELL_X1 FILLER_11_1272 ();
 FILLCELL_X4 FILLER_11_1276 ();
 FILLCELL_X4 FILLER_11_1282 ();
 FILLCELL_X16 FILLER_11_1288 ();
 FILLCELL_X8 FILLER_11_1304 ();
 FILLCELL_X2 FILLER_11_1312 ();
 FILLCELL_X1 FILLER_11_1314 ();
 FILLCELL_X8 FILLER_11_1317 ();
 FILLCELL_X1 FILLER_11_1325 ();
 FILLCELL_X4 FILLER_11_1330 ();
 FILLCELL_X4 FILLER_11_1338 ();
 FILLCELL_X4 FILLER_11_1344 ();
 FILLCELL_X32 FILLER_11_1350 ();
 FILLCELL_X32 FILLER_11_1382 ();
 FILLCELL_X32 FILLER_11_1414 ();
 FILLCELL_X32 FILLER_11_1446 ();
 FILLCELL_X32 FILLER_11_1478 ();
 FILLCELL_X32 FILLER_11_1510 ();
 FILLCELL_X4 FILLER_11_1542 ();
 FILLCELL_X32 FILLER_11_1565 ();
 FILLCELL_X32 FILLER_11_1597 ();
 FILLCELL_X32 FILLER_11_1629 ();
 FILLCELL_X32 FILLER_11_1661 ();
 FILLCELL_X8 FILLER_11_1693 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X32 FILLER_12_225 ();
 FILLCELL_X32 FILLER_12_257 ();
 FILLCELL_X32 FILLER_12_289 ();
 FILLCELL_X32 FILLER_12_321 ();
 FILLCELL_X16 FILLER_12_353 ();
 FILLCELL_X2 FILLER_12_369 ();
 FILLCELL_X4 FILLER_12_374 ();
 FILLCELL_X4 FILLER_12_384 ();
 FILLCELL_X4 FILLER_12_392 ();
 FILLCELL_X4 FILLER_12_398 ();
 FILLCELL_X4 FILLER_12_407 ();
 FILLCELL_X8 FILLER_12_424 ();
 FILLCELL_X2 FILLER_12_432 ();
 FILLCELL_X8 FILLER_12_444 ();
 FILLCELL_X2 FILLER_12_452 ();
 FILLCELL_X1 FILLER_12_454 ();
 FILLCELL_X16 FILLER_12_458 ();
 FILLCELL_X8 FILLER_12_474 ();
 FILLCELL_X4 FILLER_12_482 ();
 FILLCELL_X2 FILLER_12_486 ();
 FILLCELL_X1 FILLER_12_488 ();
 FILLCELL_X4 FILLER_12_492 ();
 FILLCELL_X4 FILLER_12_499 ();
 FILLCELL_X8 FILLER_12_506 ();
 FILLCELL_X4 FILLER_12_517 ();
 FILLCELL_X8 FILLER_12_527 ();
 FILLCELL_X2 FILLER_12_535 ();
 FILLCELL_X16 FILLER_12_541 ();
 FILLCELL_X8 FILLER_12_557 ();
 FILLCELL_X1 FILLER_12_565 ();
 FILLCELL_X4 FILLER_12_569 ();
 FILLCELL_X4 FILLER_12_577 ();
 FILLCELL_X8 FILLER_12_588 ();
 FILLCELL_X4 FILLER_12_598 ();
 FILLCELL_X4 FILLER_12_611 ();
 FILLCELL_X2 FILLER_12_615 ();
 FILLCELL_X4 FILLER_12_626 ();
 FILLCELL_X1 FILLER_12_630 ();
 FILLCELL_X4 FILLER_12_632 ();
 FILLCELL_X16 FILLER_12_645 ();
 FILLCELL_X4 FILLER_12_661 ();
 FILLCELL_X2 FILLER_12_665 ();
 FILLCELL_X4 FILLER_12_671 ();
 FILLCELL_X4 FILLER_12_679 ();
 FILLCELL_X4 FILLER_12_692 ();
 FILLCELL_X4 FILLER_12_709 ();
 FILLCELL_X4 FILLER_12_727 ();
 FILLCELL_X4 FILLER_12_735 ();
 FILLCELL_X2 FILLER_12_739 ();
 FILLCELL_X1 FILLER_12_741 ();
 FILLCELL_X8 FILLER_12_749 ();
 FILLCELL_X4 FILLER_12_764 ();
 FILLCELL_X4 FILLER_12_775 ();
 FILLCELL_X1 FILLER_12_779 ();
 FILLCELL_X8 FILLER_12_785 ();
 FILLCELL_X2 FILLER_12_793 ();
 FILLCELL_X4 FILLER_12_799 ();
 FILLCELL_X2 FILLER_12_803 ();
 FILLCELL_X1 FILLER_12_805 ();
 FILLCELL_X4 FILLER_12_809 ();
 FILLCELL_X2 FILLER_12_813 ();
 FILLCELL_X8 FILLER_12_819 ();
 FILLCELL_X4 FILLER_12_827 ();
 FILLCELL_X2 FILLER_12_831 ();
 FILLCELL_X1 FILLER_12_833 ();
 FILLCELL_X4 FILLER_12_837 ();
 FILLCELL_X16 FILLER_12_854 ();
 FILLCELL_X4 FILLER_12_870 ();
 FILLCELL_X4 FILLER_12_881 ();
 FILLCELL_X4 FILLER_12_892 ();
 FILLCELL_X4 FILLER_12_900 ();
 FILLCELL_X2 FILLER_12_904 ();
 FILLCELL_X1 FILLER_12_906 ();
 FILLCELL_X4 FILLER_12_910 ();
 FILLCELL_X4 FILLER_12_921 ();
 FILLCELL_X4 FILLER_12_928 ();
 FILLCELL_X2 FILLER_12_932 ();
 FILLCELL_X1 FILLER_12_934 ();
 FILLCELL_X8 FILLER_12_942 ();
 FILLCELL_X2 FILLER_12_950 ();
 FILLCELL_X4 FILLER_12_955 ();
 FILLCELL_X2 FILLER_12_959 ();
 FILLCELL_X4 FILLER_12_964 ();
 FILLCELL_X32 FILLER_12_971 ();
 FILLCELL_X4 FILLER_12_1003 ();
 FILLCELL_X1 FILLER_12_1007 ();
 FILLCELL_X4 FILLER_12_1015 ();
 FILLCELL_X2 FILLER_12_1019 ();
 FILLCELL_X1 FILLER_12_1021 ();
 FILLCELL_X4 FILLER_12_1027 ();
 FILLCELL_X4 FILLER_12_1035 ();
 FILLCELL_X2 FILLER_12_1039 ();
 FILLCELL_X1 FILLER_12_1041 ();
 FILLCELL_X4 FILLER_12_1049 ();
 FILLCELL_X4 FILLER_12_1060 ();
 FILLCELL_X4 FILLER_12_1071 ();
 FILLCELL_X1 FILLER_12_1075 ();
 FILLCELL_X8 FILLER_12_1079 ();
 FILLCELL_X2 FILLER_12_1087 ();
 FILLCELL_X1 FILLER_12_1089 ();
 FILLCELL_X4 FILLER_12_1094 ();
 FILLCELL_X2 FILLER_12_1098 ();
 FILLCELL_X1 FILLER_12_1100 ();
 FILLCELL_X4 FILLER_12_1105 ();
 FILLCELL_X32 FILLER_12_1114 ();
 FILLCELL_X32 FILLER_12_1146 ();
 FILLCELL_X8 FILLER_12_1178 ();
 FILLCELL_X4 FILLER_12_1186 ();
 FILLCELL_X8 FILLER_12_1197 ();
 FILLCELL_X2 FILLER_12_1205 ();
 FILLCELL_X1 FILLER_12_1207 ();
 FILLCELL_X4 FILLER_12_1212 ();
 FILLCELL_X1 FILLER_12_1216 ();
 FILLCELL_X4 FILLER_12_1226 ();
 FILLCELL_X16 FILLER_12_1237 ();
 FILLCELL_X8 FILLER_12_1253 ();
 FILLCELL_X4 FILLER_12_1261 ();
 FILLCELL_X1 FILLER_12_1265 ();
 FILLCELL_X4 FILLER_12_1270 ();
 FILLCELL_X8 FILLER_12_1288 ();
 FILLCELL_X4 FILLER_12_1307 ();
 FILLCELL_X4 FILLER_12_1322 ();
 FILLCELL_X4 FILLER_12_1330 ();
 FILLCELL_X4 FILLER_12_1338 ();
 FILLCELL_X4 FILLER_12_1349 ();
 FILLCELL_X4 FILLER_12_1357 ();
 FILLCELL_X4 FILLER_12_1364 ();
 FILLCELL_X32 FILLER_12_1370 ();
 FILLCELL_X32 FILLER_12_1402 ();
 FILLCELL_X32 FILLER_12_1434 ();
 FILLCELL_X32 FILLER_12_1466 ();
 FILLCELL_X32 FILLER_12_1498 ();
 FILLCELL_X4 FILLER_12_1530 ();
 FILLCELL_X1 FILLER_12_1534 ();
 FILLCELL_X32 FILLER_12_1539 ();
 FILLCELL_X32 FILLER_12_1571 ();
 FILLCELL_X32 FILLER_12_1603 ();
 FILLCELL_X32 FILLER_12_1635 ();
 FILLCELL_X32 FILLER_12_1667 ();
 FILLCELL_X2 FILLER_12_1699 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_225 ();
 FILLCELL_X32 FILLER_13_257 ();
 FILLCELL_X32 FILLER_13_289 ();
 FILLCELL_X32 FILLER_13_321 ();
 FILLCELL_X8 FILLER_13_353 ();
 FILLCELL_X4 FILLER_13_361 ();
 FILLCELL_X2 FILLER_13_365 ();
 FILLCELL_X1 FILLER_13_367 ();
 FILLCELL_X4 FILLER_13_372 ();
 FILLCELL_X8 FILLER_13_385 ();
 FILLCELL_X2 FILLER_13_393 ();
 FILLCELL_X1 FILLER_13_395 ();
 FILLCELL_X8 FILLER_13_405 ();
 FILLCELL_X1 FILLER_13_413 ();
 FILLCELL_X16 FILLER_13_423 ();
 FILLCELL_X4 FILLER_13_439 ();
 FILLCELL_X1 FILLER_13_443 ();
 FILLCELL_X4 FILLER_13_447 ();
 FILLCELL_X4 FILLER_13_454 ();
 FILLCELL_X8 FILLER_13_461 ();
 FILLCELL_X4 FILLER_13_469 ();
 FILLCELL_X2 FILLER_13_473 ();
 FILLCELL_X1 FILLER_13_475 ();
 FILLCELL_X4 FILLER_13_485 ();
 FILLCELL_X4 FILLER_13_493 ();
 FILLCELL_X2 FILLER_13_497 ();
 FILLCELL_X1 FILLER_13_499 ();
 FILLCELL_X4 FILLER_13_505 ();
 FILLCELL_X4 FILLER_13_512 ();
 FILLCELL_X4 FILLER_13_520 ();
 FILLCELL_X8 FILLER_13_533 ();
 FILLCELL_X2 FILLER_13_541 ();
 FILLCELL_X4 FILLER_13_549 ();
 FILLCELL_X8 FILLER_13_555 ();
 FILLCELL_X1 FILLER_13_563 ();
 FILLCELL_X4 FILLER_13_574 ();
 FILLCELL_X8 FILLER_13_587 ();
 FILLCELL_X4 FILLER_13_602 ();
 FILLCELL_X4 FILLER_13_609 ();
 FILLCELL_X8 FILLER_13_616 ();
 FILLCELL_X2 FILLER_13_624 ();
 FILLCELL_X1 FILLER_13_626 ();
 FILLCELL_X8 FILLER_13_630 ();
 FILLCELL_X4 FILLER_13_641 ();
 FILLCELL_X8 FILLER_13_655 ();
 FILLCELL_X4 FILLER_13_663 ();
 FILLCELL_X1 FILLER_13_667 ();
 FILLCELL_X4 FILLER_13_671 ();
 FILLCELL_X4 FILLER_13_678 ();
 FILLCELL_X2 FILLER_13_682 ();
 FILLCELL_X1 FILLER_13_684 ();
 FILLCELL_X16 FILLER_13_690 ();
 FILLCELL_X16 FILLER_13_711 ();
 FILLCELL_X2 FILLER_13_727 ();
 FILLCELL_X1 FILLER_13_729 ();
 FILLCELL_X8 FILLER_13_748 ();
 FILLCELL_X4 FILLER_13_756 ();
 FILLCELL_X4 FILLER_13_767 ();
 FILLCELL_X2 FILLER_13_771 ();
 FILLCELL_X4 FILLER_13_780 ();
 FILLCELL_X1 FILLER_13_784 ();
 FILLCELL_X4 FILLER_13_792 ();
 FILLCELL_X4 FILLER_13_803 ();
 FILLCELL_X16 FILLER_13_814 ();
 FILLCELL_X16 FILLER_13_837 ();
 FILLCELL_X1 FILLER_13_853 ();
 FILLCELL_X16 FILLER_13_861 ();
 FILLCELL_X4 FILLER_13_877 ();
 FILLCELL_X2 FILLER_13_881 ();
 FILLCELL_X1 FILLER_13_883 ();
 FILLCELL_X16 FILLER_13_888 ();
 FILLCELL_X8 FILLER_13_904 ();
 FILLCELL_X4 FILLER_13_918 ();
 FILLCELL_X4 FILLER_13_925 ();
 FILLCELL_X2 FILLER_13_929 ();
 FILLCELL_X1 FILLER_13_931 ();
 FILLCELL_X8 FILLER_13_945 ();
 FILLCELL_X2 FILLER_13_953 ();
 FILLCELL_X8 FILLER_13_958 ();
 FILLCELL_X4 FILLER_13_979 ();
 FILLCELL_X8 FILLER_13_986 ();
 FILLCELL_X4 FILLER_13_994 ();
 FILLCELL_X2 FILLER_13_998 ();
 FILLCELL_X1 FILLER_13_1000 ();
 FILLCELL_X4 FILLER_13_1006 ();
 FILLCELL_X2 FILLER_13_1010 ();
 FILLCELL_X1 FILLER_13_1012 ();
 FILLCELL_X8 FILLER_13_1026 ();
 FILLCELL_X2 FILLER_13_1034 ();
 FILLCELL_X8 FILLER_13_1045 ();
 FILLCELL_X1 FILLER_13_1053 ();
 FILLCELL_X8 FILLER_13_1057 ();
 FILLCELL_X4 FILLER_13_1065 ();
 FILLCELL_X16 FILLER_13_1076 ();
 FILLCELL_X8 FILLER_13_1105 ();
 FILLCELL_X2 FILLER_13_1113 ();
 FILLCELL_X1 FILLER_13_1115 ();
 FILLCELL_X4 FILLER_13_1123 ();
 FILLCELL_X4 FILLER_13_1134 ();
 FILLCELL_X4 FILLER_13_1145 ();
 FILLCELL_X4 FILLER_13_1156 ();
 FILLCELL_X4 FILLER_13_1167 ();
 FILLCELL_X2 FILLER_13_1171 ();
 FILLCELL_X1 FILLER_13_1173 ();
 FILLCELL_X4 FILLER_13_1181 ();
 FILLCELL_X4 FILLER_13_1192 ();
 FILLCELL_X8 FILLER_13_1203 ();
 FILLCELL_X16 FILLER_13_1218 ();
 FILLCELL_X2 FILLER_13_1234 ();
 FILLCELL_X4 FILLER_13_1243 ();
 FILLCELL_X8 FILLER_13_1254 ();
 FILLCELL_X1 FILLER_13_1262 ();
 FILLCELL_X4 FILLER_13_1264 ();
 FILLCELL_X4 FILLER_13_1272 ();
 FILLCELL_X8 FILLER_13_1278 ();
 FILLCELL_X1 FILLER_13_1286 ();
 FILLCELL_X4 FILLER_13_1298 ();
 FILLCELL_X2 FILLER_13_1302 ();
 FILLCELL_X4 FILLER_13_1308 ();
 FILLCELL_X4 FILLER_13_1317 ();
 FILLCELL_X4 FILLER_13_1326 ();
 FILLCELL_X8 FILLER_13_1334 ();
 FILLCELL_X4 FILLER_13_1344 ();
 FILLCELL_X4 FILLER_13_1352 ();
 FILLCELL_X32 FILLER_13_1358 ();
 FILLCELL_X32 FILLER_13_1390 ();
 FILLCELL_X32 FILLER_13_1422 ();
 FILLCELL_X32 FILLER_13_1454 ();
 FILLCELL_X32 FILLER_13_1486 ();
 FILLCELL_X32 FILLER_13_1518 ();
 FILLCELL_X32 FILLER_13_1550 ();
 FILLCELL_X32 FILLER_13_1582 ();
 FILLCELL_X32 FILLER_13_1614 ();
 FILLCELL_X32 FILLER_13_1646 ();
 FILLCELL_X16 FILLER_13_1678 ();
 FILLCELL_X4 FILLER_13_1694 ();
 FILLCELL_X2 FILLER_13_1698 ();
 FILLCELL_X1 FILLER_13_1700 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_161 ();
 FILLCELL_X32 FILLER_14_193 ();
 FILLCELL_X32 FILLER_14_225 ();
 FILLCELL_X32 FILLER_14_257 ();
 FILLCELL_X32 FILLER_14_289 ();
 FILLCELL_X32 FILLER_14_321 ();
 FILLCELL_X8 FILLER_14_353 ();
 FILLCELL_X4 FILLER_14_361 ();
 FILLCELL_X2 FILLER_14_365 ();
 FILLCELL_X1 FILLER_14_367 ();
 FILLCELL_X4 FILLER_14_372 ();
 FILLCELL_X8 FILLER_14_385 ();
 FILLCELL_X1 FILLER_14_393 ();
 FILLCELL_X4 FILLER_14_396 ();
 FILLCELL_X4 FILLER_14_403 ();
 FILLCELL_X8 FILLER_14_411 ();
 FILLCELL_X4 FILLER_14_429 ();
 FILLCELL_X4 FILLER_14_435 ();
 FILLCELL_X2 FILLER_14_439 ();
 FILLCELL_X4 FILLER_14_443 ();
 FILLCELL_X1 FILLER_14_447 ();
 FILLCELL_X4 FILLER_14_451 ();
 FILLCELL_X4 FILLER_14_460 ();
 FILLCELL_X4 FILLER_14_474 ();
 FILLCELL_X1 FILLER_14_478 ();
 FILLCELL_X4 FILLER_14_486 ();
 FILLCELL_X8 FILLER_14_497 ();
 FILLCELL_X2 FILLER_14_505 ();
 FILLCELL_X8 FILLER_14_514 ();
 FILLCELL_X2 FILLER_14_522 ();
 FILLCELL_X8 FILLER_14_530 ();
 FILLCELL_X4 FILLER_14_538 ();
 FILLCELL_X4 FILLER_14_548 ();
 FILLCELL_X16 FILLER_14_557 ();
 FILLCELL_X8 FILLER_14_573 ();
 FILLCELL_X1 FILLER_14_581 ();
 FILLCELL_X4 FILLER_14_589 ();
 FILLCELL_X2 FILLER_14_593 ();
 FILLCELL_X1 FILLER_14_595 ();
 FILLCELL_X8 FILLER_14_606 ();
 FILLCELL_X4 FILLER_14_614 ();
 FILLCELL_X2 FILLER_14_618 ();
 FILLCELL_X4 FILLER_14_627 ();
 FILLCELL_X4 FILLER_14_632 ();
 FILLCELL_X4 FILLER_14_646 ();
 FILLCELL_X4 FILLER_14_657 ();
 FILLCELL_X4 FILLER_14_668 ();
 FILLCELL_X8 FILLER_14_675 ();
 FILLCELL_X4 FILLER_14_690 ();
 FILLCELL_X2 FILLER_14_694 ();
 FILLCELL_X4 FILLER_14_703 ();
 FILLCELL_X1 FILLER_14_707 ();
 FILLCELL_X4 FILLER_14_711 ();
 FILLCELL_X8 FILLER_14_719 ();
 FILLCELL_X4 FILLER_14_730 ();
 FILLCELL_X4 FILLER_14_738 ();
 FILLCELL_X4 FILLER_14_746 ();
 FILLCELL_X4 FILLER_14_757 ();
 FILLCELL_X4 FILLER_14_768 ();
 FILLCELL_X2 FILLER_14_772 ();
 FILLCELL_X1 FILLER_14_774 ();
 FILLCELL_X4 FILLER_14_782 ();
 FILLCELL_X4 FILLER_14_789 ();
 FILLCELL_X4 FILLER_14_796 ();
 FILLCELL_X1 FILLER_14_800 ();
 FILLCELL_X4 FILLER_14_804 ();
 FILLCELL_X2 FILLER_14_808 ();
 FILLCELL_X8 FILLER_14_814 ();
 FILLCELL_X1 FILLER_14_822 ();
 FILLCELL_X4 FILLER_14_830 ();
 FILLCELL_X4 FILLER_14_841 ();
 FILLCELL_X4 FILLER_14_852 ();
 FILLCELL_X4 FILLER_14_863 ();
 FILLCELL_X8 FILLER_14_874 ();
 FILLCELL_X2 FILLER_14_882 ();
 FILLCELL_X4 FILLER_14_888 ();
 FILLCELL_X4 FILLER_14_899 ();
 FILLCELL_X4 FILLER_14_912 ();
 FILLCELL_X8 FILLER_14_919 ();
 FILLCELL_X4 FILLER_14_927 ();
 FILLCELL_X2 FILLER_14_931 ();
 FILLCELL_X1 FILLER_14_933 ();
 FILLCELL_X4 FILLER_14_937 ();
 FILLCELL_X4 FILLER_14_944 ();
 FILLCELL_X2 FILLER_14_948 ();
 FILLCELL_X8 FILLER_14_953 ();
 FILLCELL_X2 FILLER_14_961 ();
 FILLCELL_X8 FILLER_14_970 ();
 FILLCELL_X1 FILLER_14_978 ();
 FILLCELL_X4 FILLER_14_984 ();
 FILLCELL_X4 FILLER_14_997 ();
 FILLCELL_X8 FILLER_14_1014 ();
 FILLCELL_X2 FILLER_14_1022 ();
 FILLCELL_X4 FILLER_14_1028 ();
 FILLCELL_X8 FILLER_14_1035 ();
 FILLCELL_X2 FILLER_14_1043 ();
 FILLCELL_X4 FILLER_14_1052 ();
 FILLCELL_X2 FILLER_14_1056 ();
 FILLCELL_X1 FILLER_14_1058 ();
 FILLCELL_X4 FILLER_14_1072 ();
 FILLCELL_X4 FILLER_14_1083 ();
 FILLCELL_X4 FILLER_14_1090 ();
 FILLCELL_X4 FILLER_14_1101 ();
 FILLCELL_X2 FILLER_14_1105 ();
 FILLCELL_X1 FILLER_14_1107 ();
 FILLCELL_X4 FILLER_14_1112 ();
 FILLCELL_X2 FILLER_14_1116 ();
 FILLCELL_X4 FILLER_14_1125 ();
 FILLCELL_X4 FILLER_14_1136 ();
 FILLCELL_X4 FILLER_14_1147 ();
 FILLCELL_X8 FILLER_14_1158 ();
 FILLCELL_X1 FILLER_14_1166 ();
 FILLCELL_X4 FILLER_14_1174 ();
 FILLCELL_X16 FILLER_14_1185 ();
 FILLCELL_X1 FILLER_14_1201 ();
 FILLCELL_X4 FILLER_14_1209 ();
 FILLCELL_X4 FILLER_14_1220 ();
 FILLCELL_X4 FILLER_14_1231 ();
 FILLCELL_X8 FILLER_14_1242 ();
 FILLCELL_X4 FILLER_14_1259 ();
 FILLCELL_X1 FILLER_14_1263 ();
 FILLCELL_X4 FILLER_14_1266 ();
 FILLCELL_X4 FILLER_14_1274 ();
 FILLCELL_X8 FILLER_14_1282 ();
 FILLCELL_X4 FILLER_14_1290 ();
 FILLCELL_X2 FILLER_14_1294 ();
 FILLCELL_X8 FILLER_14_1301 ();
 FILLCELL_X2 FILLER_14_1309 ();
 FILLCELL_X4 FILLER_14_1314 ();
 FILLCELL_X1 FILLER_14_1318 ();
 FILLCELL_X4 FILLER_14_1324 ();
 FILLCELL_X8 FILLER_14_1332 ();
 FILLCELL_X2 FILLER_14_1340 ();
 FILLCELL_X1 FILLER_14_1342 ();
 FILLCELL_X4 FILLER_14_1345 ();
 FILLCELL_X4 FILLER_14_1353 ();
 FILLCELL_X4 FILLER_14_1361 ();
 FILLCELL_X32 FILLER_14_1368 ();
 FILLCELL_X32 FILLER_14_1400 ();
 FILLCELL_X32 FILLER_14_1432 ();
 FILLCELL_X32 FILLER_14_1464 ();
 FILLCELL_X32 FILLER_14_1496 ();
 FILLCELL_X32 FILLER_14_1528 ();
 FILLCELL_X32 FILLER_14_1560 ();
 FILLCELL_X32 FILLER_14_1592 ();
 FILLCELL_X32 FILLER_14_1624 ();
 FILLCELL_X32 FILLER_14_1656 ();
 FILLCELL_X8 FILLER_14_1688 ();
 FILLCELL_X4 FILLER_14_1696 ();
 FILLCELL_X1 FILLER_14_1700 ();
 FILLCELL_X4 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_8 ();
 FILLCELL_X32 FILLER_15_40 ();
 FILLCELL_X32 FILLER_15_72 ();
 FILLCELL_X32 FILLER_15_104 ();
 FILLCELL_X32 FILLER_15_136 ();
 FILLCELL_X32 FILLER_15_168 ();
 FILLCELL_X32 FILLER_15_200 ();
 FILLCELL_X32 FILLER_15_232 ();
 FILLCELL_X32 FILLER_15_264 ();
 FILLCELL_X32 FILLER_15_296 ();
 FILLCELL_X32 FILLER_15_328 ();
 FILLCELL_X16 FILLER_15_360 ();
 FILLCELL_X4 FILLER_15_376 ();
 FILLCELL_X4 FILLER_15_383 ();
 FILLCELL_X4 FILLER_15_389 ();
 FILLCELL_X4 FILLER_15_396 ();
 FILLCELL_X4 FILLER_15_403 ();
 FILLCELL_X4 FILLER_15_411 ();
 FILLCELL_X4 FILLER_15_418 ();
 FILLCELL_X4 FILLER_15_424 ();
 FILLCELL_X1 FILLER_15_428 ();
 FILLCELL_X4 FILLER_15_431 ();
 FILLCELL_X4 FILLER_15_444 ();
 FILLCELL_X8 FILLER_15_455 ();
 FILLCELL_X4 FILLER_15_463 ();
 FILLCELL_X2 FILLER_15_467 ();
 FILLCELL_X4 FILLER_15_476 ();
 FILLCELL_X8 FILLER_15_483 ();
 FILLCELL_X4 FILLER_15_491 ();
 FILLCELL_X2 FILLER_15_495 ();
 FILLCELL_X4 FILLER_15_502 ();
 FILLCELL_X2 FILLER_15_506 ();
 FILLCELL_X4 FILLER_15_511 ();
 FILLCELL_X4 FILLER_15_518 ();
 FILLCELL_X4 FILLER_15_526 ();
 FILLCELL_X8 FILLER_15_532 ();
 FILLCELL_X4 FILLER_15_540 ();
 FILLCELL_X1 FILLER_15_544 ();
 FILLCELL_X4 FILLER_15_548 ();
 FILLCELL_X8 FILLER_15_554 ();
 FILLCELL_X2 FILLER_15_562 ();
 FILLCELL_X4 FILLER_15_569 ();
 FILLCELL_X8 FILLER_15_575 ();
 FILLCELL_X1 FILLER_15_583 ();
 FILLCELL_X16 FILLER_15_591 ();
 FILLCELL_X4 FILLER_15_607 ();
 FILLCELL_X2 FILLER_15_611 ();
 FILLCELL_X8 FILLER_15_616 ();
 FILLCELL_X4 FILLER_15_624 ();
 FILLCELL_X1 FILLER_15_628 ();
 FILLCELL_X4 FILLER_15_636 ();
 FILLCELL_X2 FILLER_15_640 ();
 FILLCELL_X4 FILLER_15_651 ();
 FILLCELL_X8 FILLER_15_658 ();
 FILLCELL_X4 FILLER_15_666 ();
 FILLCELL_X8 FILLER_15_674 ();
 FILLCELL_X4 FILLER_15_682 ();
 FILLCELL_X2 FILLER_15_686 ();
 FILLCELL_X4 FILLER_15_695 ();
 FILLCELL_X4 FILLER_15_713 ();
 FILLCELL_X1 FILLER_15_717 ();
 FILLCELL_X4 FILLER_15_727 ();
 FILLCELL_X4 FILLER_15_738 ();
 FILLCELL_X2 FILLER_15_742 ();
 FILLCELL_X16 FILLER_15_751 ();
 FILLCELL_X8 FILLER_15_767 ();
 FILLCELL_X4 FILLER_15_782 ();
 FILLCELL_X1 FILLER_15_786 ();
 FILLCELL_X8 FILLER_15_794 ();
 FILLCELL_X4 FILLER_15_802 ();
 FILLCELL_X2 FILLER_15_806 ();
 FILLCELL_X8 FILLER_15_815 ();
 FILLCELL_X1 FILLER_15_823 ();
 FILLCELL_X16 FILLER_15_831 ();
 FILLCELL_X4 FILLER_15_847 ();
 FILLCELL_X1 FILLER_15_851 ();
 FILLCELL_X4 FILLER_15_855 ();
 FILLCELL_X8 FILLER_15_866 ();
 FILLCELL_X2 FILLER_15_874 ();
 FILLCELL_X1 FILLER_15_876 ();
 FILLCELL_X4 FILLER_15_884 ();
 FILLCELL_X8 FILLER_15_895 ();
 FILLCELL_X2 FILLER_15_903 ();
 FILLCELL_X4 FILLER_15_914 ();
 FILLCELL_X4 FILLER_15_921 ();
 FILLCELL_X2 FILLER_15_925 ();
 FILLCELL_X4 FILLER_15_934 ();
 FILLCELL_X4 FILLER_15_943 ();
 FILLCELL_X4 FILLER_15_952 ();
 FILLCELL_X16 FILLER_15_965 ();
 FILLCELL_X1 FILLER_15_981 ();
 FILLCELL_X4 FILLER_15_989 ();
 FILLCELL_X4 FILLER_15_999 ();
 FILLCELL_X2 FILLER_15_1003 ();
 FILLCELL_X1 FILLER_15_1005 ();
 FILLCELL_X4 FILLER_15_1009 ();
 FILLCELL_X1 FILLER_15_1013 ();
 FILLCELL_X4 FILLER_15_1023 ();
 FILLCELL_X4 FILLER_15_1044 ();
 FILLCELL_X4 FILLER_15_1062 ();
 FILLCELL_X4 FILLER_15_1069 ();
 FILLCELL_X2 FILLER_15_1073 ();
 FILLCELL_X1 FILLER_15_1075 ();
 FILLCELL_X4 FILLER_15_1083 ();
 FILLCELL_X8 FILLER_15_1094 ();
 FILLCELL_X2 FILLER_15_1102 ();
 FILLCELL_X1 FILLER_15_1104 ();
 FILLCELL_X4 FILLER_15_1122 ();
 FILLCELL_X8 FILLER_15_1135 ();
 FILLCELL_X4 FILLER_15_1143 ();
 FILLCELL_X1 FILLER_15_1147 ();
 FILLCELL_X16 FILLER_15_1155 ();
 FILLCELL_X8 FILLER_15_1171 ();
 FILLCELL_X4 FILLER_15_1179 ();
 FILLCELL_X1 FILLER_15_1183 ();
 FILLCELL_X8 FILLER_15_1191 ();
 FILLCELL_X1 FILLER_15_1199 ();
 FILLCELL_X8 FILLER_15_1209 ();
 FILLCELL_X4 FILLER_15_1217 ();
 FILLCELL_X1 FILLER_15_1221 ();
 FILLCELL_X8 FILLER_15_1231 ();
 FILLCELL_X1 FILLER_15_1239 ();
 FILLCELL_X4 FILLER_15_1247 ();
 FILLCELL_X4 FILLER_15_1256 ();
 FILLCELL_X2 FILLER_15_1260 ();
 FILLCELL_X1 FILLER_15_1262 ();
 FILLCELL_X8 FILLER_15_1264 ();
 FILLCELL_X2 FILLER_15_1272 ();
 FILLCELL_X4 FILLER_15_1281 ();
 FILLCELL_X4 FILLER_15_1292 ();
 FILLCELL_X4 FILLER_15_1301 ();
 FILLCELL_X4 FILLER_15_1310 ();
 FILLCELL_X4 FILLER_15_1319 ();
 FILLCELL_X4 FILLER_15_1327 ();
 FILLCELL_X16 FILLER_15_1335 ();
 FILLCELL_X2 FILLER_15_1351 ();
 FILLCELL_X4 FILLER_15_1357 ();
 FILLCELL_X32 FILLER_15_1365 ();
 FILLCELL_X32 FILLER_15_1397 ();
 FILLCELL_X32 FILLER_15_1429 ();
 FILLCELL_X32 FILLER_15_1461 ();
 FILLCELL_X32 FILLER_15_1493 ();
 FILLCELL_X8 FILLER_15_1525 ();
 FILLCELL_X4 FILLER_15_1533 ();
 FILLCELL_X2 FILLER_15_1537 ();
 FILLCELL_X1 FILLER_15_1539 ();
 FILLCELL_X4 FILLER_15_1544 ();
 FILLCELL_X2 FILLER_15_1548 ();
 FILLCELL_X1 FILLER_15_1550 ();
 FILLCELL_X32 FILLER_15_1568 ();
 FILLCELL_X32 FILLER_15_1600 ();
 FILLCELL_X32 FILLER_15_1632 ();
 FILLCELL_X32 FILLER_15_1664 ();
 FILLCELL_X4 FILLER_15_1696 ();
 FILLCELL_X1 FILLER_15_1700 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X32 FILLER_16_161 ();
 FILLCELL_X32 FILLER_16_193 ();
 FILLCELL_X32 FILLER_16_225 ();
 FILLCELL_X32 FILLER_16_257 ();
 FILLCELL_X32 FILLER_16_289 ();
 FILLCELL_X32 FILLER_16_321 ();
 FILLCELL_X16 FILLER_16_353 ();
 FILLCELL_X1 FILLER_16_369 ();
 FILLCELL_X4 FILLER_16_373 ();
 FILLCELL_X4 FILLER_16_381 ();
 FILLCELL_X2 FILLER_16_385 ();
 FILLCELL_X4 FILLER_16_392 ();
 FILLCELL_X4 FILLER_16_405 ();
 FILLCELL_X2 FILLER_16_409 ();
 FILLCELL_X4 FILLER_16_418 ();
 FILLCELL_X4 FILLER_16_431 ();
 FILLCELL_X4 FILLER_16_438 ();
 FILLCELL_X1 FILLER_16_442 ();
 FILLCELL_X4 FILLER_16_446 ();
 FILLCELL_X4 FILLER_16_459 ();
 FILLCELL_X2 FILLER_16_463 ();
 FILLCELL_X8 FILLER_16_468 ();
 FILLCELL_X1 FILLER_16_476 ();
 FILLCELL_X8 FILLER_16_486 ();
 FILLCELL_X2 FILLER_16_494 ();
 FILLCELL_X4 FILLER_16_503 ();
 FILLCELL_X2 FILLER_16_507 ();
 FILLCELL_X4 FILLER_16_516 ();
 FILLCELL_X1 FILLER_16_520 ();
 FILLCELL_X4 FILLER_16_528 ();
 FILLCELL_X4 FILLER_16_536 ();
 FILLCELL_X8 FILLER_16_543 ();
 FILLCELL_X1 FILLER_16_551 ();
 FILLCELL_X4 FILLER_16_555 ();
 FILLCELL_X4 FILLER_16_565 ();
 FILLCELL_X8 FILLER_16_579 ();
 FILLCELL_X2 FILLER_16_587 ();
 FILLCELL_X1 FILLER_16_589 ();
 FILLCELL_X4 FILLER_16_597 ();
 FILLCELL_X8 FILLER_16_608 ();
 FILLCELL_X2 FILLER_16_616 ();
 FILLCELL_X8 FILLER_16_621 ();
 FILLCELL_X2 FILLER_16_629 ();
 FILLCELL_X8 FILLER_16_632 ();
 FILLCELL_X1 FILLER_16_640 ();
 FILLCELL_X4 FILLER_16_645 ();
 FILLCELL_X4 FILLER_16_653 ();
 FILLCELL_X2 FILLER_16_657 ();
 FILLCELL_X1 FILLER_16_659 ();
 FILLCELL_X4 FILLER_16_663 ();
 FILLCELL_X8 FILLER_16_676 ();
 FILLCELL_X4 FILLER_16_684 ();
 FILLCELL_X2 FILLER_16_688 ();
 FILLCELL_X8 FILLER_16_696 ();
 FILLCELL_X8 FILLER_16_708 ();
 FILLCELL_X8 FILLER_16_719 ();
 FILLCELL_X2 FILLER_16_727 ();
 FILLCELL_X4 FILLER_16_732 ();
 FILLCELL_X8 FILLER_16_743 ();
 FILLCELL_X2 FILLER_16_751 ();
 FILLCELL_X1 FILLER_16_753 ();
 FILLCELL_X4 FILLER_16_757 ();
 FILLCELL_X4 FILLER_16_768 ();
 FILLCELL_X2 FILLER_16_772 ();
 FILLCELL_X1 FILLER_16_774 ();
 FILLCELL_X16 FILLER_16_782 ();
 FILLCELL_X1 FILLER_16_798 ();
 FILLCELL_X4 FILLER_16_806 ();
 FILLCELL_X4 FILLER_16_814 ();
 FILLCELL_X4 FILLER_16_825 ();
 FILLCELL_X8 FILLER_16_836 ();
 FILLCELL_X4 FILLER_16_844 ();
 FILLCELL_X2 FILLER_16_848 ();
 FILLCELL_X1 FILLER_16_850 ();
 FILLCELL_X32 FILLER_16_858 ();
 FILLCELL_X8 FILLER_16_894 ();
 FILLCELL_X2 FILLER_16_902 ();
 FILLCELL_X1 FILLER_16_904 ();
 FILLCELL_X8 FILLER_16_912 ();
 FILLCELL_X1 FILLER_16_920 ();
 FILLCELL_X16 FILLER_16_924 ();
 FILLCELL_X4 FILLER_16_940 ();
 FILLCELL_X2 FILLER_16_944 ();
 FILLCELL_X4 FILLER_16_949 ();
 FILLCELL_X1 FILLER_16_953 ();
 FILLCELL_X8 FILLER_16_963 ();
 FILLCELL_X4 FILLER_16_971 ();
 FILLCELL_X2 FILLER_16_975 ();
 FILLCELL_X1 FILLER_16_977 ();
 FILLCELL_X4 FILLER_16_987 ();
 FILLCELL_X4 FILLER_16_993 ();
 FILLCELL_X8 FILLER_16_1004 ();
 FILLCELL_X2 FILLER_16_1012 ();
 FILLCELL_X4 FILLER_16_1021 ();
 FILLCELL_X4 FILLER_16_1028 ();
 FILLCELL_X2 FILLER_16_1032 ();
 FILLCELL_X16 FILLER_16_1037 ();
 FILLCELL_X8 FILLER_16_1053 ();
 FILLCELL_X4 FILLER_16_1061 ();
 FILLCELL_X2 FILLER_16_1065 ();
 FILLCELL_X1 FILLER_16_1067 ();
 FILLCELL_X16 FILLER_16_1075 ();
 FILLCELL_X8 FILLER_16_1091 ();
 FILLCELL_X4 FILLER_16_1099 ();
 FILLCELL_X1 FILLER_16_1103 ();
 FILLCELL_X4 FILLER_16_1108 ();
 FILLCELL_X1 FILLER_16_1112 ();
 FILLCELL_X4 FILLER_16_1117 ();
 FILLCELL_X16 FILLER_16_1125 ();
 FILLCELL_X1 FILLER_16_1141 ();
 FILLCELL_X8 FILLER_16_1149 ();
 FILLCELL_X4 FILLER_16_1157 ();
 FILLCELL_X2 FILLER_16_1161 ();
 FILLCELL_X8 FILLER_16_1170 ();
 FILLCELL_X4 FILLER_16_1185 ();
 FILLCELL_X8 FILLER_16_1196 ();
 FILLCELL_X16 FILLER_16_1213 ();
 FILLCELL_X4 FILLER_16_1229 ();
 FILLCELL_X1 FILLER_16_1233 ();
 FILLCELL_X4 FILLER_16_1241 ();
 FILLCELL_X16 FILLER_16_1247 ();
 FILLCELL_X4 FILLER_16_1263 ();
 FILLCELL_X2 FILLER_16_1267 ();
 FILLCELL_X4 FILLER_16_1272 ();
 FILLCELL_X16 FILLER_16_1278 ();
 FILLCELL_X4 FILLER_16_1294 ();
 FILLCELL_X1 FILLER_16_1298 ();
 FILLCELL_X4 FILLER_16_1303 ();
 FILLCELL_X2 FILLER_16_1307 ();
 FILLCELL_X1 FILLER_16_1309 ();
 FILLCELL_X4 FILLER_16_1315 ();
 FILLCELL_X4 FILLER_16_1324 ();
 FILLCELL_X4 FILLER_16_1333 ();
 FILLCELL_X4 FILLER_16_1341 ();
 FILLCELL_X2 FILLER_16_1345 ();
 FILLCELL_X4 FILLER_16_1351 ();
 FILLCELL_X4 FILLER_16_1360 ();
 FILLCELL_X4 FILLER_16_1367 ();
 FILLCELL_X32 FILLER_16_1373 ();
 FILLCELL_X32 FILLER_16_1405 ();
 FILLCELL_X32 FILLER_16_1437 ();
 FILLCELL_X32 FILLER_16_1469 ();
 FILLCELL_X32 FILLER_16_1501 ();
 FILLCELL_X32 FILLER_16_1533 ();
 FILLCELL_X32 FILLER_16_1565 ();
 FILLCELL_X32 FILLER_16_1597 ();
 FILLCELL_X32 FILLER_16_1629 ();
 FILLCELL_X32 FILLER_16_1661 ();
 FILLCELL_X8 FILLER_16_1693 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X32 FILLER_17_161 ();
 FILLCELL_X32 FILLER_17_193 ();
 FILLCELL_X32 FILLER_17_225 ();
 FILLCELL_X32 FILLER_17_257 ();
 FILLCELL_X32 FILLER_17_289 ();
 FILLCELL_X32 FILLER_17_321 ();
 FILLCELL_X32 FILLER_17_353 ();
 FILLCELL_X4 FILLER_17_385 ();
 FILLCELL_X2 FILLER_17_389 ();
 FILLCELL_X4 FILLER_17_395 ();
 FILLCELL_X16 FILLER_17_403 ();
 FILLCELL_X4 FILLER_17_422 ();
 FILLCELL_X1 FILLER_17_426 ();
 FILLCELL_X8 FILLER_17_430 ();
 FILLCELL_X8 FILLER_17_445 ();
 FILLCELL_X4 FILLER_17_456 ();
 FILLCELL_X2 FILLER_17_460 ();
 FILLCELL_X1 FILLER_17_462 ();
 FILLCELL_X4 FILLER_17_470 ();
 FILLCELL_X2 FILLER_17_474 ();
 FILLCELL_X4 FILLER_17_479 ();
 FILLCELL_X4 FILLER_17_486 ();
 FILLCELL_X8 FILLER_17_493 ();
 FILLCELL_X1 FILLER_17_501 ();
 FILLCELL_X8 FILLER_17_509 ();
 FILLCELL_X4 FILLER_17_517 ();
 FILLCELL_X2 FILLER_17_521 ();
 FILLCELL_X4 FILLER_17_530 ();
 FILLCELL_X4 FILLER_17_541 ();
 FILLCELL_X4 FILLER_17_552 ();
 FILLCELL_X8 FILLER_17_562 ();
 FILLCELL_X1 FILLER_17_570 ();
 FILLCELL_X4 FILLER_17_575 ();
 FILLCELL_X4 FILLER_17_583 ();
 FILLCELL_X2 FILLER_17_587 ();
 FILLCELL_X1 FILLER_17_589 ();
 FILLCELL_X4 FILLER_17_593 ();
 FILLCELL_X2 FILLER_17_597 ();
 FILLCELL_X1 FILLER_17_599 ();
 FILLCELL_X4 FILLER_17_604 ();
 FILLCELL_X4 FILLER_17_617 ();
 FILLCELL_X4 FILLER_17_627 ();
 FILLCELL_X4 FILLER_17_638 ();
 FILLCELL_X4 FILLER_17_648 ();
 FILLCELL_X4 FILLER_17_655 ();
 FILLCELL_X4 FILLER_17_661 ();
 FILLCELL_X4 FILLER_17_672 ();
 FILLCELL_X4 FILLER_17_683 ();
 FILLCELL_X4 FILLER_17_694 ();
 FILLCELL_X4 FILLER_17_701 ();
 FILLCELL_X16 FILLER_17_708 ();
 FILLCELL_X2 FILLER_17_724 ();
 FILLCELL_X1 FILLER_17_726 ();
 FILLCELL_X4 FILLER_17_734 ();
 FILLCELL_X2 FILLER_17_738 ();
 FILLCELL_X4 FILLER_17_744 ();
 FILLCELL_X4 FILLER_17_755 ();
 FILLCELL_X2 FILLER_17_759 ();
 FILLCELL_X1 FILLER_17_761 ();
 FILLCELL_X4 FILLER_17_766 ();
 FILLCELL_X1 FILLER_17_770 ();
 FILLCELL_X4 FILLER_17_778 ();
 FILLCELL_X2 FILLER_17_782 ();
 FILLCELL_X4 FILLER_17_791 ();
 FILLCELL_X8 FILLER_17_802 ();
 FILLCELL_X2 FILLER_17_810 ();
 FILLCELL_X8 FILLER_17_819 ();
 FILLCELL_X1 FILLER_17_827 ();
 FILLCELL_X4 FILLER_17_835 ();
 FILLCELL_X4 FILLER_17_846 ();
 FILLCELL_X2 FILLER_17_850 ();
 FILLCELL_X1 FILLER_17_852 ();
 FILLCELL_X8 FILLER_17_862 ();
 FILLCELL_X1 FILLER_17_870 ();
 FILLCELL_X8 FILLER_17_874 ();
 FILLCELL_X1 FILLER_17_882 ();
 FILLCELL_X4 FILLER_17_890 ();
 FILLCELL_X4 FILLER_17_901 ();
 FILLCELL_X2 FILLER_17_905 ();
 FILLCELL_X4 FILLER_17_914 ();
 FILLCELL_X8 FILLER_17_921 ();
 FILLCELL_X1 FILLER_17_929 ();
 FILLCELL_X4 FILLER_17_940 ();
 FILLCELL_X4 FILLER_17_947 ();
 FILLCELL_X4 FILLER_17_954 ();
 FILLCELL_X4 FILLER_17_965 ();
 FILLCELL_X4 FILLER_17_973 ();
 FILLCELL_X8 FILLER_17_980 ();
 FILLCELL_X4 FILLER_17_988 ();
 FILLCELL_X2 FILLER_17_992 ();
 FILLCELL_X4 FILLER_17_1001 ();
 FILLCELL_X2 FILLER_17_1005 ();
 FILLCELL_X8 FILLER_17_1016 ();
 FILLCELL_X4 FILLER_17_1024 ();
 FILLCELL_X2 FILLER_17_1028 ();
 FILLCELL_X4 FILLER_17_1043 ();
 FILLCELL_X8 FILLER_17_1056 ();
 FILLCELL_X1 FILLER_17_1064 ();
 FILLCELL_X4 FILLER_17_1072 ();
 FILLCELL_X2 FILLER_17_1076 ();
 FILLCELL_X1 FILLER_17_1078 ();
 FILLCELL_X8 FILLER_17_1086 ();
 FILLCELL_X4 FILLER_17_1098 ();
 FILLCELL_X2 FILLER_17_1102 ();
 FILLCELL_X1 FILLER_17_1104 ();
 FILLCELL_X32 FILLER_17_1112 ();
 FILLCELL_X8 FILLER_17_1144 ();
 FILLCELL_X1 FILLER_17_1152 ();
 FILLCELL_X8 FILLER_17_1160 ();
 FILLCELL_X4 FILLER_17_1168 ();
 FILLCELL_X4 FILLER_17_1179 ();
 FILLCELL_X4 FILLER_17_1190 ();
 FILLCELL_X4 FILLER_17_1201 ();
 FILLCELL_X2 FILLER_17_1205 ();
 FILLCELL_X8 FILLER_17_1216 ();
 FILLCELL_X16 FILLER_17_1237 ();
 FILLCELL_X8 FILLER_17_1253 ();
 FILLCELL_X2 FILLER_17_1261 ();
 FILLCELL_X4 FILLER_17_1264 ();
 FILLCELL_X1 FILLER_17_1268 ();
 FILLCELL_X4 FILLER_17_1271 ();
 FILLCELL_X2 FILLER_17_1275 ();
 FILLCELL_X4 FILLER_17_1279 ();
 FILLCELL_X8 FILLER_17_1285 ();
 FILLCELL_X4 FILLER_17_1298 ();
 FILLCELL_X4 FILLER_17_1307 ();
 FILLCELL_X4 FILLER_17_1316 ();
 FILLCELL_X4 FILLER_17_1325 ();
 FILLCELL_X8 FILLER_17_1334 ();
 FILLCELL_X4 FILLER_17_1342 ();
 FILLCELL_X1 FILLER_17_1346 ();
 FILLCELL_X4 FILLER_17_1351 ();
 FILLCELL_X32 FILLER_17_1357 ();
 FILLCELL_X32 FILLER_17_1389 ();
 FILLCELL_X32 FILLER_17_1421 ();
 FILLCELL_X32 FILLER_17_1453 ();
 FILLCELL_X32 FILLER_17_1485 ();
 FILLCELL_X32 FILLER_17_1517 ();
 FILLCELL_X32 FILLER_17_1549 ();
 FILLCELL_X32 FILLER_17_1581 ();
 FILLCELL_X32 FILLER_17_1613 ();
 FILLCELL_X32 FILLER_17_1645 ();
 FILLCELL_X16 FILLER_17_1677 ();
 FILLCELL_X8 FILLER_17_1693 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X32 FILLER_18_161 ();
 FILLCELL_X32 FILLER_18_193 ();
 FILLCELL_X32 FILLER_18_225 ();
 FILLCELL_X32 FILLER_18_257 ();
 FILLCELL_X32 FILLER_18_289 ();
 FILLCELL_X32 FILLER_18_321 ();
 FILLCELL_X4 FILLER_18_353 ();
 FILLCELL_X2 FILLER_18_357 ();
 FILLCELL_X1 FILLER_18_359 ();
 FILLCELL_X8 FILLER_18_364 ();
 FILLCELL_X4 FILLER_18_376 ();
 FILLCELL_X16 FILLER_18_384 ();
 FILLCELL_X8 FILLER_18_400 ();
 FILLCELL_X1 FILLER_18_408 ();
 FILLCELL_X4 FILLER_18_418 ();
 FILLCELL_X4 FILLER_18_426 ();
 FILLCELL_X2 FILLER_18_430 ();
 FILLCELL_X1 FILLER_18_432 ();
 FILLCELL_X4 FILLER_18_442 ();
 FILLCELL_X4 FILLER_18_456 ();
 FILLCELL_X2 FILLER_18_460 ();
 FILLCELL_X4 FILLER_18_469 ();
 FILLCELL_X8 FILLER_18_480 ();
 FILLCELL_X4 FILLER_18_488 ();
 FILLCELL_X4 FILLER_18_496 ();
 FILLCELL_X8 FILLER_18_503 ();
 FILLCELL_X2 FILLER_18_511 ();
 FILLCELL_X1 FILLER_18_513 ();
 FILLCELL_X8 FILLER_18_518 ();
 FILLCELL_X4 FILLER_18_526 ();
 FILLCELL_X2 FILLER_18_530 ();
 FILLCELL_X8 FILLER_18_535 ();
 FILLCELL_X2 FILLER_18_543 ();
 FILLCELL_X4 FILLER_18_548 ();
 FILLCELL_X4 FILLER_18_555 ();
 FILLCELL_X4 FILLER_18_564 ();
 FILLCELL_X4 FILLER_18_573 ();
 FILLCELL_X4 FILLER_18_587 ();
 FILLCELL_X1 FILLER_18_591 ();
 FILLCELL_X4 FILLER_18_595 ();
 FILLCELL_X8 FILLER_18_602 ();
 FILLCELL_X1 FILLER_18_610 ();
 FILLCELL_X16 FILLER_18_614 ();
 FILLCELL_X1 FILLER_18_630 ();
 FILLCELL_X4 FILLER_18_632 ();
 FILLCELL_X4 FILLER_18_642 ();
 FILLCELL_X1 FILLER_18_646 ();
 FILLCELL_X4 FILLER_18_650 ();
 FILLCELL_X8 FILLER_18_657 ();
 FILLCELL_X4 FILLER_18_665 ();
 FILLCELL_X2 FILLER_18_669 ();
 FILLCELL_X4 FILLER_18_688 ();
 FILLCELL_X2 FILLER_18_692 ();
 FILLCELL_X1 FILLER_18_694 ();
 FILLCELL_X4 FILLER_18_702 ();
 FILLCELL_X2 FILLER_18_706 ();
 FILLCELL_X1 FILLER_18_708 ();
 FILLCELL_X8 FILLER_18_713 ();
 FILLCELL_X1 FILLER_18_721 ();
 FILLCELL_X4 FILLER_18_731 ();
 FILLCELL_X4 FILLER_18_742 ();
 FILLCELL_X4 FILLER_18_750 ();
 FILLCELL_X2 FILLER_18_754 ();
 FILLCELL_X1 FILLER_18_756 ();
 FILLCELL_X32 FILLER_18_761 ();
 FILLCELL_X16 FILLER_18_793 ();
 FILLCELL_X1 FILLER_18_809 ();
 FILLCELL_X4 FILLER_18_817 ();
 FILLCELL_X16 FILLER_18_828 ();
 FILLCELL_X2 FILLER_18_844 ();
 FILLCELL_X8 FILLER_18_853 ();
 FILLCELL_X4 FILLER_18_861 ();
 FILLCELL_X4 FILLER_18_872 ();
 FILLCELL_X1 FILLER_18_876 ();
 FILLCELL_X16 FILLER_18_880 ();
 FILLCELL_X8 FILLER_18_900 ();
 FILLCELL_X4 FILLER_18_908 ();
 FILLCELL_X2 FILLER_18_912 ();
 FILLCELL_X4 FILLER_18_917 ();
 FILLCELL_X4 FILLER_18_926 ();
 FILLCELL_X4 FILLER_18_940 ();
 FILLCELL_X2 FILLER_18_944 ();
 FILLCELL_X8 FILLER_18_953 ();
 FILLCELL_X4 FILLER_18_961 ();
 FILLCELL_X2 FILLER_18_965 ();
 FILLCELL_X4 FILLER_18_973 ();
 FILLCELL_X4 FILLER_18_982 ();
 FILLCELL_X16 FILLER_18_990 ();
 FILLCELL_X8 FILLER_18_1010 ();
 FILLCELL_X4 FILLER_18_1021 ();
 FILLCELL_X4 FILLER_18_1032 ();
 FILLCELL_X4 FILLER_18_1043 ();
 FILLCELL_X8 FILLER_18_1050 ();
 FILLCELL_X2 FILLER_18_1058 ();
 FILLCELL_X1 FILLER_18_1060 ();
 FILLCELL_X4 FILLER_18_1068 ();
 FILLCELL_X4 FILLER_18_1076 ();
 FILLCELL_X2 FILLER_18_1080 ();
 FILLCELL_X4 FILLER_18_1089 ();
 FILLCELL_X2 FILLER_18_1093 ();
 FILLCELL_X16 FILLER_18_1102 ();
 FILLCELL_X1 FILLER_18_1118 ();
 FILLCELL_X4 FILLER_18_1126 ();
 FILLCELL_X2 FILLER_18_1130 ();
 FILLCELL_X4 FILLER_18_1139 ();
 FILLCELL_X8 FILLER_18_1150 ();
 FILLCELL_X4 FILLER_18_1158 ();
 FILLCELL_X2 FILLER_18_1162 ();
 FILLCELL_X1 FILLER_18_1164 ();
 FILLCELL_X4 FILLER_18_1172 ();
 FILLCELL_X4 FILLER_18_1183 ();
 FILLCELL_X8 FILLER_18_1194 ();
 FILLCELL_X4 FILLER_18_1202 ();
 FILLCELL_X1 FILLER_18_1206 ();
 FILLCELL_X8 FILLER_18_1216 ();
 FILLCELL_X4 FILLER_18_1224 ();
 FILLCELL_X2 FILLER_18_1228 ();
 FILLCELL_X4 FILLER_18_1237 ();
 FILLCELL_X1 FILLER_18_1241 ();
 FILLCELL_X4 FILLER_18_1244 ();
 FILLCELL_X4 FILLER_18_1257 ();
 FILLCELL_X8 FILLER_18_1263 ();
 FILLCELL_X4 FILLER_18_1274 ();
 FILLCELL_X4 FILLER_18_1282 ();
 FILLCELL_X16 FILLER_18_1293 ();
 FILLCELL_X4 FILLER_18_1309 ();
 FILLCELL_X2 FILLER_18_1313 ();
 FILLCELL_X1 FILLER_18_1315 ();
 FILLCELL_X4 FILLER_18_1320 ();
 FILLCELL_X16 FILLER_18_1328 ();
 FILLCELL_X1 FILLER_18_1344 ();
 FILLCELL_X4 FILLER_18_1347 ();
 FILLCELL_X4 FILLER_18_1355 ();
 FILLCELL_X4 FILLER_18_1363 ();
 FILLCELL_X32 FILLER_18_1370 ();
 FILLCELL_X32 FILLER_18_1402 ();
 FILLCELL_X32 FILLER_18_1434 ();
 FILLCELL_X32 FILLER_18_1466 ();
 FILLCELL_X32 FILLER_18_1498 ();
 FILLCELL_X32 FILLER_18_1530 ();
 FILLCELL_X32 FILLER_18_1562 ();
 FILLCELL_X32 FILLER_18_1594 ();
 FILLCELL_X32 FILLER_18_1626 ();
 FILLCELL_X32 FILLER_18_1658 ();
 FILLCELL_X8 FILLER_18_1690 ();
 FILLCELL_X2 FILLER_18_1698 ();
 FILLCELL_X1 FILLER_18_1700 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X32 FILLER_19_193 ();
 FILLCELL_X32 FILLER_19_225 ();
 FILLCELL_X32 FILLER_19_257 ();
 FILLCELL_X32 FILLER_19_289 ();
 FILLCELL_X32 FILLER_19_321 ();
 FILLCELL_X4 FILLER_19_353 ();
 FILLCELL_X8 FILLER_19_376 ();
 FILLCELL_X4 FILLER_19_388 ();
 FILLCELL_X16 FILLER_19_396 ();
 FILLCELL_X8 FILLER_19_412 ();
 FILLCELL_X8 FILLER_19_430 ();
 FILLCELL_X4 FILLER_19_445 ();
 FILLCELL_X4 FILLER_19_459 ();
 FILLCELL_X2 FILLER_19_463 ();
 FILLCELL_X1 FILLER_19_465 ();
 FILLCELL_X4 FILLER_19_473 ();
 FILLCELL_X1 FILLER_19_477 ();
 FILLCELL_X4 FILLER_19_481 ();
 FILLCELL_X4 FILLER_19_490 ();
 FILLCELL_X4 FILLER_19_498 ();
 FILLCELL_X8 FILLER_19_505 ();
 FILLCELL_X1 FILLER_19_513 ();
 FILLCELL_X4 FILLER_19_517 ();
 FILLCELL_X8 FILLER_19_530 ();
 FILLCELL_X1 FILLER_19_538 ();
 FILLCELL_X4 FILLER_19_546 ();
 FILLCELL_X2 FILLER_19_550 ();
 FILLCELL_X1 FILLER_19_552 ();
 FILLCELL_X4 FILLER_19_555 ();
 FILLCELL_X8 FILLER_19_566 ();
 FILLCELL_X2 FILLER_19_574 ();
 FILLCELL_X1 FILLER_19_576 ();
 FILLCELL_X4 FILLER_19_590 ();
 FILLCELL_X2 FILLER_19_594 ();
 FILLCELL_X1 FILLER_19_596 ();
 FILLCELL_X4 FILLER_19_600 ();
 FILLCELL_X8 FILLER_19_606 ();
 FILLCELL_X4 FILLER_19_614 ();
 FILLCELL_X8 FILLER_19_621 ();
 FILLCELL_X4 FILLER_19_629 ();
 FILLCELL_X1 FILLER_19_633 ();
 FILLCELL_X4 FILLER_19_641 ();
 FILLCELL_X2 FILLER_19_645 ();
 FILLCELL_X1 FILLER_19_647 ();
 FILLCELL_X8 FILLER_19_651 ();
 FILLCELL_X2 FILLER_19_659 ();
 FILLCELL_X1 FILLER_19_661 ();
 FILLCELL_X16 FILLER_19_669 ();
 FILLCELL_X2 FILLER_19_685 ();
 FILLCELL_X1 FILLER_19_687 ();
 FILLCELL_X4 FILLER_19_691 ();
 FILLCELL_X4 FILLER_19_698 ();
 FILLCELL_X4 FILLER_19_706 ();
 FILLCELL_X16 FILLER_19_713 ();
 FILLCELL_X2 FILLER_19_729 ();
 FILLCELL_X1 FILLER_19_731 ();
 FILLCELL_X16 FILLER_19_736 ();
 FILLCELL_X8 FILLER_19_752 ();
 FILLCELL_X4 FILLER_19_760 ();
 FILLCELL_X8 FILLER_19_771 ();
 FILLCELL_X4 FILLER_19_779 ();
 FILLCELL_X4 FILLER_19_790 ();
 FILLCELL_X8 FILLER_19_797 ();
 FILLCELL_X2 FILLER_19_805 ();
 FILLCELL_X4 FILLER_19_811 ();
 FILLCELL_X8 FILLER_19_819 ();
 FILLCELL_X4 FILLER_19_827 ();
 FILLCELL_X2 FILLER_19_831 ();
 FILLCELL_X4 FILLER_19_840 ();
 FILLCELL_X16 FILLER_19_851 ();
 FILLCELL_X2 FILLER_19_867 ();
 FILLCELL_X1 FILLER_19_869 ();
 FILLCELL_X8 FILLER_19_874 ();
 FILLCELL_X4 FILLER_19_886 ();
 FILLCELL_X4 FILLER_19_894 ();
 FILLCELL_X1 FILLER_19_898 ();
 FILLCELL_X4 FILLER_19_902 ();
 FILLCELL_X2 FILLER_19_906 ();
 FILLCELL_X4 FILLER_19_917 ();
 FILLCELL_X8 FILLER_19_930 ();
 FILLCELL_X1 FILLER_19_938 ();
 FILLCELL_X4 FILLER_19_942 ();
 FILLCELL_X4 FILLER_19_955 ();
 FILLCELL_X8 FILLER_19_966 ();
 FILLCELL_X1 FILLER_19_974 ();
 FILLCELL_X4 FILLER_19_978 ();
 FILLCELL_X4 FILLER_19_986 ();
 FILLCELL_X8 FILLER_19_993 ();
 FILLCELL_X4 FILLER_19_1001 ();
 FILLCELL_X2 FILLER_19_1005 ();
 FILLCELL_X4 FILLER_19_1010 ();
 FILLCELL_X32 FILLER_19_1017 ();
 FILLCELL_X4 FILLER_19_1053 ();
 FILLCELL_X8 FILLER_19_1061 ();
 FILLCELL_X4 FILLER_19_1073 ();
 FILLCELL_X4 FILLER_19_1081 ();
 FILLCELL_X8 FILLER_19_1089 ();
 FILLCELL_X4 FILLER_19_1104 ();
 FILLCELL_X16 FILLER_19_1115 ();
 FILLCELL_X2 FILLER_19_1131 ();
 FILLCELL_X1 FILLER_19_1133 ();
 FILLCELL_X4 FILLER_19_1141 ();
 FILLCELL_X4 FILLER_19_1152 ();
 FILLCELL_X4 FILLER_19_1163 ();
 FILLCELL_X16 FILLER_19_1174 ();
 FILLCELL_X8 FILLER_19_1190 ();
 FILLCELL_X2 FILLER_19_1198 ();
 FILLCELL_X1 FILLER_19_1200 ();
 FILLCELL_X8 FILLER_19_1226 ();
 FILLCELL_X2 FILLER_19_1234 ();
 FILLCELL_X1 FILLER_19_1236 ();
 FILLCELL_X4 FILLER_19_1239 ();
 FILLCELL_X8 FILLER_19_1254 ();
 FILLCELL_X1 FILLER_19_1262 ();
 FILLCELL_X4 FILLER_19_1264 ();
 FILLCELL_X1 FILLER_19_1268 ();
 FILLCELL_X4 FILLER_19_1273 ();
 FILLCELL_X4 FILLER_19_1281 ();
 FILLCELL_X1 FILLER_19_1285 ();
 FILLCELL_X8 FILLER_19_1289 ();
 FILLCELL_X1 FILLER_19_1297 ();
 FILLCELL_X16 FILLER_19_1300 ();
 FILLCELL_X8 FILLER_19_1316 ();
 FILLCELL_X4 FILLER_19_1324 ();
 FILLCELL_X8 FILLER_19_1330 ();
 FILLCELL_X2 FILLER_19_1338 ();
 FILLCELL_X4 FILLER_19_1342 ();
 FILLCELL_X4 FILLER_19_1353 ();
 FILLCELL_X32 FILLER_19_1359 ();
 FILLCELL_X32 FILLER_19_1391 ();
 FILLCELL_X32 FILLER_19_1423 ();
 FILLCELL_X32 FILLER_19_1455 ();
 FILLCELL_X32 FILLER_19_1487 ();
 FILLCELL_X32 FILLER_19_1519 ();
 FILLCELL_X32 FILLER_19_1551 ();
 FILLCELL_X32 FILLER_19_1583 ();
 FILLCELL_X32 FILLER_19_1615 ();
 FILLCELL_X32 FILLER_19_1647 ();
 FILLCELL_X16 FILLER_19_1679 ();
 FILLCELL_X4 FILLER_19_1695 ();
 FILLCELL_X2 FILLER_19_1699 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X32 FILLER_20_193 ();
 FILLCELL_X32 FILLER_20_225 ();
 FILLCELL_X32 FILLER_20_257 ();
 FILLCELL_X32 FILLER_20_289 ();
 FILLCELL_X32 FILLER_20_321 ();
 FILLCELL_X16 FILLER_20_353 ();
 FILLCELL_X8 FILLER_20_388 ();
 FILLCELL_X1 FILLER_20_396 ();
 FILLCELL_X4 FILLER_20_401 ();
 FILLCELL_X4 FILLER_20_409 ();
 FILLCELL_X8 FILLER_20_415 ();
 FILLCELL_X4 FILLER_20_425 ();
 FILLCELL_X2 FILLER_20_429 ();
 FILLCELL_X1 FILLER_20_431 ();
 FILLCELL_X4 FILLER_20_435 ();
 FILLCELL_X1 FILLER_20_439 ();
 FILLCELL_X8 FILLER_20_449 ();
 FILLCELL_X4 FILLER_20_457 ();
 FILLCELL_X4 FILLER_20_464 ();
 FILLCELL_X1 FILLER_20_468 ();
 FILLCELL_X4 FILLER_20_473 ();
 FILLCELL_X4 FILLER_20_482 ();
 FILLCELL_X8 FILLER_20_492 ();
 FILLCELL_X8 FILLER_20_504 ();
 FILLCELL_X4 FILLER_20_512 ();
 FILLCELL_X1 FILLER_20_516 ();
 FILLCELL_X16 FILLER_20_524 ();
 FILLCELL_X8 FILLER_20_547 ();
 FILLCELL_X1 FILLER_20_555 ();
 FILLCELL_X4 FILLER_20_570 ();
 FILLCELL_X8 FILLER_20_585 ();
 FILLCELL_X2 FILLER_20_593 ();
 FILLCELL_X16 FILLER_20_600 ();
 FILLCELL_X2 FILLER_20_616 ();
 FILLCELL_X1 FILLER_20_618 ();
 FILLCELL_X8 FILLER_20_622 ();
 FILLCELL_X1 FILLER_20_630 ();
 FILLCELL_X8 FILLER_20_632 ();
 FILLCELL_X2 FILLER_20_640 ();
 FILLCELL_X1 FILLER_20_642 ();
 FILLCELL_X8 FILLER_20_650 ();
 FILLCELL_X2 FILLER_20_658 ();
 FILLCELL_X4 FILLER_20_667 ();
 FILLCELL_X4 FILLER_20_678 ();
 FILLCELL_X2 FILLER_20_682 ();
 FILLCELL_X4 FILLER_20_687 ();
 FILLCELL_X8 FILLER_20_700 ();
 FILLCELL_X1 FILLER_20_708 ();
 FILLCELL_X4 FILLER_20_713 ();
 FILLCELL_X1 FILLER_20_717 ();
 FILLCELL_X4 FILLER_20_722 ();
 FILLCELL_X4 FILLER_20_730 ();
 FILLCELL_X4 FILLER_20_741 ();
 FILLCELL_X4 FILLER_20_752 ();
 FILLCELL_X4 FILLER_20_763 ();
 FILLCELL_X4 FILLER_20_774 ();
 FILLCELL_X2 FILLER_20_778 ();
 FILLCELL_X4 FILLER_20_787 ();
 FILLCELL_X16 FILLER_20_798 ();
 FILLCELL_X2 FILLER_20_814 ();
 FILLCELL_X4 FILLER_20_823 ();
 FILLCELL_X8 FILLER_20_834 ();
 FILLCELL_X4 FILLER_20_842 ();
 FILLCELL_X8 FILLER_20_853 ();
 FILLCELL_X8 FILLER_20_868 ();
 FILLCELL_X2 FILLER_20_876 ();
 FILLCELL_X1 FILLER_20_878 ();
 FILLCELL_X4 FILLER_20_886 ();
 FILLCELL_X4 FILLER_20_897 ();
 FILLCELL_X4 FILLER_20_906 ();
 FILLCELL_X4 FILLER_20_915 ();
 FILLCELL_X8 FILLER_20_923 ();
 FILLCELL_X16 FILLER_20_934 ();
 FILLCELL_X2 FILLER_20_950 ();
 FILLCELL_X16 FILLER_20_955 ();
 FILLCELL_X8 FILLER_20_971 ();
 FILLCELL_X1 FILLER_20_979 ();
 FILLCELL_X4 FILLER_20_989 ();
 FILLCELL_X4 FILLER_20_1006 ();
 FILLCELL_X4 FILLER_20_1014 ();
 FILLCELL_X8 FILLER_20_1021 ();
 FILLCELL_X4 FILLER_20_1029 ();
 FILLCELL_X2 FILLER_20_1033 ();
 FILLCELL_X4 FILLER_20_1039 ();
 FILLCELL_X4 FILLER_20_1046 ();
 FILLCELL_X2 FILLER_20_1050 ();
 FILLCELL_X4 FILLER_20_1055 ();
 FILLCELL_X4 FILLER_20_1062 ();
 FILLCELL_X1 FILLER_20_1066 ();
 FILLCELL_X8 FILLER_20_1071 ();
 FILLCELL_X4 FILLER_20_1086 ();
 FILLCELL_X8 FILLER_20_1097 ();
 FILLCELL_X4 FILLER_20_1105 ();
 FILLCELL_X2 FILLER_20_1109 ();
 FILLCELL_X4 FILLER_20_1118 ();
 FILLCELL_X4 FILLER_20_1129 ();
 FILLCELL_X8 FILLER_20_1140 ();
 FILLCELL_X4 FILLER_20_1155 ();
 FILLCELL_X8 FILLER_20_1166 ();
 FILLCELL_X2 FILLER_20_1174 ();
 FILLCELL_X1 FILLER_20_1176 ();
 FILLCELL_X4 FILLER_20_1186 ();
 FILLCELL_X16 FILLER_20_1199 ();
 FILLCELL_X8 FILLER_20_1215 ();
 FILLCELL_X2 FILLER_20_1223 ();
 FILLCELL_X1 FILLER_20_1225 ();
 FILLCELL_X4 FILLER_20_1231 ();
 FILLCELL_X2 FILLER_20_1235 ();
 FILLCELL_X1 FILLER_20_1237 ();
 FILLCELL_X4 FILLER_20_1241 ();
 FILLCELL_X8 FILLER_20_1258 ();
 FILLCELL_X1 FILLER_20_1266 ();
 FILLCELL_X4 FILLER_20_1271 ();
 FILLCELL_X4 FILLER_20_1278 ();
 FILLCELL_X4 FILLER_20_1284 ();
 FILLCELL_X8 FILLER_20_1290 ();
 FILLCELL_X4 FILLER_20_1300 ();
 FILLCELL_X4 FILLER_20_1307 ();
 FILLCELL_X4 FILLER_20_1318 ();
 FILLCELL_X4 FILLER_20_1326 ();
 FILLCELL_X2 FILLER_20_1330 ();
 FILLCELL_X4 FILLER_20_1339 ();
 FILLCELL_X2 FILLER_20_1343 ();
 FILLCELL_X1 FILLER_20_1345 ();
 FILLCELL_X4 FILLER_20_1350 ();
 FILLCELL_X4 FILLER_20_1358 ();
 FILLCELL_X32 FILLER_20_1365 ();
 FILLCELL_X32 FILLER_20_1397 ();
 FILLCELL_X32 FILLER_20_1429 ();
 FILLCELL_X32 FILLER_20_1461 ();
 FILLCELL_X16 FILLER_20_1493 ();
 FILLCELL_X8 FILLER_20_1509 ();
 FILLCELL_X2 FILLER_20_1517 ();
 FILLCELL_X1 FILLER_20_1519 ();
 FILLCELL_X32 FILLER_20_1537 ();
 FILLCELL_X32 FILLER_20_1569 ();
 FILLCELL_X32 FILLER_20_1601 ();
 FILLCELL_X32 FILLER_20_1633 ();
 FILLCELL_X16 FILLER_20_1665 ();
 FILLCELL_X8 FILLER_20_1681 ();
 FILLCELL_X4 FILLER_20_1689 ();
 FILLCELL_X1 FILLER_20_1693 ();
 FILLCELL_X4 FILLER_20_1697 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X32 FILLER_21_193 ();
 FILLCELL_X32 FILLER_21_225 ();
 FILLCELL_X32 FILLER_21_257 ();
 FILLCELL_X32 FILLER_21_289 ();
 FILLCELL_X32 FILLER_21_321 ();
 FILLCELL_X32 FILLER_21_353 ();
 FILLCELL_X16 FILLER_21_385 ();
 FILLCELL_X4 FILLER_21_401 ();
 FILLCELL_X4 FILLER_21_408 ();
 FILLCELL_X32 FILLER_21_429 ();
 FILLCELL_X8 FILLER_21_465 ();
 FILLCELL_X4 FILLER_21_476 ();
 FILLCELL_X1 FILLER_21_480 ();
 FILLCELL_X4 FILLER_21_485 ();
 FILLCELL_X8 FILLER_21_492 ();
 FILLCELL_X4 FILLER_21_500 ();
 FILLCELL_X1 FILLER_21_504 ();
 FILLCELL_X4 FILLER_21_508 ();
 FILLCELL_X4 FILLER_21_521 ();
 FILLCELL_X4 FILLER_21_532 ();
 FILLCELL_X2 FILLER_21_536 ();
 FILLCELL_X1 FILLER_21_538 ();
 FILLCELL_X32 FILLER_21_543 ();
 FILLCELL_X1 FILLER_21_575 ();
 FILLCELL_X4 FILLER_21_583 ();
 FILLCELL_X4 FILLER_21_590 ();
 FILLCELL_X4 FILLER_21_599 ();
 FILLCELL_X4 FILLER_21_608 ();
 FILLCELL_X4 FILLER_21_616 ();
 FILLCELL_X4 FILLER_21_623 ();
 FILLCELL_X2 FILLER_21_627 ();
 FILLCELL_X1 FILLER_21_629 ();
 FILLCELL_X4 FILLER_21_633 ();
 FILLCELL_X4 FILLER_21_642 ();
 FILLCELL_X4 FILLER_21_649 ();
 FILLCELL_X2 FILLER_21_653 ();
 FILLCELL_X1 FILLER_21_655 ();
 FILLCELL_X4 FILLER_21_660 ();
 FILLCELL_X4 FILLER_21_667 ();
 FILLCELL_X4 FILLER_21_674 ();
 FILLCELL_X2 FILLER_21_678 ();
 FILLCELL_X1 FILLER_21_680 ();
 FILLCELL_X8 FILLER_21_685 ();
 FILLCELL_X4 FILLER_21_696 ();
 FILLCELL_X8 FILLER_21_703 ();
 FILLCELL_X8 FILLER_21_718 ();
 FILLCELL_X2 FILLER_21_726 ();
 FILLCELL_X4 FILLER_21_731 ();
 FILLCELL_X4 FILLER_21_738 ();
 FILLCELL_X8 FILLER_21_746 ();
 FILLCELL_X4 FILLER_21_754 ();
 FILLCELL_X1 FILLER_21_758 ();
 FILLCELL_X8 FILLER_21_766 ();
 FILLCELL_X2 FILLER_21_774 ();
 FILLCELL_X1 FILLER_21_776 ();
 FILLCELL_X4 FILLER_21_784 ();
 FILLCELL_X16 FILLER_21_791 ();
 FILLCELL_X1 FILLER_21_807 ();
 FILLCELL_X8 FILLER_21_815 ();
 FILLCELL_X2 FILLER_21_823 ();
 FILLCELL_X4 FILLER_21_832 ();
 FILLCELL_X2 FILLER_21_836 ();
 FILLCELL_X1 FILLER_21_838 ();
 FILLCELL_X8 FILLER_21_846 ();
 FILLCELL_X4 FILLER_21_861 ();
 FILLCELL_X8 FILLER_21_872 ();
 FILLCELL_X4 FILLER_21_887 ();
 FILLCELL_X16 FILLER_21_894 ();
 FILLCELL_X1 FILLER_21_910 ();
 FILLCELL_X4 FILLER_21_914 ();
 FILLCELL_X4 FILLER_21_921 ();
 FILLCELL_X2 FILLER_21_925 ();
 FILLCELL_X1 FILLER_21_927 ();
 FILLCELL_X16 FILLER_21_935 ();
 FILLCELL_X2 FILLER_21_951 ();
 FILLCELL_X8 FILLER_21_957 ();
 FILLCELL_X4 FILLER_21_970 ();
 FILLCELL_X4 FILLER_21_978 ();
 FILLCELL_X4 FILLER_21_985 ();
 FILLCELL_X4 FILLER_21_992 ();
 FILLCELL_X8 FILLER_21_999 ();
 FILLCELL_X1 FILLER_21_1007 ();
 FILLCELL_X4 FILLER_21_1017 ();
 FILLCELL_X4 FILLER_21_1034 ();
 FILLCELL_X4 FILLER_21_1045 ();
 FILLCELL_X8 FILLER_21_1053 ();
 FILLCELL_X4 FILLER_21_1061 ();
 FILLCELL_X4 FILLER_21_1069 ();
 FILLCELL_X4 FILLER_21_1080 ();
 FILLCELL_X8 FILLER_21_1087 ();
 FILLCELL_X4 FILLER_21_1095 ();
 FILLCELL_X1 FILLER_21_1099 ();
 FILLCELL_X8 FILLER_21_1107 ();
 FILLCELL_X4 FILLER_21_1115 ();
 FILLCELL_X1 FILLER_21_1119 ();
 FILLCELL_X8 FILLER_21_1127 ();
 FILLCELL_X2 FILLER_21_1135 ();
 FILLCELL_X4 FILLER_21_1146 ();
 FILLCELL_X8 FILLER_21_1157 ();
 FILLCELL_X4 FILLER_21_1165 ();
 FILLCELL_X1 FILLER_21_1169 ();
 FILLCELL_X4 FILLER_21_1179 ();
 FILLCELL_X16 FILLER_21_1192 ();
 FILLCELL_X1 FILLER_21_1208 ();
 FILLCELL_X4 FILLER_21_1211 ();
 FILLCELL_X8 FILLER_21_1219 ();
 FILLCELL_X4 FILLER_21_1236 ();
 FILLCELL_X8 FILLER_21_1250 ();
 FILLCELL_X4 FILLER_21_1258 ();
 FILLCELL_X1 FILLER_21_1262 ();
 FILLCELL_X4 FILLER_21_1264 ();
 FILLCELL_X4 FILLER_21_1272 ();
 FILLCELL_X8 FILLER_21_1278 ();
 FILLCELL_X4 FILLER_21_1290 ();
 FILLCELL_X4 FILLER_21_1298 ();
 FILLCELL_X4 FILLER_21_1306 ();
 FILLCELL_X4 FILLER_21_1314 ();
 FILLCELL_X1 FILLER_21_1318 ();
 FILLCELL_X4 FILLER_21_1323 ();
 FILLCELL_X4 FILLER_21_1331 ();
 FILLCELL_X1 FILLER_21_1335 ();
 FILLCELL_X4 FILLER_21_1340 ();
 FILLCELL_X4 FILLER_21_1348 ();
 FILLCELL_X32 FILLER_21_1354 ();
 FILLCELL_X32 FILLER_21_1386 ();
 FILLCELL_X32 FILLER_21_1418 ();
 FILLCELL_X32 FILLER_21_1450 ();
 FILLCELL_X32 FILLER_21_1482 ();
 FILLCELL_X32 FILLER_21_1514 ();
 FILLCELL_X32 FILLER_21_1546 ();
 FILLCELL_X32 FILLER_21_1578 ();
 FILLCELL_X32 FILLER_21_1610 ();
 FILLCELL_X32 FILLER_21_1642 ();
 FILLCELL_X16 FILLER_21_1674 ();
 FILLCELL_X8 FILLER_21_1690 ();
 FILLCELL_X2 FILLER_21_1698 ();
 FILLCELL_X1 FILLER_21_1700 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X32 FILLER_22_193 ();
 FILLCELL_X32 FILLER_22_225 ();
 FILLCELL_X32 FILLER_22_257 ();
 FILLCELL_X32 FILLER_22_289 ();
 FILLCELL_X32 FILLER_22_321 ();
 FILLCELL_X32 FILLER_22_353 ();
 FILLCELL_X16 FILLER_22_385 ();
 FILLCELL_X2 FILLER_22_401 ();
 FILLCELL_X1 FILLER_22_403 ();
 FILLCELL_X4 FILLER_22_408 ();
 FILLCELL_X8 FILLER_22_416 ();
 FILLCELL_X1 FILLER_22_424 ();
 FILLCELL_X4 FILLER_22_429 ();
 FILLCELL_X4 FILLER_22_443 ();
 FILLCELL_X2 FILLER_22_447 ();
 FILLCELL_X1 FILLER_22_449 ();
 FILLCELL_X4 FILLER_22_453 ();
 FILLCELL_X4 FILLER_22_461 ();
 FILLCELL_X4 FILLER_22_470 ();
 FILLCELL_X8 FILLER_22_479 ();
 FILLCELL_X1 FILLER_22_487 ();
 FILLCELL_X4 FILLER_22_497 ();
 FILLCELL_X4 FILLER_22_505 ();
 FILLCELL_X8 FILLER_22_516 ();
 FILLCELL_X8 FILLER_22_528 ();
 FILLCELL_X1 FILLER_22_536 ();
 FILLCELL_X8 FILLER_22_547 ();
 FILLCELL_X4 FILLER_22_555 ();
 FILLCELL_X1 FILLER_22_559 ();
 FILLCELL_X8 FILLER_22_562 ();
 FILLCELL_X4 FILLER_22_570 ();
 FILLCELL_X2 FILLER_22_574 ();
 FILLCELL_X4 FILLER_22_583 ();
 FILLCELL_X2 FILLER_22_587 ();
 FILLCELL_X1 FILLER_22_589 ();
 FILLCELL_X8 FILLER_22_594 ();
 FILLCELL_X8 FILLER_22_608 ();
 FILLCELL_X1 FILLER_22_616 ();
 FILLCELL_X4 FILLER_22_626 ();
 FILLCELL_X1 FILLER_22_630 ();
 FILLCELL_X4 FILLER_22_632 ();
 FILLCELL_X8 FILLER_22_643 ();
 FILLCELL_X8 FILLER_22_657 ();
 FILLCELL_X2 FILLER_22_665 ();
 FILLCELL_X16 FILLER_22_670 ();
 FILLCELL_X1 FILLER_22_686 ();
 FILLCELL_X4 FILLER_22_694 ();
 FILLCELL_X2 FILLER_22_698 ();
 FILLCELL_X4 FILLER_22_703 ();
 FILLCELL_X4 FILLER_22_710 ();
 FILLCELL_X4 FILLER_22_717 ();
 FILLCELL_X4 FILLER_22_724 ();
 FILLCELL_X8 FILLER_22_735 ();
 FILLCELL_X1 FILLER_22_743 ();
 FILLCELL_X4 FILLER_22_748 ();
 FILLCELL_X4 FILLER_22_759 ();
 FILLCELL_X16 FILLER_22_770 ();
 FILLCELL_X8 FILLER_22_786 ();
 FILLCELL_X2 FILLER_22_794 ();
 FILLCELL_X1 FILLER_22_796 ();
 FILLCELL_X4 FILLER_22_800 ();
 FILLCELL_X4 FILLER_22_814 ();
 FILLCELL_X4 FILLER_22_821 ();
 FILLCELL_X2 FILLER_22_825 ();
 FILLCELL_X1 FILLER_22_827 ();
 FILLCELL_X8 FILLER_22_837 ();
 FILLCELL_X4 FILLER_22_845 ();
 FILLCELL_X2 FILLER_22_849 ();
 FILLCELL_X16 FILLER_22_858 ();
 FILLCELL_X8 FILLER_22_874 ();
 FILLCELL_X2 FILLER_22_882 ();
 FILLCELL_X4 FILLER_22_891 ();
 FILLCELL_X2 FILLER_22_895 ();
 FILLCELL_X1 FILLER_22_897 ();
 FILLCELL_X4 FILLER_22_901 ();
 FILLCELL_X4 FILLER_22_909 ();
 FILLCELL_X2 FILLER_22_913 ();
 FILLCELL_X1 FILLER_22_915 ();
 FILLCELL_X8 FILLER_22_920 ();
 FILLCELL_X8 FILLER_22_934 ();
 FILLCELL_X4 FILLER_22_949 ();
 FILLCELL_X2 FILLER_22_953 ();
 FILLCELL_X4 FILLER_22_964 ();
 FILLCELL_X4 FILLER_22_974 ();
 FILLCELL_X1 FILLER_22_978 ();
 FILLCELL_X8 FILLER_22_988 ();
 FILLCELL_X1 FILLER_22_996 ();
 FILLCELL_X4 FILLER_22_1001 ();
 FILLCELL_X4 FILLER_22_1012 ();
 FILLCELL_X4 FILLER_22_1019 ();
 FILLCELL_X2 FILLER_22_1023 ();
 FILLCELL_X1 FILLER_22_1025 ();
 FILLCELL_X4 FILLER_22_1030 ();
 FILLCELL_X16 FILLER_22_1037 ();
 FILLCELL_X8 FILLER_22_1057 ();
 FILLCELL_X4 FILLER_22_1069 ();
 FILLCELL_X2 FILLER_22_1073 ();
 FILLCELL_X4 FILLER_22_1082 ();
 FILLCELL_X4 FILLER_22_1089 ();
 FILLCELL_X4 FILLER_22_1100 ();
 FILLCELL_X4 FILLER_22_1111 ();
 FILLCELL_X8 FILLER_22_1122 ();
 FILLCELL_X4 FILLER_22_1130 ();
 FILLCELL_X2 FILLER_22_1134 ();
 FILLCELL_X16 FILLER_22_1145 ();
 FILLCELL_X1 FILLER_22_1161 ();
 FILLCELL_X16 FILLER_22_1171 ();
 FILLCELL_X4 FILLER_22_1187 ();
 FILLCELL_X1 FILLER_22_1191 ();
 FILLCELL_X4 FILLER_22_1195 ();
 FILLCELL_X4 FILLER_22_1203 ();
 FILLCELL_X4 FILLER_22_1213 ();
 FILLCELL_X2 FILLER_22_1217 ();
 FILLCELL_X1 FILLER_22_1219 ();
 FILLCELL_X4 FILLER_22_1224 ();
 FILLCELL_X1 FILLER_22_1228 ();
 FILLCELL_X4 FILLER_22_1232 ();
 FILLCELL_X16 FILLER_22_1238 ();
 FILLCELL_X8 FILLER_22_1254 ();
 FILLCELL_X4 FILLER_22_1266 ();
 FILLCELL_X4 FILLER_22_1274 ();
 FILLCELL_X4 FILLER_22_1282 ();
 FILLCELL_X8 FILLER_22_1289 ();
 FILLCELL_X2 FILLER_22_1297 ();
 FILLCELL_X1 FILLER_22_1299 ();
 FILLCELL_X4 FILLER_22_1302 ();
 FILLCELL_X4 FILLER_22_1308 ();
 FILLCELL_X2 FILLER_22_1312 ();
 FILLCELL_X4 FILLER_22_1317 ();
 FILLCELL_X4 FILLER_22_1323 ();
 FILLCELL_X1 FILLER_22_1327 ();
 FILLCELL_X4 FILLER_22_1330 ();
 FILLCELL_X32 FILLER_22_1337 ();
 FILLCELL_X32 FILLER_22_1369 ();
 FILLCELL_X32 FILLER_22_1401 ();
 FILLCELL_X32 FILLER_22_1433 ();
 FILLCELL_X32 FILLER_22_1465 ();
 FILLCELL_X8 FILLER_22_1497 ();
 FILLCELL_X4 FILLER_22_1505 ();
 FILLCELL_X32 FILLER_22_1513 ();
 FILLCELL_X32 FILLER_22_1545 ();
 FILLCELL_X32 FILLER_22_1577 ();
 FILLCELL_X32 FILLER_22_1609 ();
 FILLCELL_X32 FILLER_22_1641 ();
 FILLCELL_X16 FILLER_22_1673 ();
 FILLCELL_X8 FILLER_22_1689 ();
 FILLCELL_X4 FILLER_22_1697 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X32 FILLER_23_193 ();
 FILLCELL_X32 FILLER_23_225 ();
 FILLCELL_X32 FILLER_23_257 ();
 FILLCELL_X32 FILLER_23_289 ();
 FILLCELL_X32 FILLER_23_321 ();
 FILLCELL_X16 FILLER_23_353 ();
 FILLCELL_X4 FILLER_23_369 ();
 FILLCELL_X1 FILLER_23_373 ();
 FILLCELL_X4 FILLER_23_378 ();
 FILLCELL_X16 FILLER_23_401 ();
 FILLCELL_X1 FILLER_23_417 ();
 FILLCELL_X4 FILLER_23_421 ();
 FILLCELL_X4 FILLER_23_429 ();
 FILLCELL_X4 FILLER_23_436 ();
 FILLCELL_X4 FILLER_23_450 ();
 FILLCELL_X4 FILLER_23_464 ();
 FILLCELL_X8 FILLER_23_472 ();
 FILLCELL_X4 FILLER_23_480 ();
 FILLCELL_X4 FILLER_23_491 ();
 FILLCELL_X4 FILLER_23_499 ();
 FILLCELL_X4 FILLER_23_506 ();
 FILLCELL_X2 FILLER_23_510 ();
 FILLCELL_X4 FILLER_23_522 ();
 FILLCELL_X4 FILLER_23_528 ();
 FILLCELL_X1 FILLER_23_532 ();
 FILLCELL_X8 FILLER_23_542 ();
 FILLCELL_X2 FILLER_23_550 ();
 FILLCELL_X1 FILLER_23_552 ();
 FILLCELL_X4 FILLER_23_560 ();
 FILLCELL_X4 FILLER_23_573 ();
 FILLCELL_X2 FILLER_23_577 ();
 FILLCELL_X1 FILLER_23_579 ();
 FILLCELL_X4 FILLER_23_583 ();
 FILLCELL_X4 FILLER_23_597 ();
 FILLCELL_X4 FILLER_23_605 ();
 FILLCELL_X1 FILLER_23_609 ();
 FILLCELL_X16 FILLER_23_614 ();
 FILLCELL_X2 FILLER_23_630 ();
 FILLCELL_X4 FILLER_23_641 ();
 FILLCELL_X4 FILLER_23_647 ();
 FILLCELL_X8 FILLER_23_661 ();
 FILLCELL_X1 FILLER_23_669 ();
 FILLCELL_X4 FILLER_23_673 ();
 FILLCELL_X4 FILLER_23_687 ();
 FILLCELL_X2 FILLER_23_691 ();
 FILLCELL_X4 FILLER_23_697 ();
 FILLCELL_X4 FILLER_23_708 ();
 FILLCELL_X4 FILLER_23_717 ();
 FILLCELL_X4 FILLER_23_725 ();
 FILLCELL_X4 FILLER_23_732 ();
 FILLCELL_X4 FILLER_23_740 ();
 FILLCELL_X8 FILLER_23_747 ();
 FILLCELL_X4 FILLER_23_755 ();
 FILLCELL_X2 FILLER_23_759 ();
 FILLCELL_X4 FILLER_23_768 ();
 FILLCELL_X4 FILLER_23_776 ();
 FILLCELL_X4 FILLER_23_787 ();
 FILLCELL_X4 FILLER_23_798 ();
 FILLCELL_X4 FILLER_23_807 ();
 FILLCELL_X2 FILLER_23_811 ();
 FILLCELL_X8 FILLER_23_823 ();
 FILLCELL_X1 FILLER_23_831 ();
 FILLCELL_X8 FILLER_23_841 ();
 FILLCELL_X2 FILLER_23_849 ();
 FILLCELL_X1 FILLER_23_851 ();
 FILLCELL_X8 FILLER_23_861 ();
 FILLCELL_X4 FILLER_23_869 ();
 FILLCELL_X2 FILLER_23_873 ();
 FILLCELL_X4 FILLER_23_882 ();
 FILLCELL_X2 FILLER_23_886 ();
 FILLCELL_X1 FILLER_23_888 ();
 FILLCELL_X4 FILLER_23_896 ();
 FILLCELL_X2 FILLER_23_900 ();
 FILLCELL_X1 FILLER_23_902 ();
 FILLCELL_X4 FILLER_23_907 ();
 FILLCELL_X8 FILLER_23_918 ();
 FILLCELL_X2 FILLER_23_926 ();
 FILLCELL_X1 FILLER_23_928 ();
 FILLCELL_X4 FILLER_23_932 ();
 FILLCELL_X4 FILLER_23_940 ();
 FILLCELL_X4 FILLER_23_947 ();
 FILLCELL_X2 FILLER_23_951 ();
 FILLCELL_X1 FILLER_23_953 ();
 FILLCELL_X8 FILLER_23_959 ();
 FILLCELL_X1 FILLER_23_967 ();
 FILLCELL_X8 FILLER_23_971 ();
 FILLCELL_X1 FILLER_23_979 ();
 FILLCELL_X4 FILLER_23_987 ();
 FILLCELL_X4 FILLER_23_996 ();
 FILLCELL_X8 FILLER_23_1004 ();
 FILLCELL_X2 FILLER_23_1012 ();
 FILLCELL_X4 FILLER_23_1018 ();
 FILLCELL_X2 FILLER_23_1022 ();
 FILLCELL_X4 FILLER_23_1028 ();
 FILLCELL_X8 FILLER_23_1036 ();
 FILLCELL_X2 FILLER_23_1044 ();
 FILLCELL_X1 FILLER_23_1046 ();
 FILLCELL_X4 FILLER_23_1052 ();
 FILLCELL_X4 FILLER_23_1061 ();
 FILLCELL_X16 FILLER_23_1068 ();
 FILLCELL_X4 FILLER_23_1091 ();
 FILLCELL_X16 FILLER_23_1102 ();
 FILLCELL_X4 FILLER_23_1118 ();
 FILLCELL_X1 FILLER_23_1122 ();
 FILLCELL_X16 FILLER_23_1132 ();
 FILLCELL_X4 FILLER_23_1148 ();
 FILLCELL_X2 FILLER_23_1152 ();
 FILLCELL_X4 FILLER_23_1156 ();
 FILLCELL_X4 FILLER_23_1163 ();
 FILLCELL_X4 FILLER_23_1170 ();
 FILLCELL_X2 FILLER_23_1174 ();
 FILLCELL_X8 FILLER_23_1182 ();
 FILLCELL_X1 FILLER_23_1190 ();
 FILLCELL_X4 FILLER_23_1197 ();
 FILLCELL_X8 FILLER_23_1203 ();
 FILLCELL_X2 FILLER_23_1211 ();
 FILLCELL_X8 FILLER_23_1218 ();
 FILLCELL_X2 FILLER_23_1226 ();
 FILLCELL_X1 FILLER_23_1228 ();
 FILLCELL_X4 FILLER_23_1238 ();
 FILLCELL_X16 FILLER_23_1246 ();
 FILLCELL_X1 FILLER_23_1262 ();
 FILLCELL_X4 FILLER_23_1264 ();
 FILLCELL_X4 FILLER_23_1272 ();
 FILLCELL_X4 FILLER_23_1278 ();
 FILLCELL_X2 FILLER_23_1282 ();
 FILLCELL_X4 FILLER_23_1287 ();
 FILLCELL_X4 FILLER_23_1293 ();
 FILLCELL_X4 FILLER_23_1299 ();
 FILLCELL_X2 FILLER_23_1303 ();
 FILLCELL_X8 FILLER_23_1309 ();
 FILLCELL_X4 FILLER_23_1317 ();
 FILLCELL_X2 FILLER_23_1321 ();
 FILLCELL_X1 FILLER_23_1323 ();
 FILLCELL_X4 FILLER_23_1328 ();
 FILLCELL_X2 FILLER_23_1332 ();
 FILLCELL_X4 FILLER_23_1337 ();
 FILLCELL_X32 FILLER_23_1344 ();
 FILLCELL_X32 FILLER_23_1376 ();
 FILLCELL_X32 FILLER_23_1408 ();
 FILLCELL_X32 FILLER_23_1440 ();
 FILLCELL_X32 FILLER_23_1472 ();
 FILLCELL_X32 FILLER_23_1504 ();
 FILLCELL_X32 FILLER_23_1536 ();
 FILLCELL_X32 FILLER_23_1568 ();
 FILLCELL_X32 FILLER_23_1600 ();
 FILLCELL_X32 FILLER_23_1632 ();
 FILLCELL_X32 FILLER_23_1664 ();
 FILLCELL_X4 FILLER_23_1696 ();
 FILLCELL_X1 FILLER_23_1700 ();
 FILLCELL_X4 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_8 ();
 FILLCELL_X32 FILLER_24_40 ();
 FILLCELL_X32 FILLER_24_72 ();
 FILLCELL_X32 FILLER_24_104 ();
 FILLCELL_X32 FILLER_24_136 ();
 FILLCELL_X32 FILLER_24_168 ();
 FILLCELL_X32 FILLER_24_200 ();
 FILLCELL_X32 FILLER_24_232 ();
 FILLCELL_X32 FILLER_24_264 ();
 FILLCELL_X32 FILLER_24_296 ();
 FILLCELL_X32 FILLER_24_328 ();
 FILLCELL_X32 FILLER_24_360 ();
 FILLCELL_X8 FILLER_24_392 ();
 FILLCELL_X4 FILLER_24_400 ();
 FILLCELL_X2 FILLER_24_404 ();
 FILLCELL_X8 FILLER_24_410 ();
 FILLCELL_X4 FILLER_24_418 ();
 FILLCELL_X1 FILLER_24_422 ();
 FILLCELL_X4 FILLER_24_426 ();
 FILLCELL_X4 FILLER_24_437 ();
 FILLCELL_X2 FILLER_24_441 ();
 FILLCELL_X16 FILLER_24_446 ();
 FILLCELL_X1 FILLER_24_462 ();
 FILLCELL_X8 FILLER_24_472 ();
 FILLCELL_X4 FILLER_24_480 ();
 FILLCELL_X1 FILLER_24_484 ();
 FILLCELL_X4 FILLER_24_494 ();
 FILLCELL_X4 FILLER_24_502 ();
 FILLCELL_X2 FILLER_24_506 ();
 FILLCELL_X4 FILLER_24_512 ();
 FILLCELL_X1 FILLER_24_516 ();
 FILLCELL_X4 FILLER_24_520 ();
 FILLCELL_X16 FILLER_24_527 ();
 FILLCELL_X1 FILLER_24_543 ();
 FILLCELL_X8 FILLER_24_551 ();
 FILLCELL_X1 FILLER_24_559 ();
 FILLCELL_X4 FILLER_24_570 ();
 FILLCELL_X1 FILLER_24_574 ();
 FILLCELL_X8 FILLER_24_578 ();
 FILLCELL_X4 FILLER_24_589 ();
 FILLCELL_X2 FILLER_24_593 ();
 FILLCELL_X4 FILLER_24_602 ();
 FILLCELL_X2 FILLER_24_606 ();
 FILLCELL_X4 FILLER_24_611 ();
 FILLCELL_X8 FILLER_24_618 ();
 FILLCELL_X4 FILLER_24_626 ();
 FILLCELL_X1 FILLER_24_630 ();
 FILLCELL_X4 FILLER_24_632 ();
 FILLCELL_X8 FILLER_24_643 ();
 FILLCELL_X8 FILLER_24_655 ();
 FILLCELL_X2 FILLER_24_663 ();
 FILLCELL_X1 FILLER_24_665 ();
 FILLCELL_X4 FILLER_24_676 ();
 FILLCELL_X4 FILLER_24_684 ();
 FILLCELL_X16 FILLER_24_698 ();
 FILLCELL_X1 FILLER_24_714 ();
 FILLCELL_X4 FILLER_24_718 ();
 FILLCELL_X4 FILLER_24_727 ();
 FILLCELL_X2 FILLER_24_731 ();
 FILLCELL_X1 FILLER_24_733 ();
 FILLCELL_X4 FILLER_24_741 ();
 FILLCELL_X32 FILLER_24_749 ();
 FILLCELL_X4 FILLER_24_784 ();
 FILLCELL_X2 FILLER_24_788 ();
 FILLCELL_X4 FILLER_24_799 ();
 FILLCELL_X2 FILLER_24_803 ();
 FILLCELL_X1 FILLER_24_805 ();
 FILLCELL_X4 FILLER_24_813 ();
 FILLCELL_X8 FILLER_24_819 ();
 FILLCELL_X4 FILLER_24_827 ();
 FILLCELL_X2 FILLER_24_831 ();
 FILLCELL_X1 FILLER_24_833 ();
 FILLCELL_X8 FILLER_24_844 ();
 FILLCELL_X1 FILLER_24_852 ();
 FILLCELL_X4 FILLER_24_863 ();
 FILLCELL_X4 FILLER_24_877 ();
 FILLCELL_X16 FILLER_24_884 ();
 FILLCELL_X4 FILLER_24_900 ();
 FILLCELL_X1 FILLER_24_904 ();
 FILLCELL_X4 FILLER_24_912 ();
 FILLCELL_X2 FILLER_24_916 ();
 FILLCELL_X1 FILLER_24_918 ();
 FILLCELL_X4 FILLER_24_926 ();
 FILLCELL_X1 FILLER_24_930 ();
 FILLCELL_X8 FILLER_24_944 ();
 FILLCELL_X4 FILLER_24_958 ();
 FILLCELL_X8 FILLER_24_968 ();
 FILLCELL_X1 FILLER_24_976 ();
 FILLCELL_X4 FILLER_24_986 ();
 FILLCELL_X1 FILLER_24_990 ();
 FILLCELL_X4 FILLER_24_1004 ();
 FILLCELL_X4 FILLER_24_1022 ();
 FILLCELL_X4 FILLER_24_1033 ();
 FILLCELL_X4 FILLER_24_1044 ();
 FILLCELL_X4 FILLER_24_1052 ();
 FILLCELL_X4 FILLER_24_1059 ();
 FILLCELL_X2 FILLER_24_1063 ();
 FILLCELL_X1 FILLER_24_1065 ();
 FILLCELL_X8 FILLER_24_1069 ();
 FILLCELL_X4 FILLER_24_1084 ();
 FILLCELL_X16 FILLER_24_1095 ();
 FILLCELL_X4 FILLER_24_1111 ();
 FILLCELL_X2 FILLER_24_1115 ();
 FILLCELL_X1 FILLER_24_1117 ();
 FILLCELL_X4 FILLER_24_1127 ();
 FILLCELL_X8 FILLER_24_1133 ();
 FILLCELL_X4 FILLER_24_1141 ();
 FILLCELL_X2 FILLER_24_1145 ();
 FILLCELL_X1 FILLER_24_1147 ();
 FILLCELL_X4 FILLER_24_1154 ();
 FILLCELL_X4 FILLER_24_1162 ();
 FILLCELL_X4 FILLER_24_1170 ();
 FILLCELL_X2 FILLER_24_1174 ();
 FILLCELL_X1 FILLER_24_1176 ();
 FILLCELL_X4 FILLER_24_1180 ();
 FILLCELL_X2 FILLER_24_1184 ();
 FILLCELL_X1 FILLER_24_1186 ();
 FILLCELL_X4 FILLER_24_1190 ();
 FILLCELL_X4 FILLER_24_1199 ();
 FILLCELL_X4 FILLER_24_1207 ();
 FILLCELL_X8 FILLER_24_1214 ();
 FILLCELL_X2 FILLER_24_1222 ();
 FILLCELL_X4 FILLER_24_1229 ();
 FILLCELL_X8 FILLER_24_1237 ();
 FILLCELL_X2 FILLER_24_1245 ();
 FILLCELL_X4 FILLER_24_1253 ();
 FILLCELL_X4 FILLER_24_1263 ();
 FILLCELL_X2 FILLER_24_1267 ();
 FILLCELL_X4 FILLER_24_1273 ();
 FILLCELL_X8 FILLER_24_1281 ();
 FILLCELL_X8 FILLER_24_1303 ();
 FILLCELL_X4 FILLER_24_1315 ();
 FILLCELL_X4 FILLER_24_1321 ();
 FILLCELL_X1 FILLER_24_1325 ();
 FILLCELL_X4 FILLER_24_1329 ();
 FILLCELL_X4 FILLER_24_1335 ();
 FILLCELL_X4 FILLER_24_1341 ();
 FILLCELL_X32 FILLER_24_1347 ();
 FILLCELL_X1 FILLER_24_1379 ();
 FILLCELL_X4 FILLER_24_1385 ();
 FILLCELL_X32 FILLER_24_1392 ();
 FILLCELL_X32 FILLER_24_1424 ();
 FILLCELL_X32 FILLER_24_1456 ();
 FILLCELL_X32 FILLER_24_1488 ();
 FILLCELL_X32 FILLER_24_1520 ();
 FILLCELL_X32 FILLER_24_1552 ();
 FILLCELL_X32 FILLER_24_1584 ();
 FILLCELL_X32 FILLER_24_1616 ();
 FILLCELL_X32 FILLER_24_1648 ();
 FILLCELL_X16 FILLER_24_1680 ();
 FILLCELL_X4 FILLER_24_1696 ();
 FILLCELL_X1 FILLER_24_1700 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X32 FILLER_25_193 ();
 FILLCELL_X32 FILLER_25_225 ();
 FILLCELL_X32 FILLER_25_257 ();
 FILLCELL_X32 FILLER_25_289 ();
 FILLCELL_X32 FILLER_25_321 ();
 FILLCELL_X8 FILLER_25_353 ();
 FILLCELL_X32 FILLER_25_378 ();
 FILLCELL_X16 FILLER_25_410 ();
 FILLCELL_X2 FILLER_25_426 ();
 FILLCELL_X1 FILLER_25_428 ();
 FILLCELL_X4 FILLER_25_438 ();
 FILLCELL_X2 FILLER_25_442 ();
 FILLCELL_X1 FILLER_25_444 ();
 FILLCELL_X4 FILLER_25_447 ();
 FILLCELL_X4 FILLER_25_455 ();
 FILLCELL_X8 FILLER_25_465 ();
 FILLCELL_X1 FILLER_25_473 ();
 FILLCELL_X4 FILLER_25_481 ();
 FILLCELL_X1 FILLER_25_485 ();
 FILLCELL_X8 FILLER_25_496 ();
 FILLCELL_X4 FILLER_25_504 ();
 FILLCELL_X4 FILLER_25_513 ();
 FILLCELL_X2 FILLER_25_517 ();
 FILLCELL_X1 FILLER_25_519 ();
 FILLCELL_X4 FILLER_25_523 ();
 FILLCELL_X8 FILLER_25_537 ();
 FILLCELL_X4 FILLER_25_545 ();
 FILLCELL_X1 FILLER_25_549 ();
 FILLCELL_X4 FILLER_25_554 ();
 FILLCELL_X8 FILLER_25_562 ();
 FILLCELL_X4 FILLER_25_570 ();
 FILLCELL_X2 FILLER_25_574 ();
 FILLCELL_X4 FILLER_25_585 ();
 FILLCELL_X2 FILLER_25_589 ();
 FILLCELL_X1 FILLER_25_591 ();
 FILLCELL_X4 FILLER_25_597 ();
 FILLCELL_X4 FILLER_25_606 ();
 FILLCELL_X4 FILLER_25_620 ();
 FILLCELL_X8 FILLER_25_634 ();
 FILLCELL_X1 FILLER_25_642 ();
 FILLCELL_X4 FILLER_25_648 ();
 FILLCELL_X4 FILLER_25_661 ();
 FILLCELL_X2 FILLER_25_665 ();
 FILLCELL_X4 FILLER_25_670 ();
 FILLCELL_X4 FILLER_25_677 ();
 FILLCELL_X2 FILLER_25_681 ();
 FILLCELL_X8 FILLER_25_686 ();
 FILLCELL_X8 FILLER_25_703 ();
 FILLCELL_X4 FILLER_25_715 ();
 FILLCELL_X4 FILLER_25_729 ();
 FILLCELL_X8 FILLER_25_736 ();
 FILLCELL_X4 FILLER_25_744 ();
 FILLCELL_X2 FILLER_25_748 ();
 FILLCELL_X1 FILLER_25_750 ();
 FILLCELL_X4 FILLER_25_755 ();
 FILLCELL_X2 FILLER_25_759 ();
 FILLCELL_X32 FILLER_25_770 ();
 FILLCELL_X2 FILLER_25_802 ();
 FILLCELL_X4 FILLER_25_813 ();
 FILLCELL_X2 FILLER_25_817 ();
 FILLCELL_X4 FILLER_25_823 ();
 FILLCELL_X8 FILLER_25_829 ();
 FILLCELL_X4 FILLER_25_837 ();
 FILLCELL_X1 FILLER_25_841 ();
 FILLCELL_X4 FILLER_25_851 ();
 FILLCELL_X8 FILLER_25_866 ();
 FILLCELL_X4 FILLER_25_874 ();
 FILLCELL_X16 FILLER_25_889 ();
 FILLCELL_X8 FILLER_25_905 ();
 FILLCELL_X4 FILLER_25_913 ();
 FILLCELL_X2 FILLER_25_917 ();
 FILLCELL_X1 FILLER_25_919 ();
 FILLCELL_X8 FILLER_25_927 ();
 FILLCELL_X8 FILLER_25_945 ();
 FILLCELL_X1 FILLER_25_953 ();
 FILLCELL_X4 FILLER_25_961 ();
 FILLCELL_X8 FILLER_25_968 ();
 FILLCELL_X1 FILLER_25_976 ();
 FILLCELL_X4 FILLER_25_990 ();
 FILLCELL_X16 FILLER_25_1003 ();
 FILLCELL_X8 FILLER_25_1019 ();
 FILLCELL_X4 FILLER_25_1027 ();
 FILLCELL_X1 FILLER_25_1031 ();
 FILLCELL_X4 FILLER_25_1037 ();
 FILLCELL_X8 FILLER_25_1044 ();
 FILLCELL_X2 FILLER_25_1052 ();
 FILLCELL_X4 FILLER_25_1057 ();
 FILLCELL_X8 FILLER_25_1066 ();
 FILLCELL_X8 FILLER_25_1081 ();
 FILLCELL_X4 FILLER_25_1089 ();
 FILLCELL_X1 FILLER_25_1093 ();
 FILLCELL_X4 FILLER_25_1103 ();
 FILLCELL_X4 FILLER_25_1116 ();
 FILLCELL_X1 FILLER_25_1120 ();
 FILLCELL_X8 FILLER_25_1127 ();
 FILLCELL_X4 FILLER_25_1138 ();
 FILLCELL_X4 FILLER_25_1146 ();
 FILLCELL_X2 FILLER_25_1150 ();
 FILLCELL_X4 FILLER_25_1158 ();
 FILLCELL_X4 FILLER_25_1167 ();
 FILLCELL_X4 FILLER_25_1176 ();
 FILLCELL_X4 FILLER_25_1185 ();
 FILLCELL_X4 FILLER_25_1192 ();
 FILLCELL_X8 FILLER_25_1200 ();
 FILLCELL_X4 FILLER_25_1208 ();
 FILLCELL_X2 FILLER_25_1212 ();
 FILLCELL_X4 FILLER_25_1218 ();
 FILLCELL_X2 FILLER_25_1222 ();
 FILLCELL_X1 FILLER_25_1224 ();
 FILLCELL_X8 FILLER_25_1228 ();
 FILLCELL_X1 FILLER_25_1236 ();
 FILLCELL_X4 FILLER_25_1240 ();
 FILLCELL_X2 FILLER_25_1244 ();
 FILLCELL_X8 FILLER_25_1255 ();
 FILLCELL_X16 FILLER_25_1264 ();
 FILLCELL_X4 FILLER_25_1280 ();
 FILLCELL_X2 FILLER_25_1284 ();
 FILLCELL_X1 FILLER_25_1286 ();
 FILLCELL_X4 FILLER_25_1291 ();
 FILLCELL_X4 FILLER_25_1299 ();
 FILLCELL_X2 FILLER_25_1303 ();
 FILLCELL_X1 FILLER_25_1305 ();
 FILLCELL_X4 FILLER_25_1309 ();
 FILLCELL_X4 FILLER_25_1317 ();
 FILLCELL_X1 FILLER_25_1321 ();
 FILLCELL_X4 FILLER_25_1326 ();
 FILLCELL_X4 FILLER_25_1334 ();
 FILLCELL_X32 FILLER_25_1340 ();
 FILLCELL_X32 FILLER_25_1372 ();
 FILLCELL_X32 FILLER_25_1404 ();
 FILLCELL_X32 FILLER_25_1436 ();
 FILLCELL_X32 FILLER_25_1468 ();
 FILLCELL_X32 FILLER_25_1500 ();
 FILLCELL_X32 FILLER_25_1532 ();
 FILLCELL_X32 FILLER_25_1564 ();
 FILLCELL_X32 FILLER_25_1596 ();
 FILLCELL_X32 FILLER_25_1628 ();
 FILLCELL_X32 FILLER_25_1660 ();
 FILLCELL_X8 FILLER_25_1692 ();
 FILLCELL_X1 FILLER_25_1700 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X32 FILLER_26_193 ();
 FILLCELL_X32 FILLER_26_225 ();
 FILLCELL_X32 FILLER_26_257 ();
 FILLCELL_X32 FILLER_26_289 ();
 FILLCELL_X32 FILLER_26_321 ();
 FILLCELL_X16 FILLER_26_353 ();
 FILLCELL_X8 FILLER_26_369 ();
 FILLCELL_X4 FILLER_26_396 ();
 FILLCELL_X2 FILLER_26_400 ();
 FILLCELL_X8 FILLER_26_421 ();
 FILLCELL_X2 FILLER_26_429 ();
 FILLCELL_X4 FILLER_26_435 ();
 FILLCELL_X8 FILLER_26_441 ();
 FILLCELL_X4 FILLER_26_449 ();
 FILLCELL_X8 FILLER_26_463 ();
 FILLCELL_X2 FILLER_26_471 ();
 FILLCELL_X1 FILLER_26_473 ();
 FILLCELL_X32 FILLER_26_476 ();
 FILLCELL_X1 FILLER_26_508 ();
 FILLCELL_X4 FILLER_26_513 ();
 FILLCELL_X8 FILLER_26_526 ();
 FILLCELL_X2 FILLER_26_534 ();
 FILLCELL_X4 FILLER_26_542 ();
 FILLCELL_X2 FILLER_26_546 ();
 FILLCELL_X4 FILLER_26_557 ();
 FILLCELL_X2 FILLER_26_561 ();
 FILLCELL_X1 FILLER_26_563 ();
 FILLCELL_X4 FILLER_26_574 ();
 FILLCELL_X4 FILLER_26_581 ();
 FILLCELL_X4 FILLER_26_588 ();
 FILLCELL_X4 FILLER_26_595 ();
 FILLCELL_X1 FILLER_26_599 ();
 FILLCELL_X8 FILLER_26_604 ();
 FILLCELL_X4 FILLER_26_612 ();
 FILLCELL_X2 FILLER_26_616 ();
 FILLCELL_X4 FILLER_26_627 ();
 FILLCELL_X8 FILLER_26_632 ();
 FILLCELL_X1 FILLER_26_640 ();
 FILLCELL_X4 FILLER_26_648 ();
 FILLCELL_X16 FILLER_26_655 ();
 FILLCELL_X2 FILLER_26_671 ();
 FILLCELL_X1 FILLER_26_673 ();
 FILLCELL_X8 FILLER_26_681 ();
 FILLCELL_X1 FILLER_26_689 ();
 FILLCELL_X4 FILLER_26_694 ();
 FILLCELL_X8 FILLER_26_701 ();
 FILLCELL_X2 FILLER_26_709 ();
 FILLCELL_X1 FILLER_26_711 ();
 FILLCELL_X4 FILLER_26_716 ();
 FILLCELL_X4 FILLER_26_729 ();
 FILLCELL_X4 FILLER_26_737 ();
 FILLCELL_X4 FILLER_26_743 ();
 FILLCELL_X1 FILLER_26_747 ();
 FILLCELL_X4 FILLER_26_757 ();
 FILLCELL_X2 FILLER_26_761 ();
 FILLCELL_X1 FILLER_26_763 ();
 FILLCELL_X8 FILLER_26_774 ();
 FILLCELL_X1 FILLER_26_782 ();
 FILLCELL_X8 FILLER_26_792 ();
 FILLCELL_X4 FILLER_26_800 ();
 FILLCELL_X1 FILLER_26_804 ();
 FILLCELL_X8 FILLER_26_815 ();
 FILLCELL_X4 FILLER_26_828 ();
 FILLCELL_X16 FILLER_26_841 ();
 FILLCELL_X4 FILLER_26_857 ();
 FILLCELL_X4 FILLER_26_865 ();
 FILLCELL_X1 FILLER_26_869 ();
 FILLCELL_X4 FILLER_26_874 ();
 FILLCELL_X2 FILLER_26_878 ();
 FILLCELL_X8 FILLER_26_885 ();
 FILLCELL_X1 FILLER_26_893 ();
 FILLCELL_X4 FILLER_26_905 ();
 FILLCELL_X16 FILLER_26_920 ();
 FILLCELL_X8 FILLER_26_936 ();
 FILLCELL_X4 FILLER_26_944 ();
 FILLCELL_X2 FILLER_26_948 ();
 FILLCELL_X4 FILLER_26_952 ();
 FILLCELL_X1 FILLER_26_956 ();
 FILLCELL_X4 FILLER_26_964 ();
 FILLCELL_X8 FILLER_26_974 ();
 FILLCELL_X4 FILLER_26_982 ();
 FILLCELL_X1 FILLER_26_986 ();
 FILLCELL_X16 FILLER_26_996 ();
 FILLCELL_X8 FILLER_26_1012 ();
 FILLCELL_X2 FILLER_26_1020 ();
 FILLCELL_X1 FILLER_26_1022 ();
 FILLCELL_X4 FILLER_26_1030 ();
 FILLCELL_X4 FILLER_26_1041 ();
 FILLCELL_X1 FILLER_26_1045 ();
 FILLCELL_X4 FILLER_26_1053 ();
 FILLCELL_X1 FILLER_26_1057 ();
 FILLCELL_X4 FILLER_26_1060 ();
 FILLCELL_X4 FILLER_26_1071 ();
 FILLCELL_X8 FILLER_26_1080 ();
 FILLCELL_X2 FILLER_26_1088 ();
 FILLCELL_X16 FILLER_26_1099 ();
 FILLCELL_X1 FILLER_26_1115 ();
 FILLCELL_X4 FILLER_26_1119 ();
 FILLCELL_X4 FILLER_26_1128 ();
 FILLCELL_X4 FILLER_26_1136 ();
 FILLCELL_X4 FILLER_26_1144 ();
 FILLCELL_X2 FILLER_26_1148 ();
 FILLCELL_X1 FILLER_26_1150 ();
 FILLCELL_X8 FILLER_26_1160 ();
 FILLCELL_X4 FILLER_26_1172 ();
 FILLCELL_X8 FILLER_26_1180 ();
 FILLCELL_X2 FILLER_26_1188 ();
 FILLCELL_X1 FILLER_26_1190 ();
 FILLCELL_X8 FILLER_26_1195 ();
 FILLCELL_X2 FILLER_26_1203 ();
 FILLCELL_X1 FILLER_26_1205 ();
 FILLCELL_X4 FILLER_26_1211 ();
 FILLCELL_X8 FILLER_26_1220 ();
 FILLCELL_X2 FILLER_26_1228 ();
 FILLCELL_X16 FILLER_26_1234 ();
 FILLCELL_X8 FILLER_26_1250 ();
 FILLCELL_X4 FILLER_26_1258 ();
 FILLCELL_X1 FILLER_26_1262 ();
 FILLCELL_X8 FILLER_26_1272 ();
 FILLCELL_X2 FILLER_26_1280 ();
 FILLCELL_X1 FILLER_26_1282 ();
 FILLCELL_X4 FILLER_26_1285 ();
 FILLCELL_X8 FILLER_26_1291 ();
 FILLCELL_X4 FILLER_26_1301 ();
 FILLCELL_X8 FILLER_26_1308 ();
 FILLCELL_X4 FILLER_26_1320 ();
 FILLCELL_X4 FILLER_26_1328 ();
 FILLCELL_X4 FILLER_26_1336 ();
 FILLCELL_X4 FILLER_26_1343 ();
 FILLCELL_X32 FILLER_26_1349 ();
 FILLCELL_X32 FILLER_26_1381 ();
 FILLCELL_X32 FILLER_26_1413 ();
 FILLCELL_X32 FILLER_26_1445 ();
 FILLCELL_X32 FILLER_26_1477 ();
 FILLCELL_X32 FILLER_26_1509 ();
 FILLCELL_X32 FILLER_26_1541 ();
 FILLCELL_X32 FILLER_26_1573 ();
 FILLCELL_X32 FILLER_26_1605 ();
 FILLCELL_X32 FILLER_26_1637 ();
 FILLCELL_X32 FILLER_26_1669 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X32 FILLER_27_225 ();
 FILLCELL_X32 FILLER_27_257 ();
 FILLCELL_X32 FILLER_27_289 ();
 FILLCELL_X32 FILLER_27_321 ();
 FILLCELL_X16 FILLER_27_353 ();
 FILLCELL_X1 FILLER_27_369 ();
 FILLCELL_X32 FILLER_27_374 ();
 FILLCELL_X8 FILLER_27_406 ();
 FILLCELL_X4 FILLER_27_414 ();
 FILLCELL_X2 FILLER_27_418 ();
 FILLCELL_X1 FILLER_27_420 ();
 FILLCELL_X4 FILLER_27_425 ();
 FILLCELL_X4 FILLER_27_433 ();
 FILLCELL_X4 FILLER_27_440 ();
 FILLCELL_X2 FILLER_27_444 ();
 FILLCELL_X4 FILLER_27_449 ();
 FILLCELL_X4 FILLER_27_456 ();
 FILLCELL_X4 FILLER_27_462 ();
 FILLCELL_X2 FILLER_27_466 ();
 FILLCELL_X1 FILLER_27_468 ();
 FILLCELL_X4 FILLER_27_479 ();
 FILLCELL_X16 FILLER_27_486 ();
 FILLCELL_X8 FILLER_27_506 ();
 FILLCELL_X4 FILLER_27_514 ();
 FILLCELL_X1 FILLER_27_518 ();
 FILLCELL_X8 FILLER_27_523 ();
 FILLCELL_X4 FILLER_27_531 ();
 FILLCELL_X2 FILLER_27_535 ();
 FILLCELL_X4 FILLER_27_542 ();
 FILLCELL_X4 FILLER_27_553 ();
 FILLCELL_X4 FILLER_27_560 ();
 FILLCELL_X4 FILLER_27_567 ();
 FILLCELL_X2 FILLER_27_571 ();
 FILLCELL_X1 FILLER_27_573 ();
 FILLCELL_X4 FILLER_27_583 ();
 FILLCELL_X8 FILLER_27_596 ();
 FILLCELL_X2 FILLER_27_604 ();
 FILLCELL_X8 FILLER_27_615 ();
 FILLCELL_X4 FILLER_27_623 ();
 FILLCELL_X4 FILLER_27_630 ();
 FILLCELL_X4 FILLER_27_638 ();
 FILLCELL_X2 FILLER_27_642 ();
 FILLCELL_X16 FILLER_27_649 ();
 FILLCELL_X4 FILLER_27_665 ();
 FILLCELL_X1 FILLER_27_669 ();
 FILLCELL_X4 FILLER_27_679 ();
 FILLCELL_X4 FILLER_27_690 ();
 FILLCELL_X2 FILLER_27_694 ();
 FILLCELL_X4 FILLER_27_705 ();
 FILLCELL_X4 FILLER_27_713 ();
 FILLCELL_X8 FILLER_27_720 ();
 FILLCELL_X4 FILLER_27_728 ();
 FILLCELL_X1 FILLER_27_732 ();
 FILLCELL_X4 FILLER_27_738 ();
 FILLCELL_X4 FILLER_27_745 ();
 FILLCELL_X4 FILLER_27_758 ();
 FILLCELL_X2 FILLER_27_762 ();
 FILLCELL_X4 FILLER_27_773 ();
 FILLCELL_X4 FILLER_27_781 ();
 FILLCELL_X4 FILLER_27_790 ();
 FILLCELL_X4 FILLER_27_796 ();
 FILLCELL_X4 FILLER_27_803 ();
 FILLCELL_X4 FILLER_27_811 ();
 FILLCELL_X4 FILLER_27_817 ();
 FILLCELL_X1 FILLER_27_821 ();
 FILLCELL_X8 FILLER_27_827 ();
 FILLCELL_X2 FILLER_27_835 ();
 FILLCELL_X1 FILLER_27_837 ();
 FILLCELL_X8 FILLER_27_843 ();
 FILLCELL_X2 FILLER_27_851 ();
 FILLCELL_X1 FILLER_27_853 ();
 FILLCELL_X4 FILLER_27_859 ();
 FILLCELL_X8 FILLER_27_868 ();
 FILLCELL_X2 FILLER_27_876 ();
 FILLCELL_X1 FILLER_27_878 ();
 FILLCELL_X4 FILLER_27_884 ();
 FILLCELL_X4 FILLER_27_893 ();
 FILLCELL_X4 FILLER_27_901 ();
 FILLCELL_X16 FILLER_27_916 ();
 FILLCELL_X1 FILLER_27_932 ();
 FILLCELL_X4 FILLER_27_940 ();
 FILLCELL_X8 FILLER_27_951 ();
 FILLCELL_X4 FILLER_27_959 ();
 FILLCELL_X2 FILLER_27_963 ();
 FILLCELL_X4 FILLER_27_974 ();
 FILLCELL_X2 FILLER_27_978 ();
 FILLCELL_X8 FILLER_27_984 ();
 FILLCELL_X4 FILLER_27_992 ();
 FILLCELL_X1 FILLER_27_996 ();
 FILLCELL_X4 FILLER_27_1010 ();
 FILLCELL_X4 FILLER_27_1021 ();
 FILLCELL_X8 FILLER_27_1032 ();
 FILLCELL_X2 FILLER_27_1040 ();
 FILLCELL_X8 FILLER_27_1049 ();
 FILLCELL_X1 FILLER_27_1057 ();
 FILLCELL_X4 FILLER_27_1065 ();
 FILLCELL_X2 FILLER_27_1069 ();
 FILLCELL_X4 FILLER_27_1080 ();
 FILLCELL_X2 FILLER_27_1084 ();
 FILLCELL_X1 FILLER_27_1086 ();
 FILLCELL_X8 FILLER_27_1096 ();
 FILLCELL_X4 FILLER_27_1110 ();
 FILLCELL_X4 FILLER_27_1116 ();
 FILLCELL_X1 FILLER_27_1120 ();
 FILLCELL_X4 FILLER_27_1124 ();
 FILLCELL_X32 FILLER_27_1132 ();
 FILLCELL_X16 FILLER_27_1164 ();
 FILLCELL_X2 FILLER_27_1180 ();
 FILLCELL_X1 FILLER_27_1182 ();
 FILLCELL_X8 FILLER_27_1192 ();
 FILLCELL_X4 FILLER_27_1203 ();
 FILLCELL_X4 FILLER_27_1212 ();
 FILLCELL_X8 FILLER_27_1220 ();
 FILLCELL_X4 FILLER_27_1228 ();
 FILLCELL_X1 FILLER_27_1232 ();
 FILLCELL_X4 FILLER_27_1239 ();
 FILLCELL_X4 FILLER_27_1247 ();
 FILLCELL_X2 FILLER_27_1251 ();
 FILLCELL_X4 FILLER_27_1256 ();
 FILLCELL_X2 FILLER_27_1260 ();
 FILLCELL_X1 FILLER_27_1262 ();
 FILLCELL_X4 FILLER_27_1264 ();
 FILLCELL_X4 FILLER_27_1277 ();
 FILLCELL_X4 FILLER_27_1283 ();
 FILLCELL_X4 FILLER_27_1292 ();
 FILLCELL_X8 FILLER_27_1301 ();
 FILLCELL_X1 FILLER_27_1309 ();
 FILLCELL_X4 FILLER_27_1314 ();
 FILLCELL_X4 FILLER_27_1320 ();
 FILLCELL_X4 FILLER_27_1331 ();
 FILLCELL_X32 FILLER_27_1338 ();
 FILLCELL_X16 FILLER_27_1370 ();
 FILLCELL_X8 FILLER_27_1386 ();
 FILLCELL_X2 FILLER_27_1394 ();
 FILLCELL_X32 FILLER_27_1400 ();
 FILLCELL_X32 FILLER_27_1432 ();
 FILLCELL_X32 FILLER_27_1464 ();
 FILLCELL_X32 FILLER_27_1496 ();
 FILLCELL_X16 FILLER_27_1528 ();
 FILLCELL_X4 FILLER_27_1544 ();
 FILLCELL_X2 FILLER_27_1548 ();
 FILLCELL_X8 FILLER_27_1554 ();
 FILLCELL_X4 FILLER_27_1562 ();
 FILLCELL_X32 FILLER_27_1583 ();
 FILLCELL_X32 FILLER_27_1615 ();
 FILLCELL_X32 FILLER_27_1647 ();
 FILLCELL_X16 FILLER_27_1679 ();
 FILLCELL_X4 FILLER_27_1695 ();
 FILLCELL_X2 FILLER_27_1699 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X32 FILLER_28_225 ();
 FILLCELL_X32 FILLER_28_257 ();
 FILLCELL_X32 FILLER_28_289 ();
 FILLCELL_X32 FILLER_28_321 ();
 FILLCELL_X32 FILLER_28_353 ();
 FILLCELL_X2 FILLER_28_385 ();
 FILLCELL_X1 FILLER_28_387 ();
 FILLCELL_X4 FILLER_28_392 ();
 FILLCELL_X2 FILLER_28_396 ();
 FILLCELL_X4 FILLER_28_417 ();
 FILLCELL_X4 FILLER_28_440 ();
 FILLCELL_X4 FILLER_28_450 ();
 FILLCELL_X4 FILLER_28_459 ();
 FILLCELL_X16 FILLER_28_467 ();
 FILLCELL_X4 FILLER_28_483 ();
 FILLCELL_X2 FILLER_28_487 ();
 FILLCELL_X4 FILLER_28_491 ();
 FILLCELL_X4 FILLER_28_499 ();
 FILLCELL_X4 FILLER_28_507 ();
 FILLCELL_X2 FILLER_28_511 ();
 FILLCELL_X4 FILLER_28_522 ();
 FILLCELL_X16 FILLER_28_530 ();
 FILLCELL_X1 FILLER_28_546 ();
 FILLCELL_X4 FILLER_28_556 ();
 FILLCELL_X4 FILLER_28_567 ();
 FILLCELL_X4 FILLER_28_581 ();
 FILLCELL_X16 FILLER_28_592 ();
 FILLCELL_X8 FILLER_28_608 ();
 FILLCELL_X4 FILLER_28_616 ();
 FILLCELL_X4 FILLER_28_627 ();
 FILLCELL_X4 FILLER_28_632 ();
 FILLCELL_X4 FILLER_28_649 ();
 FILLCELL_X4 FILLER_28_659 ();
 FILLCELL_X16 FILLER_28_667 ();
 FILLCELL_X4 FILLER_28_683 ();
 FILLCELL_X1 FILLER_28_687 ();
 FILLCELL_X4 FILLER_28_701 ();
 FILLCELL_X4 FILLER_28_718 ();
 FILLCELL_X4 FILLER_28_732 ();
 FILLCELL_X1 FILLER_28_736 ();
 FILLCELL_X4 FILLER_28_739 ();
 FILLCELL_X4 FILLER_28_748 ();
 FILLCELL_X8 FILLER_28_757 ();
 FILLCELL_X1 FILLER_28_765 ();
 FILLCELL_X4 FILLER_28_770 ();
 FILLCELL_X1 FILLER_28_774 ();
 FILLCELL_X4 FILLER_28_777 ();
 FILLCELL_X16 FILLER_28_784 ();
 FILLCELL_X8 FILLER_28_809 ();
 FILLCELL_X4 FILLER_28_820 ();
 FILLCELL_X4 FILLER_28_833 ();
 FILLCELL_X1 FILLER_28_837 ();
 FILLCELL_X4 FILLER_28_842 ();
 FILLCELL_X4 FILLER_28_850 ();
 FILLCELL_X4 FILLER_28_859 ();
 FILLCELL_X8 FILLER_28_868 ();
 FILLCELL_X4 FILLER_28_881 ();
 FILLCELL_X4 FILLER_28_890 ();
 FILLCELL_X4 FILLER_28_899 ();
 FILLCELL_X4 FILLER_28_908 ();
 FILLCELL_X4 FILLER_28_916 ();
 FILLCELL_X4 FILLER_28_924 ();
 FILLCELL_X2 FILLER_28_928 ();
 FILLCELL_X8 FILLER_28_936 ();
 FILLCELL_X1 FILLER_28_944 ();
 FILLCELL_X8 FILLER_28_952 ();
 FILLCELL_X1 FILLER_28_960 ();
 FILLCELL_X4 FILLER_28_968 ();
 FILLCELL_X8 FILLER_28_978 ();
 FILLCELL_X4 FILLER_28_993 ();
 FILLCELL_X4 FILLER_28_1002 ();
 FILLCELL_X2 FILLER_28_1006 ();
 FILLCELL_X1 FILLER_28_1008 ();
 FILLCELL_X8 FILLER_28_1022 ();
 FILLCELL_X4 FILLER_28_1037 ();
 FILLCELL_X16 FILLER_28_1048 ();
 FILLCELL_X4 FILLER_28_1067 ();
 FILLCELL_X8 FILLER_28_1084 ();
 FILLCELL_X4 FILLER_28_1092 ();
 FILLCELL_X2 FILLER_28_1096 ();
 FILLCELL_X8 FILLER_28_1102 ();
 FILLCELL_X1 FILLER_28_1110 ();
 FILLCELL_X4 FILLER_28_1115 ();
 FILLCELL_X4 FILLER_28_1123 ();
 FILLCELL_X4 FILLER_28_1130 ();
 FILLCELL_X1 FILLER_28_1134 ();
 FILLCELL_X8 FILLER_28_1144 ();
 FILLCELL_X2 FILLER_28_1152 ();
 FILLCELL_X4 FILLER_28_1165 ();
 FILLCELL_X8 FILLER_28_1180 ();
 FILLCELL_X4 FILLER_28_1199 ();
 FILLCELL_X8 FILLER_28_1212 ();
 FILLCELL_X4 FILLER_28_1220 ();
 FILLCELL_X1 FILLER_28_1224 ();
 FILLCELL_X4 FILLER_28_1228 ();
 FILLCELL_X2 FILLER_28_1232 ();
 FILLCELL_X1 FILLER_28_1234 ();
 FILLCELL_X4 FILLER_28_1240 ();
 FILLCELL_X1 FILLER_28_1244 ();
 FILLCELL_X4 FILLER_28_1250 ();
 FILLCELL_X4 FILLER_28_1259 ();
 FILLCELL_X1 FILLER_28_1263 ();
 FILLCELL_X4 FILLER_28_1273 ();
 FILLCELL_X4 FILLER_28_1280 ();
 FILLCELL_X4 FILLER_28_1288 ();
 FILLCELL_X4 FILLER_28_1296 ();
 FILLCELL_X4 FILLER_28_1304 ();
 FILLCELL_X4 FILLER_28_1312 ();
 FILLCELL_X4 FILLER_28_1318 ();
 FILLCELL_X32 FILLER_28_1324 ();
 FILLCELL_X32 FILLER_28_1356 ();
 FILLCELL_X4 FILLER_28_1388 ();
 FILLCELL_X1 FILLER_28_1392 ();
 FILLCELL_X32 FILLER_28_1412 ();
 FILLCELL_X32 FILLER_28_1444 ();
 FILLCELL_X32 FILLER_28_1476 ();
 FILLCELL_X32 FILLER_28_1508 ();
 FILLCELL_X4 FILLER_28_1540 ();
 FILLCELL_X1 FILLER_28_1544 ();
 FILLCELL_X32 FILLER_28_1564 ();
 FILLCELL_X32 FILLER_28_1596 ();
 FILLCELL_X32 FILLER_28_1628 ();
 FILLCELL_X32 FILLER_28_1660 ();
 FILLCELL_X8 FILLER_28_1692 ();
 FILLCELL_X1 FILLER_28_1700 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X32 FILLER_29_193 ();
 FILLCELL_X32 FILLER_29_225 ();
 FILLCELL_X32 FILLER_29_257 ();
 FILLCELL_X32 FILLER_29_289 ();
 FILLCELL_X32 FILLER_29_321 ();
 FILLCELL_X16 FILLER_29_353 ();
 FILLCELL_X8 FILLER_29_369 ();
 FILLCELL_X16 FILLER_29_396 ();
 FILLCELL_X4 FILLER_29_412 ();
 FILLCELL_X16 FILLER_29_420 ();
 FILLCELL_X4 FILLER_29_436 ();
 FILLCELL_X2 FILLER_29_440 ();
 FILLCELL_X1 FILLER_29_442 ();
 FILLCELL_X4 FILLER_29_462 ();
 FILLCELL_X4 FILLER_29_475 ();
 FILLCELL_X2 FILLER_29_479 ();
 FILLCELL_X8 FILLER_29_485 ();
 FILLCELL_X2 FILLER_29_493 ();
 FILLCELL_X1 FILLER_29_495 ();
 FILLCELL_X4 FILLER_29_506 ();
 FILLCELL_X1 FILLER_29_510 ();
 FILLCELL_X4 FILLER_29_514 ();
 FILLCELL_X4 FILLER_29_522 ();
 FILLCELL_X4 FILLER_29_530 ();
 FILLCELL_X16 FILLER_29_538 ();
 FILLCELL_X2 FILLER_29_554 ();
 FILLCELL_X4 FILLER_29_560 ();
 FILLCELL_X8 FILLER_29_567 ();
 FILLCELL_X4 FILLER_29_575 ();
 FILLCELL_X2 FILLER_29_579 ();
 FILLCELL_X1 FILLER_29_581 ();
 FILLCELL_X4 FILLER_29_584 ();
 FILLCELL_X4 FILLER_29_592 ();
 FILLCELL_X1 FILLER_29_596 ();
 FILLCELL_X4 FILLER_29_601 ();
 FILLCELL_X4 FILLER_29_609 ();
 FILLCELL_X4 FILLER_29_618 ();
 FILLCELL_X4 FILLER_29_626 ();
 FILLCELL_X4 FILLER_29_632 ();
 FILLCELL_X4 FILLER_29_639 ();
 FILLCELL_X4 FILLER_29_647 ();
 FILLCELL_X4 FILLER_29_653 ();
 FILLCELL_X8 FILLER_29_659 ();
 FILLCELL_X4 FILLER_29_667 ();
 FILLCELL_X2 FILLER_29_671 ();
 FILLCELL_X16 FILLER_29_686 ();
 FILLCELL_X4 FILLER_29_702 ();
 FILLCELL_X8 FILLER_29_710 ();
 FILLCELL_X4 FILLER_29_718 ();
 FILLCELL_X2 FILLER_29_722 ();
 FILLCELL_X1 FILLER_29_724 ();
 FILLCELL_X4 FILLER_29_732 ();
 FILLCELL_X4 FILLER_29_738 ();
 FILLCELL_X2 FILLER_29_742 ();
 FILLCELL_X1 FILLER_29_744 ();
 FILLCELL_X4 FILLER_29_749 ();
 FILLCELL_X2 FILLER_29_753 ();
 FILLCELL_X1 FILLER_29_755 ();
 FILLCELL_X8 FILLER_29_761 ();
 FILLCELL_X1 FILLER_29_769 ();
 FILLCELL_X4 FILLER_29_774 ();
 FILLCELL_X4 FILLER_29_787 ();
 FILLCELL_X1 FILLER_29_791 ();
 FILLCELL_X4 FILLER_29_796 ();
 FILLCELL_X2 FILLER_29_800 ();
 FILLCELL_X8 FILLER_29_806 ();
 FILLCELL_X4 FILLER_29_814 ();
 FILLCELL_X4 FILLER_29_820 ();
 FILLCELL_X4 FILLER_29_829 ();
 FILLCELL_X4 FILLER_29_837 ();
 FILLCELL_X4 FILLER_29_845 ();
 FILLCELL_X4 FILLER_29_854 ();
 FILLCELL_X8 FILLER_29_863 ();
 FILLCELL_X1 FILLER_29_871 ();
 FILLCELL_X4 FILLER_29_876 ();
 FILLCELL_X1 FILLER_29_880 ();
 FILLCELL_X4 FILLER_29_885 ();
 FILLCELL_X4 FILLER_29_894 ();
 FILLCELL_X4 FILLER_29_903 ();
 FILLCELL_X8 FILLER_29_911 ();
 FILLCELL_X2 FILLER_29_919 ();
 FILLCELL_X4 FILLER_29_927 ();
 FILLCELL_X1 FILLER_29_931 ();
 FILLCELL_X4 FILLER_29_941 ();
 FILLCELL_X16 FILLER_29_951 ();
 FILLCELL_X8 FILLER_29_967 ();
 FILLCELL_X4 FILLER_29_975 ();
 FILLCELL_X2 FILLER_29_979 ();
 FILLCELL_X4 FILLER_29_985 ();
 FILLCELL_X4 FILLER_29_996 ();
 FILLCELL_X2 FILLER_29_1000 ();
 FILLCELL_X16 FILLER_29_1007 ();
 FILLCELL_X8 FILLER_29_1023 ();
 FILLCELL_X2 FILLER_29_1031 ();
 FILLCELL_X4 FILLER_29_1038 ();
 FILLCELL_X8 FILLER_29_1049 ();
 FILLCELL_X4 FILLER_29_1057 ();
 FILLCELL_X1 FILLER_29_1061 ();
 FILLCELL_X8 FILLER_29_1069 ();
 FILLCELL_X4 FILLER_29_1077 ();
 FILLCELL_X2 FILLER_29_1081 ();
 FILLCELL_X1 FILLER_29_1083 ();
 FILLCELL_X4 FILLER_29_1087 ();
 FILLCELL_X4 FILLER_29_1095 ();
 FILLCELL_X4 FILLER_29_1102 ();
 FILLCELL_X2 FILLER_29_1106 ();
 FILLCELL_X4 FILLER_29_1112 ();
 FILLCELL_X8 FILLER_29_1120 ();
 FILLCELL_X2 FILLER_29_1128 ();
 FILLCELL_X4 FILLER_29_1139 ();
 FILLCELL_X16 FILLER_29_1152 ();
 FILLCELL_X1 FILLER_29_1168 ();
 FILLCELL_X4 FILLER_29_1174 ();
 FILLCELL_X4 FILLER_29_1183 ();
 FILLCELL_X8 FILLER_29_1192 ();
 FILLCELL_X2 FILLER_29_1200 ();
 FILLCELL_X1 FILLER_29_1202 ();
 FILLCELL_X4 FILLER_29_1212 ();
 FILLCELL_X4 FILLER_29_1222 ();
 FILLCELL_X4 FILLER_29_1231 ();
 FILLCELL_X4 FILLER_29_1239 ();
 FILLCELL_X4 FILLER_29_1247 ();
 FILLCELL_X8 FILLER_29_1255 ();
 FILLCELL_X4 FILLER_29_1264 ();
 FILLCELL_X4 FILLER_29_1274 ();
 FILLCELL_X32 FILLER_29_1280 ();
 FILLCELL_X32 FILLER_29_1312 ();
 FILLCELL_X32 FILLER_29_1344 ();
 FILLCELL_X32 FILLER_29_1376 ();
 FILLCELL_X32 FILLER_29_1408 ();
 FILLCELL_X32 FILLER_29_1440 ();
 FILLCELL_X32 FILLER_29_1472 ();
 FILLCELL_X2 FILLER_29_1504 ();
 FILLCELL_X16 FILLER_29_1510 ();
 FILLCELL_X4 FILLER_29_1526 ();
 FILLCELL_X2 FILLER_29_1530 ();
 FILLCELL_X32 FILLER_29_1536 ();
 FILLCELL_X2 FILLER_29_1568 ();
 FILLCELL_X1 FILLER_29_1570 ();
 FILLCELL_X32 FILLER_29_1590 ();
 FILLCELL_X32 FILLER_29_1622 ();
 FILLCELL_X32 FILLER_29_1654 ();
 FILLCELL_X8 FILLER_29_1686 ();
 FILLCELL_X4 FILLER_29_1697 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_161 ();
 FILLCELL_X32 FILLER_30_193 ();
 FILLCELL_X32 FILLER_30_225 ();
 FILLCELL_X32 FILLER_30_257 ();
 FILLCELL_X32 FILLER_30_289 ();
 FILLCELL_X32 FILLER_30_321 ();
 FILLCELL_X32 FILLER_30_353 ();
 FILLCELL_X16 FILLER_30_385 ();
 FILLCELL_X8 FILLER_30_401 ();
 FILLCELL_X2 FILLER_30_409 ();
 FILLCELL_X1 FILLER_30_411 ();
 FILLCELL_X16 FILLER_30_431 ();
 FILLCELL_X2 FILLER_30_447 ();
 FILLCELL_X4 FILLER_30_451 ();
 FILLCELL_X4 FILLER_30_460 ();
 FILLCELL_X4 FILLER_30_467 ();
 FILLCELL_X2 FILLER_30_471 ();
 FILLCELL_X16 FILLER_30_480 ();
 FILLCELL_X8 FILLER_30_496 ();
 FILLCELL_X1 FILLER_30_504 ();
 FILLCELL_X4 FILLER_30_508 ();
 FILLCELL_X4 FILLER_30_516 ();
 FILLCELL_X8 FILLER_30_522 ();
 FILLCELL_X2 FILLER_30_530 ();
 FILLCELL_X4 FILLER_30_534 ();
 FILLCELL_X1 FILLER_30_538 ();
 FILLCELL_X8 FILLER_30_543 ();
 FILLCELL_X2 FILLER_30_551 ();
 FILLCELL_X1 FILLER_30_553 ();
 FILLCELL_X8 FILLER_30_557 ();
 FILLCELL_X4 FILLER_30_565 ();
 FILLCELL_X1 FILLER_30_569 ();
 FILLCELL_X4 FILLER_30_579 ();
 FILLCELL_X1 FILLER_30_583 ();
 FILLCELL_X4 FILLER_30_587 ();
 FILLCELL_X2 FILLER_30_591 ();
 FILLCELL_X1 FILLER_30_593 ();
 FILLCELL_X4 FILLER_30_597 ();
 FILLCELL_X4 FILLER_30_611 ();
 FILLCELL_X2 FILLER_30_615 ();
 FILLCELL_X1 FILLER_30_617 ();
 FILLCELL_X4 FILLER_30_627 ();
 FILLCELL_X4 FILLER_30_632 ();
 FILLCELL_X8 FILLER_30_640 ();
 FILLCELL_X1 FILLER_30_648 ();
 FILLCELL_X4 FILLER_30_656 ();
 FILLCELL_X8 FILLER_30_673 ();
 FILLCELL_X1 FILLER_30_681 ();
 FILLCELL_X8 FILLER_30_695 ();
 FILLCELL_X8 FILLER_30_710 ();
 FILLCELL_X4 FILLER_30_718 ();
 FILLCELL_X2 FILLER_30_722 ();
 FILLCELL_X1 FILLER_30_724 ();
 FILLCELL_X8 FILLER_30_735 ();
 FILLCELL_X4 FILLER_30_745 ();
 FILLCELL_X4 FILLER_30_753 ();
 FILLCELL_X2 FILLER_30_757 ();
 FILLCELL_X4 FILLER_30_763 ();
 FILLCELL_X4 FILLER_30_771 ();
 FILLCELL_X4 FILLER_30_784 ();
 FILLCELL_X8 FILLER_30_790 ();
 FILLCELL_X4 FILLER_30_807 ();
 FILLCELL_X8 FILLER_30_815 ();
 FILLCELL_X4 FILLER_30_825 ();
 FILLCELL_X4 FILLER_30_831 ();
 FILLCELL_X16 FILLER_30_839 ();
 FILLCELL_X8 FILLER_30_855 ();
 FILLCELL_X2 FILLER_30_863 ();
 FILLCELL_X1 FILLER_30_865 ();
 FILLCELL_X16 FILLER_30_870 ();
 FILLCELL_X2 FILLER_30_886 ();
 FILLCELL_X8 FILLER_30_897 ();
 FILLCELL_X4 FILLER_30_905 ();
 FILLCELL_X8 FILLER_30_918 ();
 FILLCELL_X1 FILLER_30_926 ();
 FILLCELL_X8 FILLER_30_936 ();
 FILLCELL_X4 FILLER_30_944 ();
 FILLCELL_X4 FILLER_30_967 ();
 FILLCELL_X2 FILLER_30_971 ();
 FILLCELL_X1 FILLER_30_973 ();
 FILLCELL_X4 FILLER_30_978 ();
 FILLCELL_X4 FILLER_30_995 ();
 FILLCELL_X2 FILLER_30_999 ();
 FILLCELL_X4 FILLER_30_1008 ();
 FILLCELL_X8 FILLER_30_1016 ();
 FILLCELL_X8 FILLER_30_1031 ();
 FILLCELL_X2 FILLER_30_1039 ();
 FILLCELL_X4 FILLER_30_1050 ();
 FILLCELL_X4 FILLER_30_1063 ();
 FILLCELL_X8 FILLER_30_1070 ();
 FILLCELL_X4 FILLER_30_1082 ();
 FILLCELL_X4 FILLER_30_1092 ();
 FILLCELL_X8 FILLER_30_1099 ();
 FILLCELL_X4 FILLER_30_1107 ();
 FILLCELL_X2 FILLER_30_1111 ();
 FILLCELL_X4 FILLER_30_1119 ();
 FILLCELL_X16 FILLER_30_1126 ();
 FILLCELL_X1 FILLER_30_1142 ();
 FILLCELL_X4 FILLER_30_1154 ();
 FILLCELL_X8 FILLER_30_1169 ();
 FILLCELL_X4 FILLER_30_1186 ();
 FILLCELL_X2 FILLER_30_1190 ();
 FILLCELL_X8 FILLER_30_1196 ();
 FILLCELL_X4 FILLER_30_1210 ();
 FILLCELL_X4 FILLER_30_1218 ();
 FILLCELL_X4 FILLER_30_1226 ();
 FILLCELL_X2 FILLER_30_1230 ();
 FILLCELL_X1 FILLER_30_1232 ();
 FILLCELL_X8 FILLER_30_1235 ();
 FILLCELL_X4 FILLER_30_1243 ();
 FILLCELL_X1 FILLER_30_1247 ();
 FILLCELL_X4 FILLER_30_1252 ();
 FILLCELL_X2 FILLER_30_1256 ();
 FILLCELL_X1 FILLER_30_1258 ();
 FILLCELL_X4 FILLER_30_1264 ();
 FILLCELL_X4 FILLER_30_1277 ();
 FILLCELL_X4 FILLER_30_1286 ();
 FILLCELL_X4 FILLER_30_1294 ();
 FILLCELL_X2 FILLER_30_1298 ();
 FILLCELL_X32 FILLER_30_1302 ();
 FILLCELL_X32 FILLER_30_1334 ();
 FILLCELL_X8 FILLER_30_1366 ();
 FILLCELL_X4 FILLER_30_1374 ();
 FILLCELL_X1 FILLER_30_1378 ();
 FILLCELL_X32 FILLER_30_1383 ();
 FILLCELL_X32 FILLER_30_1415 ();
 FILLCELL_X32 FILLER_30_1447 ();
 FILLCELL_X32 FILLER_30_1479 ();
 FILLCELL_X32 FILLER_30_1511 ();
 FILLCELL_X32 FILLER_30_1543 ();
 FILLCELL_X32 FILLER_30_1575 ();
 FILLCELL_X32 FILLER_30_1607 ();
 FILLCELL_X32 FILLER_30_1639 ();
 FILLCELL_X16 FILLER_30_1671 ();
 FILLCELL_X8 FILLER_30_1687 ();
 FILLCELL_X4 FILLER_30_1695 ();
 FILLCELL_X2 FILLER_30_1699 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X32 FILLER_31_193 ();
 FILLCELL_X32 FILLER_31_225 ();
 FILLCELL_X32 FILLER_31_257 ();
 FILLCELL_X32 FILLER_31_289 ();
 FILLCELL_X32 FILLER_31_321 ();
 FILLCELL_X32 FILLER_31_353 ();
 FILLCELL_X32 FILLER_31_385 ();
 FILLCELL_X4 FILLER_31_417 ();
 FILLCELL_X2 FILLER_31_421 ();
 FILLCELL_X1 FILLER_31_423 ();
 FILLCELL_X8 FILLER_31_426 ();
 FILLCELL_X4 FILLER_31_434 ();
 FILLCELL_X2 FILLER_31_438 ();
 FILLCELL_X4 FILLER_31_443 ();
 FILLCELL_X4 FILLER_31_450 ();
 FILLCELL_X2 FILLER_31_454 ();
 FILLCELL_X1 FILLER_31_456 ();
 FILLCELL_X4 FILLER_31_462 ();
 FILLCELL_X2 FILLER_31_466 ();
 FILLCELL_X1 FILLER_31_468 ();
 FILLCELL_X4 FILLER_31_473 ();
 FILLCELL_X1 FILLER_31_477 ();
 FILLCELL_X4 FILLER_31_482 ();
 FILLCELL_X8 FILLER_31_495 ();
 FILLCELL_X16 FILLER_31_507 ();
 FILLCELL_X2 FILLER_31_523 ();
 FILLCELL_X1 FILLER_31_525 ();
 FILLCELL_X4 FILLER_31_536 ();
 FILLCELL_X4 FILLER_31_547 ();
 FILLCELL_X2 FILLER_31_551 ();
 FILLCELL_X1 FILLER_31_553 ();
 FILLCELL_X8 FILLER_31_561 ();
 FILLCELL_X4 FILLER_31_569 ();
 FILLCELL_X2 FILLER_31_573 ();
 FILLCELL_X4 FILLER_31_588 ();
 FILLCELL_X16 FILLER_31_599 ();
 FILLCELL_X8 FILLER_31_615 ();
 FILLCELL_X8 FILLER_31_627 ();
 FILLCELL_X1 FILLER_31_635 ();
 FILLCELL_X4 FILLER_31_642 ();
 FILLCELL_X4 FILLER_31_652 ();
 FILLCELL_X16 FILLER_31_661 ();
 FILLCELL_X4 FILLER_31_677 ();
 FILLCELL_X16 FILLER_31_688 ();
 FILLCELL_X2 FILLER_31_704 ();
 FILLCELL_X8 FILLER_31_708 ();
 FILLCELL_X4 FILLER_31_720 ();
 FILLCELL_X4 FILLER_31_733 ();
 FILLCELL_X8 FILLER_31_739 ();
 FILLCELL_X4 FILLER_31_751 ();
 FILLCELL_X4 FILLER_31_758 ();
 FILLCELL_X4 FILLER_31_764 ();
 FILLCELL_X1 FILLER_31_768 ();
 FILLCELL_X4 FILLER_31_774 ();
 FILLCELL_X4 FILLER_31_780 ();
 FILLCELL_X2 FILLER_31_784 ();
 FILLCELL_X1 FILLER_31_786 ();
 FILLCELL_X4 FILLER_31_789 ();
 FILLCELL_X8 FILLER_31_798 ();
 FILLCELL_X4 FILLER_31_806 ();
 FILLCELL_X2 FILLER_31_810 ();
 FILLCELL_X4 FILLER_31_814 ();
 FILLCELL_X4 FILLER_31_822 ();
 FILLCELL_X4 FILLER_31_830 ();
 FILLCELL_X4 FILLER_31_838 ();
 FILLCELL_X8 FILLER_31_851 ();
 FILLCELL_X2 FILLER_31_859 ();
 FILLCELL_X1 FILLER_31_861 ();
 FILLCELL_X8 FILLER_31_871 ();
 FILLCELL_X1 FILLER_31_879 ();
 FILLCELL_X8 FILLER_31_889 ();
 FILLCELL_X2 FILLER_31_897 ();
 FILLCELL_X1 FILLER_31_899 ();
 FILLCELL_X4 FILLER_31_910 ();
 FILLCELL_X2 FILLER_31_914 ();
 FILLCELL_X8 FILLER_31_926 ();
 FILLCELL_X4 FILLER_31_934 ();
 FILLCELL_X4 FILLER_31_947 ();
 FILLCELL_X1 FILLER_31_951 ();
 FILLCELL_X4 FILLER_31_955 ();
 FILLCELL_X8 FILLER_31_969 ();
 FILLCELL_X4 FILLER_31_977 ();
 FILLCELL_X2 FILLER_31_981 ();
 FILLCELL_X1 FILLER_31_983 ();
 FILLCELL_X4 FILLER_31_994 ();
 FILLCELL_X4 FILLER_31_1000 ();
 FILLCELL_X4 FILLER_31_1007 ();
 FILLCELL_X8 FILLER_31_1018 ();
 FILLCELL_X1 FILLER_31_1026 ();
 FILLCELL_X4 FILLER_31_1032 ();
 FILLCELL_X4 FILLER_31_1041 ();
 FILLCELL_X8 FILLER_31_1049 ();
 FILLCELL_X4 FILLER_31_1057 ();
 FILLCELL_X1 FILLER_31_1061 ();
 FILLCELL_X4 FILLER_31_1066 ();
 FILLCELL_X16 FILLER_31_1074 ();
 FILLCELL_X4 FILLER_31_1090 ();
 FILLCELL_X2 FILLER_31_1094 ();
 FILLCELL_X8 FILLER_31_1105 ();
 FILLCELL_X1 FILLER_31_1113 ();
 FILLCELL_X4 FILLER_31_1123 ();
 FILLCELL_X2 FILLER_31_1127 ();
 FILLCELL_X4 FILLER_31_1132 ();
 FILLCELL_X16 FILLER_31_1140 ();
 FILLCELL_X8 FILLER_31_1156 ();
 FILLCELL_X2 FILLER_31_1164 ();
 FILLCELL_X1 FILLER_31_1166 ();
 FILLCELL_X4 FILLER_31_1172 ();
 FILLCELL_X4 FILLER_31_1180 ();
 FILLCELL_X4 FILLER_31_1188 ();
 FILLCELL_X8 FILLER_31_1196 ();
 FILLCELL_X2 FILLER_31_1204 ();
 FILLCELL_X1 FILLER_31_1206 ();
 FILLCELL_X4 FILLER_31_1212 ();
 FILLCELL_X4 FILLER_31_1221 ();
 FILLCELL_X4 FILLER_31_1234 ();
 FILLCELL_X1 FILLER_31_1238 ();
 FILLCELL_X4 FILLER_31_1244 ();
 FILLCELL_X4 FILLER_31_1252 ();
 FILLCELL_X4 FILLER_31_1259 ();
 FILLCELL_X4 FILLER_31_1264 ();
 FILLCELL_X4 FILLER_31_1273 ();
 FILLCELL_X2 FILLER_31_1277 ();
 FILLCELL_X8 FILLER_31_1288 ();
 FILLCELL_X1 FILLER_31_1296 ();
 FILLCELL_X4 FILLER_31_1316 ();
 FILLCELL_X1 FILLER_31_1320 ();
 FILLCELL_X32 FILLER_31_1325 ();
 FILLCELL_X16 FILLER_31_1357 ();
 FILLCELL_X2 FILLER_31_1373 ();
 FILLCELL_X32 FILLER_31_1394 ();
 FILLCELL_X32 FILLER_31_1426 ();
 FILLCELL_X32 FILLER_31_1458 ();
 FILLCELL_X32 FILLER_31_1490 ();
 FILLCELL_X32 FILLER_31_1522 ();
 FILLCELL_X32 FILLER_31_1558 ();
 FILLCELL_X32 FILLER_31_1590 ();
 FILLCELL_X32 FILLER_31_1622 ();
 FILLCELL_X32 FILLER_31_1654 ();
 FILLCELL_X8 FILLER_31_1686 ();
 FILLCELL_X4 FILLER_31_1694 ();
 FILLCELL_X2 FILLER_31_1698 ();
 FILLCELL_X1 FILLER_31_1700 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X32 FILLER_32_193 ();
 FILLCELL_X32 FILLER_32_225 ();
 FILLCELL_X32 FILLER_32_257 ();
 FILLCELL_X32 FILLER_32_289 ();
 FILLCELL_X32 FILLER_32_321 ();
 FILLCELL_X32 FILLER_32_353 ();
 FILLCELL_X16 FILLER_32_385 ();
 FILLCELL_X4 FILLER_32_401 ();
 FILLCELL_X2 FILLER_32_405 ();
 FILLCELL_X1 FILLER_32_407 ();
 FILLCELL_X16 FILLER_32_412 ();
 FILLCELL_X4 FILLER_32_428 ();
 FILLCELL_X4 FILLER_32_436 ();
 FILLCELL_X1 FILLER_32_440 ();
 FILLCELL_X4 FILLER_32_445 ();
 FILLCELL_X4 FILLER_32_466 ();
 FILLCELL_X8 FILLER_32_488 ();
 FILLCELL_X4 FILLER_32_496 ();
 FILLCELL_X4 FILLER_32_509 ();
 FILLCELL_X16 FILLER_32_517 ();
 FILLCELL_X4 FILLER_32_533 ();
 FILLCELL_X1 FILLER_32_537 ();
 FILLCELL_X4 FILLER_32_541 ();
 FILLCELL_X16 FILLER_32_555 ();
 FILLCELL_X8 FILLER_32_571 ();
 FILLCELL_X2 FILLER_32_579 ();
 FILLCELL_X1 FILLER_32_581 ();
 FILLCELL_X4 FILLER_32_591 ();
 FILLCELL_X2 FILLER_32_595 ();
 FILLCELL_X1 FILLER_32_597 ();
 FILLCELL_X4 FILLER_32_600 ();
 FILLCELL_X8 FILLER_32_621 ();
 FILLCELL_X2 FILLER_32_629 ();
 FILLCELL_X4 FILLER_32_632 ();
 FILLCELL_X16 FILLER_32_639 ();
 FILLCELL_X2 FILLER_32_655 ();
 FILLCELL_X1 FILLER_32_657 ();
 FILLCELL_X4 FILLER_32_677 ();
 FILLCELL_X2 FILLER_32_681 ();
 FILLCELL_X8 FILLER_32_702 ();
 FILLCELL_X8 FILLER_32_715 ();
 FILLCELL_X1 FILLER_32_723 ();
 FILLCELL_X8 FILLER_32_731 ();
 FILLCELL_X4 FILLER_32_744 ();
 FILLCELL_X4 FILLER_32_753 ();
 FILLCELL_X16 FILLER_32_761 ();
 FILLCELL_X8 FILLER_32_777 ();
 FILLCELL_X2 FILLER_32_785 ();
 FILLCELL_X1 FILLER_32_787 ();
 FILLCELL_X4 FILLER_32_806 ();
 FILLCELL_X4 FILLER_32_816 ();
 FILLCELL_X8 FILLER_32_825 ();
 FILLCELL_X4 FILLER_32_837 ();
 FILLCELL_X4 FILLER_32_846 ();
 FILLCELL_X4 FILLER_32_855 ();
 FILLCELL_X4 FILLER_32_864 ();
 FILLCELL_X32 FILLER_32_877 ();
 FILLCELL_X8 FILLER_32_909 ();
 FILLCELL_X1 FILLER_32_917 ();
 FILLCELL_X4 FILLER_32_922 ();
 FILLCELL_X4 FILLER_32_930 ();
 FILLCELL_X2 FILLER_32_934 ();
 FILLCELL_X1 FILLER_32_936 ();
 FILLCELL_X8 FILLER_32_946 ();
 FILLCELL_X4 FILLER_32_954 ();
 FILLCELL_X1 FILLER_32_958 ();
 FILLCELL_X32 FILLER_32_963 ();
 FILLCELL_X2 FILLER_32_995 ();
 FILLCELL_X1 FILLER_32_997 ();
 FILLCELL_X4 FILLER_32_1002 ();
 FILLCELL_X32 FILLER_32_1013 ();
 FILLCELL_X8 FILLER_32_1045 ();
 FILLCELL_X4 FILLER_32_1053 ();
 FILLCELL_X4 FILLER_32_1062 ();
 FILLCELL_X4 FILLER_32_1072 ();
 FILLCELL_X4 FILLER_32_1080 ();
 FILLCELL_X1 FILLER_32_1084 ();
 FILLCELL_X8 FILLER_32_1088 ();
 FILLCELL_X4 FILLER_32_1101 ();
 FILLCELL_X8 FILLER_32_1107 ();
 FILLCELL_X4 FILLER_32_1115 ();
 FILLCELL_X2 FILLER_32_1119 ();
 FILLCELL_X1 FILLER_32_1121 ();
 FILLCELL_X4 FILLER_32_1127 ();
 FILLCELL_X8 FILLER_32_1136 ();
 FILLCELL_X1 FILLER_32_1144 ();
 FILLCELL_X4 FILLER_32_1150 ();
 FILLCELL_X2 FILLER_32_1154 ();
 FILLCELL_X4 FILLER_32_1161 ();
 FILLCELL_X4 FILLER_32_1170 ();
 FILLCELL_X4 FILLER_32_1179 ();
 FILLCELL_X4 FILLER_32_1187 ();
 FILLCELL_X2 FILLER_32_1191 ();
 FILLCELL_X1 FILLER_32_1193 ();
 FILLCELL_X8 FILLER_32_1199 ();
 FILLCELL_X2 FILLER_32_1207 ();
 FILLCELL_X8 FILLER_32_1214 ();
 FILLCELL_X2 FILLER_32_1222 ();
 FILLCELL_X1 FILLER_32_1224 ();
 FILLCELL_X8 FILLER_32_1234 ();
 FILLCELL_X4 FILLER_32_1242 ();
 FILLCELL_X8 FILLER_32_1255 ();
 FILLCELL_X1 FILLER_32_1263 ();
 FILLCELL_X8 FILLER_32_1268 ();
 FILLCELL_X4 FILLER_32_1281 ();
 FILLCELL_X2 FILLER_32_1285 ();
 FILLCELL_X1 FILLER_32_1287 ();
 FILLCELL_X4 FILLER_32_1293 ();
 FILLCELL_X4 FILLER_32_1301 ();
 FILLCELL_X2 FILLER_32_1305 ();
 FILLCELL_X1 FILLER_32_1307 ();
 FILLCELL_X8 FILLER_32_1312 ();
 FILLCELL_X4 FILLER_32_1320 ();
 FILLCELL_X2 FILLER_32_1324 ();
 FILLCELL_X1 FILLER_32_1326 ();
 FILLCELL_X32 FILLER_32_1346 ();
 FILLCELL_X32 FILLER_32_1378 ();
 FILLCELL_X32 FILLER_32_1410 ();
 FILLCELL_X32 FILLER_32_1442 ();
 FILLCELL_X32 FILLER_32_1474 ();
 FILLCELL_X32 FILLER_32_1506 ();
 FILLCELL_X16 FILLER_32_1538 ();
 FILLCELL_X8 FILLER_32_1558 ();
 FILLCELL_X2 FILLER_32_1566 ();
 FILLCELL_X32 FILLER_32_1587 ();
 FILLCELL_X32 FILLER_32_1619 ();
 FILLCELL_X32 FILLER_32_1651 ();
 FILLCELL_X16 FILLER_32_1683 ();
 FILLCELL_X2 FILLER_32_1699 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X32 FILLER_33_193 ();
 FILLCELL_X32 FILLER_33_225 ();
 FILLCELL_X32 FILLER_33_257 ();
 FILLCELL_X32 FILLER_33_289 ();
 FILLCELL_X32 FILLER_33_321 ();
 FILLCELL_X16 FILLER_33_353 ();
 FILLCELL_X8 FILLER_33_369 ();
 FILLCELL_X8 FILLER_33_402 ();
 FILLCELL_X8 FILLER_33_429 ();
 FILLCELL_X2 FILLER_33_437 ();
 FILLCELL_X4 FILLER_33_458 ();
 FILLCELL_X2 FILLER_33_462 ();
 FILLCELL_X4 FILLER_33_471 ();
 FILLCELL_X4 FILLER_33_484 ();
 FILLCELL_X2 FILLER_33_488 ();
 FILLCELL_X1 FILLER_33_490 ();
 FILLCELL_X4 FILLER_33_498 ();
 FILLCELL_X8 FILLER_33_504 ();
 FILLCELL_X2 FILLER_33_512 ();
 FILLCELL_X8 FILLER_33_523 ();
 FILLCELL_X4 FILLER_33_531 ();
 FILLCELL_X2 FILLER_33_535 ();
 FILLCELL_X8 FILLER_33_544 ();
 FILLCELL_X2 FILLER_33_552 ();
 FILLCELL_X8 FILLER_33_563 ();
 FILLCELL_X4 FILLER_33_571 ();
 FILLCELL_X4 FILLER_33_579 ();
 FILLCELL_X4 FILLER_33_587 ();
 FILLCELL_X4 FILLER_33_595 ();
 FILLCELL_X4 FILLER_33_603 ();
 FILLCELL_X4 FILLER_33_626 ();
 FILLCELL_X4 FILLER_33_649 ();
 FILLCELL_X4 FILLER_33_672 ();
 FILLCELL_X8 FILLER_33_680 ();
 FILLCELL_X2 FILLER_33_688 ();
 FILLCELL_X8 FILLER_33_709 ();
 FILLCELL_X4 FILLER_33_717 ();
 FILLCELL_X1 FILLER_33_721 ();
 FILLCELL_X4 FILLER_33_728 ();
 FILLCELL_X2 FILLER_33_732 ();
 FILLCELL_X1 FILLER_33_734 ();
 FILLCELL_X16 FILLER_33_737 ();
 FILLCELL_X8 FILLER_33_753 ();
 FILLCELL_X1 FILLER_33_761 ();
 FILLCELL_X4 FILLER_33_767 ();
 FILLCELL_X16 FILLER_33_775 ();
 FILLCELL_X2 FILLER_33_791 ();
 FILLCELL_X1 FILLER_33_793 ();
 FILLCELL_X4 FILLER_33_812 ();
 FILLCELL_X4 FILLER_33_825 ();
 FILLCELL_X2 FILLER_33_829 ();
 FILLCELL_X1 FILLER_33_831 ();
 FILLCELL_X4 FILLER_33_835 ();
 FILLCELL_X4 FILLER_33_843 ();
 FILLCELL_X4 FILLER_33_852 ();
 FILLCELL_X2 FILLER_33_856 ();
 FILLCELL_X4 FILLER_33_862 ();
 FILLCELL_X4 FILLER_33_868 ();
 FILLCELL_X2 FILLER_33_872 ();
 FILLCELL_X1 FILLER_33_874 ();
 FILLCELL_X4 FILLER_33_880 ();
 FILLCELL_X2 FILLER_33_884 ();
 FILLCELL_X4 FILLER_33_895 ();
 FILLCELL_X4 FILLER_33_909 ();
 FILLCELL_X4 FILLER_33_918 ();
 FILLCELL_X1 FILLER_33_922 ();
 FILLCELL_X8 FILLER_33_926 ();
 FILLCELL_X2 FILLER_33_934 ();
 FILLCELL_X4 FILLER_33_949 ();
 FILLCELL_X4 FILLER_33_958 ();
 FILLCELL_X4 FILLER_33_964 ();
 FILLCELL_X1 FILLER_33_968 ();
 FILLCELL_X4 FILLER_33_976 ();
 FILLCELL_X4 FILLER_33_987 ();
 FILLCELL_X8 FILLER_33_996 ();
 FILLCELL_X2 FILLER_33_1004 ();
 FILLCELL_X1 FILLER_33_1006 ();
 FILLCELL_X4 FILLER_33_1016 ();
 FILLCELL_X1 FILLER_33_1020 ();
 FILLCELL_X8 FILLER_33_1030 ();
 FILLCELL_X2 FILLER_33_1038 ();
 FILLCELL_X1 FILLER_33_1040 ();
 FILLCELL_X4 FILLER_33_1051 ();
 FILLCELL_X4 FILLER_33_1065 ();
 FILLCELL_X8 FILLER_33_1078 ();
 FILLCELL_X2 FILLER_33_1086 ();
 FILLCELL_X4 FILLER_33_1093 ();
 FILLCELL_X8 FILLER_33_1106 ();
 FILLCELL_X4 FILLER_33_1114 ();
 FILLCELL_X1 FILLER_33_1118 ();
 FILLCELL_X4 FILLER_33_1123 ();
 FILLCELL_X4 FILLER_33_1129 ();
 FILLCELL_X8 FILLER_33_1135 ();
 FILLCELL_X4 FILLER_33_1143 ();
 FILLCELL_X4 FILLER_33_1152 ();
 FILLCELL_X4 FILLER_33_1161 ();
 FILLCELL_X4 FILLER_33_1170 ();
 FILLCELL_X4 FILLER_33_1178 ();
 FILLCELL_X8 FILLER_33_1186 ();
 FILLCELL_X1 FILLER_33_1194 ();
 FILLCELL_X4 FILLER_33_1204 ();
 FILLCELL_X16 FILLER_33_1212 ();
 FILLCELL_X8 FILLER_33_1228 ();
 FILLCELL_X4 FILLER_33_1236 ();
 FILLCELL_X2 FILLER_33_1240 ();
 FILLCELL_X1 FILLER_33_1242 ();
 FILLCELL_X4 FILLER_33_1245 ();
 FILLCELL_X4 FILLER_33_1251 ();
 FILLCELL_X2 FILLER_33_1255 ();
 FILLCELL_X4 FILLER_33_1259 ();
 FILLCELL_X4 FILLER_33_1264 ();
 FILLCELL_X4 FILLER_33_1272 ();
 FILLCELL_X4 FILLER_33_1278 ();
 FILLCELL_X4 FILLER_33_1285 ();
 FILLCELL_X1 FILLER_33_1289 ();
 FILLCELL_X4 FILLER_33_1295 ();
 FILLCELL_X4 FILLER_33_1303 ();
 FILLCELL_X32 FILLER_33_1310 ();
 FILLCELL_X32 FILLER_33_1342 ();
 FILLCELL_X32 FILLER_33_1374 ();
 FILLCELL_X32 FILLER_33_1406 ();
 FILLCELL_X32 FILLER_33_1438 ();
 FILLCELL_X32 FILLER_33_1470 ();
 FILLCELL_X16 FILLER_33_1502 ();
 FILLCELL_X4 FILLER_33_1520 ();
 FILLCELL_X16 FILLER_33_1528 ();
 FILLCELL_X1 FILLER_33_1544 ();
 FILLCELL_X32 FILLER_33_1549 ();
 FILLCELL_X32 FILLER_33_1581 ();
 FILLCELL_X32 FILLER_33_1613 ();
 FILLCELL_X32 FILLER_33_1645 ();
 FILLCELL_X16 FILLER_33_1677 ();
 FILLCELL_X8 FILLER_33_1693 ();
 FILLCELL_X4 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_8 ();
 FILLCELL_X32 FILLER_34_40 ();
 FILLCELL_X32 FILLER_34_72 ();
 FILLCELL_X32 FILLER_34_104 ();
 FILLCELL_X32 FILLER_34_136 ();
 FILLCELL_X32 FILLER_34_168 ();
 FILLCELL_X32 FILLER_34_200 ();
 FILLCELL_X32 FILLER_34_232 ();
 FILLCELL_X32 FILLER_34_264 ();
 FILLCELL_X32 FILLER_34_296 ();
 FILLCELL_X32 FILLER_34_328 ();
 FILLCELL_X32 FILLER_34_360 ();
 FILLCELL_X32 FILLER_34_392 ();
 FILLCELL_X4 FILLER_34_443 ();
 FILLCELL_X1 FILLER_34_447 ();
 FILLCELL_X8 FILLER_34_452 ();
 FILLCELL_X4 FILLER_34_460 ();
 FILLCELL_X2 FILLER_34_464 ();
 FILLCELL_X4 FILLER_34_468 ();
 FILLCELL_X4 FILLER_34_475 ();
 FILLCELL_X4 FILLER_34_486 ();
 FILLCELL_X4 FILLER_34_492 ();
 FILLCELL_X4 FILLER_34_499 ();
 FILLCELL_X4 FILLER_34_508 ();
 FILLCELL_X8 FILLER_34_516 ();
 FILLCELL_X1 FILLER_34_524 ();
 FILLCELL_X4 FILLER_34_539 ();
 FILLCELL_X4 FILLER_34_552 ();
 FILLCELL_X4 FILLER_34_559 ();
 FILLCELL_X4 FILLER_34_565 ();
 FILLCELL_X2 FILLER_34_569 ();
 FILLCELL_X1 FILLER_34_571 ();
 FILLCELL_X8 FILLER_34_579 ();
 FILLCELL_X1 FILLER_34_587 ();
 FILLCELL_X4 FILLER_34_592 ();
 FILLCELL_X2 FILLER_34_596 ();
 FILLCELL_X1 FILLER_34_598 ();
 FILLCELL_X4 FILLER_34_602 ();
 FILLCELL_X1 FILLER_34_606 ();
 FILLCELL_X16 FILLER_34_612 ();
 FILLCELL_X2 FILLER_34_628 ();
 FILLCELL_X1 FILLER_34_630 ();
 FILLCELL_X16 FILLER_34_632 ();
 FILLCELL_X1 FILLER_34_648 ();
 FILLCELL_X8 FILLER_34_652 ();
 FILLCELL_X1 FILLER_34_660 ();
 FILLCELL_X8 FILLER_34_680 ();
 FILLCELL_X16 FILLER_34_707 ();
 FILLCELL_X4 FILLER_34_723 ();
 FILLCELL_X4 FILLER_34_733 ();
 FILLCELL_X2 FILLER_34_737 ();
 FILLCELL_X1 FILLER_34_739 ();
 FILLCELL_X4 FILLER_34_759 ();
 FILLCELL_X16 FILLER_34_782 ();
 FILLCELL_X8 FILLER_34_798 ();
 FILLCELL_X1 FILLER_34_806 ();
 FILLCELL_X4 FILLER_34_809 ();
 FILLCELL_X8 FILLER_34_822 ();
 FILLCELL_X4 FILLER_34_832 ();
 FILLCELL_X2 FILLER_34_836 ();
 FILLCELL_X1 FILLER_34_838 ();
 FILLCELL_X4 FILLER_34_841 ();
 FILLCELL_X4 FILLER_34_847 ();
 FILLCELL_X4 FILLER_34_855 ();
 FILLCELL_X2 FILLER_34_859 ();
 FILLCELL_X4 FILLER_34_864 ();
 FILLCELL_X2 FILLER_34_868 ();
 FILLCELL_X4 FILLER_34_874 ();
 FILLCELL_X1 FILLER_34_878 ();
 FILLCELL_X8 FILLER_34_884 ();
 FILLCELL_X2 FILLER_34_892 ();
 FILLCELL_X8 FILLER_34_903 ();
 FILLCELL_X4 FILLER_34_911 ();
 FILLCELL_X2 FILLER_34_915 ();
 FILLCELL_X1 FILLER_34_917 ();
 FILLCELL_X4 FILLER_34_920 ();
 FILLCELL_X4 FILLER_34_933 ();
 FILLCELL_X8 FILLER_34_939 ();
 FILLCELL_X4 FILLER_34_947 ();
 FILLCELL_X8 FILLER_34_953 ();
 FILLCELL_X4 FILLER_34_961 ();
 FILLCELL_X1 FILLER_34_965 ();
 FILLCELL_X4 FILLER_34_984 ();
 FILLCELL_X4 FILLER_34_991 ();
 FILLCELL_X1 FILLER_34_995 ();
 FILLCELL_X16 FILLER_34_1005 ();
 FILLCELL_X4 FILLER_34_1031 ();
 FILLCELL_X4 FILLER_34_1045 ();
 FILLCELL_X4 FILLER_34_1055 ();
 FILLCELL_X4 FILLER_34_1065 ();
 FILLCELL_X2 FILLER_34_1069 ();
 FILLCELL_X4 FILLER_34_1073 ();
 FILLCELL_X4 FILLER_34_1082 ();
 FILLCELL_X8 FILLER_34_1090 ();
 FILLCELL_X4 FILLER_34_1102 ();
 FILLCELL_X8 FILLER_34_1108 ();
 FILLCELL_X4 FILLER_34_1116 ();
 FILLCELL_X1 FILLER_34_1120 ();
 FILLCELL_X4 FILLER_34_1130 ();
 FILLCELL_X4 FILLER_34_1138 ();
 FILLCELL_X16 FILLER_34_1144 ();
 FILLCELL_X1 FILLER_34_1160 ();
 FILLCELL_X16 FILLER_34_1166 ();
 FILLCELL_X4 FILLER_34_1182 ();
 FILLCELL_X2 FILLER_34_1186 ();
 FILLCELL_X1 FILLER_34_1188 ();
 FILLCELL_X8 FILLER_34_1193 ();
 FILLCELL_X4 FILLER_34_1205 ();
 FILLCELL_X8 FILLER_34_1213 ();
 FILLCELL_X4 FILLER_34_1221 ();
 FILLCELL_X4 FILLER_34_1230 ();
 FILLCELL_X4 FILLER_34_1238 ();
 FILLCELL_X4 FILLER_34_1245 ();
 FILLCELL_X1 FILLER_34_1249 ();
 FILLCELL_X4 FILLER_34_1254 ();
 FILLCELL_X4 FILLER_34_1260 ();
 FILLCELL_X2 FILLER_34_1264 ();
 FILLCELL_X4 FILLER_34_1270 ();
 FILLCELL_X4 FILLER_34_1278 ();
 FILLCELL_X8 FILLER_34_1285 ();
 FILLCELL_X4 FILLER_34_1298 ();
 FILLCELL_X4 FILLER_34_1304 ();
 FILLCELL_X2 FILLER_34_1308 ();
 FILLCELL_X32 FILLER_34_1329 ();
 FILLCELL_X32 FILLER_34_1361 ();
 FILLCELL_X32 FILLER_34_1393 ();
 FILLCELL_X32 FILLER_34_1425 ();
 FILLCELL_X32 FILLER_34_1457 ();
 FILLCELL_X32 FILLER_34_1489 ();
 FILLCELL_X8 FILLER_34_1521 ();
 FILLCELL_X4 FILLER_34_1529 ();
 FILLCELL_X4 FILLER_34_1537 ();
 FILLCELL_X16 FILLER_34_1545 ();
 FILLCELL_X1 FILLER_34_1561 ();
 FILLCELL_X32 FILLER_34_1579 ();
 FILLCELL_X32 FILLER_34_1611 ();
 FILLCELL_X32 FILLER_34_1643 ();
 FILLCELL_X16 FILLER_34_1675 ();
 FILLCELL_X8 FILLER_34_1691 ();
 FILLCELL_X2 FILLER_34_1699 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X32 FILLER_35_161 ();
 FILLCELL_X32 FILLER_35_193 ();
 FILLCELL_X32 FILLER_35_225 ();
 FILLCELL_X32 FILLER_35_257 ();
 FILLCELL_X32 FILLER_35_289 ();
 FILLCELL_X32 FILLER_35_321 ();
 FILLCELL_X32 FILLER_35_353 ();
 FILLCELL_X32 FILLER_35_385 ();
 FILLCELL_X16 FILLER_35_417 ();
 FILLCELL_X8 FILLER_35_433 ();
 FILLCELL_X4 FILLER_35_441 ();
 FILLCELL_X16 FILLER_35_449 ();
 FILLCELL_X1 FILLER_35_465 ();
 FILLCELL_X4 FILLER_35_469 ();
 FILLCELL_X4 FILLER_35_477 ();
 FILLCELL_X4 FILLER_35_485 ();
 FILLCELL_X2 FILLER_35_489 ();
 FILLCELL_X4 FILLER_35_497 ();
 FILLCELL_X2 FILLER_35_501 ();
 FILLCELL_X4 FILLER_35_520 ();
 FILLCELL_X8 FILLER_35_531 ();
 FILLCELL_X2 FILLER_35_539 ();
 FILLCELL_X4 FILLER_35_546 ();
 FILLCELL_X8 FILLER_35_553 ();
 FILLCELL_X2 FILLER_35_561 ();
 FILLCELL_X1 FILLER_35_563 ();
 FILLCELL_X32 FILLER_35_568 ();
 FILLCELL_X1 FILLER_35_600 ();
 FILLCELL_X4 FILLER_35_620 ();
 FILLCELL_X4 FILLER_35_643 ();
 FILLCELL_X4 FILLER_35_651 ();
 FILLCELL_X8 FILLER_35_659 ();
 FILLCELL_X1 FILLER_35_667 ();
 FILLCELL_X4 FILLER_35_687 ();
 FILLCELL_X4 FILLER_35_695 ();
 FILLCELL_X1 FILLER_35_699 ();
 FILLCELL_X4 FILLER_35_719 ();
 FILLCELL_X2 FILLER_35_723 ();
 FILLCELL_X32 FILLER_35_744 ();
 FILLCELL_X32 FILLER_35_776 ();
 FILLCELL_X16 FILLER_35_808 ();
 FILLCELL_X4 FILLER_35_826 ();
 FILLCELL_X32 FILLER_35_832 ();
 FILLCELL_X4 FILLER_35_866 ();
 FILLCELL_X4 FILLER_35_875 ();
 FILLCELL_X4 FILLER_35_882 ();
 FILLCELL_X8 FILLER_35_891 ();
 FILLCELL_X1 FILLER_35_899 ();
 FILLCELL_X4 FILLER_35_909 ();
 FILLCELL_X4 FILLER_35_923 ();
 FILLCELL_X2 FILLER_35_927 ();
 FILLCELL_X1 FILLER_35_929 ();
 FILLCELL_X8 FILLER_35_940 ();
 FILLCELL_X4 FILLER_35_948 ();
 FILLCELL_X2 FILLER_35_952 ();
 FILLCELL_X1 FILLER_35_954 ();
 FILLCELL_X4 FILLER_35_964 ();
 FILLCELL_X8 FILLER_35_972 ();
 FILLCELL_X1 FILLER_35_980 ();
 FILLCELL_X4 FILLER_35_995 ();
 FILLCELL_X8 FILLER_35_1012 ();
 FILLCELL_X4 FILLER_35_1020 ();
 FILLCELL_X16 FILLER_35_1028 ();
 FILLCELL_X4 FILLER_35_1044 ();
 FILLCELL_X1 FILLER_35_1048 ();
 FILLCELL_X4 FILLER_35_1053 ();
 FILLCELL_X1 FILLER_35_1057 ();
 FILLCELL_X4 FILLER_35_1062 ();
 FILLCELL_X4 FILLER_35_1070 ();
 FILLCELL_X8 FILLER_35_1076 ();
 FILLCELL_X4 FILLER_35_1088 ();
 FILLCELL_X1 FILLER_35_1092 ();
 FILLCELL_X4 FILLER_35_1097 ();
 FILLCELL_X4 FILLER_35_1103 ();
 FILLCELL_X2 FILLER_35_1107 ();
 FILLCELL_X4 FILLER_35_1113 ();
 FILLCELL_X4 FILLER_35_1122 ();
 FILLCELL_X4 FILLER_35_1129 ();
 FILLCELL_X8 FILLER_35_1135 ();
 FILLCELL_X1 FILLER_35_1143 ();
 FILLCELL_X4 FILLER_35_1148 ();
 FILLCELL_X4 FILLER_35_1155 ();
 FILLCELL_X2 FILLER_35_1159 ();
 FILLCELL_X4 FILLER_35_1166 ();
 FILLCELL_X16 FILLER_35_1175 ();
 FILLCELL_X2 FILLER_35_1191 ();
 FILLCELL_X4 FILLER_35_1202 ();
 FILLCELL_X4 FILLER_35_1209 ();
 FILLCELL_X4 FILLER_35_1215 ();
 FILLCELL_X2 FILLER_35_1219 ();
 FILLCELL_X1 FILLER_35_1221 ();
 FILLCELL_X4 FILLER_35_1226 ();
 FILLCELL_X4 FILLER_35_1234 ();
 FILLCELL_X4 FILLER_35_1240 ();
 FILLCELL_X2 FILLER_35_1244 ();
 FILLCELL_X4 FILLER_35_1250 ();
 FILLCELL_X4 FILLER_35_1259 ();
 FILLCELL_X4 FILLER_35_1264 ();
 FILLCELL_X2 FILLER_35_1268 ();
 FILLCELL_X1 FILLER_35_1270 ();
 FILLCELL_X4 FILLER_35_1280 ();
 FILLCELL_X4 FILLER_35_1302 ();
 FILLCELL_X8 FILLER_35_1308 ();
 FILLCELL_X2 FILLER_35_1316 ();
 FILLCELL_X32 FILLER_35_1322 ();
 FILLCELL_X32 FILLER_35_1354 ();
 FILLCELL_X32 FILLER_35_1386 ();
 FILLCELL_X32 FILLER_35_1418 ();
 FILLCELL_X32 FILLER_35_1450 ();
 FILLCELL_X32 FILLER_35_1482 ();
 FILLCELL_X32 FILLER_35_1514 ();
 FILLCELL_X1 FILLER_35_1546 ();
 FILLCELL_X32 FILLER_35_1564 ();
 FILLCELL_X32 FILLER_35_1596 ();
 FILLCELL_X32 FILLER_35_1628 ();
 FILLCELL_X32 FILLER_35_1660 ();
 FILLCELL_X8 FILLER_35_1692 ();
 FILLCELL_X1 FILLER_35_1700 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X32 FILLER_36_161 ();
 FILLCELL_X32 FILLER_36_193 ();
 FILLCELL_X32 FILLER_36_225 ();
 FILLCELL_X32 FILLER_36_257 ();
 FILLCELL_X32 FILLER_36_289 ();
 FILLCELL_X32 FILLER_36_321 ();
 FILLCELL_X32 FILLER_36_353 ();
 FILLCELL_X32 FILLER_36_385 ();
 FILLCELL_X32 FILLER_36_417 ();
 FILLCELL_X16 FILLER_36_449 ();
 FILLCELL_X4 FILLER_36_465 ();
 FILLCELL_X2 FILLER_36_469 ();
 FILLCELL_X16 FILLER_36_490 ();
 FILLCELL_X4 FILLER_36_506 ();
 FILLCELL_X1 FILLER_36_510 ();
 FILLCELL_X8 FILLER_36_515 ();
 FILLCELL_X4 FILLER_36_527 ();
 FILLCELL_X4 FILLER_36_538 ();
 FILLCELL_X4 FILLER_36_545 ();
 FILLCELL_X1 FILLER_36_549 ();
 FILLCELL_X4 FILLER_36_569 ();
 FILLCELL_X8 FILLER_36_592 ();
 FILLCELL_X2 FILLER_36_600 ();
 FILLCELL_X16 FILLER_36_606 ();
 FILLCELL_X8 FILLER_36_622 ();
 FILLCELL_X1 FILLER_36_630 ();
 FILLCELL_X16 FILLER_36_632 ();
 FILLCELL_X2 FILLER_36_648 ();
 FILLCELL_X1 FILLER_36_650 ();
 FILLCELL_X8 FILLER_36_655 ();
 FILLCELL_X4 FILLER_36_663 ();
 FILLCELL_X2 FILLER_36_667 ();
 FILLCELL_X4 FILLER_36_672 ();
 FILLCELL_X2 FILLER_36_676 ();
 FILLCELL_X1 FILLER_36_678 ();
 FILLCELL_X4 FILLER_36_698 ();
 FILLCELL_X1 FILLER_36_702 ();
 FILLCELL_X16 FILLER_36_708 ();
 FILLCELL_X2 FILLER_36_724 ();
 FILLCELL_X1 FILLER_36_726 ();
 FILLCELL_X8 FILLER_36_731 ();
 FILLCELL_X2 FILLER_36_739 ();
 FILLCELL_X4 FILLER_36_745 ();
 FILLCELL_X1 FILLER_36_749 ();
 FILLCELL_X4 FILLER_36_754 ();
 FILLCELL_X8 FILLER_36_777 ();
 FILLCELL_X4 FILLER_36_785 ();
 FILLCELL_X2 FILLER_36_789 ();
 FILLCELL_X1 FILLER_36_791 ();
 FILLCELL_X4 FILLER_36_811 ();
 FILLCELL_X8 FILLER_36_834 ();
 FILLCELL_X2 FILLER_36_842 ();
 FILLCELL_X1 FILLER_36_844 ();
 FILLCELL_X8 FILLER_36_863 ();
 FILLCELL_X2 FILLER_36_871 ();
 FILLCELL_X4 FILLER_36_875 ();
 FILLCELL_X4 FILLER_36_883 ();
 FILLCELL_X2 FILLER_36_887 ();
 FILLCELL_X1 FILLER_36_889 ();
 FILLCELL_X4 FILLER_36_894 ();
 FILLCELL_X2 FILLER_36_898 ();
 FILLCELL_X1 FILLER_36_900 ();
 FILLCELL_X4 FILLER_36_906 ();
 FILLCELL_X8 FILLER_36_915 ();
 FILLCELL_X1 FILLER_36_923 ();
 FILLCELL_X4 FILLER_36_927 ();
 FILLCELL_X1 FILLER_36_931 ();
 FILLCELL_X8 FILLER_36_936 ();
 FILLCELL_X2 FILLER_36_944 ();
 FILLCELL_X4 FILLER_36_949 ();
 FILLCELL_X4 FILLER_36_957 ();
 FILLCELL_X4 FILLER_36_965 ();
 FILLCELL_X2 FILLER_36_969 ();
 FILLCELL_X1 FILLER_36_971 ();
 FILLCELL_X16 FILLER_36_976 ();
 FILLCELL_X2 FILLER_36_992 ();
 FILLCELL_X4 FILLER_36_1001 ();
 FILLCELL_X8 FILLER_36_1009 ();
 FILLCELL_X2 FILLER_36_1017 ();
 FILLCELL_X4 FILLER_36_1024 ();
 FILLCELL_X8 FILLER_36_1030 ();
 FILLCELL_X2 FILLER_36_1038 ();
 FILLCELL_X4 FILLER_36_1044 ();
 FILLCELL_X4 FILLER_36_1052 ();
 FILLCELL_X4 FILLER_36_1061 ();
 FILLCELL_X8 FILLER_36_1070 ();
 FILLCELL_X1 FILLER_36_1078 ();
 FILLCELL_X4 FILLER_36_1083 ();
 FILLCELL_X8 FILLER_36_1094 ();
 FILLCELL_X4 FILLER_36_1105 ();
 FILLCELL_X8 FILLER_36_1116 ();
 FILLCELL_X4 FILLER_36_1124 ();
 FILLCELL_X2 FILLER_36_1128 ();
 FILLCELL_X1 FILLER_36_1130 ();
 FILLCELL_X4 FILLER_36_1135 ();
 FILLCELL_X16 FILLER_36_1143 ();
 FILLCELL_X4 FILLER_36_1163 ();
 FILLCELL_X4 FILLER_36_1172 ();
 FILLCELL_X8 FILLER_36_1180 ();
 FILLCELL_X1 FILLER_36_1188 ();
 FILLCELL_X4 FILLER_36_1191 ();
 FILLCELL_X4 FILLER_36_1200 ();
 FILLCELL_X4 FILLER_36_1208 ();
 FILLCELL_X2 FILLER_36_1212 ();
 FILLCELL_X4 FILLER_36_1223 ();
 FILLCELL_X4 FILLER_36_1232 ();
 FILLCELL_X4 FILLER_36_1240 ();
 FILLCELL_X4 FILLER_36_1250 ();
 FILLCELL_X8 FILLER_36_1263 ();
 FILLCELL_X8 FILLER_36_1273 ();
 FILLCELL_X1 FILLER_36_1281 ();
 FILLCELL_X8 FILLER_36_1284 ();
 FILLCELL_X1 FILLER_36_1292 ();
 FILLCELL_X32 FILLER_36_1295 ();
 FILLCELL_X32 FILLER_36_1327 ();
 FILLCELL_X32 FILLER_36_1359 ();
 FILLCELL_X32 FILLER_36_1391 ();
 FILLCELL_X32 FILLER_36_1423 ();
 FILLCELL_X32 FILLER_36_1455 ();
 FILLCELL_X32 FILLER_36_1487 ();
 FILLCELL_X32 FILLER_36_1519 ();
 FILLCELL_X32 FILLER_36_1551 ();
 FILLCELL_X32 FILLER_36_1583 ();
 FILLCELL_X32 FILLER_36_1615 ();
 FILLCELL_X32 FILLER_36_1647 ();
 FILLCELL_X16 FILLER_36_1679 ();
 FILLCELL_X4 FILLER_36_1695 ();
 FILLCELL_X2 FILLER_36_1699 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X32 FILLER_37_161 ();
 FILLCELL_X32 FILLER_37_193 ();
 FILLCELL_X32 FILLER_37_225 ();
 FILLCELL_X32 FILLER_37_257 ();
 FILLCELL_X32 FILLER_37_289 ();
 FILLCELL_X32 FILLER_37_321 ();
 FILLCELL_X32 FILLER_37_353 ();
 FILLCELL_X32 FILLER_37_385 ();
 FILLCELL_X16 FILLER_37_417 ();
 FILLCELL_X8 FILLER_37_433 ();
 FILLCELL_X2 FILLER_37_441 ();
 FILLCELL_X8 FILLER_37_460 ();
 FILLCELL_X4 FILLER_37_468 ();
 FILLCELL_X16 FILLER_37_476 ();
 FILLCELL_X1 FILLER_37_492 ();
 FILLCELL_X16 FILLER_37_497 ();
 FILLCELL_X1 FILLER_37_513 ();
 FILLCELL_X4 FILLER_37_523 ();
 FILLCELL_X8 FILLER_37_540 ();
 FILLCELL_X4 FILLER_37_548 ();
 FILLCELL_X2 FILLER_37_552 ();
 FILLCELL_X1 FILLER_37_554 ();
 FILLCELL_X4 FILLER_37_574 ();
 FILLCELL_X4 FILLER_37_597 ();
 FILLCELL_X4 FILLER_37_620 ();
 FILLCELL_X32 FILLER_37_643 ();
 FILLCELL_X8 FILLER_37_675 ();
 FILLCELL_X4 FILLER_37_687 ();
 FILLCELL_X2 FILLER_37_691 ();
 FILLCELL_X1 FILLER_37_693 ();
 FILLCELL_X4 FILLER_37_713 ();
 FILLCELL_X4 FILLER_37_736 ();
 FILLCELL_X4 FILLER_37_759 ();
 FILLCELL_X4 FILLER_37_782 ();
 FILLCELL_X8 FILLER_37_805 ();
 FILLCELL_X1 FILLER_37_813 ();
 FILLCELL_X4 FILLER_37_833 ();
 FILLCELL_X16 FILLER_37_856 ();
 FILLCELL_X8 FILLER_37_872 ();
 FILLCELL_X4 FILLER_37_880 ();
 FILLCELL_X4 FILLER_37_886 ();
 FILLCELL_X8 FILLER_37_893 ();
 FILLCELL_X4 FILLER_37_906 ();
 FILLCELL_X4 FILLER_37_914 ();
 FILLCELL_X1 FILLER_37_918 ();
 FILLCELL_X4 FILLER_37_923 ();
 FILLCELL_X4 FILLER_37_946 ();
 FILLCELL_X2 FILLER_37_950 ();
 FILLCELL_X4 FILLER_37_956 ();
 FILLCELL_X8 FILLER_37_964 ();
 FILLCELL_X4 FILLER_37_997 ();
 FILLCELL_X2 FILLER_37_1001 ();
 FILLCELL_X4 FILLER_37_1022 ();
 FILLCELL_X2 FILLER_37_1026 ();
 FILLCELL_X1 FILLER_37_1028 ();
 FILLCELL_X4 FILLER_37_1031 ();
 FILLCELL_X4 FILLER_37_1041 ();
 FILLCELL_X4 FILLER_37_1049 ();
 FILLCELL_X1 FILLER_37_1053 ();
 FILLCELL_X4 FILLER_37_1057 ();
 FILLCELL_X4 FILLER_37_1067 ();
 FILLCELL_X16 FILLER_37_1076 ();
 FILLCELL_X2 FILLER_37_1092 ();
 FILLCELL_X1 FILLER_37_1094 ();
 FILLCELL_X4 FILLER_37_1114 ();
 FILLCELL_X8 FILLER_37_1122 ();
 FILLCELL_X4 FILLER_37_1130 ();
 FILLCELL_X1 FILLER_37_1134 ();
 FILLCELL_X4 FILLER_37_1154 ();
 FILLCELL_X4 FILLER_37_1177 ();
 FILLCELL_X8 FILLER_37_1184 ();
 FILLCELL_X2 FILLER_37_1192 ();
 FILLCELL_X4 FILLER_37_1196 ();
 FILLCELL_X2 FILLER_37_1200 ();
 FILLCELL_X8 FILLER_37_1220 ();
 FILLCELL_X4 FILLER_37_1246 ();
 FILLCELL_X4 FILLER_37_1252 ();
 FILLCELL_X4 FILLER_37_1258 ();
 FILLCELL_X1 FILLER_37_1262 ();
 FILLCELL_X4 FILLER_37_1264 ();
 FILLCELL_X4 FILLER_37_1272 ();
 FILLCELL_X4 FILLER_37_1295 ();
 FILLCELL_X32 FILLER_37_1303 ();
 FILLCELL_X4 FILLER_37_1335 ();
 FILLCELL_X2 FILLER_37_1339 ();
 FILLCELL_X8 FILLER_37_1346 ();
 FILLCELL_X4 FILLER_37_1354 ();
 FILLCELL_X2 FILLER_37_1358 ();
 FILLCELL_X32 FILLER_37_1363 ();
 FILLCELL_X32 FILLER_37_1395 ();
 FILLCELL_X32 FILLER_37_1427 ();
 FILLCELL_X16 FILLER_37_1459 ();
 FILLCELL_X2 FILLER_37_1475 ();
 FILLCELL_X1 FILLER_37_1477 ();
 FILLCELL_X4 FILLER_37_1483 ();
 FILLCELL_X32 FILLER_37_1490 ();
 FILLCELL_X32 FILLER_37_1522 ();
 FILLCELL_X32 FILLER_37_1554 ();
 FILLCELL_X32 FILLER_37_1586 ();
 FILLCELL_X32 FILLER_37_1618 ();
 FILLCELL_X32 FILLER_37_1650 ();
 FILLCELL_X16 FILLER_37_1682 ();
 FILLCELL_X2 FILLER_37_1698 ();
 FILLCELL_X1 FILLER_37_1700 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X32 FILLER_38_161 ();
 FILLCELL_X32 FILLER_38_193 ();
 FILLCELL_X32 FILLER_38_225 ();
 FILLCELL_X32 FILLER_38_257 ();
 FILLCELL_X32 FILLER_38_289 ();
 FILLCELL_X32 FILLER_38_321 ();
 FILLCELL_X16 FILLER_38_353 ();
 FILLCELL_X1 FILLER_38_369 ();
 FILLCELL_X32 FILLER_38_395 ();
 FILLCELL_X2 FILLER_38_427 ();
 FILLCELL_X1 FILLER_38_429 ();
 FILLCELL_X8 FILLER_38_434 ();
 FILLCELL_X1 FILLER_38_442 ();
 FILLCELL_X16 FILLER_38_447 ();
 FILLCELL_X4 FILLER_38_463 ();
 FILLCELL_X2 FILLER_38_467 ();
 FILLCELL_X1 FILLER_38_469 ();
 FILLCELL_X4 FILLER_38_489 ();
 FILLCELL_X1 FILLER_38_493 ();
 FILLCELL_X8 FILLER_38_513 ();
 FILLCELL_X4 FILLER_38_521 ();
 FILLCELL_X2 FILLER_38_525 ();
 FILLCELL_X1 FILLER_38_527 ();
 FILLCELL_X8 FILLER_38_531 ();
 FILLCELL_X4 FILLER_38_539 ();
 FILLCELL_X2 FILLER_38_543 ();
 FILLCELL_X16 FILLER_38_564 ();
 FILLCELL_X1 FILLER_38_580 ();
 FILLCELL_X8 FILLER_38_584 ();
 FILLCELL_X4 FILLER_38_592 ();
 FILLCELL_X2 FILLER_38_596 ();
 FILLCELL_X16 FILLER_38_601 ();
 FILLCELL_X4 FILLER_38_617 ();
 FILLCELL_X2 FILLER_38_621 ();
 FILLCELL_X4 FILLER_38_627 ();
 FILLCELL_X8 FILLER_38_632 ();
 FILLCELL_X2 FILLER_38_640 ();
 FILLCELL_X1 FILLER_38_642 ();
 FILLCELL_X4 FILLER_38_662 ();
 FILLCELL_X16 FILLER_38_670 ();
 FILLCELL_X4 FILLER_38_686 ();
 FILLCELL_X2 FILLER_38_690 ();
 FILLCELL_X4 FILLER_38_696 ();
 FILLCELL_X2 FILLER_38_700 ();
 FILLCELL_X4 FILLER_38_706 ();
 FILLCELL_X8 FILLER_38_714 ();
 FILLCELL_X8 FILLER_38_726 ();
 FILLCELL_X2 FILLER_38_734 ();
 FILLCELL_X16 FILLER_38_739 ();
 FILLCELL_X4 FILLER_38_755 ();
 FILLCELL_X4 FILLER_38_763 ();
 FILLCELL_X1 FILLER_38_767 ();
 FILLCELL_X8 FILLER_38_772 ();
 FILLCELL_X4 FILLER_38_784 ();
 FILLCELL_X8 FILLER_38_792 ();
 FILLCELL_X4 FILLER_38_800 ();
 FILLCELL_X2 FILLER_38_804 ();
 FILLCELL_X1 FILLER_38_806 ();
 FILLCELL_X32 FILLER_38_811 ();
 FILLCELL_X8 FILLER_38_843 ();
 FILLCELL_X2 FILLER_38_851 ();
 FILLCELL_X1 FILLER_38_853 ();
 FILLCELL_X16 FILLER_38_873 ();
 FILLCELL_X4 FILLER_38_889 ();
 FILLCELL_X1 FILLER_38_893 ();
 FILLCELL_X4 FILLER_38_896 ();
 FILLCELL_X4 FILLER_38_902 ();
 FILLCELL_X32 FILLER_38_908 ();
 FILLCELL_X16 FILLER_38_940 ();
 FILLCELL_X8 FILLER_38_956 ();
 FILLCELL_X32 FILLER_38_967 ();
 FILLCELL_X16 FILLER_38_999 ();
 FILLCELL_X4 FILLER_38_1015 ();
 FILLCELL_X16 FILLER_38_1023 ();
 FILLCELL_X4 FILLER_38_1042 ();
 FILLCELL_X2 FILLER_38_1046 ();
 FILLCELL_X1 FILLER_38_1048 ();
 FILLCELL_X4 FILLER_38_1051 ();
 FILLCELL_X2 FILLER_38_1055 ();
 FILLCELL_X8 FILLER_38_1059 ();
 FILLCELL_X4 FILLER_38_1067 ();
 FILLCELL_X2 FILLER_38_1071 ();
 FILLCELL_X16 FILLER_38_1092 ();
 FILLCELL_X8 FILLER_38_1108 ();
 FILLCELL_X2 FILLER_38_1116 ();
 FILLCELL_X1 FILLER_38_1118 ();
 FILLCELL_X16 FILLER_38_1138 ();
 FILLCELL_X1 FILLER_38_1154 ();
 FILLCELL_X4 FILLER_38_1158 ();
 FILLCELL_X4 FILLER_38_1164 ();
 FILLCELL_X4 FILLER_38_1170 ();
 FILLCELL_X2 FILLER_38_1174 ();
 FILLCELL_X16 FILLER_38_1195 ();
 FILLCELL_X8 FILLER_38_1211 ();
 FILLCELL_X2 FILLER_38_1219 ();
 FILLCELL_X4 FILLER_38_1223 ();
 FILLCELL_X8 FILLER_38_1246 ();
 FILLCELL_X8 FILLER_38_1273 ();
 FILLCELL_X2 FILLER_38_1281 ();
 FILLCELL_X1 FILLER_38_1283 ();
 FILLCELL_X4 FILLER_38_1287 ();
 FILLCELL_X1 FILLER_38_1291 ();
 FILLCELL_X4 FILLER_38_1311 ();
 FILLCELL_X4 FILLER_38_1334 ();
 FILLCELL_X8 FILLER_38_1357 ();
 FILLCELL_X4 FILLER_38_1368 ();
 FILLCELL_X32 FILLER_38_1375 ();
 FILLCELL_X32 FILLER_38_1407 ();
 FILLCELL_X32 FILLER_38_1439 ();
 FILLCELL_X32 FILLER_38_1471 ();
 FILLCELL_X32 FILLER_38_1503 ();
 FILLCELL_X32 FILLER_38_1535 ();
 FILLCELL_X32 FILLER_38_1567 ();
 FILLCELL_X32 FILLER_38_1599 ();
 FILLCELL_X32 FILLER_38_1631 ();
 FILLCELL_X32 FILLER_38_1663 ();
 FILLCELL_X4 FILLER_38_1695 ();
 FILLCELL_X2 FILLER_38_1699 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X32 FILLER_39_97 ();
 FILLCELL_X32 FILLER_39_129 ();
 FILLCELL_X32 FILLER_39_161 ();
 FILLCELL_X32 FILLER_39_193 ();
 FILLCELL_X32 FILLER_39_225 ();
 FILLCELL_X32 FILLER_39_257 ();
 FILLCELL_X32 FILLER_39_289 ();
 FILLCELL_X32 FILLER_39_321 ();
 FILLCELL_X32 FILLER_39_353 ();
 FILLCELL_X32 FILLER_39_385 ();
 FILLCELL_X4 FILLER_39_417 ();
 FILLCELL_X2 FILLER_39_421 ();
 FILLCELL_X1 FILLER_39_423 ();
 FILLCELL_X4 FILLER_39_443 ();
 FILLCELL_X4 FILLER_39_466 ();
 FILLCELL_X4 FILLER_39_475 ();
 FILLCELL_X4 FILLER_39_484 ();
 FILLCELL_X8 FILLER_39_491 ();
 FILLCELL_X1 FILLER_39_499 ();
 FILLCELL_X32 FILLER_39_503 ();
 FILLCELL_X4 FILLER_39_535 ();
 FILLCELL_X4 FILLER_39_542 ();
 FILLCELL_X4 FILLER_39_549 ();
 FILLCELL_X4 FILLER_39_558 ();
 FILLCELL_X4 FILLER_39_567 ();
 FILLCELL_X4 FILLER_39_575 ();
 FILLCELL_X4 FILLER_39_583 ();
 FILLCELL_X2 FILLER_39_587 ();
 FILLCELL_X8 FILLER_39_593 ();
 FILLCELL_X4 FILLER_39_601 ();
 FILLCELL_X1 FILLER_39_605 ();
 FILLCELL_X8 FILLER_39_610 ();
 FILLCELL_X2 FILLER_39_618 ();
 FILLCELL_X1 FILLER_39_620 ();
 FILLCELL_X4 FILLER_39_625 ();
 FILLCELL_X2 FILLER_39_629 ();
 FILLCELL_X4 FILLER_39_632 ();
 FILLCELL_X2 FILLER_39_636 ();
 FILLCELL_X4 FILLER_39_642 ();
 FILLCELL_X2 FILLER_39_646 ();
 FILLCELL_X16 FILLER_39_651 ();
 FILLCELL_X4 FILLER_39_667 ();
 FILLCELL_X1 FILLER_39_671 ();
 FILLCELL_X32 FILLER_39_676 ();
 FILLCELL_X4 FILLER_39_708 ();
 FILLCELL_X16 FILLER_39_715 ();
 FILLCELL_X4 FILLER_39_731 ();
 FILLCELL_X1 FILLER_39_735 ();
 FILLCELL_X4 FILLER_39_739 ();
 FILLCELL_X16 FILLER_39_747 ();
 FILLCELL_X4 FILLER_39_763 ();
 FILLCELL_X1 FILLER_39_767 ();
 FILLCELL_X32 FILLER_39_771 ();
 FILLCELL_X1 FILLER_39_803 ();
 FILLCELL_X8 FILLER_39_808 ();
 FILLCELL_X2 FILLER_39_816 ();
 FILLCELL_X4 FILLER_39_821 ();
 FILLCELL_X8 FILLER_39_829 ();
 FILLCELL_X4 FILLER_39_837 ();
 FILLCELL_X2 FILLER_39_841 ();
 FILLCELL_X8 FILLER_39_847 ();
 FILLCELL_X4 FILLER_39_855 ();
 FILLCELL_X32 FILLER_39_864 ();
 FILLCELL_X32 FILLER_39_896 ();
 FILLCELL_X4 FILLER_39_928 ();
 FILLCELL_X16 FILLER_39_937 ();
 FILLCELL_X8 FILLER_39_953 ();
 FILLCELL_X32 FILLER_39_964 ();
 FILLCELL_X8 FILLER_39_996 ();
 FILLCELL_X2 FILLER_39_1004 ();
 FILLCELL_X32 FILLER_39_1011 ();
 FILLCELL_X16 FILLER_39_1043 ();
 FILLCELL_X4 FILLER_39_1059 ();
 FILLCELL_X2 FILLER_39_1063 ();
 FILLCELL_X1 FILLER_39_1065 ();
 FILLCELL_X8 FILLER_39_1069 ();
 FILLCELL_X1 FILLER_39_1077 ();
 FILLCELL_X16 FILLER_39_1081 ();
 FILLCELL_X2 FILLER_39_1097 ();
 FILLCELL_X1 FILLER_39_1099 ();
 FILLCELL_X8 FILLER_39_1103 ();
 FILLCELL_X2 FILLER_39_1111 ();
 FILLCELL_X1 FILLER_39_1113 ();
 FILLCELL_X4 FILLER_39_1117 ();
 FILLCELL_X4 FILLER_39_1124 ();
 FILLCELL_X4 FILLER_39_1131 ();
 FILLCELL_X4 FILLER_39_1138 ();
 FILLCELL_X4 FILLER_39_1145 ();
 FILLCELL_X4 FILLER_39_1152 ();
 FILLCELL_X2 FILLER_39_1156 ();
 FILLCELL_X1 FILLER_39_1158 ();
 FILLCELL_X4 FILLER_39_1162 ();
 FILLCELL_X32 FILLER_39_1169 ();
 FILLCELL_X4 FILLER_39_1201 ();
 FILLCELL_X16 FILLER_39_1208 ();
 FILLCELL_X4 FILLER_39_1224 ();
 FILLCELL_X1 FILLER_39_1228 ();
 FILLCELL_X4 FILLER_39_1233 ();
 FILLCELL_X4 FILLER_39_1240 ();
 FILLCELL_X4 FILLER_39_1247 ();
 FILLCELL_X1 FILLER_39_1251 ();
 FILLCELL_X8 FILLER_39_1254 ();
 FILLCELL_X4 FILLER_39_1263 ();
 FILLCELL_X4 FILLER_39_1270 ();
 FILLCELL_X4 FILLER_39_1277 ();
 FILLCELL_X4 FILLER_39_1284 ();
 FILLCELL_X32 FILLER_39_1291 ();
 FILLCELL_X4 FILLER_39_1326 ();
 FILLCELL_X4 FILLER_39_1333 ();
 FILLCELL_X2 FILLER_39_1337 ();
 FILLCELL_X1 FILLER_39_1339 ();
 FILLCELL_X8 FILLER_39_1345 ();
 FILLCELL_X1 FILLER_39_1353 ();
 FILLCELL_X4 FILLER_39_1357 ();
 FILLCELL_X32 FILLER_39_1380 ();
 FILLCELL_X32 FILLER_39_1412 ();
 FILLCELL_X8 FILLER_39_1444 ();
 FILLCELL_X1 FILLER_39_1452 ();
 FILLCELL_X32 FILLER_39_1456 ();
 FILLCELL_X32 FILLER_39_1488 ();
 FILLCELL_X4 FILLER_39_1520 ();
 FILLCELL_X32 FILLER_39_1541 ();
 FILLCELL_X32 FILLER_39_1573 ();
 FILLCELL_X32 FILLER_39_1605 ();
 FILLCELL_X32 FILLER_39_1637 ();
 FILLCELL_X32 FILLER_39_1669 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X32 FILLER_40_97 ();
 FILLCELL_X32 FILLER_40_129 ();
 FILLCELL_X32 FILLER_40_161 ();
 FILLCELL_X32 FILLER_40_193 ();
 FILLCELL_X32 FILLER_40_225 ();
 FILLCELL_X32 FILLER_40_257 ();
 FILLCELL_X32 FILLER_40_289 ();
 FILLCELL_X32 FILLER_40_321 ();
 FILLCELL_X16 FILLER_40_353 ();
 FILLCELL_X8 FILLER_40_369 ();
 FILLCELL_X2 FILLER_40_377 ();
 FILLCELL_X1 FILLER_40_379 ();
 FILLCELL_X32 FILLER_40_1518 ();
 FILLCELL_X32 FILLER_40_1550 ();
 FILLCELL_X32 FILLER_40_1582 ();
 FILLCELL_X32 FILLER_40_1614 ();
 FILLCELL_X32 FILLER_40_1646 ();
 FILLCELL_X16 FILLER_40_1678 ();
 FILLCELL_X4 FILLER_40_1694 ();
 FILLCELL_X2 FILLER_40_1698 ();
 FILLCELL_X1 FILLER_40_1700 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X32 FILLER_41_97 ();
 FILLCELL_X32 FILLER_41_129 ();
 FILLCELL_X32 FILLER_41_161 ();
 FILLCELL_X32 FILLER_41_193 ();
 FILLCELL_X32 FILLER_41_225 ();
 FILLCELL_X32 FILLER_41_257 ();
 FILLCELL_X32 FILLER_41_289 ();
 FILLCELL_X32 FILLER_41_321 ();
 FILLCELL_X16 FILLER_41_353 ();
 FILLCELL_X8 FILLER_41_369 ();
 FILLCELL_X2 FILLER_41_377 ();
 FILLCELL_X1 FILLER_41_379 ();
 FILLCELL_X32 FILLER_41_1518 ();
 FILLCELL_X32 FILLER_41_1550 ();
 FILLCELL_X32 FILLER_41_1582 ();
 FILLCELL_X32 FILLER_41_1614 ();
 FILLCELL_X32 FILLER_41_1646 ();
 FILLCELL_X16 FILLER_41_1678 ();
 FILLCELL_X4 FILLER_41_1694 ();
 FILLCELL_X2 FILLER_41_1698 ();
 FILLCELL_X1 FILLER_41_1700 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X32 FILLER_42_65 ();
 FILLCELL_X32 FILLER_42_97 ();
 FILLCELL_X32 FILLER_42_129 ();
 FILLCELL_X32 FILLER_42_161 ();
 FILLCELL_X32 FILLER_42_193 ();
 FILLCELL_X32 FILLER_42_225 ();
 FILLCELL_X32 FILLER_42_257 ();
 FILLCELL_X32 FILLER_42_289 ();
 FILLCELL_X32 FILLER_42_321 ();
 FILLCELL_X16 FILLER_42_353 ();
 FILLCELL_X8 FILLER_42_369 ();
 FILLCELL_X2 FILLER_42_377 ();
 FILLCELL_X1 FILLER_42_379 ();
 FILLCELL_X4 FILLER_42_1518 ();
 FILLCELL_X32 FILLER_42_1541 ();
 FILLCELL_X32 FILLER_42_1573 ();
 FILLCELL_X32 FILLER_42_1605 ();
 FILLCELL_X32 FILLER_42_1637 ();
 FILLCELL_X32 FILLER_42_1669 ();
 FILLCELL_X4 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_9 ();
 FILLCELL_X32 FILLER_43_41 ();
 FILLCELL_X32 FILLER_43_73 ();
 FILLCELL_X32 FILLER_43_105 ();
 FILLCELL_X32 FILLER_43_137 ();
 FILLCELL_X32 FILLER_43_169 ();
 FILLCELL_X32 FILLER_43_201 ();
 FILLCELL_X32 FILLER_43_233 ();
 FILLCELL_X32 FILLER_43_265 ();
 FILLCELL_X32 FILLER_43_297 ();
 FILLCELL_X32 FILLER_43_329 ();
 FILLCELL_X16 FILLER_43_361 ();
 FILLCELL_X2 FILLER_43_377 ();
 FILLCELL_X1 FILLER_43_379 ();
 FILLCELL_X32 FILLER_43_1518 ();
 FILLCELL_X32 FILLER_43_1550 ();
 FILLCELL_X32 FILLER_43_1582 ();
 FILLCELL_X32 FILLER_43_1614 ();
 FILLCELL_X32 FILLER_43_1646 ();
 FILLCELL_X16 FILLER_43_1678 ();
 FILLCELL_X4 FILLER_43_1694 ();
 FILLCELL_X2 FILLER_43_1698 ();
 FILLCELL_X1 FILLER_43_1700 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X32 FILLER_44_33 ();
 FILLCELL_X32 FILLER_44_65 ();
 FILLCELL_X32 FILLER_44_97 ();
 FILLCELL_X32 FILLER_44_129 ();
 FILLCELL_X32 FILLER_44_161 ();
 FILLCELL_X32 FILLER_44_193 ();
 FILLCELL_X32 FILLER_44_225 ();
 FILLCELL_X32 FILLER_44_257 ();
 FILLCELL_X32 FILLER_44_289 ();
 FILLCELL_X32 FILLER_44_321 ();
 FILLCELL_X16 FILLER_44_353 ();
 FILLCELL_X8 FILLER_44_369 ();
 FILLCELL_X2 FILLER_44_377 ();
 FILLCELL_X1 FILLER_44_379 ();
 FILLCELL_X8 FILLER_44_1518 ();
 FILLCELL_X4 FILLER_44_1526 ();
 FILLCELL_X1 FILLER_44_1530 ();
 FILLCELL_X32 FILLER_44_1550 ();
 FILLCELL_X32 FILLER_44_1582 ();
 FILLCELL_X32 FILLER_44_1614 ();
 FILLCELL_X32 FILLER_44_1646 ();
 FILLCELL_X16 FILLER_44_1678 ();
 FILLCELL_X4 FILLER_44_1694 ();
 FILLCELL_X2 FILLER_44_1698 ();
 FILLCELL_X1 FILLER_44_1700 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X32 FILLER_45_33 ();
 FILLCELL_X32 FILLER_45_65 ();
 FILLCELL_X32 FILLER_45_97 ();
 FILLCELL_X32 FILLER_45_129 ();
 FILLCELL_X32 FILLER_45_161 ();
 FILLCELL_X32 FILLER_45_193 ();
 FILLCELL_X32 FILLER_45_225 ();
 FILLCELL_X32 FILLER_45_257 ();
 FILLCELL_X32 FILLER_45_289 ();
 FILLCELL_X32 FILLER_45_321 ();
 FILLCELL_X16 FILLER_45_353 ();
 FILLCELL_X8 FILLER_45_369 ();
 FILLCELL_X2 FILLER_45_377 ();
 FILLCELL_X1 FILLER_45_379 ();
 FILLCELL_X32 FILLER_45_1518 ();
 FILLCELL_X32 FILLER_45_1550 ();
 FILLCELL_X32 FILLER_45_1582 ();
 FILLCELL_X32 FILLER_45_1614 ();
 FILLCELL_X32 FILLER_45_1646 ();
 FILLCELL_X16 FILLER_45_1678 ();
 FILLCELL_X4 FILLER_45_1694 ();
 FILLCELL_X2 FILLER_45_1698 ();
 FILLCELL_X1 FILLER_45_1700 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X32 FILLER_46_33 ();
 FILLCELL_X32 FILLER_46_65 ();
 FILLCELL_X32 FILLER_46_97 ();
 FILLCELL_X32 FILLER_46_129 ();
 FILLCELL_X32 FILLER_46_161 ();
 FILLCELL_X32 FILLER_46_193 ();
 FILLCELL_X32 FILLER_46_225 ();
 FILLCELL_X32 FILLER_46_257 ();
 FILLCELL_X32 FILLER_46_289 ();
 FILLCELL_X32 FILLER_46_321 ();
 FILLCELL_X4 FILLER_46_353 ();
 FILLCELL_X4 FILLER_46_376 ();
 FILLCELL_X32 FILLER_46_1518 ();
 FILLCELL_X32 FILLER_46_1550 ();
 FILLCELL_X32 FILLER_46_1582 ();
 FILLCELL_X32 FILLER_46_1614 ();
 FILLCELL_X32 FILLER_46_1646 ();
 FILLCELL_X16 FILLER_46_1678 ();
 FILLCELL_X4 FILLER_46_1694 ();
 FILLCELL_X2 FILLER_46_1698 ();
 FILLCELL_X1 FILLER_46_1700 ();
 FILLCELL_X32 FILLER_47_1 ();
 FILLCELL_X32 FILLER_47_33 ();
 FILLCELL_X32 FILLER_47_65 ();
 FILLCELL_X32 FILLER_47_97 ();
 FILLCELL_X32 FILLER_47_129 ();
 FILLCELL_X32 FILLER_47_161 ();
 FILLCELL_X32 FILLER_47_193 ();
 FILLCELL_X32 FILLER_47_225 ();
 FILLCELL_X32 FILLER_47_257 ();
 FILLCELL_X32 FILLER_47_289 ();
 FILLCELL_X32 FILLER_47_321 ();
 FILLCELL_X16 FILLER_47_353 ();
 FILLCELL_X8 FILLER_47_369 ();
 FILLCELL_X2 FILLER_47_377 ();
 FILLCELL_X1 FILLER_47_379 ();
 FILLCELL_X4 FILLER_47_1518 ();
 FILLCELL_X32 FILLER_47_1525 ();
 FILLCELL_X32 FILLER_47_1557 ();
 FILLCELL_X32 FILLER_47_1589 ();
 FILLCELL_X32 FILLER_47_1621 ();
 FILLCELL_X32 FILLER_47_1653 ();
 FILLCELL_X8 FILLER_47_1685 ();
 FILLCELL_X1 FILLER_47_1693 ();
 FILLCELL_X4 FILLER_47_1697 ();
 FILLCELL_X32 FILLER_48_1 ();
 FILLCELL_X32 FILLER_48_33 ();
 FILLCELL_X32 FILLER_48_65 ();
 FILLCELL_X32 FILLER_48_97 ();
 FILLCELL_X32 FILLER_48_129 ();
 FILLCELL_X32 FILLER_48_161 ();
 FILLCELL_X32 FILLER_48_193 ();
 FILLCELL_X32 FILLER_48_225 ();
 FILLCELL_X32 FILLER_48_257 ();
 FILLCELL_X32 FILLER_48_289 ();
 FILLCELL_X32 FILLER_48_321 ();
 FILLCELL_X16 FILLER_48_353 ();
 FILLCELL_X8 FILLER_48_369 ();
 FILLCELL_X2 FILLER_48_377 ();
 FILLCELL_X1 FILLER_48_379 ();
 FILLCELL_X32 FILLER_48_1518 ();
 FILLCELL_X32 FILLER_48_1550 ();
 FILLCELL_X32 FILLER_48_1582 ();
 FILLCELL_X32 FILLER_48_1614 ();
 FILLCELL_X32 FILLER_48_1646 ();
 FILLCELL_X16 FILLER_48_1678 ();
 FILLCELL_X4 FILLER_48_1694 ();
 FILLCELL_X2 FILLER_48_1698 ();
 FILLCELL_X1 FILLER_48_1700 ();
 FILLCELL_X32 FILLER_49_1 ();
 FILLCELL_X32 FILLER_49_33 ();
 FILLCELL_X32 FILLER_49_65 ();
 FILLCELL_X32 FILLER_49_97 ();
 FILLCELL_X32 FILLER_49_129 ();
 FILLCELL_X32 FILLER_49_161 ();
 FILLCELL_X32 FILLER_49_193 ();
 FILLCELL_X32 FILLER_49_225 ();
 FILLCELL_X32 FILLER_49_257 ();
 FILLCELL_X32 FILLER_49_289 ();
 FILLCELL_X32 FILLER_49_321 ();
 FILLCELL_X16 FILLER_49_353 ();
 FILLCELL_X8 FILLER_49_369 ();
 FILLCELL_X2 FILLER_49_377 ();
 FILLCELL_X1 FILLER_49_379 ();
 FILLCELL_X32 FILLER_49_1518 ();
 FILLCELL_X32 FILLER_49_1550 ();
 FILLCELL_X32 FILLER_49_1582 ();
 FILLCELL_X32 FILLER_49_1614 ();
 FILLCELL_X32 FILLER_49_1646 ();
 FILLCELL_X16 FILLER_49_1678 ();
 FILLCELL_X4 FILLER_49_1694 ();
 FILLCELL_X2 FILLER_49_1698 ();
 FILLCELL_X1 FILLER_49_1700 ();
 FILLCELL_X32 FILLER_50_1 ();
 FILLCELL_X32 FILLER_50_33 ();
 FILLCELL_X32 FILLER_50_65 ();
 FILLCELL_X32 FILLER_50_97 ();
 FILLCELL_X32 FILLER_50_129 ();
 FILLCELL_X32 FILLER_50_161 ();
 FILLCELL_X32 FILLER_50_193 ();
 FILLCELL_X32 FILLER_50_225 ();
 FILLCELL_X32 FILLER_50_257 ();
 FILLCELL_X32 FILLER_50_289 ();
 FILLCELL_X32 FILLER_50_321 ();
 FILLCELL_X4 FILLER_50_353 ();
 FILLCELL_X4 FILLER_50_376 ();
 FILLCELL_X8 FILLER_50_1518 ();
 FILLCELL_X4 FILLER_50_1526 ();
 FILLCELL_X1 FILLER_50_1530 ();
 FILLCELL_X32 FILLER_50_1534 ();
 FILLCELL_X32 FILLER_50_1566 ();
 FILLCELL_X32 FILLER_50_1598 ();
 FILLCELL_X32 FILLER_50_1630 ();
 FILLCELL_X32 FILLER_50_1662 ();
 FILLCELL_X4 FILLER_50_1694 ();
 FILLCELL_X2 FILLER_50_1698 ();
 FILLCELL_X1 FILLER_50_1700 ();
 FILLCELL_X32 FILLER_51_1 ();
 FILLCELL_X32 FILLER_51_33 ();
 FILLCELL_X32 FILLER_51_65 ();
 FILLCELL_X32 FILLER_51_97 ();
 FILLCELL_X32 FILLER_51_129 ();
 FILLCELL_X32 FILLER_51_161 ();
 FILLCELL_X32 FILLER_51_193 ();
 FILLCELL_X32 FILLER_51_225 ();
 FILLCELL_X32 FILLER_51_257 ();
 FILLCELL_X32 FILLER_51_289 ();
 FILLCELL_X32 FILLER_51_321 ();
 FILLCELL_X16 FILLER_51_353 ();
 FILLCELL_X8 FILLER_51_369 ();
 FILLCELL_X2 FILLER_51_377 ();
 FILLCELL_X1 FILLER_51_379 ();
 FILLCELL_X4 FILLER_51_1518 ();
 FILLCELL_X32 FILLER_51_1541 ();
 FILLCELL_X32 FILLER_51_1573 ();
 FILLCELL_X32 FILLER_51_1605 ();
 FILLCELL_X32 FILLER_51_1637 ();
 FILLCELL_X32 FILLER_51_1669 ();
 FILLCELL_X4 FILLER_52_1 ();
 FILLCELL_X32 FILLER_52_8 ();
 FILLCELL_X32 FILLER_52_40 ();
 FILLCELL_X32 FILLER_52_72 ();
 FILLCELL_X32 FILLER_52_104 ();
 FILLCELL_X32 FILLER_52_136 ();
 FILLCELL_X32 FILLER_52_168 ();
 FILLCELL_X32 FILLER_52_200 ();
 FILLCELL_X32 FILLER_52_232 ();
 FILLCELL_X32 FILLER_52_264 ();
 FILLCELL_X32 FILLER_52_296 ();
 FILLCELL_X32 FILLER_52_328 ();
 FILLCELL_X16 FILLER_52_360 ();
 FILLCELL_X4 FILLER_52_376 ();
 FILLCELL_X4 FILLER_52_1518 ();
 FILLCELL_X32 FILLER_52_1526 ();
 FILLCELL_X32 FILLER_52_1558 ();
 FILLCELL_X32 FILLER_52_1590 ();
 FILLCELL_X32 FILLER_52_1622 ();
 FILLCELL_X32 FILLER_52_1654 ();
 FILLCELL_X8 FILLER_52_1686 ();
 FILLCELL_X4 FILLER_52_1694 ();
 FILLCELL_X2 FILLER_52_1698 ();
 FILLCELL_X1 FILLER_52_1700 ();
 FILLCELL_X32 FILLER_53_1 ();
 FILLCELL_X32 FILLER_53_33 ();
 FILLCELL_X32 FILLER_53_65 ();
 FILLCELL_X32 FILLER_53_97 ();
 FILLCELL_X32 FILLER_53_129 ();
 FILLCELL_X32 FILLER_53_161 ();
 FILLCELL_X32 FILLER_53_193 ();
 FILLCELL_X32 FILLER_53_225 ();
 FILLCELL_X32 FILLER_53_257 ();
 FILLCELL_X32 FILLER_53_289 ();
 FILLCELL_X32 FILLER_53_321 ();
 FILLCELL_X16 FILLER_53_353 ();
 FILLCELL_X8 FILLER_53_369 ();
 FILLCELL_X2 FILLER_53_377 ();
 FILLCELL_X1 FILLER_53_379 ();
 FILLCELL_X4 FILLER_53_1518 ();
 FILLCELL_X32 FILLER_53_1525 ();
 FILLCELL_X32 FILLER_53_1557 ();
 FILLCELL_X32 FILLER_53_1589 ();
 FILLCELL_X32 FILLER_53_1621 ();
 FILLCELL_X32 FILLER_53_1653 ();
 FILLCELL_X16 FILLER_53_1685 ();
 FILLCELL_X32 FILLER_54_1 ();
 FILLCELL_X32 FILLER_54_33 ();
 FILLCELL_X32 FILLER_54_65 ();
 FILLCELL_X32 FILLER_54_97 ();
 FILLCELL_X32 FILLER_54_129 ();
 FILLCELL_X32 FILLER_54_161 ();
 FILLCELL_X32 FILLER_54_193 ();
 FILLCELL_X32 FILLER_54_225 ();
 FILLCELL_X32 FILLER_54_257 ();
 FILLCELL_X32 FILLER_54_289 ();
 FILLCELL_X32 FILLER_54_321 ();
 FILLCELL_X16 FILLER_54_353 ();
 FILLCELL_X8 FILLER_54_369 ();
 FILLCELL_X2 FILLER_54_377 ();
 FILLCELL_X1 FILLER_54_379 ();
 FILLCELL_X4 FILLER_54_1518 ();
 FILLCELL_X32 FILLER_54_1527 ();
 FILLCELL_X32 FILLER_54_1559 ();
 FILLCELL_X32 FILLER_54_1591 ();
 FILLCELL_X32 FILLER_54_1623 ();
 FILLCELL_X32 FILLER_54_1655 ();
 FILLCELL_X8 FILLER_54_1687 ();
 FILLCELL_X4 FILLER_54_1695 ();
 FILLCELL_X2 FILLER_54_1699 ();
 FILLCELL_X32 FILLER_55_1 ();
 FILLCELL_X32 FILLER_55_33 ();
 FILLCELL_X32 FILLER_55_65 ();
 FILLCELL_X32 FILLER_55_97 ();
 FILLCELL_X32 FILLER_55_129 ();
 FILLCELL_X32 FILLER_55_161 ();
 FILLCELL_X32 FILLER_55_193 ();
 FILLCELL_X32 FILLER_55_225 ();
 FILLCELL_X32 FILLER_55_257 ();
 FILLCELL_X32 FILLER_55_289 ();
 FILLCELL_X32 FILLER_55_321 ();
 FILLCELL_X16 FILLER_55_353 ();
 FILLCELL_X8 FILLER_55_369 ();
 FILLCELL_X2 FILLER_55_377 ();
 FILLCELL_X1 FILLER_55_379 ();
 FILLCELL_X8 FILLER_55_1518 ();
 FILLCELL_X4 FILLER_55_1526 ();
 FILLCELL_X1 FILLER_55_1530 ();
 FILLCELL_X32 FILLER_55_1550 ();
 FILLCELL_X32 FILLER_55_1582 ();
 FILLCELL_X32 FILLER_55_1614 ();
 FILLCELL_X32 FILLER_55_1646 ();
 FILLCELL_X16 FILLER_55_1678 ();
 FILLCELL_X4 FILLER_55_1694 ();
 FILLCELL_X2 FILLER_55_1698 ();
 FILLCELL_X1 FILLER_55_1700 ();
 FILLCELL_X32 FILLER_56_1 ();
 FILLCELL_X32 FILLER_56_33 ();
 FILLCELL_X32 FILLER_56_65 ();
 FILLCELL_X32 FILLER_56_97 ();
 FILLCELL_X32 FILLER_56_129 ();
 FILLCELL_X32 FILLER_56_161 ();
 FILLCELL_X32 FILLER_56_193 ();
 FILLCELL_X32 FILLER_56_225 ();
 FILLCELL_X32 FILLER_56_257 ();
 FILLCELL_X32 FILLER_56_289 ();
 FILLCELL_X32 FILLER_56_321 ();
 FILLCELL_X16 FILLER_56_353 ();
 FILLCELL_X8 FILLER_56_369 ();
 FILLCELL_X2 FILLER_56_377 ();
 FILLCELL_X1 FILLER_56_379 ();
 FILLCELL_X32 FILLER_56_1518 ();
 FILLCELL_X32 FILLER_56_1550 ();
 FILLCELL_X32 FILLER_56_1582 ();
 FILLCELL_X32 FILLER_56_1614 ();
 FILLCELL_X32 FILLER_56_1646 ();
 FILLCELL_X16 FILLER_56_1678 ();
 FILLCELL_X4 FILLER_56_1694 ();
 FILLCELL_X2 FILLER_56_1698 ();
 FILLCELL_X1 FILLER_56_1700 ();
 FILLCELL_X32 FILLER_57_1 ();
 FILLCELL_X32 FILLER_57_33 ();
 FILLCELL_X32 FILLER_57_65 ();
 FILLCELL_X32 FILLER_57_97 ();
 FILLCELL_X32 FILLER_57_129 ();
 FILLCELL_X32 FILLER_57_161 ();
 FILLCELL_X32 FILLER_57_193 ();
 FILLCELL_X32 FILLER_57_225 ();
 FILLCELL_X32 FILLER_57_257 ();
 FILLCELL_X32 FILLER_57_289 ();
 FILLCELL_X32 FILLER_57_321 ();
 FILLCELL_X16 FILLER_57_353 ();
 FILLCELL_X8 FILLER_57_369 ();
 FILLCELL_X2 FILLER_57_377 ();
 FILLCELL_X1 FILLER_57_379 ();
 FILLCELL_X4 FILLER_57_1518 ();
 FILLCELL_X32 FILLER_57_1526 ();
 FILLCELL_X32 FILLER_57_1558 ();
 FILLCELL_X32 FILLER_57_1590 ();
 FILLCELL_X32 FILLER_57_1622 ();
 FILLCELL_X32 FILLER_57_1654 ();
 FILLCELL_X8 FILLER_57_1686 ();
 FILLCELL_X4 FILLER_57_1697 ();
 FILLCELL_X32 FILLER_58_1 ();
 FILLCELL_X32 FILLER_58_33 ();
 FILLCELL_X32 FILLER_58_65 ();
 FILLCELL_X32 FILLER_58_97 ();
 FILLCELL_X32 FILLER_58_129 ();
 FILLCELL_X32 FILLER_58_161 ();
 FILLCELL_X32 FILLER_58_193 ();
 FILLCELL_X32 FILLER_58_225 ();
 FILLCELL_X32 FILLER_58_257 ();
 FILLCELL_X32 FILLER_58_289 ();
 FILLCELL_X32 FILLER_58_321 ();
 FILLCELL_X16 FILLER_58_353 ();
 FILLCELL_X2 FILLER_58_369 ();
 FILLCELL_X4 FILLER_58_376 ();
 FILLCELL_X32 FILLER_58_1518 ();
 FILLCELL_X32 FILLER_58_1550 ();
 FILLCELL_X32 FILLER_58_1582 ();
 FILLCELL_X32 FILLER_58_1614 ();
 FILLCELL_X32 FILLER_58_1646 ();
 FILLCELL_X16 FILLER_58_1678 ();
 FILLCELL_X4 FILLER_58_1694 ();
 FILLCELL_X2 FILLER_58_1698 ();
 FILLCELL_X1 FILLER_58_1700 ();
 FILLCELL_X32 FILLER_59_1 ();
 FILLCELL_X32 FILLER_59_33 ();
 FILLCELL_X32 FILLER_59_65 ();
 FILLCELL_X32 FILLER_59_97 ();
 FILLCELL_X32 FILLER_59_129 ();
 FILLCELL_X32 FILLER_59_161 ();
 FILLCELL_X32 FILLER_59_193 ();
 FILLCELL_X32 FILLER_59_225 ();
 FILLCELL_X32 FILLER_59_257 ();
 FILLCELL_X32 FILLER_59_289 ();
 FILLCELL_X32 FILLER_59_321 ();
 FILLCELL_X16 FILLER_59_353 ();
 FILLCELL_X8 FILLER_59_369 ();
 FILLCELL_X2 FILLER_59_377 ();
 FILLCELL_X1 FILLER_59_379 ();
 FILLCELL_X4 FILLER_59_1518 ();
 FILLCELL_X32 FILLER_59_1541 ();
 FILLCELL_X32 FILLER_59_1573 ();
 FILLCELL_X32 FILLER_59_1605 ();
 FILLCELL_X32 FILLER_59_1637 ();
 FILLCELL_X32 FILLER_59_1669 ();
 FILLCELL_X32 FILLER_60_1 ();
 FILLCELL_X32 FILLER_60_33 ();
 FILLCELL_X32 FILLER_60_65 ();
 FILLCELL_X32 FILLER_60_97 ();
 FILLCELL_X32 FILLER_60_129 ();
 FILLCELL_X32 FILLER_60_161 ();
 FILLCELL_X32 FILLER_60_193 ();
 FILLCELL_X32 FILLER_60_225 ();
 FILLCELL_X32 FILLER_60_257 ();
 FILLCELL_X32 FILLER_60_289 ();
 FILLCELL_X32 FILLER_60_321 ();
 FILLCELL_X16 FILLER_60_353 ();
 FILLCELL_X2 FILLER_60_369 ();
 FILLCELL_X1 FILLER_60_371 ();
 FILLCELL_X4 FILLER_60_376 ();
 FILLCELL_X16 FILLER_60_1518 ();
 FILLCELL_X8 FILLER_60_1534 ();
 FILLCELL_X32 FILLER_60_1559 ();
 FILLCELL_X32 FILLER_60_1591 ();
 FILLCELL_X32 FILLER_60_1623 ();
 FILLCELL_X32 FILLER_60_1655 ();
 FILLCELL_X8 FILLER_60_1687 ();
 FILLCELL_X4 FILLER_60_1695 ();
 FILLCELL_X2 FILLER_60_1699 ();
 FILLCELL_X32 FILLER_61_1 ();
 FILLCELL_X32 FILLER_61_33 ();
 FILLCELL_X32 FILLER_61_65 ();
 FILLCELL_X32 FILLER_61_97 ();
 FILLCELL_X32 FILLER_61_129 ();
 FILLCELL_X32 FILLER_61_161 ();
 FILLCELL_X32 FILLER_61_193 ();
 FILLCELL_X32 FILLER_61_225 ();
 FILLCELL_X32 FILLER_61_257 ();
 FILLCELL_X32 FILLER_61_289 ();
 FILLCELL_X32 FILLER_61_321 ();
 FILLCELL_X4 FILLER_61_353 ();
 FILLCELL_X4 FILLER_61_376 ();
 FILLCELL_X4 FILLER_61_1518 ();
 FILLCELL_X32 FILLER_61_1524 ();
 FILLCELL_X32 FILLER_61_1556 ();
 FILLCELL_X32 FILLER_61_1588 ();
 FILLCELL_X32 FILLER_61_1620 ();
 FILLCELL_X32 FILLER_61_1652 ();
 FILLCELL_X16 FILLER_61_1684 ();
 FILLCELL_X1 FILLER_61_1700 ();
 FILLCELL_X4 FILLER_62_1 ();
 FILLCELL_X32 FILLER_62_12 ();
 FILLCELL_X32 FILLER_62_44 ();
 FILLCELL_X32 FILLER_62_76 ();
 FILLCELL_X32 FILLER_62_108 ();
 FILLCELL_X32 FILLER_62_140 ();
 FILLCELL_X32 FILLER_62_172 ();
 FILLCELL_X32 FILLER_62_204 ();
 FILLCELL_X32 FILLER_62_236 ();
 FILLCELL_X32 FILLER_62_268 ();
 FILLCELL_X32 FILLER_62_300 ();
 FILLCELL_X32 FILLER_62_332 ();
 FILLCELL_X4 FILLER_62_364 ();
 FILLCELL_X1 FILLER_62_368 ();
 FILLCELL_X4 FILLER_62_373 ();
 FILLCELL_X2 FILLER_62_377 ();
 FILLCELL_X1 FILLER_62_379 ();
 FILLCELL_X4 FILLER_62_1518 ();
 FILLCELL_X32 FILLER_62_1527 ();
 FILLCELL_X32 FILLER_62_1559 ();
 FILLCELL_X32 FILLER_62_1591 ();
 FILLCELL_X32 FILLER_62_1623 ();
 FILLCELL_X32 FILLER_62_1655 ();
 FILLCELL_X8 FILLER_62_1687 ();
 FILLCELL_X4 FILLER_62_1695 ();
 FILLCELL_X2 FILLER_62_1699 ();
 FILLCELL_X32 FILLER_63_1 ();
 FILLCELL_X32 FILLER_63_33 ();
 FILLCELL_X32 FILLER_63_65 ();
 FILLCELL_X32 FILLER_63_97 ();
 FILLCELL_X32 FILLER_63_129 ();
 FILLCELL_X32 FILLER_63_161 ();
 FILLCELL_X32 FILLER_63_193 ();
 FILLCELL_X32 FILLER_63_225 ();
 FILLCELL_X32 FILLER_63_257 ();
 FILLCELL_X32 FILLER_63_289 ();
 FILLCELL_X32 FILLER_63_321 ();
 FILLCELL_X16 FILLER_63_353 ();
 FILLCELL_X1 FILLER_63_369 ();
 FILLCELL_X4 FILLER_63_374 ();
 FILLCELL_X2 FILLER_63_378 ();
 FILLCELL_X32 FILLER_63_1518 ();
 FILLCELL_X32 FILLER_63_1550 ();
 FILLCELL_X32 FILLER_63_1582 ();
 FILLCELL_X32 FILLER_63_1614 ();
 FILLCELL_X32 FILLER_63_1646 ();
 FILLCELL_X16 FILLER_63_1678 ();
 FILLCELL_X4 FILLER_63_1694 ();
 FILLCELL_X2 FILLER_63_1698 ();
 FILLCELL_X1 FILLER_63_1700 ();
 FILLCELL_X32 FILLER_64_1 ();
 FILLCELL_X32 FILLER_64_33 ();
 FILLCELL_X32 FILLER_64_65 ();
 FILLCELL_X32 FILLER_64_97 ();
 FILLCELL_X32 FILLER_64_129 ();
 FILLCELL_X32 FILLER_64_161 ();
 FILLCELL_X32 FILLER_64_193 ();
 FILLCELL_X32 FILLER_64_225 ();
 FILLCELL_X32 FILLER_64_257 ();
 FILLCELL_X32 FILLER_64_289 ();
 FILLCELL_X32 FILLER_64_321 ();
 FILLCELL_X2 FILLER_64_353 ();
 FILLCELL_X1 FILLER_64_355 ();
 FILLCELL_X4 FILLER_64_375 ();
 FILLCELL_X1 FILLER_64_379 ();
 FILLCELL_X32 FILLER_64_1518 ();
 FILLCELL_X32 FILLER_64_1550 ();
 FILLCELL_X32 FILLER_64_1582 ();
 FILLCELL_X32 FILLER_64_1614 ();
 FILLCELL_X32 FILLER_64_1646 ();
 FILLCELL_X16 FILLER_64_1678 ();
 FILLCELL_X4 FILLER_64_1694 ();
 FILLCELL_X2 FILLER_64_1698 ();
 FILLCELL_X1 FILLER_64_1700 ();
 FILLCELL_X32 FILLER_65_1 ();
 FILLCELL_X32 FILLER_65_33 ();
 FILLCELL_X32 FILLER_65_65 ();
 FILLCELL_X32 FILLER_65_97 ();
 FILLCELL_X32 FILLER_65_129 ();
 FILLCELL_X32 FILLER_65_161 ();
 FILLCELL_X32 FILLER_65_193 ();
 FILLCELL_X32 FILLER_65_225 ();
 FILLCELL_X32 FILLER_65_257 ();
 FILLCELL_X32 FILLER_65_289 ();
 FILLCELL_X32 FILLER_65_321 ();
 FILLCELL_X4 FILLER_65_353 ();
 FILLCELL_X4 FILLER_65_376 ();
 FILLCELL_X32 FILLER_65_1518 ();
 FILLCELL_X32 FILLER_65_1550 ();
 FILLCELL_X32 FILLER_65_1582 ();
 FILLCELL_X32 FILLER_65_1614 ();
 FILLCELL_X32 FILLER_65_1646 ();
 FILLCELL_X16 FILLER_65_1678 ();
 FILLCELL_X4 FILLER_65_1694 ();
 FILLCELL_X2 FILLER_65_1698 ();
 FILLCELL_X1 FILLER_65_1700 ();
 FILLCELL_X32 FILLER_66_1 ();
 FILLCELL_X32 FILLER_66_33 ();
 FILLCELL_X32 FILLER_66_65 ();
 FILLCELL_X32 FILLER_66_97 ();
 FILLCELL_X32 FILLER_66_129 ();
 FILLCELL_X32 FILLER_66_161 ();
 FILLCELL_X32 FILLER_66_193 ();
 FILLCELL_X32 FILLER_66_225 ();
 FILLCELL_X32 FILLER_66_257 ();
 FILLCELL_X32 FILLER_66_289 ();
 FILLCELL_X32 FILLER_66_321 ();
 FILLCELL_X16 FILLER_66_353 ();
 FILLCELL_X4 FILLER_66_369 ();
 FILLCELL_X1 FILLER_66_373 ();
 FILLCELL_X4 FILLER_66_376 ();
 FILLCELL_X32 FILLER_66_1518 ();
 FILLCELL_X32 FILLER_66_1550 ();
 FILLCELL_X32 FILLER_66_1582 ();
 FILLCELL_X32 FILLER_66_1614 ();
 FILLCELL_X32 FILLER_66_1646 ();
 FILLCELL_X16 FILLER_66_1678 ();
 FILLCELL_X4 FILLER_66_1697 ();
 FILLCELL_X32 FILLER_67_1 ();
 FILLCELL_X32 FILLER_67_33 ();
 FILLCELL_X32 FILLER_67_65 ();
 FILLCELL_X32 FILLER_67_97 ();
 FILLCELL_X32 FILLER_67_129 ();
 FILLCELL_X32 FILLER_67_161 ();
 FILLCELL_X32 FILLER_67_193 ();
 FILLCELL_X32 FILLER_67_225 ();
 FILLCELL_X32 FILLER_67_257 ();
 FILLCELL_X32 FILLER_67_289 ();
 FILLCELL_X32 FILLER_67_321 ();
 FILLCELL_X16 FILLER_67_353 ();
 FILLCELL_X8 FILLER_67_369 ();
 FILLCELL_X2 FILLER_67_377 ();
 FILLCELL_X1 FILLER_67_379 ();
 FILLCELL_X32 FILLER_67_1518 ();
 FILLCELL_X32 FILLER_67_1550 ();
 FILLCELL_X32 FILLER_67_1582 ();
 FILLCELL_X32 FILLER_67_1614 ();
 FILLCELL_X32 FILLER_67_1646 ();
 FILLCELL_X16 FILLER_67_1678 ();
 FILLCELL_X4 FILLER_67_1694 ();
 FILLCELL_X2 FILLER_67_1698 ();
 FILLCELL_X1 FILLER_67_1700 ();
 FILLCELL_X32 FILLER_68_1 ();
 FILLCELL_X32 FILLER_68_33 ();
 FILLCELL_X32 FILLER_68_65 ();
 FILLCELL_X32 FILLER_68_97 ();
 FILLCELL_X32 FILLER_68_129 ();
 FILLCELL_X32 FILLER_68_161 ();
 FILLCELL_X32 FILLER_68_193 ();
 FILLCELL_X32 FILLER_68_225 ();
 FILLCELL_X32 FILLER_68_257 ();
 FILLCELL_X32 FILLER_68_289 ();
 FILLCELL_X32 FILLER_68_321 ();
 FILLCELL_X8 FILLER_68_353 ();
 FILLCELL_X4 FILLER_68_361 ();
 FILLCELL_X2 FILLER_68_365 ();
 FILLCELL_X8 FILLER_68_371 ();
 FILLCELL_X1 FILLER_68_379 ();
 FILLCELL_X32 FILLER_68_1518 ();
 FILLCELL_X32 FILLER_68_1550 ();
 FILLCELL_X32 FILLER_68_1582 ();
 FILLCELL_X32 FILLER_68_1614 ();
 FILLCELL_X32 FILLER_68_1646 ();
 FILLCELL_X16 FILLER_68_1678 ();
 FILLCELL_X4 FILLER_68_1694 ();
 FILLCELL_X2 FILLER_68_1698 ();
 FILLCELL_X1 FILLER_68_1700 ();
 FILLCELL_X32 FILLER_69_1 ();
 FILLCELL_X32 FILLER_69_33 ();
 FILLCELL_X32 FILLER_69_65 ();
 FILLCELL_X32 FILLER_69_97 ();
 FILLCELL_X32 FILLER_69_129 ();
 FILLCELL_X32 FILLER_69_161 ();
 FILLCELL_X32 FILLER_69_193 ();
 FILLCELL_X32 FILLER_69_225 ();
 FILLCELL_X32 FILLER_69_257 ();
 FILLCELL_X32 FILLER_69_289 ();
 FILLCELL_X32 FILLER_69_321 ();
 FILLCELL_X4 FILLER_69_353 ();
 FILLCELL_X4 FILLER_69_376 ();
 FILLCELL_X16 FILLER_69_1518 ();
 FILLCELL_X2 FILLER_69_1534 ();
 FILLCELL_X1 FILLER_69_1536 ();
 FILLCELL_X32 FILLER_69_1554 ();
 FILLCELL_X32 FILLER_69_1586 ();
 FILLCELL_X32 FILLER_69_1618 ();
 FILLCELL_X32 FILLER_69_1650 ();
 FILLCELL_X16 FILLER_69_1682 ();
 FILLCELL_X2 FILLER_69_1698 ();
 FILLCELL_X1 FILLER_69_1700 ();
 FILLCELL_X4 FILLER_70_1 ();
 FILLCELL_X32 FILLER_70_9 ();
 FILLCELL_X32 FILLER_70_41 ();
 FILLCELL_X32 FILLER_70_73 ();
 FILLCELL_X32 FILLER_70_105 ();
 FILLCELL_X32 FILLER_70_137 ();
 FILLCELL_X32 FILLER_70_169 ();
 FILLCELL_X32 FILLER_70_201 ();
 FILLCELL_X32 FILLER_70_233 ();
 FILLCELL_X32 FILLER_70_265 ();
 FILLCELL_X32 FILLER_70_297 ();
 FILLCELL_X32 FILLER_70_329 ();
 FILLCELL_X8 FILLER_70_361 ();
 FILLCELL_X1 FILLER_70_369 ();
 FILLCELL_X4 FILLER_70_374 ();
 FILLCELL_X2 FILLER_70_378 ();
 FILLCELL_X32 FILLER_70_1518 ();
 FILLCELL_X32 FILLER_70_1550 ();
 FILLCELL_X32 FILLER_70_1582 ();
 FILLCELL_X32 FILLER_70_1614 ();
 FILLCELL_X32 FILLER_70_1646 ();
 FILLCELL_X16 FILLER_70_1678 ();
 FILLCELL_X4 FILLER_70_1694 ();
 FILLCELL_X2 FILLER_70_1698 ();
 FILLCELL_X1 FILLER_70_1700 ();
 FILLCELL_X32 FILLER_71_1 ();
 FILLCELL_X32 FILLER_71_33 ();
 FILLCELL_X32 FILLER_71_65 ();
 FILLCELL_X32 FILLER_71_97 ();
 FILLCELL_X32 FILLER_71_129 ();
 FILLCELL_X32 FILLER_71_161 ();
 FILLCELL_X32 FILLER_71_193 ();
 FILLCELL_X32 FILLER_71_225 ();
 FILLCELL_X32 FILLER_71_257 ();
 FILLCELL_X32 FILLER_71_289 ();
 FILLCELL_X32 FILLER_71_321 ();
 FILLCELL_X16 FILLER_71_353 ();
 FILLCELL_X8 FILLER_71_369 ();
 FILLCELL_X2 FILLER_71_377 ();
 FILLCELL_X1 FILLER_71_379 ();
 FILLCELL_X32 FILLER_71_1518 ();
 FILLCELL_X32 FILLER_71_1550 ();
 FILLCELL_X32 FILLER_71_1582 ();
 FILLCELL_X32 FILLER_71_1614 ();
 FILLCELL_X32 FILLER_71_1646 ();
 FILLCELL_X16 FILLER_71_1678 ();
 FILLCELL_X4 FILLER_71_1694 ();
 FILLCELL_X2 FILLER_71_1698 ();
 FILLCELL_X1 FILLER_71_1700 ();
 FILLCELL_X32 FILLER_72_1 ();
 FILLCELL_X32 FILLER_72_33 ();
 FILLCELL_X32 FILLER_72_65 ();
 FILLCELL_X32 FILLER_72_97 ();
 FILLCELL_X32 FILLER_72_129 ();
 FILLCELL_X32 FILLER_72_161 ();
 FILLCELL_X32 FILLER_72_193 ();
 FILLCELL_X32 FILLER_72_225 ();
 FILLCELL_X32 FILLER_72_257 ();
 FILLCELL_X32 FILLER_72_289 ();
 FILLCELL_X32 FILLER_72_321 ();
 FILLCELL_X4 FILLER_72_353 ();
 FILLCELL_X4 FILLER_72_376 ();
 FILLCELL_X8 FILLER_72_1518 ();
 FILLCELL_X4 FILLER_72_1526 ();
 FILLCELL_X32 FILLER_72_1534 ();
 FILLCELL_X32 FILLER_72_1566 ();
 FILLCELL_X32 FILLER_72_1598 ();
 FILLCELL_X32 FILLER_72_1630 ();
 FILLCELL_X32 FILLER_72_1662 ();
 FILLCELL_X4 FILLER_72_1694 ();
 FILLCELL_X2 FILLER_72_1698 ();
 FILLCELL_X1 FILLER_72_1700 ();
 FILLCELL_X32 FILLER_73_1 ();
 FILLCELL_X32 FILLER_73_33 ();
 FILLCELL_X32 FILLER_73_65 ();
 FILLCELL_X32 FILLER_73_97 ();
 FILLCELL_X32 FILLER_73_129 ();
 FILLCELL_X32 FILLER_73_161 ();
 FILLCELL_X32 FILLER_73_193 ();
 FILLCELL_X32 FILLER_73_225 ();
 FILLCELL_X32 FILLER_73_257 ();
 FILLCELL_X32 FILLER_73_289 ();
 FILLCELL_X32 FILLER_73_321 ();
 FILLCELL_X16 FILLER_73_353 ();
 FILLCELL_X8 FILLER_73_369 ();
 FILLCELL_X2 FILLER_73_377 ();
 FILLCELL_X1 FILLER_73_379 ();
 FILLCELL_X32 FILLER_73_1518 ();
 FILLCELL_X32 FILLER_73_1550 ();
 FILLCELL_X32 FILLER_73_1582 ();
 FILLCELL_X32 FILLER_73_1614 ();
 FILLCELL_X32 FILLER_73_1646 ();
 FILLCELL_X16 FILLER_73_1678 ();
 FILLCELL_X4 FILLER_73_1694 ();
 FILLCELL_X2 FILLER_73_1698 ();
 FILLCELL_X1 FILLER_73_1700 ();
 FILLCELL_X32 FILLER_74_1 ();
 FILLCELL_X32 FILLER_74_33 ();
 FILLCELL_X32 FILLER_74_65 ();
 FILLCELL_X32 FILLER_74_97 ();
 FILLCELL_X32 FILLER_74_129 ();
 FILLCELL_X32 FILLER_74_161 ();
 FILLCELL_X32 FILLER_74_193 ();
 FILLCELL_X32 FILLER_74_225 ();
 FILLCELL_X32 FILLER_74_257 ();
 FILLCELL_X32 FILLER_74_289 ();
 FILLCELL_X32 FILLER_74_321 ();
 FILLCELL_X16 FILLER_74_353 ();
 FILLCELL_X8 FILLER_74_369 ();
 FILLCELL_X2 FILLER_74_377 ();
 FILLCELL_X1 FILLER_74_379 ();
 FILLCELL_X4 FILLER_74_1518 ();
 FILLCELL_X32 FILLER_74_1526 ();
 FILLCELL_X32 FILLER_74_1558 ();
 FILLCELL_X32 FILLER_74_1590 ();
 FILLCELL_X32 FILLER_74_1622 ();
 FILLCELL_X32 FILLER_74_1654 ();
 FILLCELL_X8 FILLER_74_1686 ();
 FILLCELL_X4 FILLER_74_1694 ();
 FILLCELL_X2 FILLER_74_1698 ();
 FILLCELL_X1 FILLER_74_1700 ();
 FILLCELL_X32 FILLER_75_1 ();
 FILLCELL_X32 FILLER_75_33 ();
 FILLCELL_X32 FILLER_75_65 ();
 FILLCELL_X32 FILLER_75_97 ();
 FILLCELL_X32 FILLER_75_129 ();
 FILLCELL_X32 FILLER_75_161 ();
 FILLCELL_X32 FILLER_75_193 ();
 FILLCELL_X32 FILLER_75_225 ();
 FILLCELL_X32 FILLER_75_257 ();
 FILLCELL_X32 FILLER_75_289 ();
 FILLCELL_X32 FILLER_75_321 ();
 FILLCELL_X16 FILLER_75_353 ();
 FILLCELL_X8 FILLER_75_369 ();
 FILLCELL_X2 FILLER_75_377 ();
 FILLCELL_X1 FILLER_75_379 ();
 FILLCELL_X32 FILLER_75_1518 ();
 FILLCELL_X32 FILLER_75_1550 ();
 FILLCELL_X32 FILLER_75_1582 ();
 FILLCELL_X32 FILLER_75_1614 ();
 FILLCELL_X32 FILLER_75_1646 ();
 FILLCELL_X16 FILLER_75_1678 ();
 FILLCELL_X4 FILLER_75_1697 ();
 FILLCELL_X32 FILLER_76_1 ();
 FILLCELL_X32 FILLER_76_33 ();
 FILLCELL_X32 FILLER_76_65 ();
 FILLCELL_X32 FILLER_76_97 ();
 FILLCELL_X32 FILLER_76_129 ();
 FILLCELL_X32 FILLER_76_161 ();
 FILLCELL_X32 FILLER_76_193 ();
 FILLCELL_X32 FILLER_76_225 ();
 FILLCELL_X32 FILLER_76_257 ();
 FILLCELL_X32 FILLER_76_289 ();
 FILLCELL_X32 FILLER_76_321 ();
 FILLCELL_X16 FILLER_76_353 ();
 FILLCELL_X4 FILLER_76_369 ();
 FILLCELL_X4 FILLER_76_376 ();
 FILLCELL_X32 FILLER_76_1518 ();
 FILLCELL_X32 FILLER_76_1550 ();
 FILLCELL_X32 FILLER_76_1582 ();
 FILLCELL_X32 FILLER_76_1614 ();
 FILLCELL_X32 FILLER_76_1646 ();
 FILLCELL_X16 FILLER_76_1678 ();
 FILLCELL_X4 FILLER_76_1694 ();
 FILLCELL_X2 FILLER_76_1698 ();
 FILLCELL_X1 FILLER_76_1700 ();
 FILLCELL_X32 FILLER_77_1 ();
 FILLCELL_X32 FILLER_77_33 ();
 FILLCELL_X32 FILLER_77_65 ();
 FILLCELL_X32 FILLER_77_97 ();
 FILLCELL_X32 FILLER_77_129 ();
 FILLCELL_X32 FILLER_77_161 ();
 FILLCELL_X32 FILLER_77_193 ();
 FILLCELL_X32 FILLER_77_225 ();
 FILLCELL_X32 FILLER_77_257 ();
 FILLCELL_X32 FILLER_77_289 ();
 FILLCELL_X32 FILLER_77_321 ();
 FILLCELL_X16 FILLER_77_353 ();
 FILLCELL_X2 FILLER_77_369 ();
 FILLCELL_X4 FILLER_77_376 ();
 FILLCELL_X32 FILLER_77_1518 ();
 FILLCELL_X32 FILLER_77_1550 ();
 FILLCELL_X32 FILLER_77_1582 ();
 FILLCELL_X32 FILLER_77_1614 ();
 FILLCELL_X32 FILLER_77_1646 ();
 FILLCELL_X16 FILLER_77_1678 ();
 FILLCELL_X4 FILLER_77_1694 ();
 FILLCELL_X2 FILLER_77_1698 ();
 FILLCELL_X1 FILLER_77_1700 ();
 FILLCELL_X32 FILLER_78_1 ();
 FILLCELL_X32 FILLER_78_33 ();
 FILLCELL_X32 FILLER_78_65 ();
 FILLCELL_X32 FILLER_78_97 ();
 FILLCELL_X32 FILLER_78_129 ();
 FILLCELL_X32 FILLER_78_161 ();
 FILLCELL_X32 FILLER_78_193 ();
 FILLCELL_X32 FILLER_78_225 ();
 FILLCELL_X32 FILLER_78_257 ();
 FILLCELL_X32 FILLER_78_289 ();
 FILLCELL_X32 FILLER_78_321 ();
 FILLCELL_X16 FILLER_78_353 ();
 FILLCELL_X8 FILLER_78_369 ();
 FILLCELL_X2 FILLER_78_377 ();
 FILLCELL_X1 FILLER_78_379 ();
 FILLCELL_X32 FILLER_78_1518 ();
 FILLCELL_X32 FILLER_78_1550 ();
 FILLCELL_X32 FILLER_78_1582 ();
 FILLCELL_X32 FILLER_78_1614 ();
 FILLCELL_X32 FILLER_78_1646 ();
 FILLCELL_X16 FILLER_78_1678 ();
 FILLCELL_X4 FILLER_78_1694 ();
 FILLCELL_X2 FILLER_78_1698 ();
 FILLCELL_X1 FILLER_78_1700 ();
 FILLCELL_X32 FILLER_79_1 ();
 FILLCELL_X32 FILLER_79_33 ();
 FILLCELL_X32 FILLER_79_65 ();
 FILLCELL_X32 FILLER_79_97 ();
 FILLCELL_X32 FILLER_79_129 ();
 FILLCELL_X32 FILLER_79_161 ();
 FILLCELL_X32 FILLER_79_193 ();
 FILLCELL_X32 FILLER_79_225 ();
 FILLCELL_X32 FILLER_79_257 ();
 FILLCELL_X32 FILLER_79_289 ();
 FILLCELL_X32 FILLER_79_321 ();
 FILLCELL_X16 FILLER_79_353 ();
 FILLCELL_X2 FILLER_79_369 ();
 FILLCELL_X4 FILLER_79_376 ();
 FILLCELL_X32 FILLER_79_1518 ();
 FILLCELL_X32 FILLER_79_1550 ();
 FILLCELL_X32 FILLER_79_1582 ();
 FILLCELL_X32 FILLER_79_1614 ();
 FILLCELL_X32 FILLER_79_1646 ();
 FILLCELL_X16 FILLER_79_1678 ();
 FILLCELL_X4 FILLER_79_1694 ();
 FILLCELL_X2 FILLER_79_1698 ();
 FILLCELL_X1 FILLER_79_1700 ();
 FILLCELL_X4 FILLER_80_1 ();
 FILLCELL_X32 FILLER_80_8 ();
 FILLCELL_X32 FILLER_80_40 ();
 FILLCELL_X32 FILLER_80_72 ();
 FILLCELL_X32 FILLER_80_104 ();
 FILLCELL_X32 FILLER_80_136 ();
 FILLCELL_X32 FILLER_80_168 ();
 FILLCELL_X32 FILLER_80_200 ();
 FILLCELL_X32 FILLER_80_232 ();
 FILLCELL_X32 FILLER_80_264 ();
 FILLCELL_X32 FILLER_80_296 ();
 FILLCELL_X32 FILLER_80_328 ();
 FILLCELL_X16 FILLER_80_360 ();
 FILLCELL_X4 FILLER_80_376 ();
 FILLCELL_X4 FILLER_80_1518 ();
 FILLCELL_X32 FILLER_80_1526 ();
 FILLCELL_X32 FILLER_80_1558 ();
 FILLCELL_X32 FILLER_80_1590 ();
 FILLCELL_X32 FILLER_80_1622 ();
 FILLCELL_X32 FILLER_80_1654 ();
 FILLCELL_X8 FILLER_80_1686 ();
 FILLCELL_X4 FILLER_80_1694 ();
 FILLCELL_X2 FILLER_80_1698 ();
 FILLCELL_X1 FILLER_80_1700 ();
 FILLCELL_X32 FILLER_81_1 ();
 FILLCELL_X32 FILLER_81_33 ();
 FILLCELL_X32 FILLER_81_65 ();
 FILLCELL_X32 FILLER_81_97 ();
 FILLCELL_X32 FILLER_81_129 ();
 FILLCELL_X32 FILLER_81_161 ();
 FILLCELL_X32 FILLER_81_193 ();
 FILLCELL_X32 FILLER_81_225 ();
 FILLCELL_X32 FILLER_81_257 ();
 FILLCELL_X32 FILLER_81_289 ();
 FILLCELL_X32 FILLER_81_321 ();
 FILLCELL_X16 FILLER_81_353 ();
 FILLCELL_X8 FILLER_81_369 ();
 FILLCELL_X2 FILLER_81_377 ();
 FILLCELL_X1 FILLER_81_379 ();
 FILLCELL_X32 FILLER_81_1518 ();
 FILLCELL_X32 FILLER_81_1550 ();
 FILLCELL_X32 FILLER_81_1582 ();
 FILLCELL_X32 FILLER_81_1614 ();
 FILLCELL_X32 FILLER_81_1646 ();
 FILLCELL_X16 FILLER_81_1678 ();
 FILLCELL_X4 FILLER_81_1694 ();
 FILLCELL_X2 FILLER_81_1698 ();
 FILLCELL_X1 FILLER_81_1700 ();
 FILLCELL_X32 FILLER_82_1 ();
 FILLCELL_X32 FILLER_82_33 ();
 FILLCELL_X32 FILLER_82_65 ();
 FILLCELL_X32 FILLER_82_97 ();
 FILLCELL_X32 FILLER_82_129 ();
 FILLCELL_X32 FILLER_82_161 ();
 FILLCELL_X32 FILLER_82_193 ();
 FILLCELL_X32 FILLER_82_225 ();
 FILLCELL_X32 FILLER_82_257 ();
 FILLCELL_X32 FILLER_82_289 ();
 FILLCELL_X32 FILLER_82_321 ();
 FILLCELL_X16 FILLER_82_353 ();
 FILLCELL_X8 FILLER_82_369 ();
 FILLCELL_X2 FILLER_82_377 ();
 FILLCELL_X1 FILLER_82_379 ();
 FILLCELL_X8 FILLER_82_1518 ();
 FILLCELL_X1 FILLER_82_1526 ();
 FILLCELL_X32 FILLER_82_1544 ();
 FILLCELL_X32 FILLER_82_1576 ();
 FILLCELL_X32 FILLER_82_1608 ();
 FILLCELL_X32 FILLER_82_1640 ();
 FILLCELL_X16 FILLER_82_1672 ();
 FILLCELL_X8 FILLER_82_1688 ();
 FILLCELL_X4 FILLER_82_1696 ();
 FILLCELL_X1 FILLER_82_1700 ();
 FILLCELL_X32 FILLER_83_1 ();
 FILLCELL_X32 FILLER_83_33 ();
 FILLCELL_X32 FILLER_83_65 ();
 FILLCELL_X32 FILLER_83_97 ();
 FILLCELL_X32 FILLER_83_129 ();
 FILLCELL_X32 FILLER_83_161 ();
 FILLCELL_X32 FILLER_83_193 ();
 FILLCELL_X32 FILLER_83_225 ();
 FILLCELL_X32 FILLER_83_257 ();
 FILLCELL_X32 FILLER_83_289 ();
 FILLCELL_X32 FILLER_83_321 ();
 FILLCELL_X16 FILLER_83_353 ();
 FILLCELL_X8 FILLER_83_369 ();
 FILLCELL_X2 FILLER_83_377 ();
 FILLCELL_X1 FILLER_83_379 ();
 FILLCELL_X32 FILLER_83_1518 ();
 FILLCELL_X32 FILLER_83_1550 ();
 FILLCELL_X32 FILLER_83_1582 ();
 FILLCELL_X32 FILLER_83_1614 ();
 FILLCELL_X32 FILLER_83_1646 ();
 FILLCELL_X16 FILLER_83_1678 ();
 FILLCELL_X4 FILLER_83_1694 ();
 FILLCELL_X2 FILLER_83_1698 ();
 FILLCELL_X1 FILLER_83_1700 ();
 FILLCELL_X32 FILLER_84_1 ();
 FILLCELL_X32 FILLER_84_33 ();
 FILLCELL_X32 FILLER_84_65 ();
 FILLCELL_X32 FILLER_84_97 ();
 FILLCELL_X32 FILLER_84_129 ();
 FILLCELL_X32 FILLER_84_161 ();
 FILLCELL_X32 FILLER_84_193 ();
 FILLCELL_X32 FILLER_84_225 ();
 FILLCELL_X32 FILLER_84_257 ();
 FILLCELL_X32 FILLER_84_289 ();
 FILLCELL_X32 FILLER_84_321 ();
 FILLCELL_X16 FILLER_84_353 ();
 FILLCELL_X8 FILLER_84_369 ();
 FILLCELL_X2 FILLER_84_377 ();
 FILLCELL_X1 FILLER_84_379 ();
 FILLCELL_X8 FILLER_84_1518 ();
 FILLCELL_X4 FILLER_84_1526 ();
 FILLCELL_X32 FILLER_84_1534 ();
 FILLCELL_X32 FILLER_84_1566 ();
 FILLCELL_X32 FILLER_84_1598 ();
 FILLCELL_X32 FILLER_84_1630 ();
 FILLCELL_X32 FILLER_84_1662 ();
 FILLCELL_X4 FILLER_84_1694 ();
 FILLCELL_X2 FILLER_84_1698 ();
 FILLCELL_X1 FILLER_84_1700 ();
 FILLCELL_X32 FILLER_85_1 ();
 FILLCELL_X32 FILLER_85_33 ();
 FILLCELL_X32 FILLER_85_65 ();
 FILLCELL_X32 FILLER_85_97 ();
 FILLCELL_X32 FILLER_85_129 ();
 FILLCELL_X32 FILLER_85_161 ();
 FILLCELL_X32 FILLER_85_193 ();
 FILLCELL_X32 FILLER_85_225 ();
 FILLCELL_X32 FILLER_85_257 ();
 FILLCELL_X32 FILLER_85_289 ();
 FILLCELL_X32 FILLER_85_321 ();
 FILLCELL_X16 FILLER_85_353 ();
 FILLCELL_X8 FILLER_85_369 ();
 FILLCELL_X2 FILLER_85_377 ();
 FILLCELL_X1 FILLER_85_379 ();
 FILLCELL_X32 FILLER_85_1518 ();
 FILLCELL_X32 FILLER_85_1550 ();
 FILLCELL_X32 FILLER_85_1582 ();
 FILLCELL_X32 FILLER_85_1614 ();
 FILLCELL_X32 FILLER_85_1646 ();
 FILLCELL_X16 FILLER_85_1678 ();
 FILLCELL_X4 FILLER_85_1697 ();
 FILLCELL_X32 FILLER_86_1 ();
 FILLCELL_X32 FILLER_86_33 ();
 FILLCELL_X32 FILLER_86_65 ();
 FILLCELL_X32 FILLER_86_97 ();
 FILLCELL_X32 FILLER_86_129 ();
 FILLCELL_X32 FILLER_86_161 ();
 FILLCELL_X32 FILLER_86_193 ();
 FILLCELL_X32 FILLER_86_225 ();
 FILLCELL_X32 FILLER_86_257 ();
 FILLCELL_X32 FILLER_86_289 ();
 FILLCELL_X32 FILLER_86_321 ();
 FILLCELL_X16 FILLER_86_353 ();
 FILLCELL_X8 FILLER_86_369 ();
 FILLCELL_X2 FILLER_86_377 ();
 FILLCELL_X1 FILLER_86_379 ();
 FILLCELL_X4 FILLER_86_1518 ();
 FILLCELL_X32 FILLER_86_1526 ();
 FILLCELL_X32 FILLER_86_1558 ();
 FILLCELL_X32 FILLER_86_1590 ();
 FILLCELL_X32 FILLER_86_1622 ();
 FILLCELL_X32 FILLER_86_1654 ();
 FILLCELL_X8 FILLER_86_1686 ();
 FILLCELL_X4 FILLER_86_1694 ();
 FILLCELL_X2 FILLER_86_1698 ();
 FILLCELL_X1 FILLER_86_1700 ();
 FILLCELL_X32 FILLER_87_1 ();
 FILLCELL_X32 FILLER_87_33 ();
 FILLCELL_X32 FILLER_87_65 ();
 FILLCELL_X32 FILLER_87_97 ();
 FILLCELL_X32 FILLER_87_129 ();
 FILLCELL_X32 FILLER_87_161 ();
 FILLCELL_X32 FILLER_87_193 ();
 FILLCELL_X32 FILLER_87_225 ();
 FILLCELL_X32 FILLER_87_257 ();
 FILLCELL_X32 FILLER_87_289 ();
 FILLCELL_X32 FILLER_87_321 ();
 FILLCELL_X16 FILLER_87_353 ();
 FILLCELL_X8 FILLER_87_369 ();
 FILLCELL_X2 FILLER_87_377 ();
 FILLCELL_X1 FILLER_87_379 ();
 FILLCELL_X4 FILLER_87_1518 ();
 FILLCELL_X32 FILLER_87_1541 ();
 FILLCELL_X32 FILLER_87_1573 ();
 FILLCELL_X32 FILLER_87_1605 ();
 FILLCELL_X32 FILLER_87_1637 ();
 FILLCELL_X32 FILLER_87_1669 ();
 FILLCELL_X32 FILLER_88_1 ();
 FILLCELL_X32 FILLER_88_33 ();
 FILLCELL_X32 FILLER_88_65 ();
 FILLCELL_X32 FILLER_88_97 ();
 FILLCELL_X32 FILLER_88_129 ();
 FILLCELL_X32 FILLER_88_161 ();
 FILLCELL_X32 FILLER_88_193 ();
 FILLCELL_X32 FILLER_88_225 ();
 FILLCELL_X32 FILLER_88_257 ();
 FILLCELL_X32 FILLER_88_289 ();
 FILLCELL_X32 FILLER_88_321 ();
 FILLCELL_X16 FILLER_88_353 ();
 FILLCELL_X8 FILLER_88_369 ();
 FILLCELL_X2 FILLER_88_377 ();
 FILLCELL_X1 FILLER_88_379 ();
 FILLCELL_X32 FILLER_88_1518 ();
 FILLCELL_X32 FILLER_88_1550 ();
 FILLCELL_X32 FILLER_88_1582 ();
 FILLCELL_X32 FILLER_88_1614 ();
 FILLCELL_X32 FILLER_88_1646 ();
 FILLCELL_X16 FILLER_88_1678 ();
 FILLCELL_X4 FILLER_88_1694 ();
 FILLCELL_X2 FILLER_88_1698 ();
 FILLCELL_X1 FILLER_88_1700 ();
 FILLCELL_X32 FILLER_89_1 ();
 FILLCELL_X32 FILLER_89_33 ();
 FILLCELL_X32 FILLER_89_65 ();
 FILLCELL_X32 FILLER_89_97 ();
 FILLCELL_X32 FILLER_89_129 ();
 FILLCELL_X32 FILLER_89_161 ();
 FILLCELL_X32 FILLER_89_193 ();
 FILLCELL_X32 FILLER_89_225 ();
 FILLCELL_X32 FILLER_89_257 ();
 FILLCELL_X32 FILLER_89_289 ();
 FILLCELL_X32 FILLER_89_321 ();
 FILLCELL_X16 FILLER_89_353 ();
 FILLCELL_X8 FILLER_89_369 ();
 FILLCELL_X2 FILLER_89_377 ();
 FILLCELL_X1 FILLER_89_379 ();
 FILLCELL_X32 FILLER_89_1518 ();
 FILLCELL_X32 FILLER_89_1550 ();
 FILLCELL_X32 FILLER_89_1582 ();
 FILLCELL_X32 FILLER_89_1614 ();
 FILLCELL_X32 FILLER_89_1646 ();
 FILLCELL_X16 FILLER_89_1678 ();
 FILLCELL_X4 FILLER_89_1694 ();
 FILLCELL_X2 FILLER_89_1698 ();
 FILLCELL_X1 FILLER_89_1700 ();
 FILLCELL_X4 FILLER_90_1 ();
 FILLCELL_X32 FILLER_90_9 ();
 FILLCELL_X32 FILLER_90_41 ();
 FILLCELL_X32 FILLER_90_73 ();
 FILLCELL_X32 FILLER_90_105 ();
 FILLCELL_X32 FILLER_90_137 ();
 FILLCELL_X32 FILLER_90_169 ();
 FILLCELL_X32 FILLER_90_201 ();
 FILLCELL_X32 FILLER_90_233 ();
 FILLCELL_X32 FILLER_90_265 ();
 FILLCELL_X32 FILLER_90_297 ();
 FILLCELL_X32 FILLER_90_329 ();
 FILLCELL_X16 FILLER_90_361 ();
 FILLCELL_X2 FILLER_90_377 ();
 FILLCELL_X1 FILLER_90_379 ();
 FILLCELL_X4 FILLER_90_1518 ();
 FILLCELL_X2 FILLER_90_1522 ();
 FILLCELL_X32 FILLER_90_1541 ();
 FILLCELL_X32 FILLER_90_1573 ();
 FILLCELL_X32 FILLER_90_1605 ();
 FILLCELL_X32 FILLER_90_1637 ();
 FILLCELL_X32 FILLER_90_1669 ();
 FILLCELL_X32 FILLER_91_1 ();
 FILLCELL_X32 FILLER_91_33 ();
 FILLCELL_X32 FILLER_91_65 ();
 FILLCELL_X32 FILLER_91_97 ();
 FILLCELL_X32 FILLER_91_129 ();
 FILLCELL_X32 FILLER_91_161 ();
 FILLCELL_X32 FILLER_91_193 ();
 FILLCELL_X32 FILLER_91_225 ();
 FILLCELL_X32 FILLER_91_257 ();
 FILLCELL_X32 FILLER_91_289 ();
 FILLCELL_X32 FILLER_91_321 ();
 FILLCELL_X16 FILLER_91_353 ();
 FILLCELL_X8 FILLER_91_369 ();
 FILLCELL_X2 FILLER_91_377 ();
 FILLCELL_X1 FILLER_91_379 ();
 FILLCELL_X32 FILLER_91_1518 ();
 FILLCELL_X32 FILLER_91_1550 ();
 FILLCELL_X32 FILLER_91_1582 ();
 FILLCELL_X32 FILLER_91_1614 ();
 FILLCELL_X32 FILLER_91_1646 ();
 FILLCELL_X16 FILLER_91_1678 ();
 FILLCELL_X4 FILLER_91_1694 ();
 FILLCELL_X2 FILLER_91_1698 ();
 FILLCELL_X1 FILLER_91_1700 ();
 FILLCELL_X32 FILLER_92_1 ();
 FILLCELL_X32 FILLER_92_33 ();
 FILLCELL_X32 FILLER_92_65 ();
 FILLCELL_X32 FILLER_92_97 ();
 FILLCELL_X32 FILLER_92_129 ();
 FILLCELL_X32 FILLER_92_161 ();
 FILLCELL_X32 FILLER_92_193 ();
 FILLCELL_X32 FILLER_92_225 ();
 FILLCELL_X32 FILLER_92_257 ();
 FILLCELL_X32 FILLER_92_289 ();
 FILLCELL_X32 FILLER_92_321 ();
 FILLCELL_X16 FILLER_92_353 ();
 FILLCELL_X8 FILLER_92_369 ();
 FILLCELL_X2 FILLER_92_377 ();
 FILLCELL_X1 FILLER_92_379 ();
 FILLCELL_X32 FILLER_92_1518 ();
 FILLCELL_X32 FILLER_92_1550 ();
 FILLCELL_X32 FILLER_92_1582 ();
 FILLCELL_X32 FILLER_92_1614 ();
 FILLCELL_X32 FILLER_92_1646 ();
 FILLCELL_X16 FILLER_92_1678 ();
 FILLCELL_X4 FILLER_92_1694 ();
 FILLCELL_X2 FILLER_92_1698 ();
 FILLCELL_X1 FILLER_92_1700 ();
 FILLCELL_X32 FILLER_93_1 ();
 FILLCELL_X32 FILLER_93_33 ();
 FILLCELL_X32 FILLER_93_65 ();
 FILLCELL_X32 FILLER_93_97 ();
 FILLCELL_X32 FILLER_93_129 ();
 FILLCELL_X32 FILLER_93_161 ();
 FILLCELL_X32 FILLER_93_193 ();
 FILLCELL_X32 FILLER_93_225 ();
 FILLCELL_X32 FILLER_93_257 ();
 FILLCELL_X32 FILLER_93_289 ();
 FILLCELL_X32 FILLER_93_321 ();
 FILLCELL_X8 FILLER_93_353 ();
 FILLCELL_X4 FILLER_93_361 ();
 FILLCELL_X2 FILLER_93_365 ();
 FILLCELL_X8 FILLER_93_371 ();
 FILLCELL_X1 FILLER_93_379 ();
 FILLCELL_X32 FILLER_93_1518 ();
 FILLCELL_X32 FILLER_93_1550 ();
 FILLCELL_X32 FILLER_93_1582 ();
 FILLCELL_X32 FILLER_93_1614 ();
 FILLCELL_X32 FILLER_93_1646 ();
 FILLCELL_X16 FILLER_93_1678 ();
 FILLCELL_X4 FILLER_93_1694 ();
 FILLCELL_X2 FILLER_93_1698 ();
 FILLCELL_X1 FILLER_93_1700 ();
 FILLCELL_X32 FILLER_94_1 ();
 FILLCELL_X32 FILLER_94_33 ();
 FILLCELL_X32 FILLER_94_65 ();
 FILLCELL_X32 FILLER_94_97 ();
 FILLCELL_X32 FILLER_94_129 ();
 FILLCELL_X32 FILLER_94_161 ();
 FILLCELL_X32 FILLER_94_193 ();
 FILLCELL_X32 FILLER_94_225 ();
 FILLCELL_X32 FILLER_94_257 ();
 FILLCELL_X32 FILLER_94_289 ();
 FILLCELL_X32 FILLER_94_321 ();
 FILLCELL_X16 FILLER_94_353 ();
 FILLCELL_X8 FILLER_94_369 ();
 FILLCELL_X2 FILLER_94_377 ();
 FILLCELL_X1 FILLER_94_379 ();
 FILLCELL_X32 FILLER_94_1518 ();
 FILLCELL_X32 FILLER_94_1550 ();
 FILLCELL_X32 FILLER_94_1582 ();
 FILLCELL_X32 FILLER_94_1614 ();
 FILLCELL_X32 FILLER_94_1646 ();
 FILLCELL_X16 FILLER_94_1678 ();
 FILLCELL_X4 FILLER_94_1697 ();
 FILLCELL_X32 FILLER_95_1 ();
 FILLCELL_X32 FILLER_95_33 ();
 FILLCELL_X32 FILLER_95_65 ();
 FILLCELL_X32 FILLER_95_97 ();
 FILLCELL_X32 FILLER_95_129 ();
 FILLCELL_X32 FILLER_95_161 ();
 FILLCELL_X32 FILLER_95_193 ();
 FILLCELL_X32 FILLER_95_225 ();
 FILLCELL_X32 FILLER_95_257 ();
 FILLCELL_X32 FILLER_95_289 ();
 FILLCELL_X32 FILLER_95_321 ();
 FILLCELL_X2 FILLER_95_353 ();
 FILLCELL_X1 FILLER_95_355 ();
 FILLCELL_X4 FILLER_95_375 ();
 FILLCELL_X1 FILLER_95_379 ();
 FILLCELL_X32 FILLER_95_1518 ();
 FILLCELL_X32 FILLER_95_1550 ();
 FILLCELL_X32 FILLER_95_1582 ();
 FILLCELL_X32 FILLER_95_1614 ();
 FILLCELL_X32 FILLER_95_1646 ();
 FILLCELL_X16 FILLER_95_1678 ();
 FILLCELL_X4 FILLER_95_1694 ();
 FILLCELL_X2 FILLER_95_1698 ();
 FILLCELL_X1 FILLER_95_1700 ();
 FILLCELL_X32 FILLER_96_1 ();
 FILLCELL_X32 FILLER_96_33 ();
 FILLCELL_X32 FILLER_96_65 ();
 FILLCELL_X32 FILLER_96_97 ();
 FILLCELL_X32 FILLER_96_129 ();
 FILLCELL_X32 FILLER_96_161 ();
 FILLCELL_X32 FILLER_96_193 ();
 FILLCELL_X32 FILLER_96_225 ();
 FILLCELL_X32 FILLER_96_257 ();
 FILLCELL_X32 FILLER_96_289 ();
 FILLCELL_X8 FILLER_96_321 ();
 FILLCELL_X4 FILLER_96_329 ();
 FILLCELL_X2 FILLER_96_333 ();
 FILLCELL_X32 FILLER_96_337 ();
 FILLCELL_X8 FILLER_96_369 ();
 FILLCELL_X2 FILLER_96_377 ();
 FILLCELL_X1 FILLER_96_379 ();
 FILLCELL_X32 FILLER_96_1518 ();
 FILLCELL_X32 FILLER_96_1550 ();
 FILLCELL_X32 FILLER_96_1582 ();
 FILLCELL_X32 FILLER_96_1614 ();
 FILLCELL_X32 FILLER_96_1646 ();
 FILLCELL_X16 FILLER_96_1678 ();
 FILLCELL_X4 FILLER_96_1694 ();
 FILLCELL_X2 FILLER_96_1698 ();
 FILLCELL_X1 FILLER_96_1700 ();
 FILLCELL_X32 FILLER_97_1 ();
 FILLCELL_X32 FILLER_97_33 ();
 FILLCELL_X32 FILLER_97_65 ();
 FILLCELL_X32 FILLER_97_97 ();
 FILLCELL_X32 FILLER_97_129 ();
 FILLCELL_X32 FILLER_97_161 ();
 FILLCELL_X32 FILLER_97_193 ();
 FILLCELL_X32 FILLER_97_225 ();
 FILLCELL_X32 FILLER_97_257 ();
 FILLCELL_X32 FILLER_97_289 ();
 FILLCELL_X8 FILLER_97_321 ();
 FILLCELL_X2 FILLER_97_329 ();
 FILLCELL_X1 FILLER_97_331 ();
 FILLCELL_X4 FILLER_97_335 ();
 FILLCELL_X4 FILLER_97_342 ();
 FILLCELL_X16 FILLER_97_349 ();
 FILLCELL_X8 FILLER_97_365 ();
 FILLCELL_X4 FILLER_97_373 ();
 FILLCELL_X2 FILLER_97_377 ();
 FILLCELL_X1 FILLER_97_379 ();
 FILLCELL_X32 FILLER_97_1518 ();
 FILLCELL_X32 FILLER_97_1550 ();
 FILLCELL_X32 FILLER_97_1582 ();
 FILLCELL_X32 FILLER_97_1614 ();
 FILLCELL_X32 FILLER_97_1646 ();
 FILLCELL_X16 FILLER_97_1678 ();
 FILLCELL_X4 FILLER_97_1694 ();
 FILLCELL_X2 FILLER_97_1698 ();
 FILLCELL_X1 FILLER_97_1700 ();
 FILLCELL_X4 FILLER_98_1 ();
 FILLCELL_X32 FILLER_98_10 ();
 FILLCELL_X32 FILLER_98_42 ();
 FILLCELL_X32 FILLER_98_74 ();
 FILLCELL_X32 FILLER_98_106 ();
 FILLCELL_X32 FILLER_98_138 ();
 FILLCELL_X32 FILLER_98_170 ();
 FILLCELL_X32 FILLER_98_202 ();
 FILLCELL_X32 FILLER_98_234 ();
 FILLCELL_X32 FILLER_98_266 ();
 FILLCELL_X4 FILLER_98_298 ();
 FILLCELL_X2 FILLER_98_302 ();
 FILLCELL_X1 FILLER_98_304 ();
 FILLCELL_X4 FILLER_98_308 ();
 FILLCELL_X4 FILLER_98_315 ();
 FILLCELL_X4 FILLER_98_336 ();
 FILLCELL_X4 FILLER_98_345 ();
 FILLCELL_X16 FILLER_98_352 ();
 FILLCELL_X8 FILLER_98_368 ();
 FILLCELL_X4 FILLER_98_376 ();
 FILLCELL_X32 FILLER_98_1518 ();
 FILLCELL_X32 FILLER_98_1550 ();
 FILLCELL_X32 FILLER_98_1582 ();
 FILLCELL_X32 FILLER_98_1614 ();
 FILLCELL_X32 FILLER_98_1646 ();
 FILLCELL_X16 FILLER_98_1678 ();
 FILLCELL_X4 FILLER_98_1694 ();
 FILLCELL_X2 FILLER_98_1698 ();
 FILLCELL_X1 FILLER_98_1700 ();
 FILLCELL_X32 FILLER_99_1 ();
 FILLCELL_X32 FILLER_99_33 ();
 FILLCELL_X32 FILLER_99_65 ();
 FILLCELL_X32 FILLER_99_97 ();
 FILLCELL_X32 FILLER_99_129 ();
 FILLCELL_X32 FILLER_99_161 ();
 FILLCELL_X32 FILLER_99_193 ();
 FILLCELL_X32 FILLER_99_225 ();
 FILLCELL_X32 FILLER_99_257 ();
 FILLCELL_X4 FILLER_99_289 ();
 FILLCELL_X2 FILLER_99_293 ();
 FILLCELL_X4 FILLER_99_314 ();
 FILLCELL_X8 FILLER_99_321 ();
 FILLCELL_X4 FILLER_99_333 ();
 FILLCELL_X4 FILLER_99_343 ();
 FILLCELL_X4 FILLER_99_351 ();
 FILLCELL_X16 FILLER_99_358 ();
 FILLCELL_X4 FILLER_99_374 ();
 FILLCELL_X2 FILLER_99_378 ();
 FILLCELL_X32 FILLER_99_1518 ();
 FILLCELL_X32 FILLER_99_1550 ();
 FILLCELL_X32 FILLER_99_1582 ();
 FILLCELL_X32 FILLER_99_1614 ();
 FILLCELL_X32 FILLER_99_1646 ();
 FILLCELL_X16 FILLER_99_1678 ();
 FILLCELL_X4 FILLER_99_1694 ();
 FILLCELL_X2 FILLER_99_1698 ();
 FILLCELL_X1 FILLER_99_1700 ();
 FILLCELL_X32 FILLER_100_1 ();
 FILLCELL_X32 FILLER_100_33 ();
 FILLCELL_X32 FILLER_100_65 ();
 FILLCELL_X32 FILLER_100_97 ();
 FILLCELL_X32 FILLER_100_129 ();
 FILLCELL_X32 FILLER_100_161 ();
 FILLCELL_X32 FILLER_100_193 ();
 FILLCELL_X32 FILLER_100_225 ();
 FILLCELL_X16 FILLER_100_257 ();
 FILLCELL_X8 FILLER_100_273 ();
 FILLCELL_X4 FILLER_100_281 ();
 FILLCELL_X4 FILLER_100_288 ();
 FILLCELL_X4 FILLER_100_295 ();
 FILLCELL_X4 FILLER_100_302 ();
 FILLCELL_X8 FILLER_100_311 ();
 FILLCELL_X1 FILLER_100_319 ();
 FILLCELL_X4 FILLER_100_324 ();
 FILLCELL_X2 FILLER_100_328 ();
 FILLCELL_X1 FILLER_100_330 ();
 FILLCELL_X4 FILLER_100_350 ();
 FILLCELL_X4 FILLER_100_359 ();
 FILLCELL_X8 FILLER_100_372 ();
 FILLCELL_X32 FILLER_100_1518 ();
 FILLCELL_X32 FILLER_100_1550 ();
 FILLCELL_X32 FILLER_100_1582 ();
 FILLCELL_X32 FILLER_100_1614 ();
 FILLCELL_X32 FILLER_100_1646 ();
 FILLCELL_X16 FILLER_100_1678 ();
 FILLCELL_X4 FILLER_100_1694 ();
 FILLCELL_X2 FILLER_100_1698 ();
 FILLCELL_X1 FILLER_100_1700 ();
 FILLCELL_X32 FILLER_101_1 ();
 FILLCELL_X32 FILLER_101_33 ();
 FILLCELL_X32 FILLER_101_65 ();
 FILLCELL_X32 FILLER_101_97 ();
 FILLCELL_X32 FILLER_101_129 ();
 FILLCELL_X32 FILLER_101_161 ();
 FILLCELL_X32 FILLER_101_193 ();
 FILLCELL_X32 FILLER_101_225 ();
 FILLCELL_X16 FILLER_101_257 ();
 FILLCELL_X4 FILLER_101_273 ();
 FILLCELL_X2 FILLER_101_277 ();
 FILLCELL_X4 FILLER_101_298 ();
 FILLCELL_X4 FILLER_101_305 ();
 FILLCELL_X2 FILLER_101_309 ();
 FILLCELL_X1 FILLER_101_311 ();
 FILLCELL_X8 FILLER_101_318 ();
 FILLCELL_X8 FILLER_101_330 ();
 FILLCELL_X4 FILLER_101_342 ();
 FILLCELL_X4 FILLER_101_350 ();
 FILLCELL_X4 FILLER_101_373 ();
 FILLCELL_X2 FILLER_101_377 ();
 FILLCELL_X1 FILLER_101_379 ();
 FILLCELL_X32 FILLER_101_1518 ();
 FILLCELL_X32 FILLER_101_1550 ();
 FILLCELL_X32 FILLER_101_1582 ();
 FILLCELL_X32 FILLER_101_1614 ();
 FILLCELL_X32 FILLER_101_1646 ();
 FILLCELL_X16 FILLER_101_1678 ();
 FILLCELL_X4 FILLER_101_1694 ();
 FILLCELL_X2 FILLER_101_1698 ();
 FILLCELL_X1 FILLER_101_1700 ();
 FILLCELL_X32 FILLER_102_1 ();
 FILLCELL_X32 FILLER_102_33 ();
 FILLCELL_X32 FILLER_102_65 ();
 FILLCELL_X32 FILLER_102_97 ();
 FILLCELL_X32 FILLER_102_129 ();
 FILLCELL_X32 FILLER_102_161 ();
 FILLCELL_X32 FILLER_102_193 ();
 FILLCELL_X32 FILLER_102_225 ();
 FILLCELL_X16 FILLER_102_257 ();
 FILLCELL_X4 FILLER_102_273 ();
 FILLCELL_X4 FILLER_102_280 ();
 FILLCELL_X4 FILLER_102_287 ();
 FILLCELL_X4 FILLER_102_296 ();
 FILLCELL_X1 FILLER_102_300 ();
 FILLCELL_X4 FILLER_102_304 ();
 FILLCELL_X4 FILLER_102_312 ();
 FILLCELL_X2 FILLER_102_316 ();
 FILLCELL_X4 FILLER_102_323 ();
 FILLCELL_X2 FILLER_102_327 ();
 FILLCELL_X4 FILLER_102_332 ();
 FILLCELL_X8 FILLER_102_341 ();
 FILLCELL_X2 FILLER_102_349 ();
 FILLCELL_X8 FILLER_102_354 ();
 FILLCELL_X8 FILLER_102_371 ();
 FILLCELL_X1 FILLER_102_379 ();
 FILLCELL_X32 FILLER_102_1518 ();
 FILLCELL_X32 FILLER_102_1550 ();
 FILLCELL_X32 FILLER_102_1582 ();
 FILLCELL_X32 FILLER_102_1614 ();
 FILLCELL_X32 FILLER_102_1646 ();
 FILLCELL_X16 FILLER_102_1678 ();
 FILLCELL_X4 FILLER_102_1694 ();
 FILLCELL_X2 FILLER_102_1698 ();
 FILLCELL_X1 FILLER_102_1700 ();
 FILLCELL_X32 FILLER_103_1 ();
 FILLCELL_X32 FILLER_103_33 ();
 FILLCELL_X32 FILLER_103_65 ();
 FILLCELL_X32 FILLER_103_97 ();
 FILLCELL_X32 FILLER_103_129 ();
 FILLCELL_X32 FILLER_103_161 ();
 FILLCELL_X32 FILLER_103_193 ();
 FILLCELL_X32 FILLER_103_225 ();
 FILLCELL_X16 FILLER_103_257 ();
 FILLCELL_X8 FILLER_103_273 ();
 FILLCELL_X4 FILLER_103_281 ();
 FILLCELL_X2 FILLER_103_285 ();
 FILLCELL_X4 FILLER_103_290 ();
 FILLCELL_X4 FILLER_103_297 ();
 FILLCELL_X4 FILLER_103_306 ();
 FILLCELL_X4 FILLER_103_316 ();
 FILLCELL_X4 FILLER_103_323 ();
 FILLCELL_X8 FILLER_103_346 ();
 FILLCELL_X2 FILLER_103_354 ();
 FILLCELL_X4 FILLER_103_360 ();
 FILLCELL_X8 FILLER_103_366 ();
 FILLCELL_X4 FILLER_103_374 ();
 FILLCELL_X2 FILLER_103_378 ();
 FILLCELL_X32 FILLER_103_1518 ();
 FILLCELL_X32 FILLER_103_1550 ();
 FILLCELL_X32 FILLER_103_1582 ();
 FILLCELL_X32 FILLER_103_1614 ();
 FILLCELL_X32 FILLER_103_1646 ();
 FILLCELL_X16 FILLER_103_1678 ();
 FILLCELL_X4 FILLER_103_1697 ();
 FILLCELL_X32 FILLER_104_1 ();
 FILLCELL_X32 FILLER_104_33 ();
 FILLCELL_X32 FILLER_104_65 ();
 FILLCELL_X32 FILLER_104_97 ();
 FILLCELL_X32 FILLER_104_129 ();
 FILLCELL_X32 FILLER_104_161 ();
 FILLCELL_X32 FILLER_104_193 ();
 FILLCELL_X32 FILLER_104_225 ();
 FILLCELL_X16 FILLER_104_257 ();
 FILLCELL_X8 FILLER_104_273 ();
 FILLCELL_X4 FILLER_104_281 ();
 FILLCELL_X4 FILLER_104_288 ();
 FILLCELL_X4 FILLER_104_297 ();
 FILLCELL_X2 FILLER_104_301 ();
 FILLCELL_X1 FILLER_104_303 ();
 FILLCELL_X8 FILLER_104_322 ();
 FILLCELL_X1 FILLER_104_330 ();
 FILLCELL_X4 FILLER_104_334 ();
 FILLCELL_X4 FILLER_104_343 ();
 FILLCELL_X4 FILLER_104_352 ();
 FILLCELL_X16 FILLER_104_360 ();
 FILLCELL_X4 FILLER_104_376 ();
 FILLCELL_X32 FILLER_104_1518 ();
 FILLCELL_X32 FILLER_104_1550 ();
 FILLCELL_X32 FILLER_104_1582 ();
 FILLCELL_X32 FILLER_104_1614 ();
 FILLCELL_X32 FILLER_104_1646 ();
 FILLCELL_X16 FILLER_104_1678 ();
 FILLCELL_X4 FILLER_104_1694 ();
 FILLCELL_X2 FILLER_104_1698 ();
 FILLCELL_X1 FILLER_104_1700 ();
 FILLCELL_X32 FILLER_105_1 ();
 FILLCELL_X32 FILLER_105_33 ();
 FILLCELL_X32 FILLER_105_65 ();
 FILLCELL_X32 FILLER_105_97 ();
 FILLCELL_X32 FILLER_105_129 ();
 FILLCELL_X32 FILLER_105_161 ();
 FILLCELL_X32 FILLER_105_193 ();
 FILLCELL_X32 FILLER_105_225 ();
 FILLCELL_X16 FILLER_105_257 ();
 FILLCELL_X4 FILLER_105_273 ();
 FILLCELL_X2 FILLER_105_277 ();
 FILLCELL_X1 FILLER_105_279 ();
 FILLCELL_X4 FILLER_105_299 ();
 FILLCELL_X2 FILLER_105_303 ();
 FILLCELL_X4 FILLER_105_310 ();
 FILLCELL_X2 FILLER_105_314 ();
 FILLCELL_X4 FILLER_105_319 ();
 FILLCELL_X4 FILLER_105_326 ();
 FILLCELL_X2 FILLER_105_330 ();
 FILLCELL_X1 FILLER_105_332 ();
 FILLCELL_X4 FILLER_105_337 ();
 FILLCELL_X4 FILLER_105_344 ();
 FILLCELL_X4 FILLER_105_351 ();
 FILLCELL_X1 FILLER_105_355 ();
 FILLCELL_X4 FILLER_105_361 ();
 FILLCELL_X8 FILLER_105_368 ();
 FILLCELL_X4 FILLER_105_376 ();
 FILLCELL_X32 FILLER_105_1518 ();
 FILLCELL_X32 FILLER_105_1550 ();
 FILLCELL_X32 FILLER_105_1582 ();
 FILLCELL_X32 FILLER_105_1614 ();
 FILLCELL_X32 FILLER_105_1646 ();
 FILLCELL_X16 FILLER_105_1678 ();
 FILLCELL_X4 FILLER_105_1694 ();
 FILLCELL_X2 FILLER_105_1698 ();
 FILLCELL_X1 FILLER_105_1700 ();
 FILLCELL_X32 FILLER_106_1 ();
 FILLCELL_X32 FILLER_106_33 ();
 FILLCELL_X32 FILLER_106_65 ();
 FILLCELL_X32 FILLER_106_97 ();
 FILLCELL_X32 FILLER_106_129 ();
 FILLCELL_X32 FILLER_106_161 ();
 FILLCELL_X32 FILLER_106_193 ();
 FILLCELL_X32 FILLER_106_225 ();
 FILLCELL_X32 FILLER_106_257 ();
 FILLCELL_X4 FILLER_106_292 ();
 FILLCELL_X4 FILLER_106_299 ();
 FILLCELL_X4 FILLER_106_306 ();
 FILLCELL_X4 FILLER_106_313 ();
 FILLCELL_X8 FILLER_106_320 ();
 FILLCELL_X4 FILLER_106_328 ();
 FILLCELL_X1 FILLER_106_332 ();
 FILLCELL_X4 FILLER_106_340 ();
 FILLCELL_X4 FILLER_106_347 ();
 FILLCELL_X1 FILLER_106_351 ();
 FILLCELL_X8 FILLER_106_371 ();
 FILLCELL_X1 FILLER_106_379 ();
 FILLCELL_X32 FILLER_106_1518 ();
 FILLCELL_X32 FILLER_106_1550 ();
 FILLCELL_X32 FILLER_106_1582 ();
 FILLCELL_X32 FILLER_106_1614 ();
 FILLCELL_X32 FILLER_106_1646 ();
 FILLCELL_X16 FILLER_106_1678 ();
 FILLCELL_X4 FILLER_106_1694 ();
 FILLCELL_X2 FILLER_106_1698 ();
 FILLCELL_X1 FILLER_106_1700 ();
 FILLCELL_X32 FILLER_107_1 ();
 FILLCELL_X32 FILLER_107_33 ();
 FILLCELL_X32 FILLER_107_65 ();
 FILLCELL_X32 FILLER_107_97 ();
 FILLCELL_X32 FILLER_107_129 ();
 FILLCELL_X32 FILLER_107_161 ();
 FILLCELL_X32 FILLER_107_193 ();
 FILLCELL_X32 FILLER_107_225 ();
 FILLCELL_X32 FILLER_107_257 ();
 FILLCELL_X4 FILLER_107_289 ();
 FILLCELL_X1 FILLER_107_293 ();
 FILLCELL_X4 FILLER_107_297 ();
 FILLCELL_X4 FILLER_107_306 ();
 FILLCELL_X4 FILLER_107_313 ();
 FILLCELL_X4 FILLER_107_321 ();
 FILLCELL_X4 FILLER_107_329 ();
 FILLCELL_X4 FILLER_107_337 ();
 FILLCELL_X1 FILLER_107_341 ();
 FILLCELL_X4 FILLER_107_344 ();
 FILLCELL_X4 FILLER_107_351 ();
 FILLCELL_X4 FILLER_107_360 ();
 FILLCELL_X1 FILLER_107_364 ();
 FILLCELL_X4 FILLER_107_368 ();
 FILLCELL_X4 FILLER_107_375 ();
 FILLCELL_X1 FILLER_107_379 ();
 FILLCELL_X32 FILLER_107_1518 ();
 FILLCELL_X32 FILLER_107_1550 ();
 FILLCELL_X32 FILLER_107_1582 ();
 FILLCELL_X32 FILLER_107_1614 ();
 FILLCELL_X32 FILLER_107_1646 ();
 FILLCELL_X16 FILLER_107_1678 ();
 FILLCELL_X4 FILLER_107_1694 ();
 FILLCELL_X2 FILLER_107_1698 ();
 FILLCELL_X1 FILLER_107_1700 ();
 FILLCELL_X4 FILLER_108_1 ();
 FILLCELL_X32 FILLER_108_8 ();
 FILLCELL_X32 FILLER_108_40 ();
 FILLCELL_X32 FILLER_108_72 ();
 FILLCELL_X32 FILLER_108_104 ();
 FILLCELL_X32 FILLER_108_136 ();
 FILLCELL_X32 FILLER_108_168 ();
 FILLCELL_X32 FILLER_108_200 ();
 FILLCELL_X32 FILLER_108_232 ();
 FILLCELL_X16 FILLER_108_264 ();
 FILLCELL_X8 FILLER_108_280 ();
 FILLCELL_X4 FILLER_108_288 ();
 FILLCELL_X8 FILLER_108_309 ();
 FILLCELL_X1 FILLER_108_317 ();
 FILLCELL_X4 FILLER_108_323 ();
 FILLCELL_X4 FILLER_108_332 ();
 FILLCELL_X4 FILLER_108_338 ();
 FILLCELL_X2 FILLER_108_342 ();
 FILLCELL_X1 FILLER_108_344 ();
 FILLCELL_X4 FILLER_108_350 ();
 FILLCELL_X2 FILLER_108_354 ();
 FILLCELL_X1 FILLER_108_356 ();
 FILLCELL_X4 FILLER_108_360 ();
 FILLCELL_X4 FILLER_108_367 ();
 FILLCELL_X2 FILLER_108_371 ();
 FILLCELL_X4 FILLER_108_376 ();
 FILLCELL_X32 FILLER_108_1518 ();
 FILLCELL_X32 FILLER_108_1550 ();
 FILLCELL_X32 FILLER_108_1582 ();
 FILLCELL_X32 FILLER_108_1614 ();
 FILLCELL_X32 FILLER_108_1646 ();
 FILLCELL_X16 FILLER_108_1678 ();
 FILLCELL_X4 FILLER_108_1694 ();
 FILLCELL_X2 FILLER_108_1698 ();
 FILLCELL_X1 FILLER_108_1700 ();
 FILLCELL_X32 FILLER_109_1 ();
 FILLCELL_X32 FILLER_109_33 ();
 FILLCELL_X32 FILLER_109_65 ();
 FILLCELL_X32 FILLER_109_97 ();
 FILLCELL_X32 FILLER_109_129 ();
 FILLCELL_X32 FILLER_109_161 ();
 FILLCELL_X32 FILLER_109_193 ();
 FILLCELL_X32 FILLER_109_225 ();
 FILLCELL_X32 FILLER_109_257 ();
 FILLCELL_X8 FILLER_109_289 ();
 FILLCELL_X4 FILLER_109_300 ();
 FILLCELL_X4 FILLER_109_307 ();
 FILLCELL_X8 FILLER_109_315 ();
 FILLCELL_X16 FILLER_109_328 ();
 FILLCELL_X1 FILLER_109_344 ();
 FILLCELL_X4 FILLER_109_348 ();
 FILLCELL_X4 FILLER_109_357 ();
 FILLCELL_X4 FILLER_109_366 ();
 FILLCELL_X1 FILLER_109_370 ();
 FILLCELL_X4 FILLER_109_373 ();
 FILLCELL_X2 FILLER_109_377 ();
 FILLCELL_X1 FILLER_109_379 ();
 FILLCELL_X32 FILLER_109_1518 ();
 FILLCELL_X32 FILLER_109_1550 ();
 FILLCELL_X32 FILLER_109_1582 ();
 FILLCELL_X32 FILLER_109_1614 ();
 FILLCELL_X32 FILLER_109_1646 ();
 FILLCELL_X16 FILLER_109_1678 ();
 FILLCELL_X4 FILLER_109_1694 ();
 FILLCELL_X2 FILLER_109_1698 ();
 FILLCELL_X1 FILLER_109_1700 ();
 FILLCELL_X32 FILLER_110_1 ();
 FILLCELL_X32 FILLER_110_33 ();
 FILLCELL_X32 FILLER_110_65 ();
 FILLCELL_X32 FILLER_110_97 ();
 FILLCELL_X32 FILLER_110_129 ();
 FILLCELL_X32 FILLER_110_161 ();
 FILLCELL_X32 FILLER_110_193 ();
 FILLCELL_X32 FILLER_110_225 ();
 FILLCELL_X32 FILLER_110_257 ();
 FILLCELL_X8 FILLER_110_289 ();
 FILLCELL_X4 FILLER_110_297 ();
 FILLCELL_X4 FILLER_110_304 ();
 FILLCELL_X8 FILLER_110_325 ();
 FILLCELL_X4 FILLER_110_337 ();
 FILLCELL_X4 FILLER_110_345 ();
 FILLCELL_X2 FILLER_110_349 ();
 FILLCELL_X4 FILLER_110_368 ();
 FILLCELL_X4 FILLER_110_376 ();
 FILLCELL_X32 FILLER_110_1518 ();
 FILLCELL_X32 FILLER_110_1550 ();
 FILLCELL_X32 FILLER_110_1582 ();
 FILLCELL_X32 FILLER_110_1614 ();
 FILLCELL_X32 FILLER_110_1646 ();
 FILLCELL_X16 FILLER_110_1678 ();
 FILLCELL_X4 FILLER_110_1694 ();
 FILLCELL_X2 FILLER_110_1698 ();
 FILLCELL_X1 FILLER_110_1700 ();
 FILLCELL_X32 FILLER_111_1 ();
 FILLCELL_X32 FILLER_111_33 ();
 FILLCELL_X32 FILLER_111_65 ();
 FILLCELL_X32 FILLER_111_97 ();
 FILLCELL_X32 FILLER_111_129 ();
 FILLCELL_X32 FILLER_111_161 ();
 FILLCELL_X32 FILLER_111_193 ();
 FILLCELL_X32 FILLER_111_225 ();
 FILLCELL_X32 FILLER_111_257 ();
 FILLCELL_X16 FILLER_111_289 ();
 FILLCELL_X4 FILLER_111_308 ();
 FILLCELL_X1 FILLER_111_312 ();
 FILLCELL_X4 FILLER_111_316 ();
 FILLCELL_X4 FILLER_111_323 ();
 FILLCELL_X4 FILLER_111_330 ();
 FILLCELL_X4 FILLER_111_339 ();
 FILLCELL_X1 FILLER_111_343 ();
 FILLCELL_X8 FILLER_111_348 ();
 FILLCELL_X1 FILLER_111_356 ();
 FILLCELL_X4 FILLER_111_360 ();
 FILLCELL_X4 FILLER_111_367 ();
 FILLCELL_X4 FILLER_111_374 ();
 FILLCELL_X2 FILLER_111_378 ();
 FILLCELL_X32 FILLER_111_1518 ();
 FILLCELL_X32 FILLER_111_1550 ();
 FILLCELL_X32 FILLER_111_1582 ();
 FILLCELL_X32 FILLER_111_1614 ();
 FILLCELL_X32 FILLER_111_1646 ();
 FILLCELL_X16 FILLER_111_1678 ();
 FILLCELL_X4 FILLER_111_1694 ();
 FILLCELL_X2 FILLER_111_1698 ();
 FILLCELL_X1 FILLER_111_1700 ();
 FILLCELL_X32 FILLER_112_1 ();
 FILLCELL_X32 FILLER_112_33 ();
 FILLCELL_X32 FILLER_112_65 ();
 FILLCELL_X32 FILLER_112_97 ();
 FILLCELL_X32 FILLER_112_129 ();
 FILLCELL_X32 FILLER_112_161 ();
 FILLCELL_X32 FILLER_112_193 ();
 FILLCELL_X32 FILLER_112_225 ();
 FILLCELL_X32 FILLER_112_257 ();
 FILLCELL_X32 FILLER_112_289 ();
 FILLCELL_X4 FILLER_112_321 ();
 FILLCELL_X8 FILLER_112_342 ();
 FILLCELL_X4 FILLER_112_354 ();
 FILLCELL_X4 FILLER_112_361 ();
 FILLCELL_X4 FILLER_112_368 ();
 FILLCELL_X1 FILLER_112_372 ();
 FILLCELL_X4 FILLER_112_376 ();
 FILLCELL_X32 FILLER_112_1518 ();
 FILLCELL_X32 FILLER_112_1550 ();
 FILLCELL_X32 FILLER_112_1582 ();
 FILLCELL_X32 FILLER_112_1614 ();
 FILLCELL_X32 FILLER_112_1646 ();
 FILLCELL_X16 FILLER_112_1678 ();
 FILLCELL_X4 FILLER_112_1694 ();
 FILLCELL_X2 FILLER_112_1698 ();
 FILLCELL_X1 FILLER_112_1700 ();
 FILLCELL_X32 FILLER_113_1 ();
 FILLCELL_X32 FILLER_113_33 ();
 FILLCELL_X32 FILLER_113_65 ();
 FILLCELL_X32 FILLER_113_97 ();
 FILLCELL_X32 FILLER_113_129 ();
 FILLCELL_X32 FILLER_113_161 ();
 FILLCELL_X32 FILLER_113_193 ();
 FILLCELL_X32 FILLER_113_225 ();
 FILLCELL_X32 FILLER_113_257 ();
 FILLCELL_X16 FILLER_113_289 ();
 FILLCELL_X8 FILLER_113_305 ();
 FILLCELL_X4 FILLER_113_313 ();
 FILLCELL_X2 FILLER_113_317 ();
 FILLCELL_X4 FILLER_113_322 ();
 FILLCELL_X4 FILLER_113_329 ();
 FILLCELL_X4 FILLER_113_336 ();
 FILLCELL_X8 FILLER_113_344 ();
 FILLCELL_X1 FILLER_113_352 ();
 FILLCELL_X4 FILLER_113_357 ();
 FILLCELL_X8 FILLER_113_370 ();
 FILLCELL_X2 FILLER_113_378 ();
 FILLCELL_X32 FILLER_113_1518 ();
 FILLCELL_X32 FILLER_113_1550 ();
 FILLCELL_X32 FILLER_113_1582 ();
 FILLCELL_X32 FILLER_113_1614 ();
 FILLCELL_X32 FILLER_113_1646 ();
 FILLCELL_X16 FILLER_113_1678 ();
 FILLCELL_X4 FILLER_113_1697 ();
 FILLCELL_X32 FILLER_114_1 ();
 FILLCELL_X32 FILLER_114_33 ();
 FILLCELL_X32 FILLER_114_65 ();
 FILLCELL_X32 FILLER_114_97 ();
 FILLCELL_X32 FILLER_114_129 ();
 FILLCELL_X32 FILLER_114_161 ();
 FILLCELL_X32 FILLER_114_193 ();
 FILLCELL_X32 FILLER_114_225 ();
 FILLCELL_X32 FILLER_114_257 ();
 FILLCELL_X32 FILLER_114_289 ();
 FILLCELL_X8 FILLER_114_321 ();
 FILLCELL_X2 FILLER_114_329 ();
 FILLCELL_X1 FILLER_114_331 ();
 FILLCELL_X4 FILLER_114_338 ();
 FILLCELL_X1 FILLER_114_342 ();
 FILLCELL_X8 FILLER_114_348 ();
 FILLCELL_X1 FILLER_114_356 ();
 FILLCELL_X4 FILLER_114_361 ();
 FILLCELL_X4 FILLER_114_368 ();
 FILLCELL_X4 FILLER_114_375 ();
 FILLCELL_X1 FILLER_114_379 ();
 FILLCELL_X32 FILLER_114_1518 ();
 FILLCELL_X32 FILLER_114_1550 ();
 FILLCELL_X32 FILLER_114_1582 ();
 FILLCELL_X32 FILLER_114_1614 ();
 FILLCELL_X32 FILLER_114_1646 ();
 FILLCELL_X16 FILLER_114_1678 ();
 FILLCELL_X4 FILLER_114_1694 ();
 FILLCELL_X2 FILLER_114_1698 ();
 FILLCELL_X1 FILLER_114_1700 ();
 FILLCELL_X32 FILLER_115_1 ();
 FILLCELL_X32 FILLER_115_33 ();
 FILLCELL_X32 FILLER_115_65 ();
 FILLCELL_X32 FILLER_115_97 ();
 FILLCELL_X32 FILLER_115_129 ();
 FILLCELL_X32 FILLER_115_161 ();
 FILLCELL_X32 FILLER_115_193 ();
 FILLCELL_X32 FILLER_115_225 ();
 FILLCELL_X32 FILLER_115_257 ();
 FILLCELL_X32 FILLER_115_289 ();
 FILLCELL_X2 FILLER_115_321 ();
 FILLCELL_X8 FILLER_115_340 ();
 FILLCELL_X2 FILLER_115_348 ();
 FILLCELL_X4 FILLER_115_356 ();
 FILLCELL_X4 FILLER_115_365 ();
 FILLCELL_X4 FILLER_115_373 ();
 FILLCELL_X2 FILLER_115_377 ();
 FILLCELL_X1 FILLER_115_379 ();
 FILLCELL_X32 FILLER_115_1518 ();
 FILLCELL_X32 FILLER_115_1550 ();
 FILLCELL_X32 FILLER_115_1582 ();
 FILLCELL_X32 FILLER_115_1614 ();
 FILLCELL_X32 FILLER_115_1646 ();
 FILLCELL_X16 FILLER_115_1678 ();
 FILLCELL_X4 FILLER_115_1694 ();
 FILLCELL_X2 FILLER_115_1698 ();
 FILLCELL_X1 FILLER_115_1700 ();
 FILLCELL_X32 FILLER_116_1 ();
 FILLCELL_X32 FILLER_116_33 ();
 FILLCELL_X32 FILLER_116_65 ();
 FILLCELL_X32 FILLER_116_97 ();
 FILLCELL_X32 FILLER_116_129 ();
 FILLCELL_X32 FILLER_116_161 ();
 FILLCELL_X32 FILLER_116_193 ();
 FILLCELL_X32 FILLER_116_225 ();
 FILLCELL_X32 FILLER_116_257 ();
 FILLCELL_X32 FILLER_116_289 ();
 FILLCELL_X1 FILLER_116_321 ();
 FILLCELL_X4 FILLER_116_324 ();
 FILLCELL_X4 FILLER_116_331 ();
 FILLCELL_X4 FILLER_116_338 ();
 FILLCELL_X4 FILLER_116_359 ();
 FILLCELL_X4 FILLER_116_366 ();
 FILLCELL_X2 FILLER_116_370 ();
 FILLCELL_X1 FILLER_116_372 ();
 FILLCELL_X4 FILLER_116_376 ();
 FILLCELL_X32 FILLER_116_1518 ();
 FILLCELL_X32 FILLER_116_1550 ();
 FILLCELL_X32 FILLER_116_1582 ();
 FILLCELL_X32 FILLER_116_1614 ();
 FILLCELL_X32 FILLER_116_1646 ();
 FILLCELL_X16 FILLER_116_1678 ();
 FILLCELL_X4 FILLER_116_1694 ();
 FILLCELL_X2 FILLER_116_1698 ();
 FILLCELL_X1 FILLER_116_1700 ();
 FILLCELL_X4 FILLER_117_1 ();
 FILLCELL_X32 FILLER_117_10 ();
 FILLCELL_X32 FILLER_117_42 ();
 FILLCELL_X32 FILLER_117_74 ();
 FILLCELL_X32 FILLER_117_106 ();
 FILLCELL_X32 FILLER_117_138 ();
 FILLCELL_X32 FILLER_117_170 ();
 FILLCELL_X32 FILLER_117_202 ();
 FILLCELL_X32 FILLER_117_234 ();
 FILLCELL_X32 FILLER_117_266 ();
 FILLCELL_X32 FILLER_117_298 ();
 FILLCELL_X4 FILLER_117_330 ();
 FILLCELL_X1 FILLER_117_334 ();
 FILLCELL_X4 FILLER_117_338 ();
 FILLCELL_X1 FILLER_117_342 ();
 FILLCELL_X4 FILLER_117_346 ();
 FILLCELL_X4 FILLER_117_367 ();
 FILLCELL_X4 FILLER_117_374 ();
 FILLCELL_X2 FILLER_117_378 ();
 FILLCELL_X32 FILLER_117_1518 ();
 FILLCELL_X32 FILLER_117_1550 ();
 FILLCELL_X32 FILLER_117_1582 ();
 FILLCELL_X32 FILLER_117_1614 ();
 FILLCELL_X32 FILLER_117_1646 ();
 FILLCELL_X16 FILLER_117_1678 ();
 FILLCELL_X4 FILLER_117_1694 ();
 FILLCELL_X2 FILLER_117_1698 ();
 FILLCELL_X1 FILLER_117_1700 ();
 FILLCELL_X32 FILLER_118_1 ();
 FILLCELL_X32 FILLER_118_33 ();
 FILLCELL_X32 FILLER_118_65 ();
 FILLCELL_X32 FILLER_118_97 ();
 FILLCELL_X32 FILLER_118_129 ();
 FILLCELL_X32 FILLER_118_161 ();
 FILLCELL_X32 FILLER_118_193 ();
 FILLCELL_X32 FILLER_118_225 ();
 FILLCELL_X32 FILLER_118_257 ();
 FILLCELL_X32 FILLER_118_289 ();
 FILLCELL_X16 FILLER_118_321 ();
 FILLCELL_X8 FILLER_118_337 ();
 FILLCELL_X4 FILLER_118_345 ();
 FILLCELL_X2 FILLER_118_349 ();
 FILLCELL_X1 FILLER_118_351 ();
 FILLCELL_X8 FILLER_118_355 ();
 FILLCELL_X1 FILLER_118_363 ();
 FILLCELL_X4 FILLER_118_367 ();
 FILLCELL_X4 FILLER_118_374 ();
 FILLCELL_X2 FILLER_118_378 ();
 FILLCELL_X32 FILLER_118_1518 ();
 FILLCELL_X32 FILLER_118_1550 ();
 FILLCELL_X32 FILLER_118_1582 ();
 FILLCELL_X32 FILLER_118_1614 ();
 FILLCELL_X32 FILLER_118_1646 ();
 FILLCELL_X16 FILLER_118_1678 ();
 FILLCELL_X4 FILLER_118_1694 ();
 FILLCELL_X2 FILLER_118_1698 ();
 FILLCELL_X1 FILLER_118_1700 ();
 FILLCELL_X32 FILLER_119_1 ();
 FILLCELL_X32 FILLER_119_33 ();
 FILLCELL_X32 FILLER_119_65 ();
 FILLCELL_X32 FILLER_119_97 ();
 FILLCELL_X32 FILLER_119_129 ();
 FILLCELL_X32 FILLER_119_161 ();
 FILLCELL_X32 FILLER_119_193 ();
 FILLCELL_X32 FILLER_119_225 ();
 FILLCELL_X32 FILLER_119_257 ();
 FILLCELL_X32 FILLER_119_289 ();
 FILLCELL_X32 FILLER_119_321 ();
 FILLCELL_X16 FILLER_119_353 ();
 FILLCELL_X8 FILLER_119_369 ();
 FILLCELL_X2 FILLER_119_377 ();
 FILLCELL_X1 FILLER_119_379 ();
 FILLCELL_X32 FILLER_119_1518 ();
 FILLCELL_X32 FILLER_119_1550 ();
 FILLCELL_X32 FILLER_119_1582 ();
 FILLCELL_X32 FILLER_119_1614 ();
 FILLCELL_X32 FILLER_119_1646 ();
 FILLCELL_X16 FILLER_119_1678 ();
 FILLCELL_X4 FILLER_119_1694 ();
 FILLCELL_X2 FILLER_119_1698 ();
 FILLCELL_X1 FILLER_119_1700 ();
 FILLCELL_X32 FILLER_120_1 ();
 FILLCELL_X32 FILLER_120_33 ();
 FILLCELL_X32 FILLER_120_65 ();
 FILLCELL_X32 FILLER_120_97 ();
 FILLCELL_X32 FILLER_120_129 ();
 FILLCELL_X32 FILLER_120_161 ();
 FILLCELL_X32 FILLER_120_193 ();
 FILLCELL_X32 FILLER_120_225 ();
 FILLCELL_X32 FILLER_120_257 ();
 FILLCELL_X32 FILLER_120_289 ();
 FILLCELL_X32 FILLER_120_321 ();
 FILLCELL_X4 FILLER_120_353 ();
 FILLCELL_X2 FILLER_120_357 ();
 FILLCELL_X4 FILLER_120_362 ();
 FILLCELL_X4 FILLER_120_369 ();
 FILLCELL_X4 FILLER_120_376 ();
 FILLCELL_X32 FILLER_120_1518 ();
 FILLCELL_X32 FILLER_120_1550 ();
 FILLCELL_X32 FILLER_120_1582 ();
 FILLCELL_X32 FILLER_120_1614 ();
 FILLCELL_X32 FILLER_120_1646 ();
 FILLCELL_X16 FILLER_120_1678 ();
 FILLCELL_X4 FILLER_120_1694 ();
 FILLCELL_X2 FILLER_120_1698 ();
 FILLCELL_X1 FILLER_120_1700 ();
 FILLCELL_X32 FILLER_121_1 ();
 FILLCELL_X32 FILLER_121_33 ();
 FILLCELL_X32 FILLER_121_65 ();
 FILLCELL_X32 FILLER_121_97 ();
 FILLCELL_X32 FILLER_121_129 ();
 FILLCELL_X32 FILLER_121_161 ();
 FILLCELL_X32 FILLER_121_193 ();
 FILLCELL_X32 FILLER_121_225 ();
 FILLCELL_X32 FILLER_121_257 ();
 FILLCELL_X32 FILLER_121_289 ();
 FILLCELL_X32 FILLER_121_321 ();
 FILLCELL_X16 FILLER_121_353 ();
 FILLCELL_X4 FILLER_121_369 ();
 FILLCELL_X4 FILLER_121_376 ();
 FILLCELL_X32 FILLER_121_1518 ();
 FILLCELL_X32 FILLER_121_1550 ();
 FILLCELL_X32 FILLER_121_1582 ();
 FILLCELL_X32 FILLER_121_1614 ();
 FILLCELL_X32 FILLER_121_1646 ();
 FILLCELL_X16 FILLER_121_1678 ();
 FILLCELL_X4 FILLER_121_1694 ();
 FILLCELL_X2 FILLER_121_1698 ();
 FILLCELL_X1 FILLER_121_1700 ();
 FILLCELL_X32 FILLER_122_1 ();
 FILLCELL_X32 FILLER_122_33 ();
 FILLCELL_X32 FILLER_122_65 ();
 FILLCELL_X32 FILLER_122_97 ();
 FILLCELL_X32 FILLER_122_129 ();
 FILLCELL_X32 FILLER_122_161 ();
 FILLCELL_X32 FILLER_122_193 ();
 FILLCELL_X32 FILLER_122_225 ();
 FILLCELL_X32 FILLER_122_257 ();
 FILLCELL_X32 FILLER_122_289 ();
 FILLCELL_X32 FILLER_122_321 ();
 FILLCELL_X16 FILLER_122_353 ();
 FILLCELL_X8 FILLER_122_369 ();
 FILLCELL_X2 FILLER_122_377 ();
 FILLCELL_X1 FILLER_122_379 ();
 FILLCELL_X32 FILLER_122_1518 ();
 FILLCELL_X32 FILLER_122_1550 ();
 FILLCELL_X32 FILLER_122_1582 ();
 FILLCELL_X32 FILLER_122_1614 ();
 FILLCELL_X32 FILLER_122_1646 ();
 FILLCELL_X8 FILLER_122_1678 ();
 FILLCELL_X4 FILLER_122_1686 ();
 FILLCELL_X2 FILLER_122_1690 ();
 FILLCELL_X1 FILLER_122_1692 ();
 FILLCELL_X4 FILLER_122_1697 ();
 FILLCELL_X32 FILLER_123_1 ();
 FILLCELL_X32 FILLER_123_33 ();
 FILLCELL_X32 FILLER_123_65 ();
 FILLCELL_X32 FILLER_123_97 ();
 FILLCELL_X32 FILLER_123_129 ();
 FILLCELL_X32 FILLER_123_161 ();
 FILLCELL_X32 FILLER_123_193 ();
 FILLCELL_X32 FILLER_123_225 ();
 FILLCELL_X32 FILLER_123_257 ();
 FILLCELL_X32 FILLER_123_289 ();
 FILLCELL_X32 FILLER_123_321 ();
 FILLCELL_X8 FILLER_123_353 ();
 FILLCELL_X4 FILLER_123_361 ();
 FILLCELL_X1 FILLER_123_365 ();
 FILLCELL_X4 FILLER_123_369 ();
 FILLCELL_X4 FILLER_123_376 ();
 FILLCELL_X32 FILLER_123_1518 ();
 FILLCELL_X32 FILLER_123_1550 ();
 FILLCELL_X32 FILLER_123_1582 ();
 FILLCELL_X32 FILLER_123_1614 ();
 FILLCELL_X32 FILLER_123_1646 ();
 FILLCELL_X16 FILLER_123_1678 ();
 FILLCELL_X4 FILLER_123_1694 ();
 FILLCELL_X2 FILLER_123_1698 ();
 FILLCELL_X1 FILLER_123_1700 ();
 FILLCELL_X32 FILLER_124_1 ();
 FILLCELL_X32 FILLER_124_33 ();
 FILLCELL_X32 FILLER_124_65 ();
 FILLCELL_X32 FILLER_124_97 ();
 FILLCELL_X32 FILLER_124_129 ();
 FILLCELL_X32 FILLER_124_161 ();
 FILLCELL_X32 FILLER_124_193 ();
 FILLCELL_X32 FILLER_124_225 ();
 FILLCELL_X32 FILLER_124_257 ();
 FILLCELL_X32 FILLER_124_289 ();
 FILLCELL_X32 FILLER_124_321 ();
 FILLCELL_X16 FILLER_124_353 ();
 FILLCELL_X8 FILLER_124_369 ();
 FILLCELL_X2 FILLER_124_377 ();
 FILLCELL_X1 FILLER_124_379 ();
 FILLCELL_X32 FILLER_124_1518 ();
 FILLCELL_X32 FILLER_124_1550 ();
 FILLCELL_X32 FILLER_124_1582 ();
 FILLCELL_X32 FILLER_124_1614 ();
 FILLCELL_X32 FILLER_124_1646 ();
 FILLCELL_X16 FILLER_124_1678 ();
 FILLCELL_X4 FILLER_124_1694 ();
 FILLCELL_X2 FILLER_124_1698 ();
 FILLCELL_X1 FILLER_124_1700 ();
 FILLCELL_X32 FILLER_125_1 ();
 FILLCELL_X32 FILLER_125_33 ();
 FILLCELL_X32 FILLER_125_65 ();
 FILLCELL_X32 FILLER_125_97 ();
 FILLCELL_X32 FILLER_125_129 ();
 FILLCELL_X32 FILLER_125_161 ();
 FILLCELL_X32 FILLER_125_193 ();
 FILLCELL_X32 FILLER_125_225 ();
 FILLCELL_X32 FILLER_125_257 ();
 FILLCELL_X32 FILLER_125_289 ();
 FILLCELL_X32 FILLER_125_321 ();
 FILLCELL_X16 FILLER_125_353 ();
 FILLCELL_X8 FILLER_125_369 ();
 FILLCELL_X2 FILLER_125_377 ();
 FILLCELL_X1 FILLER_125_379 ();
 FILLCELL_X32 FILLER_125_1518 ();
 FILLCELL_X32 FILLER_125_1550 ();
 FILLCELL_X32 FILLER_125_1582 ();
 FILLCELL_X32 FILLER_125_1614 ();
 FILLCELL_X32 FILLER_125_1646 ();
 FILLCELL_X16 FILLER_125_1678 ();
 FILLCELL_X4 FILLER_125_1694 ();
 FILLCELL_X2 FILLER_125_1698 ();
 FILLCELL_X1 FILLER_125_1700 ();
 FILLCELL_X4 FILLER_126_1 ();
 FILLCELL_X32 FILLER_126_8 ();
 FILLCELL_X32 FILLER_126_40 ();
 FILLCELL_X32 FILLER_126_72 ();
 FILLCELL_X32 FILLER_126_104 ();
 FILLCELL_X32 FILLER_126_136 ();
 FILLCELL_X32 FILLER_126_168 ();
 FILLCELL_X32 FILLER_126_200 ();
 FILLCELL_X32 FILLER_126_232 ();
 FILLCELL_X32 FILLER_126_264 ();
 FILLCELL_X32 FILLER_126_296 ();
 FILLCELL_X32 FILLER_126_328 ();
 FILLCELL_X8 FILLER_126_360 ();
 FILLCELL_X4 FILLER_126_368 ();
 FILLCELL_X1 FILLER_126_372 ();
 FILLCELL_X4 FILLER_126_376 ();
 FILLCELL_X32 FILLER_126_1518 ();
 FILLCELL_X32 FILLER_126_1550 ();
 FILLCELL_X32 FILLER_126_1582 ();
 FILLCELL_X32 FILLER_126_1614 ();
 FILLCELL_X32 FILLER_126_1646 ();
 FILLCELL_X16 FILLER_126_1678 ();
 FILLCELL_X4 FILLER_126_1694 ();
 FILLCELL_X2 FILLER_126_1698 ();
 FILLCELL_X1 FILLER_126_1700 ();
 FILLCELL_X32 FILLER_127_1 ();
 FILLCELL_X32 FILLER_127_33 ();
 FILLCELL_X32 FILLER_127_65 ();
 FILLCELL_X32 FILLER_127_97 ();
 FILLCELL_X32 FILLER_127_129 ();
 FILLCELL_X32 FILLER_127_161 ();
 FILLCELL_X32 FILLER_127_193 ();
 FILLCELL_X32 FILLER_127_225 ();
 FILLCELL_X32 FILLER_127_257 ();
 FILLCELL_X32 FILLER_127_289 ();
 FILLCELL_X32 FILLER_127_321 ();
 FILLCELL_X16 FILLER_127_353 ();
 FILLCELL_X8 FILLER_127_369 ();
 FILLCELL_X2 FILLER_127_377 ();
 FILLCELL_X1 FILLER_127_379 ();
 FILLCELL_X32 FILLER_127_1518 ();
 FILLCELL_X32 FILLER_127_1550 ();
 FILLCELL_X32 FILLER_127_1582 ();
 FILLCELL_X32 FILLER_127_1614 ();
 FILLCELL_X32 FILLER_127_1646 ();
 FILLCELL_X16 FILLER_127_1678 ();
 FILLCELL_X4 FILLER_127_1694 ();
 FILLCELL_X2 FILLER_127_1698 ();
 FILLCELL_X1 FILLER_127_1700 ();
 FILLCELL_X32 FILLER_128_1 ();
 FILLCELL_X32 FILLER_128_33 ();
 FILLCELL_X32 FILLER_128_65 ();
 FILLCELL_X32 FILLER_128_97 ();
 FILLCELL_X32 FILLER_128_129 ();
 FILLCELL_X32 FILLER_128_161 ();
 FILLCELL_X32 FILLER_128_193 ();
 FILLCELL_X32 FILLER_128_225 ();
 FILLCELL_X32 FILLER_128_257 ();
 FILLCELL_X32 FILLER_128_289 ();
 FILLCELL_X32 FILLER_128_321 ();
 FILLCELL_X16 FILLER_128_353 ();
 FILLCELL_X8 FILLER_128_369 ();
 FILLCELL_X2 FILLER_128_377 ();
 FILLCELL_X1 FILLER_128_379 ();
 FILLCELL_X32 FILLER_128_1518 ();
 FILLCELL_X32 FILLER_128_1550 ();
 FILLCELL_X32 FILLER_128_1582 ();
 FILLCELL_X32 FILLER_128_1614 ();
 FILLCELL_X32 FILLER_128_1646 ();
 FILLCELL_X16 FILLER_128_1678 ();
 FILLCELL_X4 FILLER_128_1694 ();
 FILLCELL_X2 FILLER_128_1698 ();
 FILLCELL_X1 FILLER_128_1700 ();
 FILLCELL_X32 FILLER_129_1 ();
 FILLCELL_X32 FILLER_129_33 ();
 FILLCELL_X32 FILLER_129_65 ();
 FILLCELL_X32 FILLER_129_97 ();
 FILLCELL_X32 FILLER_129_129 ();
 FILLCELL_X32 FILLER_129_161 ();
 FILLCELL_X32 FILLER_129_193 ();
 FILLCELL_X32 FILLER_129_225 ();
 FILLCELL_X32 FILLER_129_257 ();
 FILLCELL_X32 FILLER_129_289 ();
 FILLCELL_X32 FILLER_129_321 ();
 FILLCELL_X16 FILLER_129_353 ();
 FILLCELL_X8 FILLER_129_369 ();
 FILLCELL_X2 FILLER_129_377 ();
 FILLCELL_X1 FILLER_129_379 ();
 FILLCELL_X32 FILLER_129_1518 ();
 FILLCELL_X32 FILLER_129_1550 ();
 FILLCELL_X32 FILLER_129_1582 ();
 FILLCELL_X32 FILLER_129_1614 ();
 FILLCELL_X32 FILLER_129_1646 ();
 FILLCELL_X16 FILLER_129_1678 ();
 FILLCELL_X4 FILLER_129_1694 ();
 FILLCELL_X2 FILLER_129_1698 ();
 FILLCELL_X1 FILLER_129_1700 ();
 FILLCELL_X32 FILLER_130_1 ();
 FILLCELL_X32 FILLER_130_33 ();
 FILLCELL_X32 FILLER_130_65 ();
 FILLCELL_X32 FILLER_130_97 ();
 FILLCELL_X32 FILLER_130_129 ();
 FILLCELL_X32 FILLER_130_161 ();
 FILLCELL_X32 FILLER_130_193 ();
 FILLCELL_X32 FILLER_130_225 ();
 FILLCELL_X32 FILLER_130_257 ();
 FILLCELL_X32 FILLER_130_289 ();
 FILLCELL_X32 FILLER_130_321 ();
 FILLCELL_X16 FILLER_130_353 ();
 FILLCELL_X8 FILLER_130_369 ();
 FILLCELL_X2 FILLER_130_377 ();
 FILLCELL_X1 FILLER_130_379 ();
 FILLCELL_X32 FILLER_130_1518 ();
 FILLCELL_X32 FILLER_130_1550 ();
 FILLCELL_X32 FILLER_130_1582 ();
 FILLCELL_X32 FILLER_130_1614 ();
 FILLCELL_X32 FILLER_130_1646 ();
 FILLCELL_X16 FILLER_130_1678 ();
 FILLCELL_X4 FILLER_130_1694 ();
 FILLCELL_X2 FILLER_130_1698 ();
 FILLCELL_X1 FILLER_130_1700 ();
 FILLCELL_X32 FILLER_131_1 ();
 FILLCELL_X32 FILLER_131_33 ();
 FILLCELL_X32 FILLER_131_65 ();
 FILLCELL_X32 FILLER_131_97 ();
 FILLCELL_X32 FILLER_131_129 ();
 FILLCELL_X32 FILLER_131_161 ();
 FILLCELL_X32 FILLER_131_193 ();
 FILLCELL_X32 FILLER_131_225 ();
 FILLCELL_X32 FILLER_131_257 ();
 FILLCELL_X32 FILLER_131_289 ();
 FILLCELL_X32 FILLER_131_321 ();
 FILLCELL_X16 FILLER_131_353 ();
 FILLCELL_X8 FILLER_131_369 ();
 FILLCELL_X2 FILLER_131_377 ();
 FILLCELL_X1 FILLER_131_379 ();
 FILLCELL_X32 FILLER_131_1518 ();
 FILLCELL_X32 FILLER_131_1550 ();
 FILLCELL_X32 FILLER_131_1582 ();
 FILLCELL_X32 FILLER_131_1614 ();
 FILLCELL_X32 FILLER_131_1646 ();
 FILLCELL_X16 FILLER_131_1678 ();
 FILLCELL_X4 FILLER_131_1697 ();
 FILLCELL_X32 FILLER_132_1 ();
 FILLCELL_X32 FILLER_132_33 ();
 FILLCELL_X32 FILLER_132_65 ();
 FILLCELL_X32 FILLER_132_97 ();
 FILLCELL_X32 FILLER_132_129 ();
 FILLCELL_X32 FILLER_132_161 ();
 FILLCELL_X32 FILLER_132_193 ();
 FILLCELL_X32 FILLER_132_225 ();
 FILLCELL_X32 FILLER_132_257 ();
 FILLCELL_X32 FILLER_132_289 ();
 FILLCELL_X32 FILLER_132_321 ();
 FILLCELL_X16 FILLER_132_353 ();
 FILLCELL_X8 FILLER_132_369 ();
 FILLCELL_X2 FILLER_132_377 ();
 FILLCELL_X1 FILLER_132_379 ();
 FILLCELL_X32 FILLER_132_1518 ();
 FILLCELL_X32 FILLER_132_1550 ();
 FILLCELL_X32 FILLER_132_1582 ();
 FILLCELL_X32 FILLER_132_1614 ();
 FILLCELL_X32 FILLER_132_1646 ();
 FILLCELL_X16 FILLER_132_1678 ();
 FILLCELL_X4 FILLER_132_1694 ();
 FILLCELL_X2 FILLER_132_1698 ();
 FILLCELL_X1 FILLER_132_1700 ();
 FILLCELL_X32 FILLER_133_1 ();
 FILLCELL_X32 FILLER_133_33 ();
 FILLCELL_X32 FILLER_133_65 ();
 FILLCELL_X32 FILLER_133_97 ();
 FILLCELL_X32 FILLER_133_129 ();
 FILLCELL_X32 FILLER_133_161 ();
 FILLCELL_X32 FILLER_133_193 ();
 FILLCELL_X32 FILLER_133_225 ();
 FILLCELL_X32 FILLER_133_257 ();
 FILLCELL_X32 FILLER_133_289 ();
 FILLCELL_X32 FILLER_133_321 ();
 FILLCELL_X16 FILLER_133_353 ();
 FILLCELL_X8 FILLER_133_369 ();
 FILLCELL_X2 FILLER_133_377 ();
 FILLCELL_X1 FILLER_133_379 ();
 FILLCELL_X32 FILLER_133_1518 ();
 FILLCELL_X32 FILLER_133_1550 ();
 FILLCELL_X32 FILLER_133_1582 ();
 FILLCELL_X32 FILLER_133_1614 ();
 FILLCELL_X32 FILLER_133_1646 ();
 FILLCELL_X16 FILLER_133_1678 ();
 FILLCELL_X4 FILLER_133_1694 ();
 FILLCELL_X2 FILLER_133_1698 ();
 FILLCELL_X1 FILLER_133_1700 ();
 FILLCELL_X32 FILLER_134_1 ();
 FILLCELL_X32 FILLER_134_33 ();
 FILLCELL_X32 FILLER_134_65 ();
 FILLCELL_X32 FILLER_134_97 ();
 FILLCELL_X32 FILLER_134_129 ();
 FILLCELL_X32 FILLER_134_161 ();
 FILLCELL_X32 FILLER_134_193 ();
 FILLCELL_X32 FILLER_134_225 ();
 FILLCELL_X32 FILLER_134_257 ();
 FILLCELL_X32 FILLER_134_289 ();
 FILLCELL_X32 FILLER_134_321 ();
 FILLCELL_X16 FILLER_134_353 ();
 FILLCELL_X8 FILLER_134_369 ();
 FILLCELL_X2 FILLER_134_377 ();
 FILLCELL_X1 FILLER_134_379 ();
 FILLCELL_X32 FILLER_134_1518 ();
 FILLCELL_X32 FILLER_134_1550 ();
 FILLCELL_X32 FILLER_134_1582 ();
 FILLCELL_X32 FILLER_134_1614 ();
 FILLCELL_X32 FILLER_134_1646 ();
 FILLCELL_X16 FILLER_134_1678 ();
 FILLCELL_X4 FILLER_134_1694 ();
 FILLCELL_X2 FILLER_134_1698 ();
 FILLCELL_X1 FILLER_134_1700 ();
 FILLCELL_X32 FILLER_135_1 ();
 FILLCELL_X32 FILLER_135_33 ();
 FILLCELL_X32 FILLER_135_65 ();
 FILLCELL_X32 FILLER_135_97 ();
 FILLCELL_X32 FILLER_135_129 ();
 FILLCELL_X32 FILLER_135_161 ();
 FILLCELL_X32 FILLER_135_193 ();
 FILLCELL_X32 FILLER_135_225 ();
 FILLCELL_X32 FILLER_135_257 ();
 FILLCELL_X32 FILLER_135_289 ();
 FILLCELL_X32 FILLER_135_321 ();
 FILLCELL_X16 FILLER_135_353 ();
 FILLCELL_X8 FILLER_135_369 ();
 FILLCELL_X2 FILLER_135_377 ();
 FILLCELL_X1 FILLER_135_379 ();
 FILLCELL_X32 FILLER_135_1518 ();
 FILLCELL_X32 FILLER_135_1550 ();
 FILLCELL_X32 FILLER_135_1582 ();
 FILLCELL_X32 FILLER_135_1614 ();
 FILLCELL_X32 FILLER_135_1646 ();
 FILLCELL_X16 FILLER_135_1678 ();
 FILLCELL_X4 FILLER_135_1694 ();
 FILLCELL_X2 FILLER_135_1698 ();
 FILLCELL_X1 FILLER_135_1700 ();
 FILLCELL_X4 FILLER_136_1 ();
 FILLCELL_X32 FILLER_136_8 ();
 FILLCELL_X32 FILLER_136_40 ();
 FILLCELL_X32 FILLER_136_72 ();
 FILLCELL_X32 FILLER_136_104 ();
 FILLCELL_X32 FILLER_136_136 ();
 FILLCELL_X32 FILLER_136_168 ();
 FILLCELL_X32 FILLER_136_200 ();
 FILLCELL_X32 FILLER_136_232 ();
 FILLCELL_X32 FILLER_136_264 ();
 FILLCELL_X32 FILLER_136_296 ();
 FILLCELL_X32 FILLER_136_328 ();
 FILLCELL_X16 FILLER_136_360 ();
 FILLCELL_X4 FILLER_136_376 ();
 FILLCELL_X32 FILLER_136_1518 ();
 FILLCELL_X4 FILLER_136_1550 ();
 FILLCELL_X2 FILLER_136_1554 ();
 FILLCELL_X32 FILLER_136_1561 ();
 FILLCELL_X32 FILLER_136_1593 ();
 FILLCELL_X32 FILLER_136_1625 ();
 FILLCELL_X32 FILLER_136_1657 ();
 FILLCELL_X8 FILLER_136_1689 ();
 FILLCELL_X4 FILLER_136_1697 ();
 FILLCELL_X32 FILLER_137_1 ();
 FILLCELL_X32 FILLER_137_33 ();
 FILLCELL_X32 FILLER_137_65 ();
 FILLCELL_X32 FILLER_137_97 ();
 FILLCELL_X32 FILLER_137_129 ();
 FILLCELL_X32 FILLER_137_161 ();
 FILLCELL_X32 FILLER_137_193 ();
 FILLCELL_X32 FILLER_137_225 ();
 FILLCELL_X32 FILLER_137_257 ();
 FILLCELL_X32 FILLER_137_289 ();
 FILLCELL_X32 FILLER_137_321 ();
 FILLCELL_X16 FILLER_137_353 ();
 FILLCELL_X8 FILLER_137_369 ();
 FILLCELL_X2 FILLER_137_377 ();
 FILLCELL_X1 FILLER_137_379 ();
 FILLCELL_X32 FILLER_137_1518 ();
 FILLCELL_X32 FILLER_137_1550 ();
 FILLCELL_X32 FILLER_137_1582 ();
 FILLCELL_X32 FILLER_137_1614 ();
 FILLCELL_X32 FILLER_137_1646 ();
 FILLCELL_X16 FILLER_137_1678 ();
 FILLCELL_X4 FILLER_137_1694 ();
 FILLCELL_X2 FILLER_137_1698 ();
 FILLCELL_X1 FILLER_137_1700 ();
 FILLCELL_X32 FILLER_138_1 ();
 FILLCELL_X32 FILLER_138_33 ();
 FILLCELL_X32 FILLER_138_65 ();
 FILLCELL_X32 FILLER_138_97 ();
 FILLCELL_X32 FILLER_138_129 ();
 FILLCELL_X32 FILLER_138_161 ();
 FILLCELL_X32 FILLER_138_193 ();
 FILLCELL_X32 FILLER_138_225 ();
 FILLCELL_X32 FILLER_138_257 ();
 FILLCELL_X32 FILLER_138_289 ();
 FILLCELL_X32 FILLER_138_321 ();
 FILLCELL_X16 FILLER_138_353 ();
 FILLCELL_X8 FILLER_138_369 ();
 FILLCELL_X2 FILLER_138_377 ();
 FILLCELL_X1 FILLER_138_379 ();
 FILLCELL_X32 FILLER_138_1518 ();
 FILLCELL_X32 FILLER_138_1550 ();
 FILLCELL_X32 FILLER_138_1582 ();
 FILLCELL_X32 FILLER_138_1614 ();
 FILLCELL_X32 FILLER_138_1646 ();
 FILLCELL_X16 FILLER_138_1678 ();
 FILLCELL_X4 FILLER_138_1694 ();
 FILLCELL_X2 FILLER_138_1698 ();
 FILLCELL_X1 FILLER_138_1700 ();
 FILLCELL_X32 FILLER_139_1 ();
 FILLCELL_X32 FILLER_139_33 ();
 FILLCELL_X32 FILLER_139_65 ();
 FILLCELL_X32 FILLER_139_97 ();
 FILLCELL_X32 FILLER_139_129 ();
 FILLCELL_X32 FILLER_139_161 ();
 FILLCELL_X32 FILLER_139_193 ();
 FILLCELL_X32 FILLER_139_225 ();
 FILLCELL_X32 FILLER_139_257 ();
 FILLCELL_X32 FILLER_139_289 ();
 FILLCELL_X32 FILLER_139_321 ();
 FILLCELL_X16 FILLER_139_353 ();
 FILLCELL_X8 FILLER_139_369 ();
 FILLCELL_X2 FILLER_139_377 ();
 FILLCELL_X1 FILLER_139_379 ();
 FILLCELL_X32 FILLER_139_1518 ();
 FILLCELL_X32 FILLER_139_1550 ();
 FILLCELL_X32 FILLER_139_1582 ();
 FILLCELL_X32 FILLER_139_1614 ();
 FILLCELL_X32 FILLER_139_1646 ();
 FILLCELL_X16 FILLER_139_1678 ();
 FILLCELL_X4 FILLER_139_1694 ();
 FILLCELL_X2 FILLER_139_1698 ();
 FILLCELL_X1 FILLER_139_1700 ();
 FILLCELL_X32 FILLER_140_1 ();
 FILLCELL_X32 FILLER_140_33 ();
 FILLCELL_X32 FILLER_140_65 ();
 FILLCELL_X32 FILLER_140_97 ();
 FILLCELL_X32 FILLER_140_129 ();
 FILLCELL_X32 FILLER_140_161 ();
 FILLCELL_X32 FILLER_140_193 ();
 FILLCELL_X32 FILLER_140_225 ();
 FILLCELL_X32 FILLER_140_257 ();
 FILLCELL_X32 FILLER_140_289 ();
 FILLCELL_X32 FILLER_140_321 ();
 FILLCELL_X16 FILLER_140_353 ();
 FILLCELL_X8 FILLER_140_369 ();
 FILLCELL_X2 FILLER_140_377 ();
 FILLCELL_X1 FILLER_140_379 ();
 FILLCELL_X32 FILLER_140_1518 ();
 FILLCELL_X32 FILLER_140_1550 ();
 FILLCELL_X32 FILLER_140_1582 ();
 FILLCELL_X32 FILLER_140_1614 ();
 FILLCELL_X32 FILLER_140_1646 ();
 FILLCELL_X16 FILLER_140_1678 ();
 FILLCELL_X4 FILLER_140_1697 ();
 FILLCELL_X32 FILLER_141_1 ();
 FILLCELL_X32 FILLER_141_33 ();
 FILLCELL_X32 FILLER_141_65 ();
 FILLCELL_X32 FILLER_141_97 ();
 FILLCELL_X32 FILLER_141_129 ();
 FILLCELL_X32 FILLER_141_161 ();
 FILLCELL_X32 FILLER_141_193 ();
 FILLCELL_X32 FILLER_141_225 ();
 FILLCELL_X32 FILLER_141_257 ();
 FILLCELL_X32 FILLER_141_289 ();
 FILLCELL_X32 FILLER_141_321 ();
 FILLCELL_X16 FILLER_141_353 ();
 FILLCELL_X8 FILLER_141_369 ();
 FILLCELL_X2 FILLER_141_377 ();
 FILLCELL_X1 FILLER_141_379 ();
 FILLCELL_X32 FILLER_141_1518 ();
 FILLCELL_X32 FILLER_141_1550 ();
 FILLCELL_X32 FILLER_141_1582 ();
 FILLCELL_X32 FILLER_141_1614 ();
 FILLCELL_X32 FILLER_141_1646 ();
 FILLCELL_X16 FILLER_141_1678 ();
 FILLCELL_X4 FILLER_141_1694 ();
 FILLCELL_X2 FILLER_141_1698 ();
 FILLCELL_X1 FILLER_141_1700 ();
 FILLCELL_X32 FILLER_142_1 ();
 FILLCELL_X32 FILLER_142_33 ();
 FILLCELL_X32 FILLER_142_65 ();
 FILLCELL_X32 FILLER_142_97 ();
 FILLCELL_X32 FILLER_142_129 ();
 FILLCELL_X32 FILLER_142_161 ();
 FILLCELL_X32 FILLER_142_193 ();
 FILLCELL_X32 FILLER_142_225 ();
 FILLCELL_X32 FILLER_142_257 ();
 FILLCELL_X32 FILLER_142_289 ();
 FILLCELL_X32 FILLER_142_321 ();
 FILLCELL_X16 FILLER_142_353 ();
 FILLCELL_X8 FILLER_142_369 ();
 FILLCELL_X2 FILLER_142_377 ();
 FILLCELL_X1 FILLER_142_379 ();
 FILLCELL_X32 FILLER_142_1518 ();
 FILLCELL_X32 FILLER_142_1550 ();
 FILLCELL_X32 FILLER_142_1582 ();
 FILLCELL_X32 FILLER_142_1614 ();
 FILLCELL_X32 FILLER_142_1646 ();
 FILLCELL_X16 FILLER_142_1678 ();
 FILLCELL_X4 FILLER_142_1694 ();
 FILLCELL_X2 FILLER_142_1698 ();
 FILLCELL_X1 FILLER_142_1700 ();
 FILLCELL_X32 FILLER_143_1 ();
 FILLCELL_X32 FILLER_143_33 ();
 FILLCELL_X32 FILLER_143_65 ();
 FILLCELL_X32 FILLER_143_97 ();
 FILLCELL_X32 FILLER_143_129 ();
 FILLCELL_X32 FILLER_143_161 ();
 FILLCELL_X32 FILLER_143_193 ();
 FILLCELL_X32 FILLER_143_225 ();
 FILLCELL_X32 FILLER_143_257 ();
 FILLCELL_X32 FILLER_143_289 ();
 FILLCELL_X32 FILLER_143_321 ();
 FILLCELL_X16 FILLER_143_353 ();
 FILLCELL_X8 FILLER_143_369 ();
 FILLCELL_X2 FILLER_143_377 ();
 FILLCELL_X1 FILLER_143_379 ();
 FILLCELL_X32 FILLER_143_1518 ();
 FILLCELL_X32 FILLER_143_1550 ();
 FILLCELL_X32 FILLER_143_1582 ();
 FILLCELL_X32 FILLER_143_1614 ();
 FILLCELL_X32 FILLER_143_1646 ();
 FILLCELL_X16 FILLER_143_1678 ();
 FILLCELL_X4 FILLER_143_1694 ();
 FILLCELL_X2 FILLER_143_1698 ();
 FILLCELL_X1 FILLER_143_1700 ();
 FILLCELL_X32 FILLER_144_1 ();
 FILLCELL_X32 FILLER_144_33 ();
 FILLCELL_X32 FILLER_144_65 ();
 FILLCELL_X32 FILLER_144_97 ();
 FILLCELL_X32 FILLER_144_129 ();
 FILLCELL_X32 FILLER_144_161 ();
 FILLCELL_X32 FILLER_144_193 ();
 FILLCELL_X32 FILLER_144_225 ();
 FILLCELL_X32 FILLER_144_257 ();
 FILLCELL_X32 FILLER_144_289 ();
 FILLCELL_X32 FILLER_144_321 ();
 FILLCELL_X16 FILLER_144_353 ();
 FILLCELL_X8 FILLER_144_369 ();
 FILLCELL_X2 FILLER_144_377 ();
 FILLCELL_X1 FILLER_144_379 ();
 FILLCELL_X32 FILLER_144_1518 ();
 FILLCELL_X32 FILLER_144_1550 ();
 FILLCELL_X32 FILLER_144_1582 ();
 FILLCELL_X32 FILLER_144_1614 ();
 FILLCELL_X32 FILLER_144_1646 ();
 FILLCELL_X16 FILLER_144_1678 ();
 FILLCELL_X4 FILLER_144_1694 ();
 FILLCELL_X2 FILLER_144_1698 ();
 FILLCELL_X1 FILLER_144_1700 ();
 FILLCELL_X4 FILLER_145_1 ();
 FILLCELL_X32 FILLER_145_10 ();
 FILLCELL_X32 FILLER_145_42 ();
 FILLCELL_X32 FILLER_145_74 ();
 FILLCELL_X32 FILLER_145_106 ();
 FILLCELL_X32 FILLER_145_138 ();
 FILLCELL_X32 FILLER_145_170 ();
 FILLCELL_X32 FILLER_145_202 ();
 FILLCELL_X32 FILLER_145_234 ();
 FILLCELL_X32 FILLER_145_266 ();
 FILLCELL_X32 FILLER_145_298 ();
 FILLCELL_X32 FILLER_145_330 ();
 FILLCELL_X16 FILLER_145_362 ();
 FILLCELL_X2 FILLER_145_378 ();
 FILLCELL_X32 FILLER_145_1518 ();
 FILLCELL_X32 FILLER_145_1550 ();
 FILLCELL_X32 FILLER_145_1582 ();
 FILLCELL_X32 FILLER_145_1614 ();
 FILLCELL_X32 FILLER_145_1646 ();
 FILLCELL_X16 FILLER_145_1678 ();
 FILLCELL_X4 FILLER_145_1694 ();
 FILLCELL_X2 FILLER_145_1698 ();
 FILLCELL_X1 FILLER_145_1700 ();
 FILLCELL_X32 FILLER_146_1 ();
 FILLCELL_X32 FILLER_146_33 ();
 FILLCELL_X32 FILLER_146_65 ();
 FILLCELL_X32 FILLER_146_97 ();
 FILLCELL_X32 FILLER_146_129 ();
 FILLCELL_X32 FILLER_146_161 ();
 FILLCELL_X32 FILLER_146_193 ();
 FILLCELL_X32 FILLER_146_225 ();
 FILLCELL_X32 FILLER_146_257 ();
 FILLCELL_X32 FILLER_146_289 ();
 FILLCELL_X32 FILLER_146_321 ();
 FILLCELL_X16 FILLER_146_353 ();
 FILLCELL_X8 FILLER_146_369 ();
 FILLCELL_X2 FILLER_146_377 ();
 FILLCELL_X1 FILLER_146_379 ();
 FILLCELL_X32 FILLER_146_1518 ();
 FILLCELL_X32 FILLER_146_1550 ();
 FILLCELL_X32 FILLER_146_1582 ();
 FILLCELL_X32 FILLER_146_1614 ();
 FILLCELL_X32 FILLER_146_1646 ();
 FILLCELL_X16 FILLER_146_1678 ();
 FILLCELL_X4 FILLER_146_1694 ();
 FILLCELL_X2 FILLER_146_1698 ();
 FILLCELL_X1 FILLER_146_1700 ();
 FILLCELL_X32 FILLER_147_1 ();
 FILLCELL_X32 FILLER_147_33 ();
 FILLCELL_X32 FILLER_147_65 ();
 FILLCELL_X32 FILLER_147_97 ();
 FILLCELL_X32 FILLER_147_129 ();
 FILLCELL_X32 FILLER_147_161 ();
 FILLCELL_X32 FILLER_147_193 ();
 FILLCELL_X32 FILLER_147_225 ();
 FILLCELL_X32 FILLER_147_257 ();
 FILLCELL_X32 FILLER_147_289 ();
 FILLCELL_X32 FILLER_147_321 ();
 FILLCELL_X16 FILLER_147_353 ();
 FILLCELL_X8 FILLER_147_369 ();
 FILLCELL_X2 FILLER_147_377 ();
 FILLCELL_X1 FILLER_147_379 ();
 FILLCELL_X32 FILLER_147_1518 ();
 FILLCELL_X32 FILLER_147_1550 ();
 FILLCELL_X32 FILLER_147_1582 ();
 FILLCELL_X32 FILLER_147_1614 ();
 FILLCELL_X32 FILLER_147_1646 ();
 FILLCELL_X16 FILLER_147_1678 ();
 FILLCELL_X4 FILLER_147_1694 ();
 FILLCELL_X2 FILLER_147_1698 ();
 FILLCELL_X1 FILLER_147_1700 ();
 FILLCELL_X32 FILLER_148_1 ();
 FILLCELL_X32 FILLER_148_33 ();
 FILLCELL_X32 FILLER_148_65 ();
 FILLCELL_X32 FILLER_148_97 ();
 FILLCELL_X32 FILLER_148_129 ();
 FILLCELL_X32 FILLER_148_161 ();
 FILLCELL_X32 FILLER_148_193 ();
 FILLCELL_X32 FILLER_148_225 ();
 FILLCELL_X32 FILLER_148_257 ();
 FILLCELL_X32 FILLER_148_289 ();
 FILLCELL_X32 FILLER_148_321 ();
 FILLCELL_X16 FILLER_148_353 ();
 FILLCELL_X8 FILLER_148_369 ();
 FILLCELL_X2 FILLER_148_377 ();
 FILLCELL_X1 FILLER_148_379 ();
 FILLCELL_X32 FILLER_148_1518 ();
 FILLCELL_X32 FILLER_148_1550 ();
 FILLCELL_X32 FILLER_148_1582 ();
 FILLCELL_X32 FILLER_148_1614 ();
 FILLCELL_X32 FILLER_148_1646 ();
 FILLCELL_X16 FILLER_148_1678 ();
 FILLCELL_X4 FILLER_148_1694 ();
 FILLCELL_X2 FILLER_148_1698 ();
 FILLCELL_X1 FILLER_148_1700 ();
 FILLCELL_X32 FILLER_149_1 ();
 FILLCELL_X32 FILLER_149_33 ();
 FILLCELL_X32 FILLER_149_65 ();
 FILLCELL_X32 FILLER_149_97 ();
 FILLCELL_X32 FILLER_149_129 ();
 FILLCELL_X32 FILLER_149_161 ();
 FILLCELL_X32 FILLER_149_193 ();
 FILLCELL_X32 FILLER_149_225 ();
 FILLCELL_X32 FILLER_149_257 ();
 FILLCELL_X32 FILLER_149_289 ();
 FILLCELL_X32 FILLER_149_321 ();
 FILLCELL_X16 FILLER_149_353 ();
 FILLCELL_X8 FILLER_149_369 ();
 FILLCELL_X2 FILLER_149_377 ();
 FILLCELL_X1 FILLER_149_379 ();
 FILLCELL_X32 FILLER_149_1518 ();
 FILLCELL_X32 FILLER_149_1550 ();
 FILLCELL_X32 FILLER_149_1582 ();
 FILLCELL_X32 FILLER_149_1614 ();
 FILLCELL_X32 FILLER_149_1646 ();
 FILLCELL_X16 FILLER_149_1678 ();
 FILLCELL_X4 FILLER_149_1694 ();
 FILLCELL_X2 FILLER_149_1698 ();
 FILLCELL_X1 FILLER_149_1700 ();
 FILLCELL_X32 FILLER_150_1 ();
 FILLCELL_X32 FILLER_150_33 ();
 FILLCELL_X32 FILLER_150_65 ();
 FILLCELL_X32 FILLER_150_97 ();
 FILLCELL_X32 FILLER_150_129 ();
 FILLCELL_X32 FILLER_150_161 ();
 FILLCELL_X32 FILLER_150_193 ();
 FILLCELL_X32 FILLER_150_225 ();
 FILLCELL_X32 FILLER_150_257 ();
 FILLCELL_X32 FILLER_150_289 ();
 FILLCELL_X32 FILLER_150_321 ();
 FILLCELL_X16 FILLER_150_353 ();
 FILLCELL_X8 FILLER_150_369 ();
 FILLCELL_X2 FILLER_150_377 ();
 FILLCELL_X1 FILLER_150_379 ();
 FILLCELL_X32 FILLER_150_1518 ();
 FILLCELL_X32 FILLER_150_1550 ();
 FILLCELL_X32 FILLER_150_1582 ();
 FILLCELL_X32 FILLER_150_1614 ();
 FILLCELL_X32 FILLER_150_1646 ();
 FILLCELL_X16 FILLER_150_1678 ();
 FILLCELL_X4 FILLER_150_1697 ();
 FILLCELL_X32 FILLER_151_1 ();
 FILLCELL_X32 FILLER_151_33 ();
 FILLCELL_X32 FILLER_151_65 ();
 FILLCELL_X32 FILLER_151_97 ();
 FILLCELL_X32 FILLER_151_129 ();
 FILLCELL_X32 FILLER_151_161 ();
 FILLCELL_X32 FILLER_151_193 ();
 FILLCELL_X32 FILLER_151_225 ();
 FILLCELL_X32 FILLER_151_257 ();
 FILLCELL_X32 FILLER_151_289 ();
 FILLCELL_X32 FILLER_151_321 ();
 FILLCELL_X16 FILLER_151_353 ();
 FILLCELL_X8 FILLER_151_369 ();
 FILLCELL_X2 FILLER_151_377 ();
 FILLCELL_X1 FILLER_151_379 ();
 FILLCELL_X32 FILLER_151_1518 ();
 FILLCELL_X32 FILLER_151_1550 ();
 FILLCELL_X32 FILLER_151_1582 ();
 FILLCELL_X32 FILLER_151_1614 ();
 FILLCELL_X32 FILLER_151_1646 ();
 FILLCELL_X16 FILLER_151_1678 ();
 FILLCELL_X4 FILLER_151_1694 ();
 FILLCELL_X2 FILLER_151_1698 ();
 FILLCELL_X1 FILLER_151_1700 ();
 FILLCELL_X32 FILLER_152_1 ();
 FILLCELL_X32 FILLER_152_33 ();
 FILLCELL_X32 FILLER_152_65 ();
 FILLCELL_X32 FILLER_152_97 ();
 FILLCELL_X32 FILLER_152_129 ();
 FILLCELL_X32 FILLER_152_161 ();
 FILLCELL_X32 FILLER_152_193 ();
 FILLCELL_X32 FILLER_152_225 ();
 FILLCELL_X32 FILLER_152_257 ();
 FILLCELL_X32 FILLER_152_289 ();
 FILLCELL_X32 FILLER_152_321 ();
 FILLCELL_X16 FILLER_152_353 ();
 FILLCELL_X8 FILLER_152_369 ();
 FILLCELL_X2 FILLER_152_377 ();
 FILLCELL_X1 FILLER_152_379 ();
 FILLCELL_X32 FILLER_152_1518 ();
 FILLCELL_X32 FILLER_152_1550 ();
 FILLCELL_X32 FILLER_152_1582 ();
 FILLCELL_X32 FILLER_152_1614 ();
 FILLCELL_X32 FILLER_152_1646 ();
 FILLCELL_X16 FILLER_152_1678 ();
 FILLCELL_X4 FILLER_152_1694 ();
 FILLCELL_X2 FILLER_152_1698 ();
 FILLCELL_X1 FILLER_152_1700 ();
 FILLCELL_X32 FILLER_153_1 ();
 FILLCELL_X32 FILLER_153_33 ();
 FILLCELL_X32 FILLER_153_65 ();
 FILLCELL_X32 FILLER_153_97 ();
 FILLCELL_X32 FILLER_153_129 ();
 FILLCELL_X32 FILLER_153_161 ();
 FILLCELL_X32 FILLER_153_193 ();
 FILLCELL_X32 FILLER_153_225 ();
 FILLCELL_X32 FILLER_153_257 ();
 FILLCELL_X32 FILLER_153_289 ();
 FILLCELL_X32 FILLER_153_321 ();
 FILLCELL_X16 FILLER_153_353 ();
 FILLCELL_X8 FILLER_153_369 ();
 FILLCELL_X2 FILLER_153_377 ();
 FILLCELL_X1 FILLER_153_379 ();
 FILLCELL_X32 FILLER_153_1518 ();
 FILLCELL_X32 FILLER_153_1550 ();
 FILLCELL_X32 FILLER_153_1582 ();
 FILLCELL_X32 FILLER_153_1614 ();
 FILLCELL_X32 FILLER_153_1646 ();
 FILLCELL_X16 FILLER_153_1678 ();
 FILLCELL_X4 FILLER_153_1694 ();
 FILLCELL_X2 FILLER_153_1698 ();
 FILLCELL_X1 FILLER_153_1700 ();
 FILLCELL_X4 FILLER_154_1 ();
 FILLCELL_X32 FILLER_154_12 ();
 FILLCELL_X32 FILLER_154_44 ();
 FILLCELL_X32 FILLER_154_76 ();
 FILLCELL_X32 FILLER_154_108 ();
 FILLCELL_X32 FILLER_154_140 ();
 FILLCELL_X32 FILLER_154_172 ();
 FILLCELL_X32 FILLER_154_204 ();
 FILLCELL_X32 FILLER_154_236 ();
 FILLCELL_X32 FILLER_154_268 ();
 FILLCELL_X32 FILLER_154_300 ();
 FILLCELL_X32 FILLER_154_332 ();
 FILLCELL_X16 FILLER_154_364 ();
 FILLCELL_X32 FILLER_154_1518 ();
 FILLCELL_X32 FILLER_154_1550 ();
 FILLCELL_X32 FILLER_154_1582 ();
 FILLCELL_X32 FILLER_154_1614 ();
 FILLCELL_X32 FILLER_154_1646 ();
 FILLCELL_X16 FILLER_154_1678 ();
 FILLCELL_X4 FILLER_154_1694 ();
 FILLCELL_X2 FILLER_154_1698 ();
 FILLCELL_X1 FILLER_154_1700 ();
 FILLCELL_X32 FILLER_155_1 ();
 FILLCELL_X32 FILLER_155_33 ();
 FILLCELL_X32 FILLER_155_65 ();
 FILLCELL_X32 FILLER_155_97 ();
 FILLCELL_X32 FILLER_155_129 ();
 FILLCELL_X32 FILLER_155_161 ();
 FILLCELL_X32 FILLER_155_193 ();
 FILLCELL_X32 FILLER_155_225 ();
 FILLCELL_X32 FILLER_155_257 ();
 FILLCELL_X32 FILLER_155_289 ();
 FILLCELL_X32 FILLER_155_321 ();
 FILLCELL_X16 FILLER_155_353 ();
 FILLCELL_X8 FILLER_155_369 ();
 FILLCELL_X2 FILLER_155_377 ();
 FILLCELL_X1 FILLER_155_379 ();
 FILLCELL_X32 FILLER_155_1518 ();
 FILLCELL_X32 FILLER_155_1550 ();
 FILLCELL_X32 FILLER_155_1582 ();
 FILLCELL_X32 FILLER_155_1614 ();
 FILLCELL_X32 FILLER_155_1646 ();
 FILLCELL_X16 FILLER_155_1678 ();
 FILLCELL_X4 FILLER_155_1694 ();
 FILLCELL_X2 FILLER_155_1698 ();
 FILLCELL_X1 FILLER_155_1700 ();
 FILLCELL_X32 FILLER_156_1 ();
 FILLCELL_X32 FILLER_156_33 ();
 FILLCELL_X32 FILLER_156_65 ();
 FILLCELL_X32 FILLER_156_97 ();
 FILLCELL_X32 FILLER_156_129 ();
 FILLCELL_X32 FILLER_156_161 ();
 FILLCELL_X32 FILLER_156_193 ();
 FILLCELL_X32 FILLER_156_225 ();
 FILLCELL_X32 FILLER_156_257 ();
 FILLCELL_X32 FILLER_156_289 ();
 FILLCELL_X32 FILLER_156_321 ();
 FILLCELL_X16 FILLER_156_353 ();
 FILLCELL_X8 FILLER_156_369 ();
 FILLCELL_X2 FILLER_156_377 ();
 FILLCELL_X1 FILLER_156_379 ();
 FILLCELL_X32 FILLER_156_1518 ();
 FILLCELL_X32 FILLER_156_1550 ();
 FILLCELL_X32 FILLER_156_1582 ();
 FILLCELL_X32 FILLER_156_1614 ();
 FILLCELL_X32 FILLER_156_1646 ();
 FILLCELL_X16 FILLER_156_1678 ();
 FILLCELL_X4 FILLER_156_1694 ();
 FILLCELL_X2 FILLER_156_1698 ();
 FILLCELL_X1 FILLER_156_1700 ();
 FILLCELL_X32 FILLER_157_1 ();
 FILLCELL_X32 FILLER_157_33 ();
 FILLCELL_X32 FILLER_157_65 ();
 FILLCELL_X32 FILLER_157_97 ();
 FILLCELL_X32 FILLER_157_129 ();
 FILLCELL_X32 FILLER_157_161 ();
 FILLCELL_X32 FILLER_157_193 ();
 FILLCELL_X32 FILLER_157_225 ();
 FILLCELL_X32 FILLER_157_257 ();
 FILLCELL_X32 FILLER_157_289 ();
 FILLCELL_X32 FILLER_157_321 ();
 FILLCELL_X16 FILLER_157_353 ();
 FILLCELL_X8 FILLER_157_369 ();
 FILLCELL_X2 FILLER_157_377 ();
 FILLCELL_X1 FILLER_157_379 ();
 FILLCELL_X32 FILLER_157_1518 ();
 FILLCELL_X32 FILLER_157_1550 ();
 FILLCELL_X32 FILLER_157_1582 ();
 FILLCELL_X32 FILLER_157_1614 ();
 FILLCELL_X32 FILLER_157_1646 ();
 FILLCELL_X16 FILLER_157_1678 ();
 FILLCELL_X4 FILLER_157_1694 ();
 FILLCELL_X2 FILLER_157_1698 ();
 FILLCELL_X1 FILLER_157_1700 ();
 FILLCELL_X32 FILLER_158_1 ();
 FILLCELL_X32 FILLER_158_33 ();
 FILLCELL_X32 FILLER_158_65 ();
 FILLCELL_X32 FILLER_158_97 ();
 FILLCELL_X32 FILLER_158_129 ();
 FILLCELL_X32 FILLER_158_161 ();
 FILLCELL_X32 FILLER_158_193 ();
 FILLCELL_X32 FILLER_158_225 ();
 FILLCELL_X32 FILLER_158_257 ();
 FILLCELL_X32 FILLER_158_289 ();
 FILLCELL_X32 FILLER_158_321 ();
 FILLCELL_X16 FILLER_158_353 ();
 FILLCELL_X8 FILLER_158_369 ();
 FILLCELL_X2 FILLER_158_377 ();
 FILLCELL_X1 FILLER_158_379 ();
 FILLCELL_X32 FILLER_158_1518 ();
 FILLCELL_X32 FILLER_158_1550 ();
 FILLCELL_X32 FILLER_158_1582 ();
 FILLCELL_X32 FILLER_158_1614 ();
 FILLCELL_X32 FILLER_158_1646 ();
 FILLCELL_X16 FILLER_158_1678 ();
 FILLCELL_X4 FILLER_158_1694 ();
 FILLCELL_X2 FILLER_158_1698 ();
 FILLCELL_X1 FILLER_158_1700 ();
 FILLCELL_X32 FILLER_159_1 ();
 FILLCELL_X32 FILLER_159_33 ();
 FILLCELL_X32 FILLER_159_65 ();
 FILLCELL_X32 FILLER_159_97 ();
 FILLCELL_X32 FILLER_159_129 ();
 FILLCELL_X32 FILLER_159_161 ();
 FILLCELL_X32 FILLER_159_193 ();
 FILLCELL_X32 FILLER_159_225 ();
 FILLCELL_X32 FILLER_159_257 ();
 FILLCELL_X32 FILLER_159_289 ();
 FILLCELL_X32 FILLER_159_321 ();
 FILLCELL_X16 FILLER_159_353 ();
 FILLCELL_X8 FILLER_159_369 ();
 FILLCELL_X2 FILLER_159_377 ();
 FILLCELL_X1 FILLER_159_379 ();
 FILLCELL_X32 FILLER_159_1518 ();
 FILLCELL_X32 FILLER_159_1550 ();
 FILLCELL_X32 FILLER_159_1582 ();
 FILLCELL_X32 FILLER_159_1614 ();
 FILLCELL_X32 FILLER_159_1646 ();
 FILLCELL_X16 FILLER_159_1678 ();
 FILLCELL_X4 FILLER_159_1697 ();
 FILLCELL_X32 FILLER_160_1 ();
 FILLCELL_X32 FILLER_160_33 ();
 FILLCELL_X32 FILLER_160_65 ();
 FILLCELL_X32 FILLER_160_97 ();
 FILLCELL_X32 FILLER_160_129 ();
 FILLCELL_X32 FILLER_160_161 ();
 FILLCELL_X32 FILLER_160_193 ();
 FILLCELL_X32 FILLER_160_225 ();
 FILLCELL_X32 FILLER_160_257 ();
 FILLCELL_X32 FILLER_160_289 ();
 FILLCELL_X32 FILLER_160_321 ();
 FILLCELL_X16 FILLER_160_353 ();
 FILLCELL_X8 FILLER_160_369 ();
 FILLCELL_X2 FILLER_160_377 ();
 FILLCELL_X1 FILLER_160_379 ();
 FILLCELL_X32 FILLER_160_1518 ();
 FILLCELL_X32 FILLER_160_1550 ();
 FILLCELL_X32 FILLER_160_1582 ();
 FILLCELL_X32 FILLER_160_1614 ();
 FILLCELL_X32 FILLER_160_1646 ();
 FILLCELL_X16 FILLER_160_1678 ();
 FILLCELL_X4 FILLER_160_1694 ();
 FILLCELL_X2 FILLER_160_1698 ();
 FILLCELL_X1 FILLER_160_1700 ();
 FILLCELL_X32 FILLER_161_1 ();
 FILLCELL_X32 FILLER_161_33 ();
 FILLCELL_X32 FILLER_161_65 ();
 FILLCELL_X32 FILLER_161_97 ();
 FILLCELL_X32 FILLER_161_129 ();
 FILLCELL_X32 FILLER_161_161 ();
 FILLCELL_X32 FILLER_161_193 ();
 FILLCELL_X32 FILLER_161_225 ();
 FILLCELL_X32 FILLER_161_257 ();
 FILLCELL_X32 FILLER_161_289 ();
 FILLCELL_X32 FILLER_161_321 ();
 FILLCELL_X16 FILLER_161_353 ();
 FILLCELL_X8 FILLER_161_369 ();
 FILLCELL_X2 FILLER_161_377 ();
 FILLCELL_X1 FILLER_161_379 ();
 FILLCELL_X32 FILLER_161_1518 ();
 FILLCELL_X32 FILLER_161_1550 ();
 FILLCELL_X32 FILLER_161_1582 ();
 FILLCELL_X32 FILLER_161_1614 ();
 FILLCELL_X32 FILLER_161_1646 ();
 FILLCELL_X16 FILLER_161_1678 ();
 FILLCELL_X4 FILLER_161_1694 ();
 FILLCELL_X2 FILLER_161_1698 ();
 FILLCELL_X1 FILLER_161_1700 ();
 FILLCELL_X32 FILLER_162_1 ();
 FILLCELL_X32 FILLER_162_33 ();
 FILLCELL_X32 FILLER_162_65 ();
 FILLCELL_X32 FILLER_162_97 ();
 FILLCELL_X32 FILLER_162_129 ();
 FILLCELL_X32 FILLER_162_161 ();
 FILLCELL_X32 FILLER_162_193 ();
 FILLCELL_X32 FILLER_162_225 ();
 FILLCELL_X32 FILLER_162_257 ();
 FILLCELL_X32 FILLER_162_289 ();
 FILLCELL_X32 FILLER_162_321 ();
 FILLCELL_X16 FILLER_162_353 ();
 FILLCELL_X8 FILLER_162_369 ();
 FILLCELL_X2 FILLER_162_377 ();
 FILLCELL_X1 FILLER_162_379 ();
 FILLCELL_X32 FILLER_162_1518 ();
 FILLCELL_X32 FILLER_162_1550 ();
 FILLCELL_X32 FILLER_162_1582 ();
 FILLCELL_X32 FILLER_162_1614 ();
 FILLCELL_X32 FILLER_162_1646 ();
 FILLCELL_X16 FILLER_162_1678 ();
 FILLCELL_X4 FILLER_162_1694 ();
 FILLCELL_X2 FILLER_162_1698 ();
 FILLCELL_X1 FILLER_162_1700 ();
 FILLCELL_X4 FILLER_163_1 ();
 FILLCELL_X32 FILLER_163_8 ();
 FILLCELL_X32 FILLER_163_40 ();
 FILLCELL_X32 FILLER_163_72 ();
 FILLCELL_X32 FILLER_163_104 ();
 FILLCELL_X32 FILLER_163_136 ();
 FILLCELL_X32 FILLER_163_168 ();
 FILLCELL_X32 FILLER_163_200 ();
 FILLCELL_X32 FILLER_163_232 ();
 FILLCELL_X32 FILLER_163_264 ();
 FILLCELL_X32 FILLER_163_296 ();
 FILLCELL_X32 FILLER_163_328 ();
 FILLCELL_X16 FILLER_163_360 ();
 FILLCELL_X4 FILLER_163_376 ();
 FILLCELL_X32 FILLER_163_1518 ();
 FILLCELL_X32 FILLER_163_1550 ();
 FILLCELL_X32 FILLER_163_1582 ();
 FILLCELL_X32 FILLER_163_1614 ();
 FILLCELL_X32 FILLER_163_1646 ();
 FILLCELL_X16 FILLER_163_1678 ();
 FILLCELL_X4 FILLER_163_1694 ();
 FILLCELL_X2 FILLER_163_1698 ();
 FILLCELL_X1 FILLER_163_1700 ();
 FILLCELL_X32 FILLER_164_1 ();
 FILLCELL_X32 FILLER_164_33 ();
 FILLCELL_X32 FILLER_164_65 ();
 FILLCELL_X32 FILLER_164_97 ();
 FILLCELL_X32 FILLER_164_129 ();
 FILLCELL_X32 FILLER_164_161 ();
 FILLCELL_X32 FILLER_164_193 ();
 FILLCELL_X32 FILLER_164_225 ();
 FILLCELL_X32 FILLER_164_257 ();
 FILLCELL_X32 FILLER_164_289 ();
 FILLCELL_X32 FILLER_164_321 ();
 FILLCELL_X16 FILLER_164_353 ();
 FILLCELL_X8 FILLER_164_369 ();
 FILLCELL_X2 FILLER_164_377 ();
 FILLCELL_X1 FILLER_164_379 ();
 FILLCELL_X32 FILLER_164_1518 ();
 FILLCELL_X32 FILLER_164_1550 ();
 FILLCELL_X32 FILLER_164_1582 ();
 FILLCELL_X32 FILLER_164_1614 ();
 FILLCELL_X32 FILLER_164_1646 ();
 FILLCELL_X16 FILLER_164_1678 ();
 FILLCELL_X4 FILLER_164_1694 ();
 FILLCELL_X2 FILLER_164_1698 ();
 FILLCELL_X1 FILLER_164_1700 ();
 FILLCELL_X32 FILLER_165_1 ();
 FILLCELL_X32 FILLER_165_33 ();
 FILLCELL_X32 FILLER_165_65 ();
 FILLCELL_X32 FILLER_165_97 ();
 FILLCELL_X32 FILLER_165_129 ();
 FILLCELL_X32 FILLER_165_161 ();
 FILLCELL_X32 FILLER_165_193 ();
 FILLCELL_X32 FILLER_165_225 ();
 FILLCELL_X32 FILLER_165_257 ();
 FILLCELL_X32 FILLER_165_289 ();
 FILLCELL_X32 FILLER_165_321 ();
 FILLCELL_X16 FILLER_165_353 ();
 FILLCELL_X8 FILLER_165_369 ();
 FILLCELL_X2 FILLER_165_377 ();
 FILLCELL_X1 FILLER_165_379 ();
 FILLCELL_X32 FILLER_165_1518 ();
 FILLCELL_X32 FILLER_165_1550 ();
 FILLCELL_X32 FILLER_165_1582 ();
 FILLCELL_X32 FILLER_165_1614 ();
 FILLCELL_X32 FILLER_165_1646 ();
 FILLCELL_X16 FILLER_165_1678 ();
 FILLCELL_X4 FILLER_165_1694 ();
 FILLCELL_X2 FILLER_165_1698 ();
 FILLCELL_X1 FILLER_165_1700 ();
 FILLCELL_X32 FILLER_166_1 ();
 FILLCELL_X32 FILLER_166_33 ();
 FILLCELL_X32 FILLER_166_65 ();
 FILLCELL_X32 FILLER_166_97 ();
 FILLCELL_X32 FILLER_166_129 ();
 FILLCELL_X32 FILLER_166_161 ();
 FILLCELL_X32 FILLER_166_193 ();
 FILLCELL_X32 FILLER_166_225 ();
 FILLCELL_X32 FILLER_166_257 ();
 FILLCELL_X32 FILLER_166_289 ();
 FILLCELL_X32 FILLER_166_321 ();
 FILLCELL_X16 FILLER_166_353 ();
 FILLCELL_X8 FILLER_166_369 ();
 FILLCELL_X2 FILLER_166_377 ();
 FILLCELL_X1 FILLER_166_379 ();
 FILLCELL_X32 FILLER_166_1518 ();
 FILLCELL_X32 FILLER_166_1550 ();
 FILLCELL_X32 FILLER_166_1582 ();
 FILLCELL_X32 FILLER_166_1614 ();
 FILLCELL_X32 FILLER_166_1646 ();
 FILLCELL_X16 FILLER_166_1678 ();
 FILLCELL_X4 FILLER_166_1694 ();
 FILLCELL_X2 FILLER_166_1698 ();
 FILLCELL_X1 FILLER_166_1700 ();
 FILLCELL_X32 FILLER_167_1 ();
 FILLCELL_X32 FILLER_167_33 ();
 FILLCELL_X32 FILLER_167_65 ();
 FILLCELL_X32 FILLER_167_97 ();
 FILLCELL_X32 FILLER_167_129 ();
 FILLCELL_X32 FILLER_167_161 ();
 FILLCELL_X32 FILLER_167_193 ();
 FILLCELL_X32 FILLER_167_225 ();
 FILLCELL_X32 FILLER_167_257 ();
 FILLCELL_X32 FILLER_167_289 ();
 FILLCELL_X32 FILLER_167_321 ();
 FILLCELL_X16 FILLER_167_353 ();
 FILLCELL_X8 FILLER_167_369 ();
 FILLCELL_X2 FILLER_167_377 ();
 FILLCELL_X1 FILLER_167_379 ();
 FILLCELL_X32 FILLER_167_1518 ();
 FILLCELL_X32 FILLER_167_1550 ();
 FILLCELL_X32 FILLER_167_1582 ();
 FILLCELL_X32 FILLER_167_1614 ();
 FILLCELL_X32 FILLER_167_1646 ();
 FILLCELL_X16 FILLER_167_1678 ();
 FILLCELL_X4 FILLER_167_1694 ();
 FILLCELL_X2 FILLER_167_1698 ();
 FILLCELL_X1 FILLER_167_1700 ();
 FILLCELL_X32 FILLER_168_1 ();
 FILLCELL_X32 FILLER_168_33 ();
 FILLCELL_X32 FILLER_168_65 ();
 FILLCELL_X32 FILLER_168_97 ();
 FILLCELL_X32 FILLER_168_129 ();
 FILLCELL_X32 FILLER_168_161 ();
 FILLCELL_X32 FILLER_168_193 ();
 FILLCELL_X32 FILLER_168_225 ();
 FILLCELL_X32 FILLER_168_257 ();
 FILLCELL_X32 FILLER_168_289 ();
 FILLCELL_X32 FILLER_168_321 ();
 FILLCELL_X16 FILLER_168_353 ();
 FILLCELL_X8 FILLER_168_369 ();
 FILLCELL_X2 FILLER_168_377 ();
 FILLCELL_X1 FILLER_168_379 ();
 FILLCELL_X32 FILLER_168_1518 ();
 FILLCELL_X32 FILLER_168_1550 ();
 FILLCELL_X32 FILLER_168_1582 ();
 FILLCELL_X32 FILLER_168_1614 ();
 FILLCELL_X32 FILLER_168_1646 ();
 FILLCELL_X8 FILLER_168_1678 ();
 FILLCELL_X4 FILLER_168_1686 ();
 FILLCELL_X2 FILLER_168_1690 ();
 FILLCELL_X4 FILLER_168_1697 ();
 FILLCELL_X32 FILLER_169_1 ();
 FILLCELL_X32 FILLER_169_33 ();
 FILLCELL_X32 FILLER_169_65 ();
 FILLCELL_X32 FILLER_169_97 ();
 FILLCELL_X32 FILLER_169_129 ();
 FILLCELL_X32 FILLER_169_161 ();
 FILLCELL_X32 FILLER_169_193 ();
 FILLCELL_X32 FILLER_169_225 ();
 FILLCELL_X32 FILLER_169_257 ();
 FILLCELL_X32 FILLER_169_289 ();
 FILLCELL_X32 FILLER_169_321 ();
 FILLCELL_X16 FILLER_169_353 ();
 FILLCELL_X8 FILLER_169_369 ();
 FILLCELL_X2 FILLER_169_377 ();
 FILLCELL_X1 FILLER_169_379 ();
 FILLCELL_X32 FILLER_169_1518 ();
 FILLCELL_X32 FILLER_169_1550 ();
 FILLCELL_X32 FILLER_169_1582 ();
 FILLCELL_X32 FILLER_169_1614 ();
 FILLCELL_X32 FILLER_169_1646 ();
 FILLCELL_X16 FILLER_169_1678 ();
 FILLCELL_X4 FILLER_169_1694 ();
 FILLCELL_X2 FILLER_169_1698 ();
 FILLCELL_X1 FILLER_169_1700 ();
 FILLCELL_X32 FILLER_170_1 ();
 FILLCELL_X32 FILLER_170_33 ();
 FILLCELL_X32 FILLER_170_65 ();
 FILLCELL_X32 FILLER_170_97 ();
 FILLCELL_X32 FILLER_170_129 ();
 FILLCELL_X32 FILLER_170_161 ();
 FILLCELL_X32 FILLER_170_193 ();
 FILLCELL_X32 FILLER_170_225 ();
 FILLCELL_X32 FILLER_170_257 ();
 FILLCELL_X32 FILLER_170_289 ();
 FILLCELL_X32 FILLER_170_321 ();
 FILLCELL_X16 FILLER_170_353 ();
 FILLCELL_X8 FILLER_170_369 ();
 FILLCELL_X2 FILLER_170_377 ();
 FILLCELL_X1 FILLER_170_379 ();
 FILLCELL_X32 FILLER_170_1518 ();
 FILLCELL_X32 FILLER_170_1550 ();
 FILLCELL_X32 FILLER_170_1582 ();
 FILLCELL_X32 FILLER_170_1614 ();
 FILLCELL_X32 FILLER_170_1646 ();
 FILLCELL_X16 FILLER_170_1678 ();
 FILLCELL_X4 FILLER_170_1694 ();
 FILLCELL_X2 FILLER_170_1698 ();
 FILLCELL_X1 FILLER_170_1700 ();
 FILLCELL_X32 FILLER_171_1 ();
 FILLCELL_X32 FILLER_171_33 ();
 FILLCELL_X32 FILLER_171_65 ();
 FILLCELL_X32 FILLER_171_97 ();
 FILLCELL_X32 FILLER_171_129 ();
 FILLCELL_X32 FILLER_171_161 ();
 FILLCELL_X32 FILLER_171_193 ();
 FILLCELL_X32 FILLER_171_225 ();
 FILLCELL_X32 FILLER_171_257 ();
 FILLCELL_X32 FILLER_171_289 ();
 FILLCELL_X32 FILLER_171_321 ();
 FILLCELL_X16 FILLER_171_353 ();
 FILLCELL_X8 FILLER_171_369 ();
 FILLCELL_X2 FILLER_171_377 ();
 FILLCELL_X1 FILLER_171_379 ();
 FILLCELL_X32 FILLER_171_1518 ();
 FILLCELL_X32 FILLER_171_1550 ();
 FILLCELL_X32 FILLER_171_1582 ();
 FILLCELL_X32 FILLER_171_1614 ();
 FILLCELL_X32 FILLER_171_1646 ();
 FILLCELL_X16 FILLER_171_1678 ();
 FILLCELL_X4 FILLER_171_1694 ();
 FILLCELL_X2 FILLER_171_1698 ();
 FILLCELL_X1 FILLER_171_1700 ();
 FILLCELL_X32 FILLER_172_1 ();
 FILLCELL_X32 FILLER_172_33 ();
 FILLCELL_X32 FILLER_172_65 ();
 FILLCELL_X32 FILLER_172_97 ();
 FILLCELL_X32 FILLER_172_129 ();
 FILLCELL_X32 FILLER_172_161 ();
 FILLCELL_X32 FILLER_172_193 ();
 FILLCELL_X32 FILLER_172_225 ();
 FILLCELL_X32 FILLER_172_257 ();
 FILLCELL_X32 FILLER_172_289 ();
 FILLCELL_X32 FILLER_172_321 ();
 FILLCELL_X16 FILLER_172_353 ();
 FILLCELL_X8 FILLER_172_369 ();
 FILLCELL_X2 FILLER_172_377 ();
 FILLCELL_X1 FILLER_172_379 ();
 FILLCELL_X32 FILLER_172_1518 ();
 FILLCELL_X32 FILLER_172_1550 ();
 FILLCELL_X32 FILLER_172_1582 ();
 FILLCELL_X32 FILLER_172_1614 ();
 FILLCELL_X32 FILLER_172_1646 ();
 FILLCELL_X16 FILLER_172_1678 ();
 FILLCELL_X4 FILLER_172_1694 ();
 FILLCELL_X2 FILLER_172_1698 ();
 FILLCELL_X1 FILLER_172_1700 ();
 FILLCELL_X4 FILLER_173_1 ();
 FILLCELL_X32 FILLER_173_10 ();
 FILLCELL_X32 FILLER_173_42 ();
 FILLCELL_X32 FILLER_173_74 ();
 FILLCELL_X32 FILLER_173_106 ();
 FILLCELL_X32 FILLER_173_138 ();
 FILLCELL_X32 FILLER_173_170 ();
 FILLCELL_X32 FILLER_173_202 ();
 FILLCELL_X32 FILLER_173_234 ();
 FILLCELL_X32 FILLER_173_266 ();
 FILLCELL_X32 FILLER_173_298 ();
 FILLCELL_X32 FILLER_173_330 ();
 FILLCELL_X16 FILLER_173_362 ();
 FILLCELL_X2 FILLER_173_378 ();
 FILLCELL_X32 FILLER_173_1518 ();
 FILLCELL_X32 FILLER_173_1550 ();
 FILLCELL_X32 FILLER_173_1582 ();
 FILLCELL_X32 FILLER_173_1614 ();
 FILLCELL_X32 FILLER_173_1646 ();
 FILLCELL_X16 FILLER_173_1678 ();
 FILLCELL_X4 FILLER_173_1694 ();
 FILLCELL_X2 FILLER_173_1698 ();
 FILLCELL_X1 FILLER_173_1700 ();
 FILLCELL_X32 FILLER_174_1 ();
 FILLCELL_X32 FILLER_174_33 ();
 FILLCELL_X32 FILLER_174_65 ();
 FILLCELL_X32 FILLER_174_97 ();
 FILLCELL_X32 FILLER_174_129 ();
 FILLCELL_X32 FILLER_174_161 ();
 FILLCELL_X32 FILLER_174_193 ();
 FILLCELL_X32 FILLER_174_225 ();
 FILLCELL_X32 FILLER_174_257 ();
 FILLCELL_X32 FILLER_174_289 ();
 FILLCELL_X32 FILLER_174_321 ();
 FILLCELL_X16 FILLER_174_353 ();
 FILLCELL_X8 FILLER_174_369 ();
 FILLCELL_X2 FILLER_174_377 ();
 FILLCELL_X1 FILLER_174_379 ();
 FILLCELL_X32 FILLER_174_1518 ();
 FILLCELL_X32 FILLER_174_1550 ();
 FILLCELL_X32 FILLER_174_1582 ();
 FILLCELL_X32 FILLER_174_1614 ();
 FILLCELL_X32 FILLER_174_1646 ();
 FILLCELL_X16 FILLER_174_1678 ();
 FILLCELL_X4 FILLER_174_1694 ();
 FILLCELL_X2 FILLER_174_1698 ();
 FILLCELL_X1 FILLER_174_1700 ();
 FILLCELL_X32 FILLER_175_1 ();
 FILLCELL_X32 FILLER_175_33 ();
 FILLCELL_X32 FILLER_175_65 ();
 FILLCELL_X32 FILLER_175_97 ();
 FILLCELL_X32 FILLER_175_129 ();
 FILLCELL_X32 FILLER_175_161 ();
 FILLCELL_X32 FILLER_175_193 ();
 FILLCELL_X32 FILLER_175_225 ();
 FILLCELL_X32 FILLER_175_257 ();
 FILLCELL_X32 FILLER_175_289 ();
 FILLCELL_X32 FILLER_175_321 ();
 FILLCELL_X16 FILLER_175_353 ();
 FILLCELL_X8 FILLER_175_369 ();
 FILLCELL_X2 FILLER_175_377 ();
 FILLCELL_X1 FILLER_175_379 ();
 FILLCELL_X32 FILLER_175_1518 ();
 FILLCELL_X32 FILLER_175_1550 ();
 FILLCELL_X32 FILLER_175_1582 ();
 FILLCELL_X32 FILLER_175_1614 ();
 FILLCELL_X32 FILLER_175_1646 ();
 FILLCELL_X16 FILLER_175_1678 ();
 FILLCELL_X4 FILLER_175_1694 ();
 FILLCELL_X2 FILLER_175_1698 ();
 FILLCELL_X1 FILLER_175_1700 ();
 FILLCELL_X32 FILLER_176_1 ();
 FILLCELL_X32 FILLER_176_33 ();
 FILLCELL_X32 FILLER_176_65 ();
 FILLCELL_X32 FILLER_176_97 ();
 FILLCELL_X32 FILLER_176_129 ();
 FILLCELL_X32 FILLER_176_161 ();
 FILLCELL_X32 FILLER_176_193 ();
 FILLCELL_X32 FILLER_176_225 ();
 FILLCELL_X32 FILLER_176_257 ();
 FILLCELL_X32 FILLER_176_289 ();
 FILLCELL_X32 FILLER_176_321 ();
 FILLCELL_X16 FILLER_176_353 ();
 FILLCELL_X8 FILLER_176_369 ();
 FILLCELL_X2 FILLER_176_377 ();
 FILLCELL_X1 FILLER_176_379 ();
 FILLCELL_X32 FILLER_176_1518 ();
 FILLCELL_X32 FILLER_176_1550 ();
 FILLCELL_X32 FILLER_176_1582 ();
 FILLCELL_X32 FILLER_176_1614 ();
 FILLCELL_X32 FILLER_176_1646 ();
 FILLCELL_X16 FILLER_176_1678 ();
 FILLCELL_X4 FILLER_176_1694 ();
 FILLCELL_X2 FILLER_176_1698 ();
 FILLCELL_X1 FILLER_176_1700 ();
 FILLCELL_X32 FILLER_177_1 ();
 FILLCELL_X32 FILLER_177_33 ();
 FILLCELL_X32 FILLER_177_65 ();
 FILLCELL_X32 FILLER_177_97 ();
 FILLCELL_X32 FILLER_177_129 ();
 FILLCELL_X32 FILLER_177_161 ();
 FILLCELL_X32 FILLER_177_193 ();
 FILLCELL_X32 FILLER_177_225 ();
 FILLCELL_X32 FILLER_177_257 ();
 FILLCELL_X32 FILLER_177_289 ();
 FILLCELL_X32 FILLER_177_321 ();
 FILLCELL_X16 FILLER_177_353 ();
 FILLCELL_X8 FILLER_177_369 ();
 FILLCELL_X2 FILLER_177_377 ();
 FILLCELL_X1 FILLER_177_379 ();
 FILLCELL_X32 FILLER_177_1518 ();
 FILLCELL_X32 FILLER_177_1550 ();
 FILLCELL_X32 FILLER_177_1582 ();
 FILLCELL_X32 FILLER_177_1614 ();
 FILLCELL_X32 FILLER_177_1646 ();
 FILLCELL_X16 FILLER_177_1678 ();
 FILLCELL_X4 FILLER_177_1694 ();
 FILLCELL_X2 FILLER_177_1698 ();
 FILLCELL_X1 FILLER_177_1700 ();
 FILLCELL_X32 FILLER_178_1 ();
 FILLCELL_X32 FILLER_178_33 ();
 FILLCELL_X32 FILLER_178_65 ();
 FILLCELL_X32 FILLER_178_97 ();
 FILLCELL_X32 FILLER_178_129 ();
 FILLCELL_X32 FILLER_178_161 ();
 FILLCELL_X32 FILLER_178_193 ();
 FILLCELL_X32 FILLER_178_225 ();
 FILLCELL_X32 FILLER_178_257 ();
 FILLCELL_X32 FILLER_178_289 ();
 FILLCELL_X32 FILLER_178_321 ();
 FILLCELL_X16 FILLER_178_353 ();
 FILLCELL_X8 FILLER_178_369 ();
 FILLCELL_X2 FILLER_178_377 ();
 FILLCELL_X1 FILLER_178_379 ();
 FILLCELL_X32 FILLER_178_1518 ();
 FILLCELL_X32 FILLER_178_1550 ();
 FILLCELL_X32 FILLER_178_1582 ();
 FILLCELL_X32 FILLER_178_1614 ();
 FILLCELL_X32 FILLER_178_1646 ();
 FILLCELL_X16 FILLER_178_1678 ();
 FILLCELL_X4 FILLER_178_1697 ();
 FILLCELL_X32 FILLER_179_1 ();
 FILLCELL_X32 FILLER_179_33 ();
 FILLCELL_X32 FILLER_179_65 ();
 FILLCELL_X32 FILLER_179_97 ();
 FILLCELL_X32 FILLER_179_129 ();
 FILLCELL_X32 FILLER_179_161 ();
 FILLCELL_X32 FILLER_179_193 ();
 FILLCELL_X32 FILLER_179_225 ();
 FILLCELL_X32 FILLER_179_257 ();
 FILLCELL_X32 FILLER_179_289 ();
 FILLCELL_X32 FILLER_179_321 ();
 FILLCELL_X16 FILLER_179_353 ();
 FILLCELL_X8 FILLER_179_369 ();
 FILLCELL_X2 FILLER_179_377 ();
 FILLCELL_X1 FILLER_179_379 ();
 FILLCELL_X32 FILLER_179_1518 ();
 FILLCELL_X32 FILLER_179_1550 ();
 FILLCELL_X32 FILLER_179_1582 ();
 FILLCELL_X32 FILLER_179_1614 ();
 FILLCELL_X32 FILLER_179_1646 ();
 FILLCELL_X16 FILLER_179_1678 ();
 FILLCELL_X4 FILLER_179_1694 ();
 FILLCELL_X2 FILLER_179_1698 ();
 FILLCELL_X1 FILLER_179_1700 ();
 FILLCELL_X32 FILLER_180_1 ();
 FILLCELL_X32 FILLER_180_33 ();
 FILLCELL_X32 FILLER_180_65 ();
 FILLCELL_X32 FILLER_180_97 ();
 FILLCELL_X32 FILLER_180_129 ();
 FILLCELL_X32 FILLER_180_161 ();
 FILLCELL_X32 FILLER_180_193 ();
 FILLCELL_X32 FILLER_180_225 ();
 FILLCELL_X32 FILLER_180_257 ();
 FILLCELL_X32 FILLER_180_289 ();
 FILLCELL_X32 FILLER_180_321 ();
 FILLCELL_X16 FILLER_180_353 ();
 FILLCELL_X8 FILLER_180_369 ();
 FILLCELL_X2 FILLER_180_377 ();
 FILLCELL_X1 FILLER_180_379 ();
 FILLCELL_X32 FILLER_180_1518 ();
 FILLCELL_X32 FILLER_180_1550 ();
 FILLCELL_X32 FILLER_180_1582 ();
 FILLCELL_X32 FILLER_180_1614 ();
 FILLCELL_X32 FILLER_180_1646 ();
 FILLCELL_X16 FILLER_180_1678 ();
 FILLCELL_X4 FILLER_180_1694 ();
 FILLCELL_X2 FILLER_180_1698 ();
 FILLCELL_X1 FILLER_180_1700 ();
 FILLCELL_X32 FILLER_181_1 ();
 FILLCELL_X32 FILLER_181_33 ();
 FILLCELL_X32 FILLER_181_65 ();
 FILLCELL_X32 FILLER_181_97 ();
 FILLCELL_X32 FILLER_181_129 ();
 FILLCELL_X32 FILLER_181_161 ();
 FILLCELL_X32 FILLER_181_193 ();
 FILLCELL_X32 FILLER_181_225 ();
 FILLCELL_X32 FILLER_181_257 ();
 FILLCELL_X32 FILLER_181_289 ();
 FILLCELL_X32 FILLER_181_321 ();
 FILLCELL_X16 FILLER_181_353 ();
 FILLCELL_X8 FILLER_181_369 ();
 FILLCELL_X2 FILLER_181_377 ();
 FILLCELL_X1 FILLER_181_379 ();
 FILLCELL_X32 FILLER_181_1518 ();
 FILLCELL_X32 FILLER_181_1550 ();
 FILLCELL_X32 FILLER_181_1582 ();
 FILLCELL_X32 FILLER_181_1614 ();
 FILLCELL_X32 FILLER_181_1646 ();
 FILLCELL_X16 FILLER_181_1678 ();
 FILLCELL_X4 FILLER_181_1694 ();
 FILLCELL_X2 FILLER_181_1698 ();
 FILLCELL_X1 FILLER_181_1700 ();
 FILLCELL_X4 FILLER_182_1 ();
 FILLCELL_X32 FILLER_182_12 ();
 FILLCELL_X32 FILLER_182_44 ();
 FILLCELL_X32 FILLER_182_76 ();
 FILLCELL_X32 FILLER_182_108 ();
 FILLCELL_X32 FILLER_182_140 ();
 FILLCELL_X32 FILLER_182_172 ();
 FILLCELL_X32 FILLER_182_204 ();
 FILLCELL_X32 FILLER_182_236 ();
 FILLCELL_X32 FILLER_182_268 ();
 FILLCELL_X32 FILLER_182_300 ();
 FILLCELL_X32 FILLER_182_332 ();
 FILLCELL_X16 FILLER_182_364 ();
 FILLCELL_X32 FILLER_182_1518 ();
 FILLCELL_X32 FILLER_182_1550 ();
 FILLCELL_X32 FILLER_182_1582 ();
 FILLCELL_X32 FILLER_182_1614 ();
 FILLCELL_X32 FILLER_182_1646 ();
 FILLCELL_X16 FILLER_182_1678 ();
 FILLCELL_X4 FILLER_182_1694 ();
 FILLCELL_X2 FILLER_182_1698 ();
 FILLCELL_X1 FILLER_182_1700 ();
 FILLCELL_X32 FILLER_183_1 ();
 FILLCELL_X32 FILLER_183_33 ();
 FILLCELL_X32 FILLER_183_65 ();
 FILLCELL_X32 FILLER_183_97 ();
 FILLCELL_X32 FILLER_183_129 ();
 FILLCELL_X32 FILLER_183_161 ();
 FILLCELL_X32 FILLER_183_193 ();
 FILLCELL_X32 FILLER_183_225 ();
 FILLCELL_X32 FILLER_183_257 ();
 FILLCELL_X32 FILLER_183_289 ();
 FILLCELL_X32 FILLER_183_321 ();
 FILLCELL_X16 FILLER_183_353 ();
 FILLCELL_X8 FILLER_183_369 ();
 FILLCELL_X2 FILLER_183_377 ();
 FILLCELL_X1 FILLER_183_379 ();
 FILLCELL_X32 FILLER_183_1518 ();
 FILLCELL_X32 FILLER_183_1550 ();
 FILLCELL_X32 FILLER_183_1582 ();
 FILLCELL_X32 FILLER_183_1614 ();
 FILLCELL_X32 FILLER_183_1646 ();
 FILLCELL_X16 FILLER_183_1678 ();
 FILLCELL_X4 FILLER_183_1694 ();
 FILLCELL_X2 FILLER_183_1698 ();
 FILLCELL_X1 FILLER_183_1700 ();
 FILLCELL_X32 FILLER_184_1 ();
 FILLCELL_X32 FILLER_184_33 ();
 FILLCELL_X32 FILLER_184_65 ();
 FILLCELL_X32 FILLER_184_97 ();
 FILLCELL_X32 FILLER_184_129 ();
 FILLCELL_X32 FILLER_184_161 ();
 FILLCELL_X32 FILLER_184_193 ();
 FILLCELL_X32 FILLER_184_225 ();
 FILLCELL_X32 FILLER_184_257 ();
 FILLCELL_X32 FILLER_184_289 ();
 FILLCELL_X32 FILLER_184_321 ();
 FILLCELL_X16 FILLER_184_353 ();
 FILLCELL_X8 FILLER_184_369 ();
 FILLCELL_X2 FILLER_184_377 ();
 FILLCELL_X1 FILLER_184_379 ();
 FILLCELL_X32 FILLER_184_1518 ();
 FILLCELL_X32 FILLER_184_1550 ();
 FILLCELL_X32 FILLER_184_1582 ();
 FILLCELL_X32 FILLER_184_1614 ();
 FILLCELL_X32 FILLER_184_1646 ();
 FILLCELL_X16 FILLER_184_1678 ();
 FILLCELL_X4 FILLER_184_1694 ();
 FILLCELL_X2 FILLER_184_1698 ();
 FILLCELL_X1 FILLER_184_1700 ();
 FILLCELL_X32 FILLER_185_1 ();
 FILLCELL_X32 FILLER_185_33 ();
 FILLCELL_X32 FILLER_185_65 ();
 FILLCELL_X32 FILLER_185_97 ();
 FILLCELL_X32 FILLER_185_129 ();
 FILLCELL_X32 FILLER_185_161 ();
 FILLCELL_X32 FILLER_185_193 ();
 FILLCELL_X32 FILLER_185_225 ();
 FILLCELL_X32 FILLER_185_257 ();
 FILLCELL_X32 FILLER_185_289 ();
 FILLCELL_X32 FILLER_185_321 ();
 FILLCELL_X16 FILLER_185_353 ();
 FILLCELL_X8 FILLER_185_369 ();
 FILLCELL_X2 FILLER_185_377 ();
 FILLCELL_X1 FILLER_185_379 ();
 FILLCELL_X32 FILLER_185_1518 ();
 FILLCELL_X32 FILLER_185_1550 ();
 FILLCELL_X32 FILLER_185_1582 ();
 FILLCELL_X32 FILLER_185_1614 ();
 FILLCELL_X32 FILLER_185_1646 ();
 FILLCELL_X16 FILLER_185_1678 ();
 FILLCELL_X4 FILLER_185_1694 ();
 FILLCELL_X2 FILLER_185_1698 ();
 FILLCELL_X1 FILLER_185_1700 ();
 FILLCELL_X32 FILLER_186_1 ();
 FILLCELL_X32 FILLER_186_33 ();
 FILLCELL_X32 FILLER_186_65 ();
 FILLCELL_X32 FILLER_186_97 ();
 FILLCELL_X32 FILLER_186_129 ();
 FILLCELL_X32 FILLER_186_161 ();
 FILLCELL_X32 FILLER_186_193 ();
 FILLCELL_X32 FILLER_186_225 ();
 FILLCELL_X32 FILLER_186_257 ();
 FILLCELL_X32 FILLER_186_289 ();
 FILLCELL_X32 FILLER_186_321 ();
 FILLCELL_X16 FILLER_186_353 ();
 FILLCELL_X8 FILLER_186_369 ();
 FILLCELL_X2 FILLER_186_377 ();
 FILLCELL_X1 FILLER_186_379 ();
 FILLCELL_X32 FILLER_186_1518 ();
 FILLCELL_X32 FILLER_186_1550 ();
 FILLCELL_X32 FILLER_186_1582 ();
 FILLCELL_X32 FILLER_186_1614 ();
 FILLCELL_X32 FILLER_186_1646 ();
 FILLCELL_X16 FILLER_186_1678 ();
 FILLCELL_X4 FILLER_186_1697 ();
 FILLCELL_X32 FILLER_187_1 ();
 FILLCELL_X32 FILLER_187_33 ();
 FILLCELL_X32 FILLER_187_65 ();
 FILLCELL_X32 FILLER_187_97 ();
 FILLCELL_X32 FILLER_187_129 ();
 FILLCELL_X32 FILLER_187_161 ();
 FILLCELL_X32 FILLER_187_193 ();
 FILLCELL_X32 FILLER_187_225 ();
 FILLCELL_X32 FILLER_187_257 ();
 FILLCELL_X32 FILLER_187_289 ();
 FILLCELL_X32 FILLER_187_321 ();
 FILLCELL_X16 FILLER_187_353 ();
 FILLCELL_X8 FILLER_187_369 ();
 FILLCELL_X2 FILLER_187_377 ();
 FILLCELL_X1 FILLER_187_379 ();
 FILLCELL_X32 FILLER_187_1518 ();
 FILLCELL_X32 FILLER_187_1550 ();
 FILLCELL_X32 FILLER_187_1582 ();
 FILLCELL_X32 FILLER_187_1614 ();
 FILLCELL_X32 FILLER_187_1646 ();
 FILLCELL_X16 FILLER_187_1678 ();
 FILLCELL_X4 FILLER_187_1694 ();
 FILLCELL_X2 FILLER_187_1698 ();
 FILLCELL_X1 FILLER_187_1700 ();
 FILLCELL_X32 FILLER_188_1 ();
 FILLCELL_X32 FILLER_188_33 ();
 FILLCELL_X32 FILLER_188_65 ();
 FILLCELL_X32 FILLER_188_97 ();
 FILLCELL_X32 FILLER_188_129 ();
 FILLCELL_X32 FILLER_188_161 ();
 FILLCELL_X32 FILLER_188_193 ();
 FILLCELL_X32 FILLER_188_225 ();
 FILLCELL_X32 FILLER_188_257 ();
 FILLCELL_X32 FILLER_188_289 ();
 FILLCELL_X32 FILLER_188_321 ();
 FILLCELL_X16 FILLER_188_353 ();
 FILLCELL_X8 FILLER_188_369 ();
 FILLCELL_X2 FILLER_188_377 ();
 FILLCELL_X1 FILLER_188_379 ();
 FILLCELL_X32 FILLER_188_1518 ();
 FILLCELL_X32 FILLER_188_1550 ();
 FILLCELL_X32 FILLER_188_1582 ();
 FILLCELL_X32 FILLER_188_1614 ();
 FILLCELL_X32 FILLER_188_1646 ();
 FILLCELL_X16 FILLER_188_1678 ();
 FILLCELL_X4 FILLER_188_1694 ();
 FILLCELL_X2 FILLER_188_1698 ();
 FILLCELL_X1 FILLER_188_1700 ();
 FILLCELL_X32 FILLER_189_1 ();
 FILLCELL_X32 FILLER_189_33 ();
 FILLCELL_X32 FILLER_189_65 ();
 FILLCELL_X32 FILLER_189_97 ();
 FILLCELL_X32 FILLER_189_129 ();
 FILLCELL_X32 FILLER_189_161 ();
 FILLCELL_X32 FILLER_189_193 ();
 FILLCELL_X32 FILLER_189_225 ();
 FILLCELL_X32 FILLER_189_257 ();
 FILLCELL_X32 FILLER_189_289 ();
 FILLCELL_X32 FILLER_189_321 ();
 FILLCELL_X16 FILLER_189_353 ();
 FILLCELL_X8 FILLER_189_369 ();
 FILLCELL_X2 FILLER_189_377 ();
 FILLCELL_X1 FILLER_189_379 ();
 FILLCELL_X32 FILLER_189_1518 ();
 FILLCELL_X32 FILLER_189_1550 ();
 FILLCELL_X32 FILLER_189_1582 ();
 FILLCELL_X32 FILLER_189_1614 ();
 FILLCELL_X32 FILLER_189_1646 ();
 FILLCELL_X16 FILLER_189_1678 ();
 FILLCELL_X4 FILLER_189_1694 ();
 FILLCELL_X2 FILLER_189_1698 ();
 FILLCELL_X1 FILLER_189_1700 ();
 FILLCELL_X32 FILLER_190_1 ();
 FILLCELL_X32 FILLER_190_33 ();
 FILLCELL_X32 FILLER_190_65 ();
 FILLCELL_X32 FILLER_190_97 ();
 FILLCELL_X32 FILLER_190_129 ();
 FILLCELL_X32 FILLER_190_161 ();
 FILLCELL_X32 FILLER_190_193 ();
 FILLCELL_X32 FILLER_190_225 ();
 FILLCELL_X32 FILLER_190_257 ();
 FILLCELL_X32 FILLER_190_289 ();
 FILLCELL_X32 FILLER_190_321 ();
 FILLCELL_X16 FILLER_190_353 ();
 FILLCELL_X8 FILLER_190_369 ();
 FILLCELL_X2 FILLER_190_377 ();
 FILLCELL_X1 FILLER_190_379 ();
 FILLCELL_X32 FILLER_190_1518 ();
 FILLCELL_X32 FILLER_190_1550 ();
 FILLCELL_X32 FILLER_190_1582 ();
 FILLCELL_X32 FILLER_190_1614 ();
 FILLCELL_X32 FILLER_190_1646 ();
 FILLCELL_X16 FILLER_190_1678 ();
 FILLCELL_X4 FILLER_190_1694 ();
 FILLCELL_X2 FILLER_190_1698 ();
 FILLCELL_X1 FILLER_190_1700 ();
 FILLCELL_X4 FILLER_191_1 ();
 FILLCELL_X32 FILLER_191_8 ();
 FILLCELL_X32 FILLER_191_40 ();
 FILLCELL_X32 FILLER_191_72 ();
 FILLCELL_X32 FILLER_191_104 ();
 FILLCELL_X32 FILLER_191_136 ();
 FILLCELL_X32 FILLER_191_168 ();
 FILLCELL_X32 FILLER_191_200 ();
 FILLCELL_X32 FILLER_191_232 ();
 FILLCELL_X32 FILLER_191_264 ();
 FILLCELL_X32 FILLER_191_296 ();
 FILLCELL_X32 FILLER_191_328 ();
 FILLCELL_X16 FILLER_191_360 ();
 FILLCELL_X4 FILLER_191_376 ();
 FILLCELL_X32 FILLER_191_1518 ();
 FILLCELL_X32 FILLER_191_1550 ();
 FILLCELL_X32 FILLER_191_1582 ();
 FILLCELL_X32 FILLER_191_1614 ();
 FILLCELL_X32 FILLER_191_1646 ();
 FILLCELL_X16 FILLER_191_1678 ();
 FILLCELL_X4 FILLER_191_1694 ();
 FILLCELL_X2 FILLER_191_1698 ();
 FILLCELL_X1 FILLER_191_1700 ();
 FILLCELL_X32 FILLER_192_1 ();
 FILLCELL_X32 FILLER_192_33 ();
 FILLCELL_X32 FILLER_192_65 ();
 FILLCELL_X32 FILLER_192_97 ();
 FILLCELL_X32 FILLER_192_129 ();
 FILLCELL_X32 FILLER_192_161 ();
 FILLCELL_X32 FILLER_192_193 ();
 FILLCELL_X32 FILLER_192_225 ();
 FILLCELL_X32 FILLER_192_257 ();
 FILLCELL_X32 FILLER_192_289 ();
 FILLCELL_X32 FILLER_192_321 ();
 FILLCELL_X16 FILLER_192_353 ();
 FILLCELL_X8 FILLER_192_369 ();
 FILLCELL_X2 FILLER_192_377 ();
 FILLCELL_X1 FILLER_192_379 ();
 FILLCELL_X32 FILLER_192_1518 ();
 FILLCELL_X32 FILLER_192_1550 ();
 FILLCELL_X32 FILLER_192_1582 ();
 FILLCELL_X32 FILLER_192_1614 ();
 FILLCELL_X32 FILLER_192_1646 ();
 FILLCELL_X16 FILLER_192_1678 ();
 FILLCELL_X4 FILLER_192_1694 ();
 FILLCELL_X2 FILLER_192_1698 ();
 FILLCELL_X1 FILLER_192_1700 ();
 FILLCELL_X32 FILLER_193_1 ();
 FILLCELL_X32 FILLER_193_33 ();
 FILLCELL_X32 FILLER_193_65 ();
 FILLCELL_X32 FILLER_193_97 ();
 FILLCELL_X32 FILLER_193_129 ();
 FILLCELL_X32 FILLER_193_161 ();
 FILLCELL_X32 FILLER_193_193 ();
 FILLCELL_X32 FILLER_193_225 ();
 FILLCELL_X32 FILLER_193_257 ();
 FILLCELL_X32 FILLER_193_289 ();
 FILLCELL_X32 FILLER_193_321 ();
 FILLCELL_X16 FILLER_193_353 ();
 FILLCELL_X8 FILLER_193_369 ();
 FILLCELL_X2 FILLER_193_377 ();
 FILLCELL_X1 FILLER_193_379 ();
 FILLCELL_X32 FILLER_193_1518 ();
 FILLCELL_X32 FILLER_193_1550 ();
 FILLCELL_X32 FILLER_193_1582 ();
 FILLCELL_X32 FILLER_193_1614 ();
 FILLCELL_X32 FILLER_193_1646 ();
 FILLCELL_X16 FILLER_193_1678 ();
 FILLCELL_X4 FILLER_193_1694 ();
 FILLCELL_X2 FILLER_193_1698 ();
 FILLCELL_X1 FILLER_193_1700 ();
 FILLCELL_X32 FILLER_194_1 ();
 FILLCELL_X32 FILLER_194_33 ();
 FILLCELL_X32 FILLER_194_65 ();
 FILLCELL_X32 FILLER_194_97 ();
 FILLCELL_X32 FILLER_194_129 ();
 FILLCELL_X32 FILLER_194_161 ();
 FILLCELL_X32 FILLER_194_193 ();
 FILLCELL_X32 FILLER_194_225 ();
 FILLCELL_X32 FILLER_194_257 ();
 FILLCELL_X32 FILLER_194_289 ();
 FILLCELL_X32 FILLER_194_321 ();
 FILLCELL_X16 FILLER_194_353 ();
 FILLCELL_X8 FILLER_194_369 ();
 FILLCELL_X2 FILLER_194_377 ();
 FILLCELL_X1 FILLER_194_379 ();
 FILLCELL_X32 FILLER_194_1518 ();
 FILLCELL_X32 FILLER_194_1550 ();
 FILLCELL_X32 FILLER_194_1582 ();
 FILLCELL_X32 FILLER_194_1614 ();
 FILLCELL_X32 FILLER_194_1646 ();
 FILLCELL_X16 FILLER_194_1678 ();
 FILLCELL_X4 FILLER_194_1694 ();
 FILLCELL_X2 FILLER_194_1698 ();
 FILLCELL_X1 FILLER_194_1700 ();
 FILLCELL_X32 FILLER_195_1 ();
 FILLCELL_X32 FILLER_195_33 ();
 FILLCELL_X32 FILLER_195_65 ();
 FILLCELL_X32 FILLER_195_97 ();
 FILLCELL_X32 FILLER_195_129 ();
 FILLCELL_X32 FILLER_195_161 ();
 FILLCELL_X32 FILLER_195_193 ();
 FILLCELL_X32 FILLER_195_225 ();
 FILLCELL_X32 FILLER_195_257 ();
 FILLCELL_X32 FILLER_195_289 ();
 FILLCELL_X32 FILLER_195_321 ();
 FILLCELL_X16 FILLER_195_353 ();
 FILLCELL_X8 FILLER_195_369 ();
 FILLCELL_X2 FILLER_195_377 ();
 FILLCELL_X1 FILLER_195_379 ();
 FILLCELL_X32 FILLER_195_1518 ();
 FILLCELL_X32 FILLER_195_1550 ();
 FILLCELL_X32 FILLER_195_1582 ();
 FILLCELL_X32 FILLER_195_1614 ();
 FILLCELL_X32 FILLER_195_1646 ();
 FILLCELL_X16 FILLER_195_1678 ();
 FILLCELL_X4 FILLER_195_1694 ();
 FILLCELL_X2 FILLER_195_1698 ();
 FILLCELL_X1 FILLER_195_1700 ();
 FILLCELL_X32 FILLER_196_1 ();
 FILLCELL_X32 FILLER_196_33 ();
 FILLCELL_X32 FILLER_196_65 ();
 FILLCELL_X32 FILLER_196_97 ();
 FILLCELL_X32 FILLER_196_129 ();
 FILLCELL_X32 FILLER_196_161 ();
 FILLCELL_X32 FILLER_196_193 ();
 FILLCELL_X32 FILLER_196_225 ();
 FILLCELL_X32 FILLER_196_257 ();
 FILLCELL_X32 FILLER_196_289 ();
 FILLCELL_X32 FILLER_196_321 ();
 FILLCELL_X16 FILLER_196_353 ();
 FILLCELL_X8 FILLER_196_369 ();
 FILLCELL_X2 FILLER_196_377 ();
 FILLCELL_X1 FILLER_196_379 ();
 FILLCELL_X32 FILLER_196_1518 ();
 FILLCELL_X32 FILLER_196_1550 ();
 FILLCELL_X32 FILLER_196_1582 ();
 FILLCELL_X32 FILLER_196_1614 ();
 FILLCELL_X32 FILLER_196_1646 ();
 FILLCELL_X16 FILLER_196_1678 ();
 FILLCELL_X4 FILLER_196_1697 ();
 FILLCELL_X32 FILLER_197_1 ();
 FILLCELL_X32 FILLER_197_33 ();
 FILLCELL_X32 FILLER_197_65 ();
 FILLCELL_X32 FILLER_197_97 ();
 FILLCELL_X32 FILLER_197_129 ();
 FILLCELL_X32 FILLER_197_161 ();
 FILLCELL_X32 FILLER_197_193 ();
 FILLCELL_X32 FILLER_197_225 ();
 FILLCELL_X32 FILLER_197_257 ();
 FILLCELL_X32 FILLER_197_289 ();
 FILLCELL_X32 FILLER_197_321 ();
 FILLCELL_X16 FILLER_197_353 ();
 FILLCELL_X8 FILLER_197_369 ();
 FILLCELL_X2 FILLER_197_377 ();
 FILLCELL_X1 FILLER_197_379 ();
 FILLCELL_X32 FILLER_197_1518 ();
 FILLCELL_X32 FILLER_197_1550 ();
 FILLCELL_X32 FILLER_197_1582 ();
 FILLCELL_X32 FILLER_197_1614 ();
 FILLCELL_X32 FILLER_197_1646 ();
 FILLCELL_X16 FILLER_197_1678 ();
 FILLCELL_X4 FILLER_197_1694 ();
 FILLCELL_X2 FILLER_197_1698 ();
 FILLCELL_X1 FILLER_197_1700 ();
 FILLCELL_X32 FILLER_198_1 ();
 FILLCELL_X32 FILLER_198_33 ();
 FILLCELL_X32 FILLER_198_65 ();
 FILLCELL_X32 FILLER_198_97 ();
 FILLCELL_X32 FILLER_198_129 ();
 FILLCELL_X32 FILLER_198_161 ();
 FILLCELL_X32 FILLER_198_193 ();
 FILLCELL_X32 FILLER_198_225 ();
 FILLCELL_X32 FILLER_198_257 ();
 FILLCELL_X32 FILLER_198_289 ();
 FILLCELL_X32 FILLER_198_321 ();
 FILLCELL_X16 FILLER_198_353 ();
 FILLCELL_X8 FILLER_198_369 ();
 FILLCELL_X2 FILLER_198_377 ();
 FILLCELL_X1 FILLER_198_379 ();
 FILLCELL_X32 FILLER_198_1518 ();
 FILLCELL_X32 FILLER_198_1550 ();
 FILLCELL_X32 FILLER_198_1582 ();
 FILLCELL_X32 FILLER_198_1614 ();
 FILLCELL_X32 FILLER_198_1646 ();
 FILLCELL_X16 FILLER_198_1678 ();
 FILLCELL_X4 FILLER_198_1694 ();
 FILLCELL_X2 FILLER_198_1698 ();
 FILLCELL_X1 FILLER_198_1700 ();
 FILLCELL_X32 FILLER_199_1 ();
 FILLCELL_X32 FILLER_199_33 ();
 FILLCELL_X32 FILLER_199_65 ();
 FILLCELL_X32 FILLER_199_97 ();
 FILLCELL_X32 FILLER_199_129 ();
 FILLCELL_X32 FILLER_199_161 ();
 FILLCELL_X32 FILLER_199_193 ();
 FILLCELL_X32 FILLER_199_225 ();
 FILLCELL_X32 FILLER_199_257 ();
 FILLCELL_X32 FILLER_199_289 ();
 FILLCELL_X32 FILLER_199_321 ();
 FILLCELL_X16 FILLER_199_353 ();
 FILLCELL_X8 FILLER_199_369 ();
 FILLCELL_X2 FILLER_199_377 ();
 FILLCELL_X1 FILLER_199_379 ();
 FILLCELL_X32 FILLER_199_1518 ();
 FILLCELL_X32 FILLER_199_1550 ();
 FILLCELL_X32 FILLER_199_1582 ();
 FILLCELL_X32 FILLER_199_1614 ();
 FILLCELL_X32 FILLER_199_1646 ();
 FILLCELL_X16 FILLER_199_1678 ();
 FILLCELL_X4 FILLER_199_1694 ();
 FILLCELL_X2 FILLER_199_1698 ();
 FILLCELL_X1 FILLER_199_1700 ();
 FILLCELL_X32 FILLER_200_1 ();
 FILLCELL_X32 FILLER_200_33 ();
 FILLCELL_X32 FILLER_200_65 ();
 FILLCELL_X32 FILLER_200_97 ();
 FILLCELL_X32 FILLER_200_129 ();
 FILLCELL_X32 FILLER_200_161 ();
 FILLCELL_X32 FILLER_200_193 ();
 FILLCELL_X32 FILLER_200_225 ();
 FILLCELL_X32 FILLER_200_257 ();
 FILLCELL_X32 FILLER_200_289 ();
 FILLCELL_X32 FILLER_200_321 ();
 FILLCELL_X16 FILLER_200_353 ();
 FILLCELL_X8 FILLER_200_369 ();
 FILLCELL_X2 FILLER_200_377 ();
 FILLCELL_X1 FILLER_200_379 ();
 FILLCELL_X32 FILLER_200_1518 ();
 FILLCELL_X32 FILLER_200_1550 ();
 FILLCELL_X32 FILLER_200_1582 ();
 FILLCELL_X32 FILLER_200_1614 ();
 FILLCELL_X32 FILLER_200_1646 ();
 FILLCELL_X16 FILLER_200_1678 ();
 FILLCELL_X4 FILLER_200_1694 ();
 FILLCELL_X2 FILLER_200_1698 ();
 FILLCELL_X1 FILLER_200_1700 ();
 FILLCELL_X4 FILLER_201_1 ();
 FILLCELL_X32 FILLER_201_54 ();
 FILLCELL_X32 FILLER_201_86 ();
 FILLCELL_X32 FILLER_201_118 ();
 FILLCELL_X32 FILLER_201_150 ();
 FILLCELL_X32 FILLER_201_182 ();
 FILLCELL_X32 FILLER_201_214 ();
 FILLCELL_X32 FILLER_201_246 ();
 FILLCELL_X32 FILLER_201_278 ();
 FILLCELL_X32 FILLER_201_310 ();
 FILLCELL_X32 FILLER_201_342 ();
 FILLCELL_X4 FILLER_201_374 ();
 FILLCELL_X2 FILLER_201_378 ();
 FILLCELL_X32 FILLER_201_1518 ();
 FILLCELL_X32 FILLER_201_1550 ();
 FILLCELL_X32 FILLER_201_1582 ();
 FILLCELL_X32 FILLER_201_1614 ();
 FILLCELL_X32 FILLER_201_1646 ();
 FILLCELL_X16 FILLER_201_1678 ();
 FILLCELL_X4 FILLER_201_1694 ();
 FILLCELL_X2 FILLER_201_1698 ();
 FILLCELL_X1 FILLER_201_1700 ();
 FILLCELL_X32 FILLER_202_1 ();
 FILLCELL_X32 FILLER_202_33 ();
 FILLCELL_X32 FILLER_202_65 ();
 FILLCELL_X32 FILLER_202_97 ();
 FILLCELL_X32 FILLER_202_129 ();
 FILLCELL_X32 FILLER_202_161 ();
 FILLCELL_X32 FILLER_202_193 ();
 FILLCELL_X32 FILLER_202_225 ();
 FILLCELL_X32 FILLER_202_257 ();
 FILLCELL_X32 FILLER_202_289 ();
 FILLCELL_X32 FILLER_202_321 ();
 FILLCELL_X16 FILLER_202_353 ();
 FILLCELL_X8 FILLER_202_369 ();
 FILLCELL_X2 FILLER_202_377 ();
 FILLCELL_X1 FILLER_202_379 ();
 FILLCELL_X32 FILLER_202_1518 ();
 FILLCELL_X32 FILLER_202_1550 ();
 FILLCELL_X32 FILLER_202_1582 ();
 FILLCELL_X32 FILLER_202_1614 ();
 FILLCELL_X32 FILLER_202_1646 ();
 FILLCELL_X16 FILLER_202_1678 ();
 FILLCELL_X4 FILLER_202_1694 ();
 FILLCELL_X2 FILLER_202_1698 ();
 FILLCELL_X1 FILLER_202_1700 ();
 FILLCELL_X32 FILLER_203_1 ();
 FILLCELL_X32 FILLER_203_33 ();
 FILLCELL_X32 FILLER_203_65 ();
 FILLCELL_X32 FILLER_203_97 ();
 FILLCELL_X32 FILLER_203_129 ();
 FILLCELL_X32 FILLER_203_161 ();
 FILLCELL_X32 FILLER_203_193 ();
 FILLCELL_X32 FILLER_203_225 ();
 FILLCELL_X32 FILLER_203_257 ();
 FILLCELL_X32 FILLER_203_289 ();
 FILLCELL_X32 FILLER_203_321 ();
 FILLCELL_X16 FILLER_203_353 ();
 FILLCELL_X8 FILLER_203_369 ();
 FILLCELL_X2 FILLER_203_377 ();
 FILLCELL_X1 FILLER_203_379 ();
 FILLCELL_X32 FILLER_203_1518 ();
 FILLCELL_X32 FILLER_203_1550 ();
 FILLCELL_X32 FILLER_203_1582 ();
 FILLCELL_X32 FILLER_203_1614 ();
 FILLCELL_X32 FILLER_203_1646 ();
 FILLCELL_X16 FILLER_203_1678 ();
 FILLCELL_X4 FILLER_203_1694 ();
 FILLCELL_X2 FILLER_203_1698 ();
 FILLCELL_X1 FILLER_203_1700 ();
 FILLCELL_X32 FILLER_204_1 ();
 FILLCELL_X32 FILLER_204_33 ();
 FILLCELL_X32 FILLER_204_65 ();
 FILLCELL_X32 FILLER_204_97 ();
 FILLCELL_X32 FILLER_204_129 ();
 FILLCELL_X32 FILLER_204_161 ();
 FILLCELL_X32 FILLER_204_193 ();
 FILLCELL_X32 FILLER_204_225 ();
 FILLCELL_X32 FILLER_204_257 ();
 FILLCELL_X32 FILLER_204_289 ();
 FILLCELL_X32 FILLER_204_321 ();
 FILLCELL_X16 FILLER_204_353 ();
 FILLCELL_X8 FILLER_204_369 ();
 FILLCELL_X2 FILLER_204_377 ();
 FILLCELL_X1 FILLER_204_379 ();
 FILLCELL_X32 FILLER_204_1518 ();
 FILLCELL_X32 FILLER_204_1550 ();
 FILLCELL_X32 FILLER_204_1582 ();
 FILLCELL_X32 FILLER_204_1614 ();
 FILLCELL_X32 FILLER_204_1646 ();
 FILLCELL_X16 FILLER_204_1678 ();
 FILLCELL_X4 FILLER_204_1694 ();
 FILLCELL_X2 FILLER_204_1698 ();
 FILLCELL_X1 FILLER_204_1700 ();
 FILLCELL_X32 FILLER_205_1 ();
 FILLCELL_X32 FILLER_205_33 ();
 FILLCELL_X32 FILLER_205_65 ();
 FILLCELL_X32 FILLER_205_97 ();
 FILLCELL_X32 FILLER_205_129 ();
 FILLCELL_X32 FILLER_205_161 ();
 FILLCELL_X32 FILLER_205_193 ();
 FILLCELL_X32 FILLER_205_225 ();
 FILLCELL_X32 FILLER_205_257 ();
 FILLCELL_X32 FILLER_205_289 ();
 FILLCELL_X32 FILLER_205_321 ();
 FILLCELL_X16 FILLER_205_353 ();
 FILLCELL_X8 FILLER_205_369 ();
 FILLCELL_X2 FILLER_205_377 ();
 FILLCELL_X1 FILLER_205_379 ();
 FILLCELL_X32 FILLER_205_1518 ();
 FILLCELL_X32 FILLER_205_1550 ();
 FILLCELL_X32 FILLER_205_1582 ();
 FILLCELL_X32 FILLER_205_1614 ();
 FILLCELL_X32 FILLER_205_1646 ();
 FILLCELL_X16 FILLER_205_1678 ();
 FILLCELL_X4 FILLER_205_1694 ();
 FILLCELL_X2 FILLER_205_1698 ();
 FILLCELL_X1 FILLER_205_1700 ();
 FILLCELL_X32 FILLER_206_1 ();
 FILLCELL_X32 FILLER_206_33 ();
 FILLCELL_X32 FILLER_206_65 ();
 FILLCELL_X32 FILLER_206_97 ();
 FILLCELL_X32 FILLER_206_129 ();
 FILLCELL_X32 FILLER_206_161 ();
 FILLCELL_X32 FILLER_206_193 ();
 FILLCELL_X32 FILLER_206_225 ();
 FILLCELL_X32 FILLER_206_257 ();
 FILLCELL_X32 FILLER_206_289 ();
 FILLCELL_X32 FILLER_206_321 ();
 FILLCELL_X16 FILLER_206_353 ();
 FILLCELL_X8 FILLER_206_369 ();
 FILLCELL_X2 FILLER_206_377 ();
 FILLCELL_X1 FILLER_206_379 ();
 FILLCELL_X32 FILLER_206_1518 ();
 FILLCELL_X32 FILLER_206_1550 ();
 FILLCELL_X32 FILLER_206_1582 ();
 FILLCELL_X32 FILLER_206_1614 ();
 FILLCELL_X32 FILLER_206_1646 ();
 FILLCELL_X8 FILLER_206_1678 ();
 FILLCELL_X4 FILLER_206_1686 ();
 FILLCELL_X2 FILLER_206_1690 ();
 FILLCELL_X4 FILLER_206_1697 ();
 FILLCELL_X32 FILLER_207_1 ();
 FILLCELL_X32 FILLER_207_33 ();
 FILLCELL_X32 FILLER_207_65 ();
 FILLCELL_X32 FILLER_207_97 ();
 FILLCELL_X32 FILLER_207_129 ();
 FILLCELL_X32 FILLER_207_161 ();
 FILLCELL_X32 FILLER_207_193 ();
 FILLCELL_X32 FILLER_207_225 ();
 FILLCELL_X32 FILLER_207_257 ();
 FILLCELL_X32 FILLER_207_289 ();
 FILLCELL_X32 FILLER_207_321 ();
 FILLCELL_X16 FILLER_207_353 ();
 FILLCELL_X8 FILLER_207_369 ();
 FILLCELL_X2 FILLER_207_377 ();
 FILLCELL_X1 FILLER_207_379 ();
 FILLCELL_X32 FILLER_207_1518 ();
 FILLCELL_X32 FILLER_207_1550 ();
 FILLCELL_X32 FILLER_207_1582 ();
 FILLCELL_X32 FILLER_207_1614 ();
 FILLCELL_X32 FILLER_207_1646 ();
 FILLCELL_X16 FILLER_207_1678 ();
 FILLCELL_X4 FILLER_207_1694 ();
 FILLCELL_X2 FILLER_207_1698 ();
 FILLCELL_X1 FILLER_207_1700 ();
 FILLCELL_X32 FILLER_208_1 ();
 FILLCELL_X32 FILLER_208_33 ();
 FILLCELL_X32 FILLER_208_65 ();
 FILLCELL_X32 FILLER_208_97 ();
 FILLCELL_X32 FILLER_208_129 ();
 FILLCELL_X32 FILLER_208_161 ();
 FILLCELL_X32 FILLER_208_193 ();
 FILLCELL_X32 FILLER_208_225 ();
 FILLCELL_X32 FILLER_208_257 ();
 FILLCELL_X32 FILLER_208_289 ();
 FILLCELL_X32 FILLER_208_321 ();
 FILLCELL_X32 FILLER_208_353 ();
 FILLCELL_X32 FILLER_208_385 ();
 FILLCELL_X32 FILLER_208_417 ();
 FILLCELL_X32 FILLER_208_449 ();
 FILLCELL_X32 FILLER_208_481 ();
 FILLCELL_X32 FILLER_208_513 ();
 FILLCELL_X32 FILLER_208_545 ();
 FILLCELL_X32 FILLER_208_577 ();
 FILLCELL_X16 FILLER_208_609 ();
 FILLCELL_X4 FILLER_208_625 ();
 FILLCELL_X2 FILLER_208_629 ();
 FILLCELL_X32 FILLER_208_632 ();
 FILLCELL_X32 FILLER_208_664 ();
 FILLCELL_X32 FILLER_208_696 ();
 FILLCELL_X32 FILLER_208_728 ();
 FILLCELL_X32 FILLER_208_760 ();
 FILLCELL_X32 FILLER_208_792 ();
 FILLCELL_X32 FILLER_208_824 ();
 FILLCELL_X32 FILLER_208_856 ();
 FILLCELL_X32 FILLER_208_888 ();
 FILLCELL_X32 FILLER_208_920 ();
 FILLCELL_X32 FILLER_208_952 ();
 FILLCELL_X32 FILLER_208_984 ();
 FILLCELL_X32 FILLER_208_1016 ();
 FILLCELL_X16 FILLER_208_1048 ();
 FILLCELL_X8 FILLER_208_1064 ();
 FILLCELL_X4 FILLER_208_1072 ();
 FILLCELL_X32 FILLER_208_1081 ();
 FILLCELL_X32 FILLER_208_1113 ();
 FILLCELL_X32 FILLER_208_1145 ();
 FILLCELL_X32 FILLER_208_1177 ();
 FILLCELL_X32 FILLER_208_1209 ();
 FILLCELL_X16 FILLER_208_1241 ();
 FILLCELL_X4 FILLER_208_1257 ();
 FILLCELL_X1 FILLER_208_1261 ();
 FILLCELL_X32 FILLER_208_1263 ();
 FILLCELL_X32 FILLER_208_1295 ();
 FILLCELL_X32 FILLER_208_1327 ();
 FILLCELL_X32 FILLER_208_1359 ();
 FILLCELL_X32 FILLER_208_1391 ();
 FILLCELL_X32 FILLER_208_1423 ();
 FILLCELL_X32 FILLER_208_1455 ();
 FILLCELL_X32 FILLER_208_1487 ();
 FILLCELL_X32 FILLER_208_1519 ();
 FILLCELL_X32 FILLER_208_1551 ();
 FILLCELL_X32 FILLER_208_1583 ();
 FILLCELL_X32 FILLER_208_1615 ();
 FILLCELL_X32 FILLER_208_1647 ();
 FILLCELL_X16 FILLER_208_1679 ();
 FILLCELL_X4 FILLER_208_1695 ();
 FILLCELL_X2 FILLER_208_1699 ();
 FILLCELL_X32 FILLER_209_1 ();
 FILLCELL_X32 FILLER_209_33 ();
 FILLCELL_X32 FILLER_209_65 ();
 FILLCELL_X32 FILLER_209_97 ();
 FILLCELL_X32 FILLER_209_129 ();
 FILLCELL_X32 FILLER_209_161 ();
 FILLCELL_X32 FILLER_209_193 ();
 FILLCELL_X32 FILLER_209_225 ();
 FILLCELL_X32 FILLER_209_257 ();
 FILLCELL_X32 FILLER_209_289 ();
 FILLCELL_X32 FILLER_209_321 ();
 FILLCELL_X32 FILLER_209_353 ();
 FILLCELL_X32 FILLER_209_385 ();
 FILLCELL_X32 FILLER_209_417 ();
 FILLCELL_X32 FILLER_209_449 ();
 FILLCELL_X32 FILLER_209_481 ();
 FILLCELL_X32 FILLER_209_513 ();
 FILLCELL_X32 FILLER_209_545 ();
 FILLCELL_X32 FILLER_209_577 ();
 FILLCELL_X32 FILLER_209_609 ();
 FILLCELL_X32 FILLER_209_641 ();
 FILLCELL_X32 FILLER_209_673 ();
 FILLCELL_X32 FILLER_209_705 ();
 FILLCELL_X32 FILLER_209_737 ();
 FILLCELL_X32 FILLER_209_769 ();
 FILLCELL_X32 FILLER_209_801 ();
 FILLCELL_X32 FILLER_209_833 ();
 FILLCELL_X32 FILLER_209_865 ();
 FILLCELL_X32 FILLER_209_897 ();
 FILLCELL_X32 FILLER_209_929 ();
 FILLCELL_X32 FILLER_209_961 ();
 FILLCELL_X32 FILLER_209_993 ();
 FILLCELL_X32 FILLER_209_1025 ();
 FILLCELL_X32 FILLER_209_1057 ();
 FILLCELL_X32 FILLER_209_1089 ();
 FILLCELL_X32 FILLER_209_1121 ();
 FILLCELL_X32 FILLER_209_1153 ();
 FILLCELL_X32 FILLER_209_1185 ();
 FILLCELL_X32 FILLER_209_1217 ();
 FILLCELL_X8 FILLER_209_1249 ();
 FILLCELL_X4 FILLER_209_1257 ();
 FILLCELL_X2 FILLER_209_1261 ();
 FILLCELL_X32 FILLER_209_1264 ();
 FILLCELL_X32 FILLER_209_1296 ();
 FILLCELL_X32 FILLER_209_1328 ();
 FILLCELL_X32 FILLER_209_1360 ();
 FILLCELL_X32 FILLER_209_1392 ();
 FILLCELL_X32 FILLER_209_1424 ();
 FILLCELL_X32 FILLER_209_1456 ();
 FILLCELL_X32 FILLER_209_1488 ();
 FILLCELL_X32 FILLER_209_1520 ();
 FILLCELL_X32 FILLER_209_1552 ();
 FILLCELL_X32 FILLER_209_1584 ();
 FILLCELL_X32 FILLER_209_1616 ();
 FILLCELL_X32 FILLER_209_1648 ();
 FILLCELL_X16 FILLER_209_1680 ();
 FILLCELL_X4 FILLER_209_1696 ();
 FILLCELL_X1 FILLER_209_1700 ();
 FILLCELL_X4 FILLER_210_1 ();
 FILLCELL_X32 FILLER_210_10 ();
 FILLCELL_X32 FILLER_210_42 ();
 FILLCELL_X32 FILLER_210_74 ();
 FILLCELL_X32 FILLER_210_106 ();
 FILLCELL_X32 FILLER_210_138 ();
 FILLCELL_X32 FILLER_210_170 ();
 FILLCELL_X32 FILLER_210_202 ();
 FILLCELL_X32 FILLER_210_234 ();
 FILLCELL_X32 FILLER_210_266 ();
 FILLCELL_X32 FILLER_210_298 ();
 FILLCELL_X32 FILLER_210_330 ();
 FILLCELL_X32 FILLER_210_362 ();
 FILLCELL_X32 FILLER_210_394 ();
 FILLCELL_X32 FILLER_210_426 ();
 FILLCELL_X32 FILLER_210_458 ();
 FILLCELL_X32 FILLER_210_490 ();
 FILLCELL_X32 FILLER_210_522 ();
 FILLCELL_X32 FILLER_210_554 ();
 FILLCELL_X32 FILLER_210_586 ();
 FILLCELL_X8 FILLER_210_618 ();
 FILLCELL_X4 FILLER_210_626 ();
 FILLCELL_X1 FILLER_210_630 ();
 FILLCELL_X32 FILLER_210_632 ();
 FILLCELL_X32 FILLER_210_664 ();
 FILLCELL_X32 FILLER_210_696 ();
 FILLCELL_X32 FILLER_210_728 ();
 FILLCELL_X32 FILLER_210_760 ();
 FILLCELL_X32 FILLER_210_792 ();
 FILLCELL_X32 FILLER_210_824 ();
 FILLCELL_X32 FILLER_210_856 ();
 FILLCELL_X32 FILLER_210_888 ();
 FILLCELL_X32 FILLER_210_920 ();
 FILLCELL_X32 FILLER_210_952 ();
 FILLCELL_X32 FILLER_210_984 ();
 FILLCELL_X32 FILLER_210_1016 ();
 FILLCELL_X32 FILLER_210_1048 ();
 FILLCELL_X32 FILLER_210_1080 ();
 FILLCELL_X32 FILLER_210_1112 ();
 FILLCELL_X32 FILLER_210_1144 ();
 FILLCELL_X32 FILLER_210_1176 ();
 FILLCELL_X32 FILLER_210_1208 ();
 FILLCELL_X32 FILLER_210_1240 ();
 FILLCELL_X32 FILLER_210_1272 ();
 FILLCELL_X32 FILLER_210_1304 ();
 FILLCELL_X32 FILLER_210_1336 ();
 FILLCELL_X32 FILLER_210_1368 ();
 FILLCELL_X32 FILLER_210_1400 ();
 FILLCELL_X32 FILLER_210_1432 ();
 FILLCELL_X32 FILLER_210_1464 ();
 FILLCELL_X32 FILLER_210_1496 ();
 FILLCELL_X32 FILLER_210_1528 ();
 FILLCELL_X32 FILLER_210_1560 ();
 FILLCELL_X32 FILLER_210_1592 ();
 FILLCELL_X32 FILLER_210_1624 ();
 FILLCELL_X32 FILLER_210_1656 ();
 FILLCELL_X8 FILLER_210_1688 ();
 FILLCELL_X4 FILLER_210_1696 ();
 FILLCELL_X1 FILLER_210_1700 ();
 FILLCELL_X32 FILLER_211_1 ();
 FILLCELL_X32 FILLER_211_33 ();
 FILLCELL_X32 FILLER_211_65 ();
 FILLCELL_X32 FILLER_211_97 ();
 FILLCELL_X32 FILLER_211_129 ();
 FILLCELL_X32 FILLER_211_161 ();
 FILLCELL_X32 FILLER_211_193 ();
 FILLCELL_X32 FILLER_211_225 ();
 FILLCELL_X32 FILLER_211_257 ();
 FILLCELL_X32 FILLER_211_289 ();
 FILLCELL_X32 FILLER_211_321 ();
 FILLCELL_X32 FILLER_211_353 ();
 FILLCELL_X32 FILLER_211_385 ();
 FILLCELL_X32 FILLER_211_417 ();
 FILLCELL_X32 FILLER_211_449 ();
 FILLCELL_X32 FILLER_211_481 ();
 FILLCELL_X32 FILLER_211_513 ();
 FILLCELL_X32 FILLER_211_545 ();
 FILLCELL_X32 FILLER_211_577 ();
 FILLCELL_X32 FILLER_211_609 ();
 FILLCELL_X32 FILLER_211_641 ();
 FILLCELL_X32 FILLER_211_673 ();
 FILLCELL_X32 FILLER_211_705 ();
 FILLCELL_X32 FILLER_211_737 ();
 FILLCELL_X32 FILLER_211_769 ();
 FILLCELL_X32 FILLER_211_801 ();
 FILLCELL_X32 FILLER_211_833 ();
 FILLCELL_X32 FILLER_211_865 ();
 FILLCELL_X32 FILLER_211_897 ();
 FILLCELL_X32 FILLER_211_929 ();
 FILLCELL_X32 FILLER_211_961 ();
 FILLCELL_X32 FILLER_211_993 ();
 FILLCELL_X32 FILLER_211_1025 ();
 FILLCELL_X32 FILLER_211_1057 ();
 FILLCELL_X32 FILLER_211_1089 ();
 FILLCELL_X32 FILLER_211_1121 ();
 FILLCELL_X32 FILLER_211_1153 ();
 FILLCELL_X32 FILLER_211_1185 ();
 FILLCELL_X32 FILLER_211_1217 ();
 FILLCELL_X8 FILLER_211_1249 ();
 FILLCELL_X4 FILLER_211_1257 ();
 FILLCELL_X2 FILLER_211_1261 ();
 FILLCELL_X32 FILLER_211_1264 ();
 FILLCELL_X32 FILLER_211_1296 ();
 FILLCELL_X32 FILLER_211_1328 ();
 FILLCELL_X32 FILLER_211_1360 ();
 FILLCELL_X32 FILLER_211_1392 ();
 FILLCELL_X32 FILLER_211_1424 ();
 FILLCELL_X32 FILLER_211_1456 ();
 FILLCELL_X32 FILLER_211_1488 ();
 FILLCELL_X32 FILLER_211_1520 ();
 FILLCELL_X32 FILLER_211_1552 ();
 FILLCELL_X32 FILLER_211_1584 ();
 FILLCELL_X32 FILLER_211_1616 ();
 FILLCELL_X32 FILLER_211_1648 ();
 FILLCELL_X16 FILLER_211_1680 ();
 FILLCELL_X4 FILLER_211_1696 ();
 FILLCELL_X1 FILLER_211_1700 ();
 FILLCELL_X32 FILLER_212_1 ();
 FILLCELL_X32 FILLER_212_33 ();
 FILLCELL_X32 FILLER_212_65 ();
 FILLCELL_X32 FILLER_212_97 ();
 FILLCELL_X32 FILLER_212_129 ();
 FILLCELL_X32 FILLER_212_161 ();
 FILLCELL_X32 FILLER_212_193 ();
 FILLCELL_X32 FILLER_212_225 ();
 FILLCELL_X32 FILLER_212_257 ();
 FILLCELL_X32 FILLER_212_289 ();
 FILLCELL_X32 FILLER_212_321 ();
 FILLCELL_X32 FILLER_212_353 ();
 FILLCELL_X32 FILLER_212_385 ();
 FILLCELL_X32 FILLER_212_417 ();
 FILLCELL_X32 FILLER_212_449 ();
 FILLCELL_X32 FILLER_212_481 ();
 FILLCELL_X32 FILLER_212_513 ();
 FILLCELL_X32 FILLER_212_545 ();
 FILLCELL_X32 FILLER_212_577 ();
 FILLCELL_X16 FILLER_212_609 ();
 FILLCELL_X4 FILLER_212_625 ();
 FILLCELL_X2 FILLER_212_629 ();
 FILLCELL_X32 FILLER_212_632 ();
 FILLCELL_X32 FILLER_212_664 ();
 FILLCELL_X32 FILLER_212_696 ();
 FILLCELL_X32 FILLER_212_728 ();
 FILLCELL_X32 FILLER_212_760 ();
 FILLCELL_X32 FILLER_212_792 ();
 FILLCELL_X32 FILLER_212_824 ();
 FILLCELL_X32 FILLER_212_856 ();
 FILLCELL_X32 FILLER_212_888 ();
 FILLCELL_X32 FILLER_212_920 ();
 FILLCELL_X32 FILLER_212_952 ();
 FILLCELL_X32 FILLER_212_984 ();
 FILLCELL_X32 FILLER_212_1016 ();
 FILLCELL_X32 FILLER_212_1048 ();
 FILLCELL_X32 FILLER_212_1080 ();
 FILLCELL_X32 FILLER_212_1112 ();
 FILLCELL_X32 FILLER_212_1144 ();
 FILLCELL_X32 FILLER_212_1176 ();
 FILLCELL_X32 FILLER_212_1208 ();
 FILLCELL_X32 FILLER_212_1240 ();
 FILLCELL_X32 FILLER_212_1272 ();
 FILLCELL_X32 FILLER_212_1304 ();
 FILLCELL_X32 FILLER_212_1336 ();
 FILLCELL_X32 FILLER_212_1368 ();
 FILLCELL_X32 FILLER_212_1400 ();
 FILLCELL_X32 FILLER_212_1432 ();
 FILLCELL_X32 FILLER_212_1464 ();
 FILLCELL_X32 FILLER_212_1496 ();
 FILLCELL_X32 FILLER_212_1528 ();
 FILLCELL_X32 FILLER_212_1560 ();
 FILLCELL_X32 FILLER_212_1592 ();
 FILLCELL_X32 FILLER_212_1624 ();
 FILLCELL_X32 FILLER_212_1656 ();
 FILLCELL_X8 FILLER_212_1688 ();
 FILLCELL_X4 FILLER_212_1696 ();
 FILLCELL_X1 FILLER_212_1700 ();
 FILLCELL_X32 FILLER_213_1 ();
 FILLCELL_X32 FILLER_213_33 ();
 FILLCELL_X32 FILLER_213_65 ();
 FILLCELL_X32 FILLER_213_97 ();
 FILLCELL_X32 FILLER_213_129 ();
 FILLCELL_X32 FILLER_213_161 ();
 FILLCELL_X32 FILLER_213_193 ();
 FILLCELL_X32 FILLER_213_225 ();
 FILLCELL_X32 FILLER_213_257 ();
 FILLCELL_X32 FILLER_213_289 ();
 FILLCELL_X32 FILLER_213_321 ();
 FILLCELL_X32 FILLER_213_353 ();
 FILLCELL_X32 FILLER_213_385 ();
 FILLCELL_X32 FILLER_213_417 ();
 FILLCELL_X32 FILLER_213_449 ();
 FILLCELL_X32 FILLER_213_481 ();
 FILLCELL_X32 FILLER_213_513 ();
 FILLCELL_X32 FILLER_213_545 ();
 FILLCELL_X32 FILLER_213_577 ();
 FILLCELL_X32 FILLER_213_609 ();
 FILLCELL_X32 FILLER_213_641 ();
 FILLCELL_X32 FILLER_213_673 ();
 FILLCELL_X32 FILLER_213_705 ();
 FILLCELL_X32 FILLER_213_737 ();
 FILLCELL_X32 FILLER_213_769 ();
 FILLCELL_X32 FILLER_213_801 ();
 FILLCELL_X32 FILLER_213_833 ();
 FILLCELL_X32 FILLER_213_865 ();
 FILLCELL_X32 FILLER_213_897 ();
 FILLCELL_X32 FILLER_213_929 ();
 FILLCELL_X32 FILLER_213_961 ();
 FILLCELL_X32 FILLER_213_993 ();
 FILLCELL_X32 FILLER_213_1025 ();
 FILLCELL_X32 FILLER_213_1057 ();
 FILLCELL_X32 FILLER_213_1089 ();
 FILLCELL_X32 FILLER_213_1121 ();
 FILLCELL_X32 FILLER_213_1153 ();
 FILLCELL_X32 FILLER_213_1185 ();
 FILLCELL_X32 FILLER_213_1217 ();
 FILLCELL_X8 FILLER_213_1249 ();
 FILLCELL_X4 FILLER_213_1257 ();
 FILLCELL_X2 FILLER_213_1261 ();
 FILLCELL_X32 FILLER_213_1264 ();
 FILLCELL_X32 FILLER_213_1296 ();
 FILLCELL_X32 FILLER_213_1328 ();
 FILLCELL_X32 FILLER_213_1360 ();
 FILLCELL_X32 FILLER_213_1392 ();
 FILLCELL_X32 FILLER_213_1424 ();
 FILLCELL_X32 FILLER_213_1456 ();
 FILLCELL_X32 FILLER_213_1488 ();
 FILLCELL_X32 FILLER_213_1520 ();
 FILLCELL_X32 FILLER_213_1552 ();
 FILLCELL_X32 FILLER_213_1584 ();
 FILLCELL_X32 FILLER_213_1616 ();
 FILLCELL_X32 FILLER_213_1648 ();
 FILLCELL_X16 FILLER_213_1680 ();
 FILLCELL_X4 FILLER_213_1696 ();
 FILLCELL_X1 FILLER_213_1700 ();
 FILLCELL_X32 FILLER_214_1 ();
 FILLCELL_X32 FILLER_214_33 ();
 FILLCELL_X32 FILLER_214_65 ();
 FILLCELL_X32 FILLER_214_97 ();
 FILLCELL_X32 FILLER_214_129 ();
 FILLCELL_X32 FILLER_214_161 ();
 FILLCELL_X32 FILLER_214_193 ();
 FILLCELL_X32 FILLER_214_225 ();
 FILLCELL_X32 FILLER_214_257 ();
 FILLCELL_X32 FILLER_214_289 ();
 FILLCELL_X32 FILLER_214_321 ();
 FILLCELL_X32 FILLER_214_353 ();
 FILLCELL_X32 FILLER_214_385 ();
 FILLCELL_X32 FILLER_214_417 ();
 FILLCELL_X32 FILLER_214_449 ();
 FILLCELL_X32 FILLER_214_481 ();
 FILLCELL_X32 FILLER_214_513 ();
 FILLCELL_X32 FILLER_214_545 ();
 FILLCELL_X32 FILLER_214_577 ();
 FILLCELL_X16 FILLER_214_609 ();
 FILLCELL_X4 FILLER_214_625 ();
 FILLCELL_X2 FILLER_214_629 ();
 FILLCELL_X32 FILLER_214_632 ();
 FILLCELL_X32 FILLER_214_664 ();
 FILLCELL_X32 FILLER_214_696 ();
 FILLCELL_X32 FILLER_214_728 ();
 FILLCELL_X32 FILLER_214_760 ();
 FILLCELL_X32 FILLER_214_792 ();
 FILLCELL_X32 FILLER_214_824 ();
 FILLCELL_X32 FILLER_214_856 ();
 FILLCELL_X32 FILLER_214_888 ();
 FILLCELL_X32 FILLER_214_920 ();
 FILLCELL_X32 FILLER_214_952 ();
 FILLCELL_X32 FILLER_214_984 ();
 FILLCELL_X32 FILLER_214_1016 ();
 FILLCELL_X32 FILLER_214_1048 ();
 FILLCELL_X32 FILLER_214_1080 ();
 FILLCELL_X32 FILLER_214_1112 ();
 FILLCELL_X32 FILLER_214_1144 ();
 FILLCELL_X32 FILLER_214_1176 ();
 FILLCELL_X32 FILLER_214_1208 ();
 FILLCELL_X32 FILLER_214_1240 ();
 FILLCELL_X32 FILLER_214_1272 ();
 FILLCELL_X32 FILLER_214_1304 ();
 FILLCELL_X32 FILLER_214_1336 ();
 FILLCELL_X32 FILLER_214_1368 ();
 FILLCELL_X32 FILLER_214_1400 ();
 FILLCELL_X32 FILLER_214_1432 ();
 FILLCELL_X32 FILLER_214_1464 ();
 FILLCELL_X32 FILLER_214_1496 ();
 FILLCELL_X32 FILLER_214_1528 ();
 FILLCELL_X32 FILLER_214_1560 ();
 FILLCELL_X32 FILLER_214_1592 ();
 FILLCELL_X32 FILLER_214_1624 ();
 FILLCELL_X32 FILLER_214_1656 ();
 FILLCELL_X4 FILLER_214_1688 ();
 FILLCELL_X4 FILLER_214_1697 ();
 FILLCELL_X32 FILLER_215_1 ();
 FILLCELL_X32 FILLER_215_33 ();
 FILLCELL_X32 FILLER_215_65 ();
 FILLCELL_X32 FILLER_215_97 ();
 FILLCELL_X32 FILLER_215_129 ();
 FILLCELL_X32 FILLER_215_161 ();
 FILLCELL_X32 FILLER_215_193 ();
 FILLCELL_X32 FILLER_215_225 ();
 FILLCELL_X32 FILLER_215_257 ();
 FILLCELL_X32 FILLER_215_289 ();
 FILLCELL_X32 FILLER_215_321 ();
 FILLCELL_X32 FILLER_215_353 ();
 FILLCELL_X32 FILLER_215_385 ();
 FILLCELL_X32 FILLER_215_417 ();
 FILLCELL_X32 FILLER_215_449 ();
 FILLCELL_X32 FILLER_215_481 ();
 FILLCELL_X32 FILLER_215_513 ();
 FILLCELL_X32 FILLER_215_545 ();
 FILLCELL_X32 FILLER_215_577 ();
 FILLCELL_X32 FILLER_215_609 ();
 FILLCELL_X32 FILLER_215_641 ();
 FILLCELL_X32 FILLER_215_673 ();
 FILLCELL_X32 FILLER_215_705 ();
 FILLCELL_X32 FILLER_215_737 ();
 FILLCELL_X32 FILLER_215_769 ();
 FILLCELL_X32 FILLER_215_801 ();
 FILLCELL_X32 FILLER_215_833 ();
 FILLCELL_X32 FILLER_215_865 ();
 FILLCELL_X32 FILLER_215_897 ();
 FILLCELL_X32 FILLER_215_929 ();
 FILLCELL_X32 FILLER_215_961 ();
 FILLCELL_X32 FILLER_215_993 ();
 FILLCELL_X32 FILLER_215_1025 ();
 FILLCELL_X32 FILLER_215_1057 ();
 FILLCELL_X32 FILLER_215_1089 ();
 FILLCELL_X32 FILLER_215_1121 ();
 FILLCELL_X32 FILLER_215_1153 ();
 FILLCELL_X32 FILLER_215_1185 ();
 FILLCELL_X32 FILLER_215_1217 ();
 FILLCELL_X8 FILLER_215_1249 ();
 FILLCELL_X4 FILLER_215_1257 ();
 FILLCELL_X2 FILLER_215_1261 ();
 FILLCELL_X32 FILLER_215_1264 ();
 FILLCELL_X32 FILLER_215_1296 ();
 FILLCELL_X32 FILLER_215_1328 ();
 FILLCELL_X32 FILLER_215_1360 ();
 FILLCELL_X32 FILLER_215_1392 ();
 FILLCELL_X32 FILLER_215_1424 ();
 FILLCELL_X32 FILLER_215_1456 ();
 FILLCELL_X32 FILLER_215_1488 ();
 FILLCELL_X32 FILLER_215_1520 ();
 FILLCELL_X32 FILLER_215_1552 ();
 FILLCELL_X32 FILLER_215_1584 ();
 FILLCELL_X32 FILLER_215_1616 ();
 FILLCELL_X32 FILLER_215_1648 ();
 FILLCELL_X16 FILLER_215_1680 ();
 FILLCELL_X4 FILLER_215_1696 ();
 FILLCELL_X1 FILLER_215_1700 ();
 FILLCELL_X32 FILLER_216_1 ();
 FILLCELL_X32 FILLER_216_33 ();
 FILLCELL_X32 FILLER_216_65 ();
 FILLCELL_X32 FILLER_216_97 ();
 FILLCELL_X32 FILLER_216_129 ();
 FILLCELL_X32 FILLER_216_161 ();
 FILLCELL_X32 FILLER_216_193 ();
 FILLCELL_X32 FILLER_216_225 ();
 FILLCELL_X32 FILLER_216_257 ();
 FILLCELL_X32 FILLER_216_289 ();
 FILLCELL_X32 FILLER_216_321 ();
 FILLCELL_X32 FILLER_216_353 ();
 FILLCELL_X32 FILLER_216_385 ();
 FILLCELL_X32 FILLER_216_417 ();
 FILLCELL_X32 FILLER_216_449 ();
 FILLCELL_X32 FILLER_216_481 ();
 FILLCELL_X32 FILLER_216_513 ();
 FILLCELL_X32 FILLER_216_545 ();
 FILLCELL_X32 FILLER_216_577 ();
 FILLCELL_X16 FILLER_216_609 ();
 FILLCELL_X4 FILLER_216_625 ();
 FILLCELL_X2 FILLER_216_629 ();
 FILLCELL_X32 FILLER_216_632 ();
 FILLCELL_X32 FILLER_216_664 ();
 FILLCELL_X32 FILLER_216_696 ();
 FILLCELL_X32 FILLER_216_728 ();
 FILLCELL_X32 FILLER_216_760 ();
 FILLCELL_X32 FILLER_216_792 ();
 FILLCELL_X32 FILLER_216_824 ();
 FILLCELL_X32 FILLER_216_856 ();
 FILLCELL_X32 FILLER_216_888 ();
 FILLCELL_X32 FILLER_216_920 ();
 FILLCELL_X32 FILLER_216_952 ();
 FILLCELL_X32 FILLER_216_984 ();
 FILLCELL_X32 FILLER_216_1016 ();
 FILLCELL_X32 FILLER_216_1048 ();
 FILLCELL_X32 FILLER_216_1080 ();
 FILLCELL_X32 FILLER_216_1112 ();
 FILLCELL_X32 FILLER_216_1144 ();
 FILLCELL_X32 FILLER_216_1176 ();
 FILLCELL_X32 FILLER_216_1208 ();
 FILLCELL_X32 FILLER_216_1240 ();
 FILLCELL_X32 FILLER_216_1272 ();
 FILLCELL_X32 FILLER_216_1304 ();
 FILLCELL_X32 FILLER_216_1336 ();
 FILLCELL_X32 FILLER_216_1368 ();
 FILLCELL_X32 FILLER_216_1400 ();
 FILLCELL_X32 FILLER_216_1432 ();
 FILLCELL_X32 FILLER_216_1464 ();
 FILLCELL_X32 FILLER_216_1496 ();
 FILLCELL_X32 FILLER_216_1528 ();
 FILLCELL_X32 FILLER_216_1560 ();
 FILLCELL_X32 FILLER_216_1592 ();
 FILLCELL_X32 FILLER_216_1624 ();
 FILLCELL_X32 FILLER_216_1656 ();
 FILLCELL_X8 FILLER_216_1688 ();
 FILLCELL_X4 FILLER_216_1696 ();
 FILLCELL_X1 FILLER_216_1700 ();
 FILLCELL_X32 FILLER_217_1 ();
 FILLCELL_X32 FILLER_217_33 ();
 FILLCELL_X32 FILLER_217_65 ();
 FILLCELL_X32 FILLER_217_97 ();
 FILLCELL_X32 FILLER_217_129 ();
 FILLCELL_X32 FILLER_217_161 ();
 FILLCELL_X32 FILLER_217_193 ();
 FILLCELL_X32 FILLER_217_225 ();
 FILLCELL_X32 FILLER_217_257 ();
 FILLCELL_X32 FILLER_217_289 ();
 FILLCELL_X32 FILLER_217_321 ();
 FILLCELL_X32 FILLER_217_353 ();
 FILLCELL_X32 FILLER_217_385 ();
 FILLCELL_X32 FILLER_217_417 ();
 FILLCELL_X32 FILLER_217_449 ();
 FILLCELL_X32 FILLER_217_481 ();
 FILLCELL_X32 FILLER_217_513 ();
 FILLCELL_X32 FILLER_217_545 ();
 FILLCELL_X32 FILLER_217_577 ();
 FILLCELL_X32 FILLER_217_609 ();
 FILLCELL_X32 FILLER_217_641 ();
 FILLCELL_X32 FILLER_217_673 ();
 FILLCELL_X32 FILLER_217_705 ();
 FILLCELL_X32 FILLER_217_737 ();
 FILLCELL_X32 FILLER_217_769 ();
 FILLCELL_X32 FILLER_217_801 ();
 FILLCELL_X32 FILLER_217_833 ();
 FILLCELL_X32 FILLER_217_865 ();
 FILLCELL_X32 FILLER_217_897 ();
 FILLCELL_X32 FILLER_217_929 ();
 FILLCELL_X32 FILLER_217_961 ();
 FILLCELL_X32 FILLER_217_993 ();
 FILLCELL_X32 FILLER_217_1025 ();
 FILLCELL_X32 FILLER_217_1057 ();
 FILLCELL_X32 FILLER_217_1089 ();
 FILLCELL_X32 FILLER_217_1121 ();
 FILLCELL_X32 FILLER_217_1153 ();
 FILLCELL_X32 FILLER_217_1185 ();
 FILLCELL_X32 FILLER_217_1217 ();
 FILLCELL_X8 FILLER_217_1249 ();
 FILLCELL_X4 FILLER_217_1257 ();
 FILLCELL_X2 FILLER_217_1261 ();
 FILLCELL_X32 FILLER_217_1264 ();
 FILLCELL_X32 FILLER_217_1296 ();
 FILLCELL_X32 FILLER_217_1328 ();
 FILLCELL_X32 FILLER_217_1360 ();
 FILLCELL_X32 FILLER_217_1392 ();
 FILLCELL_X32 FILLER_217_1424 ();
 FILLCELL_X32 FILLER_217_1456 ();
 FILLCELL_X32 FILLER_217_1488 ();
 FILLCELL_X32 FILLER_217_1520 ();
 FILLCELL_X32 FILLER_217_1552 ();
 FILLCELL_X32 FILLER_217_1584 ();
 FILLCELL_X32 FILLER_217_1616 ();
 FILLCELL_X32 FILLER_217_1648 ();
 FILLCELL_X16 FILLER_217_1680 ();
 FILLCELL_X4 FILLER_217_1696 ();
 FILLCELL_X1 FILLER_217_1700 ();
 FILLCELL_X32 FILLER_218_1 ();
 FILLCELL_X32 FILLER_218_33 ();
 FILLCELL_X32 FILLER_218_65 ();
 FILLCELL_X32 FILLER_218_97 ();
 FILLCELL_X32 FILLER_218_129 ();
 FILLCELL_X32 FILLER_218_161 ();
 FILLCELL_X32 FILLER_218_193 ();
 FILLCELL_X32 FILLER_218_225 ();
 FILLCELL_X32 FILLER_218_257 ();
 FILLCELL_X32 FILLER_218_289 ();
 FILLCELL_X32 FILLER_218_321 ();
 FILLCELL_X32 FILLER_218_353 ();
 FILLCELL_X32 FILLER_218_385 ();
 FILLCELL_X32 FILLER_218_417 ();
 FILLCELL_X32 FILLER_218_449 ();
 FILLCELL_X32 FILLER_218_481 ();
 FILLCELL_X32 FILLER_218_513 ();
 FILLCELL_X32 FILLER_218_545 ();
 FILLCELL_X32 FILLER_218_577 ();
 FILLCELL_X16 FILLER_218_609 ();
 FILLCELL_X4 FILLER_218_625 ();
 FILLCELL_X2 FILLER_218_629 ();
 FILLCELL_X32 FILLER_218_632 ();
 FILLCELL_X32 FILLER_218_664 ();
 FILLCELL_X32 FILLER_218_696 ();
 FILLCELL_X32 FILLER_218_728 ();
 FILLCELL_X32 FILLER_218_760 ();
 FILLCELL_X32 FILLER_218_792 ();
 FILLCELL_X32 FILLER_218_824 ();
 FILLCELL_X32 FILLER_218_856 ();
 FILLCELL_X32 FILLER_218_888 ();
 FILLCELL_X32 FILLER_218_920 ();
 FILLCELL_X32 FILLER_218_952 ();
 FILLCELL_X32 FILLER_218_984 ();
 FILLCELL_X32 FILLER_218_1016 ();
 FILLCELL_X32 FILLER_218_1048 ();
 FILLCELL_X32 FILLER_218_1080 ();
 FILLCELL_X32 FILLER_218_1112 ();
 FILLCELL_X32 FILLER_218_1144 ();
 FILLCELL_X32 FILLER_218_1176 ();
 FILLCELL_X32 FILLER_218_1208 ();
 FILLCELL_X32 FILLER_218_1240 ();
 FILLCELL_X32 FILLER_218_1272 ();
 FILLCELL_X32 FILLER_218_1304 ();
 FILLCELL_X32 FILLER_218_1336 ();
 FILLCELL_X32 FILLER_218_1368 ();
 FILLCELL_X32 FILLER_218_1400 ();
 FILLCELL_X32 FILLER_218_1432 ();
 FILLCELL_X32 FILLER_218_1464 ();
 FILLCELL_X32 FILLER_218_1496 ();
 FILLCELL_X32 FILLER_218_1528 ();
 FILLCELL_X32 FILLER_218_1560 ();
 FILLCELL_X32 FILLER_218_1592 ();
 FILLCELL_X32 FILLER_218_1624 ();
 FILLCELL_X32 FILLER_218_1656 ();
 FILLCELL_X8 FILLER_218_1688 ();
 FILLCELL_X4 FILLER_218_1696 ();
 FILLCELL_X1 FILLER_218_1700 ();
 FILLCELL_X4 FILLER_219_1 ();
 FILLCELL_X32 FILLER_219_12 ();
 FILLCELL_X32 FILLER_219_44 ();
 FILLCELL_X32 FILLER_219_76 ();
 FILLCELL_X32 FILLER_219_108 ();
 FILLCELL_X32 FILLER_219_140 ();
 FILLCELL_X32 FILLER_219_172 ();
 FILLCELL_X32 FILLER_219_204 ();
 FILLCELL_X32 FILLER_219_236 ();
 FILLCELL_X32 FILLER_219_268 ();
 FILLCELL_X32 FILLER_219_300 ();
 FILLCELL_X32 FILLER_219_332 ();
 FILLCELL_X32 FILLER_219_364 ();
 FILLCELL_X32 FILLER_219_396 ();
 FILLCELL_X32 FILLER_219_428 ();
 FILLCELL_X32 FILLER_219_460 ();
 FILLCELL_X32 FILLER_219_492 ();
 FILLCELL_X32 FILLER_219_524 ();
 FILLCELL_X32 FILLER_219_556 ();
 FILLCELL_X32 FILLER_219_588 ();
 FILLCELL_X32 FILLER_219_620 ();
 FILLCELL_X32 FILLER_219_652 ();
 FILLCELL_X32 FILLER_219_684 ();
 FILLCELL_X32 FILLER_219_716 ();
 FILLCELL_X32 FILLER_219_748 ();
 FILLCELL_X32 FILLER_219_780 ();
 FILLCELL_X32 FILLER_219_812 ();
 FILLCELL_X32 FILLER_219_844 ();
 FILLCELL_X32 FILLER_219_876 ();
 FILLCELL_X32 FILLER_219_908 ();
 FILLCELL_X32 FILLER_219_940 ();
 FILLCELL_X32 FILLER_219_972 ();
 FILLCELL_X32 FILLER_219_1004 ();
 FILLCELL_X32 FILLER_219_1036 ();
 FILLCELL_X32 FILLER_219_1068 ();
 FILLCELL_X32 FILLER_219_1100 ();
 FILLCELL_X32 FILLER_219_1132 ();
 FILLCELL_X32 FILLER_219_1164 ();
 FILLCELL_X32 FILLER_219_1196 ();
 FILLCELL_X32 FILLER_219_1228 ();
 FILLCELL_X2 FILLER_219_1260 ();
 FILLCELL_X1 FILLER_219_1262 ();
 FILLCELL_X32 FILLER_219_1264 ();
 FILLCELL_X32 FILLER_219_1296 ();
 FILLCELL_X32 FILLER_219_1328 ();
 FILLCELL_X32 FILLER_219_1360 ();
 FILLCELL_X32 FILLER_219_1392 ();
 FILLCELL_X32 FILLER_219_1424 ();
 FILLCELL_X32 FILLER_219_1456 ();
 FILLCELL_X32 FILLER_219_1488 ();
 FILLCELL_X32 FILLER_219_1520 ();
 FILLCELL_X32 FILLER_219_1552 ();
 FILLCELL_X32 FILLER_219_1584 ();
 FILLCELL_X32 FILLER_219_1616 ();
 FILLCELL_X32 FILLER_219_1648 ();
 FILLCELL_X16 FILLER_219_1680 ();
 FILLCELL_X4 FILLER_219_1696 ();
 FILLCELL_X1 FILLER_219_1700 ();
 FILLCELL_X32 FILLER_220_1 ();
 FILLCELL_X32 FILLER_220_33 ();
 FILLCELL_X32 FILLER_220_65 ();
 FILLCELL_X32 FILLER_220_97 ();
 FILLCELL_X32 FILLER_220_129 ();
 FILLCELL_X32 FILLER_220_161 ();
 FILLCELL_X32 FILLER_220_193 ();
 FILLCELL_X32 FILLER_220_225 ();
 FILLCELL_X32 FILLER_220_257 ();
 FILLCELL_X32 FILLER_220_289 ();
 FILLCELL_X32 FILLER_220_321 ();
 FILLCELL_X32 FILLER_220_353 ();
 FILLCELL_X32 FILLER_220_385 ();
 FILLCELL_X32 FILLER_220_417 ();
 FILLCELL_X32 FILLER_220_449 ();
 FILLCELL_X32 FILLER_220_481 ();
 FILLCELL_X32 FILLER_220_513 ();
 FILLCELL_X32 FILLER_220_545 ();
 FILLCELL_X32 FILLER_220_577 ();
 FILLCELL_X16 FILLER_220_609 ();
 FILLCELL_X4 FILLER_220_625 ();
 FILLCELL_X2 FILLER_220_629 ();
 FILLCELL_X32 FILLER_220_632 ();
 FILLCELL_X32 FILLER_220_664 ();
 FILLCELL_X32 FILLER_220_696 ();
 FILLCELL_X32 FILLER_220_728 ();
 FILLCELL_X32 FILLER_220_760 ();
 FILLCELL_X32 FILLER_220_792 ();
 FILLCELL_X32 FILLER_220_824 ();
 FILLCELL_X32 FILLER_220_856 ();
 FILLCELL_X32 FILLER_220_888 ();
 FILLCELL_X32 FILLER_220_920 ();
 FILLCELL_X32 FILLER_220_952 ();
 FILLCELL_X32 FILLER_220_984 ();
 FILLCELL_X32 FILLER_220_1016 ();
 FILLCELL_X32 FILLER_220_1048 ();
 FILLCELL_X32 FILLER_220_1080 ();
 FILLCELL_X32 FILLER_220_1112 ();
 FILLCELL_X32 FILLER_220_1144 ();
 FILLCELL_X32 FILLER_220_1176 ();
 FILLCELL_X32 FILLER_220_1208 ();
 FILLCELL_X32 FILLER_220_1240 ();
 FILLCELL_X32 FILLER_220_1272 ();
 FILLCELL_X32 FILLER_220_1304 ();
 FILLCELL_X32 FILLER_220_1336 ();
 FILLCELL_X32 FILLER_220_1368 ();
 FILLCELL_X32 FILLER_220_1400 ();
 FILLCELL_X32 FILLER_220_1432 ();
 FILLCELL_X32 FILLER_220_1464 ();
 FILLCELL_X32 FILLER_220_1496 ();
 FILLCELL_X32 FILLER_220_1528 ();
 FILLCELL_X32 FILLER_220_1560 ();
 FILLCELL_X32 FILLER_220_1592 ();
 FILLCELL_X32 FILLER_220_1624 ();
 FILLCELL_X32 FILLER_220_1656 ();
 FILLCELL_X8 FILLER_220_1688 ();
 FILLCELL_X4 FILLER_220_1696 ();
 FILLCELL_X1 FILLER_220_1700 ();
 FILLCELL_X32 FILLER_221_1 ();
 FILLCELL_X32 FILLER_221_33 ();
 FILLCELL_X32 FILLER_221_65 ();
 FILLCELL_X32 FILLER_221_97 ();
 FILLCELL_X32 FILLER_221_129 ();
 FILLCELL_X32 FILLER_221_161 ();
 FILLCELL_X32 FILLER_221_193 ();
 FILLCELL_X32 FILLER_221_225 ();
 FILLCELL_X32 FILLER_221_257 ();
 FILLCELL_X32 FILLER_221_289 ();
 FILLCELL_X32 FILLER_221_321 ();
 FILLCELL_X32 FILLER_221_353 ();
 FILLCELL_X32 FILLER_221_385 ();
 FILLCELL_X32 FILLER_221_417 ();
 FILLCELL_X32 FILLER_221_449 ();
 FILLCELL_X32 FILLER_221_481 ();
 FILLCELL_X32 FILLER_221_513 ();
 FILLCELL_X32 FILLER_221_545 ();
 FILLCELL_X32 FILLER_221_577 ();
 FILLCELL_X32 FILLER_221_609 ();
 FILLCELL_X32 FILLER_221_641 ();
 FILLCELL_X32 FILLER_221_673 ();
 FILLCELL_X32 FILLER_221_705 ();
 FILLCELL_X32 FILLER_221_737 ();
 FILLCELL_X32 FILLER_221_769 ();
 FILLCELL_X32 FILLER_221_801 ();
 FILLCELL_X32 FILLER_221_833 ();
 FILLCELL_X32 FILLER_221_865 ();
 FILLCELL_X32 FILLER_221_897 ();
 FILLCELL_X32 FILLER_221_929 ();
 FILLCELL_X32 FILLER_221_961 ();
 FILLCELL_X32 FILLER_221_993 ();
 FILLCELL_X32 FILLER_221_1025 ();
 FILLCELL_X32 FILLER_221_1057 ();
 FILLCELL_X32 FILLER_221_1089 ();
 FILLCELL_X32 FILLER_221_1121 ();
 FILLCELL_X32 FILLER_221_1153 ();
 FILLCELL_X32 FILLER_221_1185 ();
 FILLCELL_X32 FILLER_221_1217 ();
 FILLCELL_X8 FILLER_221_1249 ();
 FILLCELL_X4 FILLER_221_1257 ();
 FILLCELL_X2 FILLER_221_1261 ();
 FILLCELL_X32 FILLER_221_1264 ();
 FILLCELL_X32 FILLER_221_1296 ();
 FILLCELL_X32 FILLER_221_1328 ();
 FILLCELL_X32 FILLER_221_1360 ();
 FILLCELL_X32 FILLER_221_1392 ();
 FILLCELL_X32 FILLER_221_1424 ();
 FILLCELL_X32 FILLER_221_1456 ();
 FILLCELL_X32 FILLER_221_1488 ();
 FILLCELL_X32 FILLER_221_1520 ();
 FILLCELL_X32 FILLER_221_1552 ();
 FILLCELL_X32 FILLER_221_1584 ();
 FILLCELL_X32 FILLER_221_1616 ();
 FILLCELL_X32 FILLER_221_1648 ();
 FILLCELL_X16 FILLER_221_1680 ();
 FILLCELL_X4 FILLER_221_1696 ();
 FILLCELL_X1 FILLER_221_1700 ();
 FILLCELL_X32 FILLER_222_1 ();
 FILLCELL_X32 FILLER_222_33 ();
 FILLCELL_X32 FILLER_222_65 ();
 FILLCELL_X32 FILLER_222_97 ();
 FILLCELL_X32 FILLER_222_129 ();
 FILLCELL_X32 FILLER_222_161 ();
 FILLCELL_X32 FILLER_222_193 ();
 FILLCELL_X32 FILLER_222_225 ();
 FILLCELL_X32 FILLER_222_257 ();
 FILLCELL_X32 FILLER_222_289 ();
 FILLCELL_X32 FILLER_222_321 ();
 FILLCELL_X32 FILLER_222_353 ();
 FILLCELL_X32 FILLER_222_385 ();
 FILLCELL_X32 FILLER_222_417 ();
 FILLCELL_X32 FILLER_222_449 ();
 FILLCELL_X32 FILLER_222_481 ();
 FILLCELL_X32 FILLER_222_513 ();
 FILLCELL_X32 FILLER_222_545 ();
 FILLCELL_X32 FILLER_222_577 ();
 FILLCELL_X16 FILLER_222_609 ();
 FILLCELL_X4 FILLER_222_625 ();
 FILLCELL_X2 FILLER_222_629 ();
 FILLCELL_X32 FILLER_222_632 ();
 FILLCELL_X32 FILLER_222_664 ();
 FILLCELL_X32 FILLER_222_696 ();
 FILLCELL_X32 FILLER_222_728 ();
 FILLCELL_X32 FILLER_222_760 ();
 FILLCELL_X32 FILLER_222_792 ();
 FILLCELL_X32 FILLER_222_824 ();
 FILLCELL_X32 FILLER_222_856 ();
 FILLCELL_X32 FILLER_222_888 ();
 FILLCELL_X32 FILLER_222_920 ();
 FILLCELL_X32 FILLER_222_952 ();
 FILLCELL_X32 FILLER_222_984 ();
 FILLCELL_X32 FILLER_222_1016 ();
 FILLCELL_X32 FILLER_222_1048 ();
 FILLCELL_X32 FILLER_222_1080 ();
 FILLCELL_X32 FILLER_222_1112 ();
 FILLCELL_X32 FILLER_222_1144 ();
 FILLCELL_X32 FILLER_222_1176 ();
 FILLCELL_X32 FILLER_222_1208 ();
 FILLCELL_X32 FILLER_222_1240 ();
 FILLCELL_X32 FILLER_222_1272 ();
 FILLCELL_X32 FILLER_222_1304 ();
 FILLCELL_X32 FILLER_222_1336 ();
 FILLCELL_X32 FILLER_222_1368 ();
 FILLCELL_X32 FILLER_222_1400 ();
 FILLCELL_X32 FILLER_222_1432 ();
 FILLCELL_X32 FILLER_222_1464 ();
 FILLCELL_X32 FILLER_222_1496 ();
 FILLCELL_X32 FILLER_222_1528 ();
 FILLCELL_X32 FILLER_222_1560 ();
 FILLCELL_X32 FILLER_222_1592 ();
 FILLCELL_X32 FILLER_222_1624 ();
 FILLCELL_X32 FILLER_222_1656 ();
 FILLCELL_X8 FILLER_222_1688 ();
 FILLCELL_X4 FILLER_222_1696 ();
 FILLCELL_X1 FILLER_222_1700 ();
 FILLCELL_X32 FILLER_223_1 ();
 FILLCELL_X32 FILLER_223_33 ();
 FILLCELL_X32 FILLER_223_65 ();
 FILLCELL_X32 FILLER_223_97 ();
 FILLCELL_X32 FILLER_223_129 ();
 FILLCELL_X32 FILLER_223_161 ();
 FILLCELL_X32 FILLER_223_193 ();
 FILLCELL_X32 FILLER_223_225 ();
 FILLCELL_X32 FILLER_223_257 ();
 FILLCELL_X32 FILLER_223_289 ();
 FILLCELL_X32 FILLER_223_321 ();
 FILLCELL_X32 FILLER_223_353 ();
 FILLCELL_X32 FILLER_223_385 ();
 FILLCELL_X32 FILLER_223_417 ();
 FILLCELL_X32 FILLER_223_449 ();
 FILLCELL_X32 FILLER_223_481 ();
 FILLCELL_X32 FILLER_223_513 ();
 FILLCELL_X32 FILLER_223_545 ();
 FILLCELL_X32 FILLER_223_577 ();
 FILLCELL_X32 FILLER_223_609 ();
 FILLCELL_X32 FILLER_223_641 ();
 FILLCELL_X32 FILLER_223_673 ();
 FILLCELL_X32 FILLER_223_705 ();
 FILLCELL_X32 FILLER_223_737 ();
 FILLCELL_X32 FILLER_223_769 ();
 FILLCELL_X32 FILLER_223_801 ();
 FILLCELL_X32 FILLER_223_833 ();
 FILLCELL_X32 FILLER_223_865 ();
 FILLCELL_X32 FILLER_223_897 ();
 FILLCELL_X32 FILLER_223_929 ();
 FILLCELL_X32 FILLER_223_961 ();
 FILLCELL_X32 FILLER_223_993 ();
 FILLCELL_X32 FILLER_223_1025 ();
 FILLCELL_X32 FILLER_223_1057 ();
 FILLCELL_X32 FILLER_223_1089 ();
 FILLCELL_X32 FILLER_223_1121 ();
 FILLCELL_X32 FILLER_223_1153 ();
 FILLCELL_X32 FILLER_223_1185 ();
 FILLCELL_X32 FILLER_223_1217 ();
 FILLCELL_X8 FILLER_223_1249 ();
 FILLCELL_X4 FILLER_223_1257 ();
 FILLCELL_X2 FILLER_223_1261 ();
 FILLCELL_X32 FILLER_223_1264 ();
 FILLCELL_X32 FILLER_223_1296 ();
 FILLCELL_X32 FILLER_223_1328 ();
 FILLCELL_X32 FILLER_223_1360 ();
 FILLCELL_X32 FILLER_223_1392 ();
 FILLCELL_X32 FILLER_223_1424 ();
 FILLCELL_X32 FILLER_223_1456 ();
 FILLCELL_X32 FILLER_223_1488 ();
 FILLCELL_X32 FILLER_223_1520 ();
 FILLCELL_X32 FILLER_223_1552 ();
 FILLCELL_X32 FILLER_223_1584 ();
 FILLCELL_X32 FILLER_223_1616 ();
 FILLCELL_X32 FILLER_223_1648 ();
 FILLCELL_X16 FILLER_223_1680 ();
 FILLCELL_X4 FILLER_223_1696 ();
 FILLCELL_X1 FILLER_223_1700 ();
 FILLCELL_X32 FILLER_224_1 ();
 FILLCELL_X32 FILLER_224_33 ();
 FILLCELL_X32 FILLER_224_65 ();
 FILLCELL_X32 FILLER_224_97 ();
 FILLCELL_X32 FILLER_224_129 ();
 FILLCELL_X32 FILLER_224_161 ();
 FILLCELL_X32 FILLER_224_193 ();
 FILLCELL_X32 FILLER_224_225 ();
 FILLCELL_X32 FILLER_224_257 ();
 FILLCELL_X32 FILLER_224_289 ();
 FILLCELL_X32 FILLER_224_321 ();
 FILLCELL_X32 FILLER_224_353 ();
 FILLCELL_X32 FILLER_224_385 ();
 FILLCELL_X32 FILLER_224_417 ();
 FILLCELL_X32 FILLER_224_449 ();
 FILLCELL_X32 FILLER_224_481 ();
 FILLCELL_X32 FILLER_224_513 ();
 FILLCELL_X32 FILLER_224_545 ();
 FILLCELL_X32 FILLER_224_577 ();
 FILLCELL_X16 FILLER_224_609 ();
 FILLCELL_X4 FILLER_224_625 ();
 FILLCELL_X2 FILLER_224_629 ();
 FILLCELL_X32 FILLER_224_632 ();
 FILLCELL_X32 FILLER_224_664 ();
 FILLCELL_X32 FILLER_224_696 ();
 FILLCELL_X32 FILLER_224_728 ();
 FILLCELL_X32 FILLER_224_760 ();
 FILLCELL_X32 FILLER_224_792 ();
 FILLCELL_X32 FILLER_224_824 ();
 FILLCELL_X32 FILLER_224_856 ();
 FILLCELL_X32 FILLER_224_888 ();
 FILLCELL_X32 FILLER_224_920 ();
 FILLCELL_X32 FILLER_224_952 ();
 FILLCELL_X32 FILLER_224_984 ();
 FILLCELL_X32 FILLER_224_1016 ();
 FILLCELL_X32 FILLER_224_1048 ();
 FILLCELL_X32 FILLER_224_1080 ();
 FILLCELL_X32 FILLER_224_1112 ();
 FILLCELL_X32 FILLER_224_1144 ();
 FILLCELL_X32 FILLER_224_1176 ();
 FILLCELL_X32 FILLER_224_1208 ();
 FILLCELL_X32 FILLER_224_1240 ();
 FILLCELL_X32 FILLER_224_1272 ();
 FILLCELL_X32 FILLER_224_1304 ();
 FILLCELL_X32 FILLER_224_1336 ();
 FILLCELL_X32 FILLER_224_1368 ();
 FILLCELL_X32 FILLER_224_1400 ();
 FILLCELL_X32 FILLER_224_1432 ();
 FILLCELL_X32 FILLER_224_1464 ();
 FILLCELL_X32 FILLER_224_1496 ();
 FILLCELL_X32 FILLER_224_1528 ();
 FILLCELL_X32 FILLER_224_1560 ();
 FILLCELL_X32 FILLER_224_1592 ();
 FILLCELL_X32 FILLER_224_1624 ();
 FILLCELL_X32 FILLER_224_1656 ();
 FILLCELL_X2 FILLER_224_1688 ();
 FILLCELL_X4 FILLER_224_1697 ();
 FILLCELL_X32 FILLER_225_1 ();
 FILLCELL_X32 FILLER_225_33 ();
 FILLCELL_X32 FILLER_225_65 ();
 FILLCELL_X32 FILLER_225_97 ();
 FILLCELL_X32 FILLER_225_129 ();
 FILLCELL_X32 FILLER_225_161 ();
 FILLCELL_X32 FILLER_225_193 ();
 FILLCELL_X32 FILLER_225_225 ();
 FILLCELL_X32 FILLER_225_257 ();
 FILLCELL_X32 FILLER_225_289 ();
 FILLCELL_X32 FILLER_225_321 ();
 FILLCELL_X32 FILLER_225_353 ();
 FILLCELL_X32 FILLER_225_385 ();
 FILLCELL_X32 FILLER_225_417 ();
 FILLCELL_X32 FILLER_225_449 ();
 FILLCELL_X32 FILLER_225_481 ();
 FILLCELL_X32 FILLER_225_513 ();
 FILLCELL_X32 FILLER_225_545 ();
 FILLCELL_X32 FILLER_225_577 ();
 FILLCELL_X32 FILLER_225_609 ();
 FILLCELL_X32 FILLER_225_641 ();
 FILLCELL_X32 FILLER_225_673 ();
 FILLCELL_X32 FILLER_225_705 ();
 FILLCELL_X32 FILLER_225_737 ();
 FILLCELL_X32 FILLER_225_769 ();
 FILLCELL_X32 FILLER_225_801 ();
 FILLCELL_X32 FILLER_225_833 ();
 FILLCELL_X32 FILLER_225_865 ();
 FILLCELL_X32 FILLER_225_897 ();
 FILLCELL_X32 FILLER_225_929 ();
 FILLCELL_X32 FILLER_225_961 ();
 FILLCELL_X32 FILLER_225_993 ();
 FILLCELL_X32 FILLER_225_1025 ();
 FILLCELL_X32 FILLER_225_1057 ();
 FILLCELL_X32 FILLER_225_1089 ();
 FILLCELL_X32 FILLER_225_1121 ();
 FILLCELL_X32 FILLER_225_1153 ();
 FILLCELL_X32 FILLER_225_1185 ();
 FILLCELL_X32 FILLER_225_1217 ();
 FILLCELL_X8 FILLER_225_1249 ();
 FILLCELL_X4 FILLER_225_1257 ();
 FILLCELL_X2 FILLER_225_1261 ();
 FILLCELL_X32 FILLER_225_1264 ();
 FILLCELL_X32 FILLER_225_1296 ();
 FILLCELL_X32 FILLER_225_1328 ();
 FILLCELL_X32 FILLER_225_1360 ();
 FILLCELL_X32 FILLER_225_1392 ();
 FILLCELL_X32 FILLER_225_1424 ();
 FILLCELL_X32 FILLER_225_1456 ();
 FILLCELL_X32 FILLER_225_1488 ();
 FILLCELL_X32 FILLER_225_1520 ();
 FILLCELL_X32 FILLER_225_1552 ();
 FILLCELL_X32 FILLER_225_1584 ();
 FILLCELL_X32 FILLER_225_1616 ();
 FILLCELL_X32 FILLER_225_1648 ();
 FILLCELL_X16 FILLER_225_1680 ();
 FILLCELL_X4 FILLER_225_1696 ();
 FILLCELL_X1 FILLER_225_1700 ();
 FILLCELL_X32 FILLER_226_1 ();
 FILLCELL_X32 FILLER_226_33 ();
 FILLCELL_X32 FILLER_226_65 ();
 FILLCELL_X32 FILLER_226_97 ();
 FILLCELL_X32 FILLER_226_129 ();
 FILLCELL_X32 FILLER_226_161 ();
 FILLCELL_X32 FILLER_226_193 ();
 FILLCELL_X32 FILLER_226_225 ();
 FILLCELL_X32 FILLER_226_257 ();
 FILLCELL_X32 FILLER_226_289 ();
 FILLCELL_X32 FILLER_226_321 ();
 FILLCELL_X32 FILLER_226_353 ();
 FILLCELL_X32 FILLER_226_385 ();
 FILLCELL_X32 FILLER_226_417 ();
 FILLCELL_X32 FILLER_226_449 ();
 FILLCELL_X32 FILLER_226_481 ();
 FILLCELL_X32 FILLER_226_513 ();
 FILLCELL_X32 FILLER_226_545 ();
 FILLCELL_X32 FILLER_226_577 ();
 FILLCELL_X16 FILLER_226_609 ();
 FILLCELL_X4 FILLER_226_625 ();
 FILLCELL_X2 FILLER_226_629 ();
 FILLCELL_X32 FILLER_226_632 ();
 FILLCELL_X32 FILLER_226_664 ();
 FILLCELL_X32 FILLER_226_696 ();
 FILLCELL_X32 FILLER_226_728 ();
 FILLCELL_X32 FILLER_226_760 ();
 FILLCELL_X32 FILLER_226_792 ();
 FILLCELL_X32 FILLER_226_824 ();
 FILLCELL_X32 FILLER_226_856 ();
 FILLCELL_X32 FILLER_226_888 ();
 FILLCELL_X32 FILLER_226_920 ();
 FILLCELL_X32 FILLER_226_952 ();
 FILLCELL_X32 FILLER_226_984 ();
 FILLCELL_X32 FILLER_226_1016 ();
 FILLCELL_X32 FILLER_226_1048 ();
 FILLCELL_X32 FILLER_226_1080 ();
 FILLCELL_X32 FILLER_226_1112 ();
 FILLCELL_X32 FILLER_226_1144 ();
 FILLCELL_X32 FILLER_226_1176 ();
 FILLCELL_X32 FILLER_226_1208 ();
 FILLCELL_X32 FILLER_226_1240 ();
 FILLCELL_X32 FILLER_226_1272 ();
 FILLCELL_X32 FILLER_226_1304 ();
 FILLCELL_X32 FILLER_226_1336 ();
 FILLCELL_X32 FILLER_226_1368 ();
 FILLCELL_X32 FILLER_226_1400 ();
 FILLCELL_X32 FILLER_226_1432 ();
 FILLCELL_X32 FILLER_226_1464 ();
 FILLCELL_X32 FILLER_226_1496 ();
 FILLCELL_X32 FILLER_226_1528 ();
 FILLCELL_X32 FILLER_226_1560 ();
 FILLCELL_X32 FILLER_226_1592 ();
 FILLCELL_X32 FILLER_226_1624 ();
 FILLCELL_X32 FILLER_226_1656 ();
 FILLCELL_X8 FILLER_226_1688 ();
 FILLCELL_X4 FILLER_226_1696 ();
 FILLCELL_X1 FILLER_226_1700 ();
 FILLCELL_X32 FILLER_227_1 ();
 FILLCELL_X32 FILLER_227_33 ();
 FILLCELL_X32 FILLER_227_65 ();
 FILLCELL_X32 FILLER_227_97 ();
 FILLCELL_X32 FILLER_227_129 ();
 FILLCELL_X32 FILLER_227_161 ();
 FILLCELL_X32 FILLER_227_193 ();
 FILLCELL_X32 FILLER_227_225 ();
 FILLCELL_X32 FILLER_227_257 ();
 FILLCELL_X32 FILLER_227_289 ();
 FILLCELL_X32 FILLER_227_321 ();
 FILLCELL_X32 FILLER_227_353 ();
 FILLCELL_X32 FILLER_227_385 ();
 FILLCELL_X32 FILLER_227_417 ();
 FILLCELL_X32 FILLER_227_449 ();
 FILLCELL_X32 FILLER_227_481 ();
 FILLCELL_X32 FILLER_227_513 ();
 FILLCELL_X32 FILLER_227_545 ();
 FILLCELL_X32 FILLER_227_577 ();
 FILLCELL_X32 FILLER_227_609 ();
 FILLCELL_X32 FILLER_227_641 ();
 FILLCELL_X32 FILLER_227_673 ();
 FILLCELL_X32 FILLER_227_705 ();
 FILLCELL_X32 FILLER_227_737 ();
 FILLCELL_X32 FILLER_227_769 ();
 FILLCELL_X32 FILLER_227_801 ();
 FILLCELL_X32 FILLER_227_833 ();
 FILLCELL_X32 FILLER_227_865 ();
 FILLCELL_X32 FILLER_227_897 ();
 FILLCELL_X32 FILLER_227_929 ();
 FILLCELL_X32 FILLER_227_961 ();
 FILLCELL_X32 FILLER_227_993 ();
 FILLCELL_X32 FILLER_227_1025 ();
 FILLCELL_X32 FILLER_227_1057 ();
 FILLCELL_X32 FILLER_227_1089 ();
 FILLCELL_X32 FILLER_227_1121 ();
 FILLCELL_X32 FILLER_227_1153 ();
 FILLCELL_X32 FILLER_227_1185 ();
 FILLCELL_X32 FILLER_227_1217 ();
 FILLCELL_X8 FILLER_227_1249 ();
 FILLCELL_X4 FILLER_227_1257 ();
 FILLCELL_X2 FILLER_227_1261 ();
 FILLCELL_X32 FILLER_227_1264 ();
 FILLCELL_X32 FILLER_227_1296 ();
 FILLCELL_X32 FILLER_227_1328 ();
 FILLCELL_X32 FILLER_227_1360 ();
 FILLCELL_X32 FILLER_227_1392 ();
 FILLCELL_X32 FILLER_227_1424 ();
 FILLCELL_X32 FILLER_227_1456 ();
 FILLCELL_X32 FILLER_227_1488 ();
 FILLCELL_X32 FILLER_227_1520 ();
 FILLCELL_X32 FILLER_227_1552 ();
 FILLCELL_X32 FILLER_227_1584 ();
 FILLCELL_X32 FILLER_227_1616 ();
 FILLCELL_X32 FILLER_227_1648 ();
 FILLCELL_X16 FILLER_227_1680 ();
 FILLCELL_X4 FILLER_227_1696 ();
 FILLCELL_X1 FILLER_227_1700 ();
 FILLCELL_X4 FILLER_228_1 ();
 FILLCELL_X32 FILLER_228_8 ();
 FILLCELL_X32 FILLER_228_40 ();
 FILLCELL_X32 FILLER_228_72 ();
 FILLCELL_X32 FILLER_228_104 ();
 FILLCELL_X32 FILLER_228_136 ();
 FILLCELL_X32 FILLER_228_168 ();
 FILLCELL_X32 FILLER_228_200 ();
 FILLCELL_X32 FILLER_228_232 ();
 FILLCELL_X32 FILLER_228_264 ();
 FILLCELL_X32 FILLER_228_296 ();
 FILLCELL_X32 FILLER_228_328 ();
 FILLCELL_X32 FILLER_228_360 ();
 FILLCELL_X32 FILLER_228_392 ();
 FILLCELL_X32 FILLER_228_424 ();
 FILLCELL_X32 FILLER_228_456 ();
 FILLCELL_X32 FILLER_228_488 ();
 FILLCELL_X32 FILLER_228_520 ();
 FILLCELL_X32 FILLER_228_552 ();
 FILLCELL_X32 FILLER_228_584 ();
 FILLCELL_X8 FILLER_228_616 ();
 FILLCELL_X4 FILLER_228_624 ();
 FILLCELL_X2 FILLER_228_628 ();
 FILLCELL_X1 FILLER_228_630 ();
 FILLCELL_X32 FILLER_228_632 ();
 FILLCELL_X32 FILLER_228_664 ();
 FILLCELL_X32 FILLER_228_696 ();
 FILLCELL_X32 FILLER_228_728 ();
 FILLCELL_X32 FILLER_228_760 ();
 FILLCELL_X32 FILLER_228_792 ();
 FILLCELL_X32 FILLER_228_824 ();
 FILLCELL_X32 FILLER_228_856 ();
 FILLCELL_X32 FILLER_228_888 ();
 FILLCELL_X32 FILLER_228_920 ();
 FILLCELL_X32 FILLER_228_952 ();
 FILLCELL_X32 FILLER_228_984 ();
 FILLCELL_X32 FILLER_228_1016 ();
 FILLCELL_X32 FILLER_228_1048 ();
 FILLCELL_X32 FILLER_228_1080 ();
 FILLCELL_X32 FILLER_228_1112 ();
 FILLCELL_X32 FILLER_228_1144 ();
 FILLCELL_X32 FILLER_228_1176 ();
 FILLCELL_X32 FILLER_228_1208 ();
 FILLCELL_X32 FILLER_228_1240 ();
 FILLCELL_X32 FILLER_228_1272 ();
 FILLCELL_X32 FILLER_228_1304 ();
 FILLCELL_X32 FILLER_228_1336 ();
 FILLCELL_X32 FILLER_228_1368 ();
 FILLCELL_X32 FILLER_228_1400 ();
 FILLCELL_X32 FILLER_228_1432 ();
 FILLCELL_X32 FILLER_228_1464 ();
 FILLCELL_X32 FILLER_228_1496 ();
 FILLCELL_X32 FILLER_228_1528 ();
 FILLCELL_X32 FILLER_228_1560 ();
 FILLCELL_X32 FILLER_228_1592 ();
 FILLCELL_X32 FILLER_228_1624 ();
 FILLCELL_X32 FILLER_228_1656 ();
 FILLCELL_X8 FILLER_228_1688 ();
 FILLCELL_X4 FILLER_228_1696 ();
 FILLCELL_X1 FILLER_228_1700 ();
 FILLCELL_X8 FILLER_229_1 ();
 FILLCELL_X32 FILLER_229_12 ();
 FILLCELL_X32 FILLER_229_44 ();
 FILLCELL_X4 FILLER_229_76 ();
 FILLCELL_X32 FILLER_229_83 ();
 FILLCELL_X32 FILLER_229_115 ();
 FILLCELL_X2 FILLER_229_147 ();
 FILLCELL_X1 FILLER_229_149 ();
 FILLCELL_X32 FILLER_229_153 ();
 FILLCELL_X16 FILLER_229_185 ();
 FILLCELL_X8 FILLER_229_201 ();
 FILLCELL_X4 FILLER_229_209 ();
 FILLCELL_X2 FILLER_229_213 ();
 FILLCELL_X32 FILLER_229_218 ();
 FILLCELL_X32 FILLER_229_250 ();
 FILLCELL_X4 FILLER_229_282 ();
 FILLCELL_X32 FILLER_229_289 ();
 FILLCELL_X16 FILLER_229_321 ();
 FILLCELL_X8 FILLER_229_337 ();
 FILLCELL_X4 FILLER_229_345 ();
 FILLCELL_X2 FILLER_229_349 ();
 FILLCELL_X32 FILLER_229_354 ();
 FILLCELL_X32 FILLER_229_386 ();
 FILLCELL_X4 FILLER_229_418 ();
 FILLCELL_X32 FILLER_229_425 ();
 FILLCELL_X32 FILLER_229_457 ();
 FILLCELL_X2 FILLER_229_489 ();
 FILLCELL_X1 FILLER_229_491 ();
 FILLCELL_X32 FILLER_229_495 ();
 FILLCELL_X16 FILLER_229_527 ();
 FILLCELL_X8 FILLER_229_543 ();
 FILLCELL_X4 FILLER_229_551 ();
 FILLCELL_X2 FILLER_229_555 ();
 FILLCELL_X32 FILLER_229_564 ();
 FILLCELL_X32 FILLER_229_596 ();
 FILLCELL_X2 FILLER_229_628 ();
 FILLCELL_X1 FILLER_229_630 ();
 FILLCELL_X4 FILLER_229_632 ();
 FILLCELL_X32 FILLER_229_643 ();
 FILLCELL_X16 FILLER_229_675 ();
 FILLCELL_X2 FILLER_229_691 ();
 FILLCELL_X32 FILLER_229_696 ();
 FILLCELL_X32 FILLER_229_728 ();
 FILLCELL_X2 FILLER_229_760 ();
 FILLCELL_X1 FILLER_229_762 ();
 FILLCELL_X32 FILLER_229_770 ();
 FILLCELL_X32 FILLER_229_802 ();
 FILLCELL_X32 FILLER_229_837 ();
 FILLCELL_X16 FILLER_229_869 ();
 FILLCELL_X8 FILLER_229_885 ();
 FILLCELL_X4 FILLER_229_893 ();
 FILLCELL_X2 FILLER_229_897 ();
 FILLCELL_X32 FILLER_229_902 ();
 FILLCELL_X32 FILLER_229_934 ();
 FILLCELL_X4 FILLER_229_966 ();
 FILLCELL_X32 FILLER_229_977 ();
 FILLCELL_X16 FILLER_229_1009 ();
 FILLCELL_X8 FILLER_229_1025 ();
 FILLCELL_X2 FILLER_229_1033 ();
 FILLCELL_X32 FILLER_229_1042 ();
 FILLCELL_X16 FILLER_229_1074 ();
 FILLCELL_X8 FILLER_229_1090 ();
 FILLCELL_X4 FILLER_229_1098 ();
 FILLCELL_X2 FILLER_229_1102 ();
 FILLCELL_X1 FILLER_229_1104 ();
 FILLCELL_X32 FILLER_229_1108 ();
 FILLCELL_X32 FILLER_229_1140 ();
 FILLCELL_X4 FILLER_229_1172 ();
 FILLCELL_X32 FILLER_229_1179 ();
 FILLCELL_X16 FILLER_229_1211 ();
 FILLCELL_X8 FILLER_229_1227 ();
 FILLCELL_X4 FILLER_229_1235 ();
 FILLCELL_X2 FILLER_229_1239 ();
 FILLCELL_X16 FILLER_229_1244 ();
 FILLCELL_X2 FILLER_229_1260 ();
 FILLCELL_X32 FILLER_229_1263 ();
 FILLCELL_X16 FILLER_229_1295 ();
 FILLCELL_X1 FILLER_229_1311 ();
 FILLCELL_X32 FILLER_229_1315 ();
 FILLCELL_X16 FILLER_229_1347 ();
 FILLCELL_X8 FILLER_229_1363 ();
 FILLCELL_X4 FILLER_229_1371 ();
 FILLCELL_X1 FILLER_229_1375 ();
 FILLCELL_X32 FILLER_229_1379 ();
 FILLCELL_X32 FILLER_229_1411 ();
 FILLCELL_X4 FILLER_229_1443 ();
 FILLCELL_X32 FILLER_229_1450 ();
 FILLCELL_X32 FILLER_229_1482 ();
 FILLCELL_X4 FILLER_229_1514 ();
 FILLCELL_X32 FILLER_229_1521 ();
 FILLCELL_X16 FILLER_229_1553 ();
 FILLCELL_X8 FILLER_229_1569 ();
 FILLCELL_X4 FILLER_229_1577 ();
 FILLCELL_X2 FILLER_229_1581 ();
 FILLCELL_X32 FILLER_229_1586 ();
 FILLCELL_X32 FILLER_229_1618 ();
 FILLCELL_X4 FILLER_229_1650 ();
 FILLCELL_X32 FILLER_229_1661 ();
 FILLCELL_X1 FILLER_229_1693 ();
 FILLCELL_X4 FILLER_229_1697 ();
 assign init_done = curr_state[1];
 assign valid_out = valid_reg_out;
endmodule
