module sram_multiplier_system (clk,
    init_done,
    init_enable,
    pe_ce,
    rst_n,
    valid_out,
    data_in,
    data_out);
 input clk;
 output init_done;
 input init_enable;
 input pe_ce;
 input rst_n;
 output valid_out;
 input [7:0] data_in;
 output [15:0] data_out;

 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire u_multiplier_pp_0 ;
 wire u_multiplier_pp_14 ;
 wire net46;
 wire u_multiplier_STAGE1__016_ ;
 wire u_multiplier_STAGE1__017_ ;
 wire u_multiplier_STAGE1__018_ ;
 wire u_multiplier_STAGE1__019_ ;
 wire u_multiplier_STAGE1__020_ ;
 wire u_multiplier_STAGE1__021_ ;
 wire u_multiplier_STAGE1__022_ ;
 wire u_multiplier_STAGE1__023_ ;
 wire u_multiplier_STAGE1__024_ ;
 wire u_multiplier_STAGE1__025_ ;
 wire u_multiplier_STAGE1__026_ ;
 wire u_multiplier_STAGE1__027_ ;
 wire u_multiplier_STAGE1__028_ ;
 wire u_multiplier_STAGE1__029_ ;
 wire u_multiplier_STAGE1__030_ ;
 wire u_multiplier_STAGE1__031_ ;
 wire u_multiplier_STAGE1__032_ ;
 wire u_multiplier_STAGE1__033_ ;
 wire u_multiplier_STAGE1__034_ ;
 wire u_multiplier_STAGE1__035_ ;
 wire u_multiplier_STAGE1__036_ ;
 wire u_multiplier_STAGE1__037_ ;
 wire u_multiplier_STAGE1__038_ ;
 wire u_multiplier_STAGE1__039_ ;
 wire u_multiplier_STAGE1__040_ ;
 wire u_multiplier_STAGE1__041_ ;
 wire u_multiplier_STAGE1__042_ ;
 wire u_multiplier_STAGE1__043_ ;
 wire u_multiplier_STAGE1__044_ ;
 wire u_multiplier_STAGE1__045_ ;
 wire u_multiplier_STAGE1__046_ ;
 wire u_multiplier_STAGE1__047_ ;
 wire u_multiplier_STAGE1__048_ ;
 wire u_multiplier_STAGE1__049_ ;
 wire u_multiplier_STAGE1__050_ ;
 wire u_multiplier_STAGE1__051_ ;
 wire u_multiplier_STAGE1__052_ ;
 wire u_multiplier_STAGE1__053_ ;
 wire u_multiplier_STAGE1__054_ ;
 wire u_multiplier_STAGE1_pp_10_c2 ;
 wire u_multiplier_STAGE1_pp_5_c2 ;
 wire u_multiplier_STAGE1_pp_6_c2 ;
 wire u_multiplier_STAGE1_pp_7_c2 ;
 wire u_multiplier_STAGE1_pp_7_c4 ;
 wire u_multiplier_STAGE1_pp_8_c2 ;
 wire u_multiplier_STAGE1_pp_8_c4 ;
 wire u_multiplier_STAGE1_pp_9_c2 ;
 wire net52;
 wire u_multiplier_STAGE1_E_4_2_pp_10__08_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_10__09_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_10__10_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_10__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_10__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_10__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_10__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_5__08_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_5__09_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_5__10_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_5__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_5__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_5__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_5__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_6__08_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_6__09_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_6__10_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_6__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_6__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_6__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_6__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_7_1__08_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_7_1__09_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_7_1__10_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_7_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_7_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_7_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_7_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_7_2__08_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_7_2__09_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_7_2__10_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_7_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_7_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_7_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_7_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_8_1__08_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_8_1__09_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_8_1__10_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_8_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_8_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_8_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_8_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_8_2__08_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_8_2__09_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_8_2__10_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_8_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_8_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_8_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_8_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_9_1__08_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_9_1__09_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_9_1__10_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_9_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_9_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_9_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_9_1__14_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_11__05_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_11__06_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_11__07_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_11__08_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_9__05_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_9__06_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_9__07_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_9__08_ ;
 wire u_multiplier_STAGE2_pp_10_c1 ;
 wire u_multiplier_STAGE2_pp_10_c2 ;
 wire u_multiplier_STAGE2_pp_10_s ;
 wire u_multiplier_STAGE2_pp_11_c1 ;
 wire u_multiplier_STAGE2_pp_11_c2 ;
 wire u_multiplier_STAGE2_pp_11_s ;
 wire u_multiplier_STAGE2_pp_12_c1 ;
 wire u_multiplier_STAGE2_pp_12_c2 ;
 wire u_multiplier_STAGE2_pp_12_s ;
 wire u_multiplier_STAGE2_pp_13_c ;
 wire u_multiplier_STAGE2_pp_13_s ;
 wire u_multiplier_STAGE2_pp_2_c ;
 wire u_multiplier_STAGE2_pp_2_s ;
 wire u_multiplier_STAGE2_pp_3_c1 ;
 wire u_multiplier_STAGE2_pp_3_c2 ;
 wire u_multiplier_STAGE2_pp_3_s ;
 wire u_multiplier_STAGE2_pp_4_c1 ;
 wire u_multiplier_STAGE2_pp_4_c2 ;
 wire u_multiplier_STAGE2_pp_4_s ;
 wire u_multiplier_STAGE2_pp_5_c1 ;
 wire u_multiplier_STAGE2_pp_5_c2 ;
 wire u_multiplier_STAGE2_pp_5_s ;
 wire u_multiplier_STAGE2_pp_6_c1 ;
 wire u_multiplier_STAGE2_pp_6_c2 ;
 wire u_multiplier_STAGE2_pp_6_s ;
 wire u_multiplier_STAGE2_pp_7_c1 ;
 wire u_multiplier_STAGE2_pp_7_c2 ;
 wire u_multiplier_STAGE2_pp_7_s ;
 wire u_multiplier_STAGE2_pp_8_c1 ;
 wire u_multiplier_STAGE2_pp_8_c2 ;
 wire u_multiplier_STAGE2_pp_8_s ;
 wire u_multiplier_STAGE2_pp_9_c1 ;
 wire u_multiplier_STAGE2_pp_9_c2 ;
 wire u_multiplier_STAGE2_pp_9_s ;
 wire net65;
 wire u_multiplier_STAGE2_E_4_2_pp_10__08_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_10__09_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_10__10_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_10__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_10__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_10__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_10__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_11__08_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_11__09_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_11__10_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_11__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_11__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_11__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_11__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_12__08_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_12__09_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_12__10_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_12__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_12__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_12__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_12__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_3__08_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_3__09_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_3__10_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_4__08_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_4__09_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_4__10_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_5__08_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_5__09_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_5__10_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_5__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_5__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_5__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_5__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_6__08_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_6__09_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_6__10_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_6__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_6__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_6__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_6__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_7__08_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_7__09_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_7__10_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_7__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_7__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_7__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_7__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_8__08_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_8__09_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_8__10_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_8__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_8__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_8__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_8__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_9__08_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_9__09_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_9__10_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_9__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_9__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_9__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp_9__14_ ;
 wire u_multiplier_STAGE2_Final_add_Cout ;
 wire u_multiplier_STAGE2_Final_add_c1 ;
 wire u_multiplier_STAGE2_Final_add_c2 ;
 wire u_multiplier_STAGE2_Final_add_c3 ;
 wire u_multiplier_STAGE2_Final_add_cla1__14_ ;
 wire u_multiplier_STAGE2_Final_add_cla1__15_ ;
 wire u_multiplier_STAGE2_Final_add_cla1__16_ ;
 wire u_multiplier_STAGE2_Final_add_cla1__17_ ;
 wire u_multiplier_STAGE2_Final_add_cla1__18_ ;
 wire u_multiplier_STAGE2_Final_add_cla1__19_ ;
 wire u_multiplier_STAGE2_Final_add_cla1__20_ ;
 wire u_multiplier_STAGE2_Final_add_cla1__21_ ;
 wire u_multiplier_STAGE2_Final_add_cla1__22_ ;
 wire u_multiplier_STAGE2_Final_add_cla1__23_ ;
 wire u_multiplier_STAGE2_Final_add_cla1__24_ ;
 wire u_multiplier_STAGE2_Final_add_cla1__25_ ;
 wire u_multiplier_STAGE2_Final_add_cla1__26_ ;
 wire u_multiplier_STAGE2_Final_add_cla1__27_ ;
 wire u_multiplier_STAGE2_Final_add_cla1__28_ ;
 wire u_multiplier_STAGE2_Final_add_cla2__14_ ;
 wire u_multiplier_STAGE2_Final_add_cla2__15_ ;
 wire u_multiplier_STAGE2_Final_add_cla2__16_ ;
 wire u_multiplier_STAGE2_Final_add_cla2__17_ ;
 wire u_multiplier_STAGE2_Final_add_cla2__18_ ;
 wire u_multiplier_STAGE2_Final_add_cla2__19_ ;
 wire u_multiplier_STAGE2_Final_add_cla2__20_ ;
 wire u_multiplier_STAGE2_Final_add_cla2__21_ ;
 wire u_multiplier_STAGE2_Final_add_cla2__22_ ;
 wire u_multiplier_STAGE2_Final_add_cla2__23_ ;
 wire u_multiplier_STAGE2_Final_add_cla2__24_ ;
 wire u_multiplier_STAGE2_Final_add_cla2__25_ ;
 wire u_multiplier_STAGE2_Final_add_cla2__26_ ;
 wire u_multiplier_STAGE2_Final_add_cla2__27_ ;
 wire u_multiplier_STAGE2_Final_add_cla2__28_ ;
 wire u_multiplier_STAGE2_Final_add_cla3__14_ ;
 wire u_multiplier_STAGE2_Final_add_cla3__15_ ;
 wire u_multiplier_STAGE2_Final_add_cla3__16_ ;
 wire u_multiplier_STAGE2_Final_add_cla3__17_ ;
 wire u_multiplier_STAGE2_Final_add_cla3__18_ ;
 wire u_multiplier_STAGE2_Final_add_cla3__19_ ;
 wire u_multiplier_STAGE2_Final_add_cla3__20_ ;
 wire u_multiplier_STAGE2_Final_add_cla3__21_ ;
 wire u_multiplier_STAGE2_Final_add_cla3__22_ ;
 wire u_multiplier_STAGE2_Final_add_cla3__23_ ;
 wire u_multiplier_STAGE2_Final_add_cla3__24_ ;
 wire u_multiplier_STAGE2_Final_add_cla3__25_ ;
 wire u_multiplier_STAGE2_Final_add_cla3__26_ ;
 wire u_multiplier_STAGE2_Final_add_cla3__27_ ;
 wire u_multiplier_STAGE2_Final_add_cla3__28_ ;
 wire u_multiplier_STAGE2_Final_add_cla4__14_ ;
 wire u_multiplier_STAGE2_Final_add_cla4__15_ ;
 wire u_multiplier_STAGE2_Final_add_cla4__16_ ;
 wire u_multiplier_STAGE2_Final_add_cla4__17_ ;
 wire u_multiplier_STAGE2_Final_add_cla4__18_ ;
 wire u_multiplier_STAGE2_Final_add_cla4__19_ ;
 wire u_multiplier_STAGE2_Final_add_cla4__20_ ;
 wire u_multiplier_STAGE2_Final_add_cla4__21_ ;
 wire u_multiplier_STAGE2_Final_add_cla4__22_ ;
 wire u_multiplier_STAGE2_Final_add_cla4__23_ ;
 wire u_multiplier_STAGE2_Final_add_cla4__24_ ;
 wire u_multiplier_STAGE2_Final_add_cla4__25_ ;
 wire u_multiplier_STAGE2_Final_add_cla4__26_ ;
 wire u_multiplier_STAGE2_Final_add_cla4__27_ ;
 wire u_multiplier_STAGE2_Final_add_cla4__28_ ;
 wire u_multiplier_STAGE2_Full_adder_pp_13__05_ ;
 wire u_multiplier_STAGE2_Full_adder_pp_13__06_ ;
 wire u_multiplier_STAGE2_Full_adder_pp_13__07_ ;
 wire u_multiplier_STAGE2_Full_adder_pp_13__08_ ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire valid_reg_out;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire [3:0] addr_ptr;
 wire [2:0] curr_state;
 wire [7:0] data_in_reg;
 wire [3:0] init_count;
 wire [15:0] product;
 wire [7:0] sram_rdata;
 wire [7:0] sram_rdata_reg;
 wire [15:0] u_multiplier_approx ;
 wire [1:0] u_multiplier_pp_1 ;
 wire [3:0] u_multiplier_pp_10 ;
 wire [3:0] u_multiplier_pp_11 ;
 wire [3:0] u_multiplier_pp_12 ;
 wire [1:0] u_multiplier_pp_13 ;
 wire [2:0] u_multiplier_pp_2 ;
 wire [3:0] u_multiplier_pp_3 ;
 wire [3:0] u_multiplier_pp_4 ;
 wire [3:0] u_multiplier_pp_5 ;
 wire [3:0] u_multiplier_pp_6 ;
 wire [3:0] u_multiplier_pp_7 ;
 wire [3:0] u_multiplier_pp_8 ;
 wire [3:0] u_multiplier_pp_9 ;

 INV_X1 _279_ (.A(net10),
    .ZN(_050_));
 INV_X1 _280_ (.A(addr_ptr[3]),
    .ZN(_081_));
 INV_X1 _281_ (.A(net101),
    .ZN(_082_));
 INV_X1 _282_ (.A(init_count[2]),
    .ZN(_083_));
 NAND2_X2 _283_ (.A1(_050_),
    .A2(net11),
    .ZN(_084_));
 NAND2_X1 _284_ (.A1(init_count[3]),
    .A2(init_count[2]),
    .ZN(_085_));
 NAND2_X1 _285_ (.A1(init_count[1]),
    .A2(init_count[0]),
    .ZN(_086_));
 NAND4_X1 _286_ (.A1(init_count[1]),
    .A2(init_count[0]),
    .A3(init_count[3]),
    .A4(init_count[2]),
    .ZN(_087_));
 AND2_X1 _287_ (.A1(curr_state[2]),
    .A2(_087_),
    .ZN(_088_));
 AND2_X2 _288_ (.A1(net10),
    .A2(net11),
    .ZN(_089_));
 NAND2_X1 _289_ (.A1(net10),
    .A2(net11),
    .ZN(_090_));
 OAI21_X1 _290_ (.A(_089_),
    .B1(_088_),
    .B2(net12),
    .ZN(_091_));
 NAND2_X1 _291_ (.A1(addr_ptr[0]),
    .A2(addr_ptr[1]),
    .ZN(_092_));
 XOR2_X1 _292_ (.A(addr_ptr[2]),
    .B(_092_),
    .Z(_093_));
 OAI22_X1 _293_ (.A1(net65),
    .A2(_084_),
    .B1(_091_),
    .B2(_093_),
    .ZN(_008_));
 AND4_X1 _294_ (.A1(addr_ptr[2]),
    .A2(net10),
    .A3(addr_ptr[0]),
    .A4(addr_ptr[1]),
    .ZN(_094_));
 OAI21_X1 _295_ (.A(_094_),
    .B1(_088_),
    .B2(_081_),
    .ZN(_095_));
 NOR3_X1 _296_ (.A1(net12),
    .A2(_050_),
    .A3(_088_),
    .ZN(_096_));
 NAND2_X1 _297_ (.A1(_082_),
    .A2(_094_),
    .ZN(_097_));
 NAND2_X1 _298_ (.A1(net11),
    .A2(_097_),
    .ZN(_098_));
 AOI211_X1 _299_ (.A(_096_),
    .B(_098_),
    .C1(net102),
    .C2(_095_),
    .ZN(_009_));
 NAND2_X1 _300_ (.A1(net116),
    .A2(net11),
    .ZN(_051_));
 AND2_X4 _301_ (.A1(net12),
    .A2(net11),
    .ZN(_046_));
 INV_X1 _302_ (.A(_046_),
    .ZN(_099_));
 NAND2_X1 _303_ (.A1(net116),
    .A2(_089_),
    .ZN(_100_));
 OAI21_X1 _304_ (.A(_099_),
    .B1(_100_),
    .B2(_087_),
    .ZN(_048_));
 NAND2_X1 _305_ (.A1(_088_),
    .A2(_089_),
    .ZN(_101_));
 NAND3_X1 _306_ (.A1(net9),
    .A2(net107),
    .A3(_089_),
    .ZN(_102_));
 OAI211_X1 _307_ (.A(_101_),
    .B(net108),
    .C1(net10),
    .C2(_051_),
    .ZN(_049_));
 AOI22_X1 _308_ (.A1(net11),
    .A2(net69),
    .B1(_089_),
    .B2(net9),
    .ZN(_047_));
 AND2_X1 _309_ (.A1(net11),
    .A2(sram_rdata[0]),
    .ZN(_038_));
 AND2_X1 _310_ (.A1(net11),
    .A2(sram_rdata[1]),
    .ZN(_039_));
 AND2_X1 _311_ (.A1(net11),
    .A2(sram_rdata[2]),
    .ZN(_040_));
 AND2_X1 _312_ (.A1(net11),
    .A2(sram_rdata[3]),
    .ZN(_041_));
 AND2_X1 _313_ (.A1(net11),
    .A2(sram_rdata[4]),
    .ZN(_042_));
 AND2_X1 _314_ (.A1(net11),
    .A2(sram_rdata[5]),
    .ZN(_043_));
 AND2_X1 _315_ (.A1(net11),
    .A2(sram_rdata[6]),
    .ZN(_044_));
 AND2_X1 _316_ (.A1(net11),
    .A2(sram_rdata[7]),
    .ZN(_045_));
 AND2_X1 _317_ (.A1(product[0]),
    .A2(_046_),
    .ZN(_018_));
 AND2_X1 _318_ (.A1(product[1]),
    .A2(_046_),
    .ZN(_025_));
 AND2_X1 _319_ (.A1(product[2]),
    .A2(_046_),
    .ZN(_026_));
 AND2_X1 _320_ (.A1(product[3]),
    .A2(_046_),
    .ZN(_027_));
 AND2_X1 _321_ (.A1(product[4]),
    .A2(_046_),
    .ZN(_028_));
 AND2_X1 _322_ (.A1(product[5]),
    .A2(_046_),
    .ZN(_029_));
 AND2_X1 _323_ (.A1(product[6]),
    .A2(_046_),
    .ZN(_030_));
 AND2_X1 _324_ (.A1(product[7]),
    .A2(_046_),
    .ZN(_031_));
 AND2_X1 _325_ (.A1(product[8]),
    .A2(_046_),
    .ZN(_032_));
 AND2_X1 _326_ (.A1(product[9]),
    .A2(_046_),
    .ZN(_033_));
 AND2_X1 _327_ (.A1(product[10]),
    .A2(_046_),
    .ZN(_019_));
 AND2_X1 _328_ (.A1(product[11]),
    .A2(_046_),
    .ZN(_020_));
 AND2_X1 _329_ (.A1(product[12]),
    .A2(_046_),
    .ZN(_021_));
 AND2_X1 _330_ (.A1(product[13]),
    .A2(_046_),
    .ZN(_022_));
 AND2_X1 _331_ (.A1(product[14]),
    .A2(_046_),
    .ZN(_023_));
 AND2_X1 _332_ (.A1(product[15]),
    .A2(_046_),
    .ZN(_024_));
 AND2_X1 _333_ (.A1(net11),
    .A2(net1),
    .ZN(_010_));
 AND2_X1 _334_ (.A1(net11),
    .A2(net2),
    .ZN(_011_));
 AND2_X1 _335_ (.A1(net11),
    .A2(net3),
    .ZN(_012_));
 AND2_X1 _336_ (.A1(net11),
    .A2(net4),
    .ZN(_013_));
 AND2_X1 _337_ (.A1(net11),
    .A2(net5),
    .ZN(_014_));
 AND2_X1 _338_ (.A1(net11),
    .A2(net6),
    .ZN(_015_));
 AND2_X1 _339_ (.A1(net11),
    .A2(net7),
    .ZN(_016_));
 AND2_X1 _340_ (.A1(net11),
    .A2(net8),
    .ZN(_017_));
 OAI21_X1 _341_ (.A(init_count[0]),
    .B1(_267_),
    .B2(_085_),
    .ZN(_103_));
 AOI22_X1 _342_ (.A1(net12),
    .A2(init_count[0]),
    .B1(_103_),
    .B2(curr_state[2]),
    .ZN(_104_));
 OAI22_X1 _343_ (.A1(net99),
    .A2(_084_),
    .B1(_090_),
    .B2(_104_),
    .ZN(_034_));
 NAND3_X1 _344_ (.A1(init_count[1]),
    .A2(init_count[0]),
    .A3(_085_),
    .ZN(_105_));
 OAI21_X1 _345_ (.A(curr_state[2]),
    .B1(init_count[1]),
    .B2(init_count[0]),
    .ZN(_106_));
 INV_X1 _346_ (.A(_106_),
    .ZN(_107_));
 AOI22_X1 _347_ (.A1(net12),
    .A2(init_count[1]),
    .B1(_105_),
    .B2(_107_),
    .ZN(_108_));
 OAI22_X1 _348_ (.A1(net105),
    .A2(_084_),
    .B1(_090_),
    .B2(_108_),
    .ZN(_035_));
 OR3_X1 _349_ (.A1(init_count[3]),
    .A2(_083_),
    .A3(_086_),
    .ZN(_109_));
 AOI21_X1 _350_ (.A(net12),
    .B1(_109_),
    .B2(curr_state[2]),
    .ZN(_110_));
 AND3_X1 _351_ (.A1(curr_state[2]),
    .A2(init_count[1]),
    .A3(init_count[0]),
    .ZN(_111_));
 OAI21_X1 _352_ (.A(_089_),
    .B1(_111_),
    .B2(init_count[2]),
    .ZN(_112_));
 OAI22_X1 _353_ (.A1(net96),
    .A2(_084_),
    .B1(_110_),
    .B2(_112_),
    .ZN(_036_));
 OAI21_X1 _354_ (.A(net92),
    .B1(_086_),
    .B2(_268_),
    .ZN(_113_));
 AOI22_X1 _355_ (.A1(net12),
    .A2(init_count[3]),
    .B1(_113_),
    .B2(curr_state[2]),
    .ZN(_114_));
 OAI22_X1 _356_ (.A1(net93),
    .A2(_084_),
    .B1(_090_),
    .B2(_114_),
    .ZN(_037_));
 NAND3_X1 _357_ (.A1(net88),
    .A2(_088_),
    .A3(_089_),
    .ZN(_115_));
 NAND2_X1 _358_ (.A1(net10),
    .A2(_046_),
    .ZN(_116_));
 OAI221_X1 _359_ (.A(net89),
    .B1(_116_),
    .B2(addr_ptr[0]),
    .C1(net79),
    .C2(_084_),
    .ZN(_006_));
 XNOR2_X1 _360_ (.A(addr_ptr[0]),
    .B(addr_ptr[1]),
    .ZN(_117_));
 OAI22_X1 _361_ (.A1(net67),
    .A2(_084_),
    .B1(_091_),
    .B2(_117_),
    .ZN(_007_));
 DFF_X1 _362_ (.D(net70),
    .CK(clknet_2_1__leaf_clk),
    .Q(curr_state[0]),
    .QN(_226_));
 DFF_X2 _363_ (.D(net117),
    .CK(clknet_2_1__leaf_clk),
    .Q(net12),
    .QN(_227_));
 DFF_X2 _364_ (.D(net109),
    .CK(clknet_2_1__leaf_clk),
    .Q(curr_state[2]),
    .QN(_228_));
 DFF_X1 _365_ (.D(_018_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net13),
    .QN(_229_));
 DFF_X2 _366_ (.D(_025_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net20),
    .QN(_230_));
 DFF_X1 _367_ (.D(_026_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net21),
    .QN(_231_));
 DFF_X2 _368_ (.D(_027_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net22),
    .QN(_232_));
 DFF_X1 _369_ (.D(_028_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net23),
    .QN(_233_));
 DFF_X1 _370_ (.D(_029_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net24),
    .QN(_234_));
 DFF_X1 _371_ (.D(_030_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net25),
    .QN(_235_));
 DFF_X1 _372_ (.D(_031_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net26),
    .QN(_236_));
 DFF_X1 _373_ (.D(_032_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net27),
    .QN(_237_));
 DFF_X2 _374_ (.D(_033_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net28),
    .QN(_238_));
 DFF_X1 _375_ (.D(_019_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net14),
    .QN(_239_));
 DFF_X2 _376_ (.D(_020_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net15),
    .QN(_240_));
 DFF_X1 _377_ (.D(_021_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net16),
    .QN(_241_));
 DFF_X1 _378_ (.D(_022_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net17),
    .QN(_242_));
 DFF_X2 _379_ (.D(_023_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net18),
    .QN(_243_));
 DFF_X1 _380_ (.D(_024_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net19),
    .QN(_244_));
 DFF_X2 _381_ (.D(_010_),
    .CK(clknet_2_0__leaf_clk),
    .Q(data_in_reg[0]),
    .QN(_245_));
 DFF_X2 _382_ (.D(_011_),
    .CK(clknet_2_0__leaf_clk),
    .Q(data_in_reg[1]),
    .QN(_246_));
 DFF_X2 _383_ (.D(_012_),
    .CK(clknet_2_2__leaf_clk),
    .Q(data_in_reg[2]),
    .QN(_247_));
 DFF_X2 _384_ (.D(_013_),
    .CK(clknet_2_0__leaf_clk),
    .Q(data_in_reg[3]),
    .QN(_248_));
 DFF_X2 _385_ (.D(_014_),
    .CK(clknet_2_2__leaf_clk),
    .Q(data_in_reg[4]),
    .QN(_249_));
 DFF_X2 _386_ (.D(_015_),
    .CK(clknet_2_2__leaf_clk),
    .Q(data_in_reg[5]),
    .QN(_250_));
 DFF_X2 _387_ (.D(_016_),
    .CK(clknet_2_2__leaf_clk),
    .Q(data_in_reg[6]),
    .QN(_251_));
 DFF_X2 _388_ (.D(_017_),
    .CK(clknet_2_0__leaf_clk),
    .Q(data_in_reg[7]),
    .QN(_252_));
 DFF_X2 _389_ (.D(_038_),
    .CK(clknet_2_0__leaf_clk),
    .Q(sram_rdata_reg[0]),
    .QN(_253_));
 DFF_X2 _390_ (.D(_039_),
    .CK(clknet_2_0__leaf_clk),
    .Q(sram_rdata_reg[1]),
    .QN(_254_));
 DFF_X2 _391_ (.D(_040_),
    .CK(clknet_2_2__leaf_clk),
    .Q(sram_rdata_reg[2]),
    .QN(_255_));
 DFF_X2 _392_ (.D(_041_),
    .CK(clknet_2_2__leaf_clk),
    .Q(sram_rdata_reg[3]),
    .QN(_256_));
 DFF_X2 _393_ (.D(_042_),
    .CK(clknet_2_2__leaf_clk),
    .Q(sram_rdata_reg[4]),
    .QN(_257_));
 DFF_X2 _394_ (.D(_043_),
    .CK(clknet_2_2__leaf_clk),
    .Q(sram_rdata_reg[5]),
    .QN(_258_));
 DFF_X2 _395_ (.D(_044_),
    .CK(clknet_2_2__leaf_clk),
    .Q(sram_rdata_reg[6]),
    .QN(_259_));
 DFF_X1 _396_ (.D(_045_),
    .CK(clknet_2_3__leaf_clk),
    .Q(sram_rdata_reg[7]),
    .QN(_260_));
 DFF_X1 _397_ (.D(_046_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net29),
    .QN(_261_));
 DFF_X2 _398_ (.D(net90),
    .CK(clknet_2_1__leaf_clk),
    .Q(addr_ptr[0]),
    .QN(_262_));
 DFF_X1 _399_ (.D(net68),
    .CK(clknet_2_1__leaf_clk),
    .Q(addr_ptr[1]),
    .QN(_263_));
 DFF_X1 _400_ (.D(net66),
    .CK(clknet_2_1__leaf_clk),
    .Q(addr_ptr[2]),
    .QN(_264_));
 DFF_X1 _401_ (.D(net103),
    .CK(clknet_2_1__leaf_clk),
    .Q(addr_ptr[3]),
    .QN(_265_));
 DFF_X2 _402_ (.D(net100),
    .CK(clknet_2_1__leaf_clk),
    .Q(init_count[0]),
    .QN(_266_));
 DFF_X2 _403_ (.D(net106),
    .CK(clknet_2_1__leaf_clk),
    .Q(init_count[1]),
    .QN(_267_));
 DFF_X1 _404_ (.D(net97),
    .CK(clknet_2_1__leaf_clk),
    .Q(init_count[2]),
    .QN(_268_));
 DFF_X1 _405_ (.D(net94),
    .CK(clknet_2_1__leaf_clk),
    .Q(init_count[3]),
    .QN(_269_));
 SRAM_6T_CORE_16x8_MC_TB sram_inst (.ce_in(_050_),
    .we_in(_051_),
    .clk(clknet_2_0__leaf_clk),
    .addr_in({net113,
    net78,
    net111,
    net80}),
    .rd_out({sram_rdata[7],
    sram_rdata[6],
    sram_rdata[5],
    sram_rdata[4],
    sram_rdata[3],
    sram_rdata[2],
    sram_rdata[1],
    sram_rdata[0]}),
    .wd_in({net81,
    net82,
    net83,
    net84,
    net91,
    net87,
    net86,
    net85}));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_10__18_  (.A(u_multiplier_STAGE1_pp_9_c2 ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_10__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_10__19_  (.A1(u_multiplier_STAGE1__050_ ),
    .A2(u_multiplier_STAGE1__049_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_10__08_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_10__20_  (.A(u_multiplier_STAGE1__050_ ),
    .B(u_multiplier_STAGE1__049_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_10__09_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_10__21_  (.A1(u_multiplier_STAGE1__051_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_10__09_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_10__10_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_10__22_  (.A(u_multiplier_STAGE1__051_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_10__09_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_10__11_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_10__23_  (.A1(u_multiplier_STAGE1__052_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_10__11_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_10__12_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_10__24_  (.A(u_multiplier_STAGE1__052_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_10__11_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_10__13_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_10__25_  (.A(u_multiplier_STAGE1_pp_9_c2 ),
    .B(u_multiplier_STAGE1_E_4_2_pp_10__13_ ),
    .ZN(u_multiplier_pp_10 [3]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_10__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_10__08_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_10__10_ ),
    .ZN(u_multiplier_STAGE1_pp_10_c2 ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_10__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_10__12_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_10__13_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_10__14_ ),
    .ZN(u_multiplier_pp_11 [0]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_5__18_  (.A(net46),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_5__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_5__19_  (.A1(u_multiplier_STAGE1__019_ ),
    .A2(u_multiplier_STAGE1__018_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_5__08_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_5__20_  (.A(u_multiplier_STAGE1__019_ ),
    .B(u_multiplier_STAGE1__018_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_5__09_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_5__21_  (.A1(u_multiplier_STAGE1__020_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_5__09_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_5__10_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_5__22_  (.A(u_multiplier_STAGE1__020_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_5__09_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_5__11_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_5__23_  (.A1(u_multiplier_STAGE1__021_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_5__11_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_5__12_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_5__24_  (.A(u_multiplier_STAGE1__021_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_5__11_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_5__13_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_5__25_  (.A(net47),
    .B(u_multiplier_STAGE1_E_4_2_pp_5__13_ ),
    .ZN(u_multiplier_pp_5 [0]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_5__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_5__08_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_5__10_ ),
    .ZN(u_multiplier_STAGE1_pp_5_c2 ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_5__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_5__12_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_5__13_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_5__14_ ),
    .ZN(u_multiplier_pp_6 [3]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_6__18_  (.A(u_multiplier_STAGE1_pp_5_c2 ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_6__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_6__19_  (.A1(u_multiplier_STAGE1__023_ ),
    .A2(u_multiplier_STAGE1__022_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_6__08_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_6__20_  (.A(u_multiplier_STAGE1__023_ ),
    .B(u_multiplier_STAGE1__022_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_6__09_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_6__21_  (.A1(u_multiplier_STAGE1__024_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_6__09_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_6__10_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_6__22_  (.A(u_multiplier_STAGE1__024_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_6__09_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_6__11_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_6__23_  (.A1(u_multiplier_STAGE1__025_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_6__11_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_6__12_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_6__24_  (.A(u_multiplier_STAGE1__025_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_6__11_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_6__13_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_6__25_  (.A(u_multiplier_STAGE1_pp_5_c2 ),
    .B(u_multiplier_STAGE1_E_4_2_pp_6__13_ ),
    .ZN(u_multiplier_pp_6 [0]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_6__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_6__08_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_6__10_ ),
    .ZN(u_multiplier_STAGE1_pp_6_c2 ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_6__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_6__12_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_6__13_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_6__14_ ),
    .ZN(u_multiplier_pp_7 [2]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_7_1__18_  (.A(u_multiplier_STAGE1_pp_6_c2 ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_7_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_7_1__19_  (.A1(u_multiplier_STAGE1__029_ ),
    .A2(u_multiplier_STAGE1__028_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_7_1__08_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_7_1__20_  (.A(u_multiplier_STAGE1__029_ ),
    .B(u_multiplier_STAGE1__028_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_7_1__09_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_7_1__21_  (.A1(u_multiplier_STAGE1__030_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_7_1__09_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_7_1__10_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_7_1__22_  (.A(u_multiplier_STAGE1__030_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_7_1__09_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_7_1__11_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_7_1__23_  (.A1(u_multiplier_STAGE1__031_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_7_1__11_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_7_1__12_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_7_1__24_  (.A(u_multiplier_STAGE1__031_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_7_1__11_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_7_1__13_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_7_1__25_  (.A(u_multiplier_STAGE1_pp_6_c2 ),
    .B(u_multiplier_STAGE1_E_4_2_pp_7_1__13_ ),
    .ZN(u_multiplier_pp_7 [0]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_7_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_7_1__08_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_7_1__10_ ),
    .ZN(u_multiplier_STAGE1_pp_7_c2 ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_7_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_7_1__12_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_7_1__13_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_7_1__14_ ),
    .ZN(u_multiplier_pp_8 [2]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_7_2__18_  (.A(net48),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_7_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_7_2__19_  (.A1(u_multiplier_STAGE1__033_ ),
    .A2(u_multiplier_STAGE1__032_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_7_2__08_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_7_2__20_  (.A(u_multiplier_STAGE1__033_ ),
    .B(u_multiplier_STAGE1__032_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_7_2__09_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_7_2__21_  (.A1(u_multiplier_STAGE1__034_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_7_2__09_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_7_2__10_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_7_2__22_  (.A(u_multiplier_STAGE1__034_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_7_2__09_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_7_2__11_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_7_2__23_  (.A1(u_multiplier_STAGE1__035_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_7_2__11_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_7_2__12_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_7_2__24_  (.A(u_multiplier_STAGE1__035_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_7_2__11_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_7_2__13_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_7_2__25_  (.A(net49),
    .B(u_multiplier_STAGE1_E_4_2_pp_7_2__13_ ),
    .ZN(u_multiplier_pp_7 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_7_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_7_2__08_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_7_2__10_ ),
    .ZN(u_multiplier_STAGE1_pp_7_c4 ));
 OAI21_X1 u_multiplier_STAGE1_E_4_2_pp_7_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_7_2__12_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_7_2__13_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_7_2__14_ ),
    .ZN(u_multiplier_pp_8 [3]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_8_1__18_  (.A(u_multiplier_STAGE1_pp_7_c2 ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_8_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_8_1__19_  (.A1(u_multiplier_STAGE1__037_ ),
    .A2(u_multiplier_STAGE1__036_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_8_1__08_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_8_1__20_  (.A(u_multiplier_STAGE1__037_ ),
    .B(u_multiplier_STAGE1__036_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_8_1__09_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_8_1__21_  (.A1(u_multiplier_STAGE1__038_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_8_1__09_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_8_1__10_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_8_1__22_  (.A(u_multiplier_STAGE1__038_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_8_1__09_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_8_1__11_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_8_1__23_  (.A1(u_multiplier_STAGE1__039_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_8_1__11_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_8_1__12_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_8_1__24_  (.A(u_multiplier_STAGE1__039_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_8_1__11_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_8_1__13_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_8_1__25_  (.A(u_multiplier_STAGE1_pp_7_c2 ),
    .B(u_multiplier_STAGE1_E_4_2_pp_8_1__13_ ),
    .ZN(u_multiplier_pp_8 [0]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_8_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_8_1__08_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_8_1__10_ ),
    .ZN(u_multiplier_STAGE1_pp_8_c2 ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_8_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_8_1__12_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_8_1__13_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_8_1__14_ ),
    .ZN(u_multiplier_pp_9 [2]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_8_2__18_  (.A(net50),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_8_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_8_2__19_  (.A1(u_multiplier_STAGE1__041_ ),
    .A2(u_multiplier_STAGE1__040_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_8_2__08_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_8_2__20_  (.A(u_multiplier_STAGE1__041_ ),
    .B(u_multiplier_STAGE1__040_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_8_2__09_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_8_2__21_  (.A1(u_multiplier_STAGE1__042_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_8_2__09_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_8_2__10_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_8_2__22_  (.A(u_multiplier_STAGE1__042_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_8_2__09_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_8_2__11_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_8_2__23_  (.A1(u_multiplier_STAGE1_pp_7_c4 ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_8_2__11_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_8_2__12_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_8_2__24_  (.A(u_multiplier_STAGE1_pp_7_c4 ),
    .B(u_multiplier_STAGE1_E_4_2_pp_8_2__11_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_8_2__13_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_8_2__25_  (.A(net51),
    .B(u_multiplier_STAGE1_E_4_2_pp_8_2__13_ ),
    .ZN(u_multiplier_pp_8 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_8_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_8_2__08_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_8_2__10_ ),
    .ZN(u_multiplier_STAGE1_pp_8_c4 ));
 OAI21_X1 u_multiplier_STAGE1_E_4_2_pp_8_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_8_2__12_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_8_2__13_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_8_2__14_ ),
    .ZN(u_multiplier_pp_9 [3]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_9_1__18_  (.A(u_multiplier_STAGE1_pp_8_c2 ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_9_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_9_1__19_  (.A1(u_multiplier_STAGE1__044_ ),
    .A2(u_multiplier_STAGE1__043_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_9_1__08_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_9_1__20_  (.A(u_multiplier_STAGE1__044_ ),
    .B(u_multiplier_STAGE1__043_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_9_1__09_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_9_1__21_  (.A1(u_multiplier_STAGE1__045_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_9_1__09_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_9_1__10_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_9_1__22_  (.A(u_multiplier_STAGE1__045_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_9_1__09_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_9_1__11_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_9_1__23_  (.A1(u_multiplier_STAGE1__046_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_9_1__11_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_9_1__12_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_9_1__24_  (.A(u_multiplier_STAGE1__046_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_9_1__11_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_9_1__13_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_9_1__25_  (.A(u_multiplier_STAGE1_pp_8_c2 ),
    .B(u_multiplier_STAGE1_E_4_2_pp_9_1__13_ ),
    .ZN(u_multiplier_pp_9 [0]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_9_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_9_1__08_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_9_1__10_ ),
    .ZN(u_multiplier_STAGE1_pp_9_c2 ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_9_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_9_1__12_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_9_1__13_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_9_1__14_ ),
    .ZN(u_multiplier_pp_10 [1]));
 INV_X1 u_multiplier_STAGE1_Full_adder_pp_11__12_  (.A(u_multiplier_STAGE1_pp_10_c2 ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_11__05_ ));
 NAND3_X1 u_multiplier_STAGE1_Full_adder_pp_11__13_  (.A1(u_multiplier_STAGE1__054_ ),
    .A2(u_multiplier_STAGE1__053_ ),
    .A3(u_multiplier_STAGE1_pp_10_c2 ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_11__06_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_11__14_  (.A1(u_multiplier_STAGE1__054_ ),
    .A2(u_multiplier_STAGE1__053_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_11__07_ ));
 AOI21_X1 u_multiplier_STAGE1_Full_adder_pp_11__15_  (.A(u_multiplier_STAGE1_pp_10_c2 ),
    .B1(u_multiplier_STAGE1__053_ ),
    .B2(u_multiplier_STAGE1__054_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_11__08_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_11__16_  (.A1(u_multiplier_STAGE1_Full_adder_pp_11__07_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_11__08_ ),
    .ZN(u_multiplier_pp_12 [0]));
 AOI22_X4 u_multiplier_STAGE1_Full_adder_pp_11__17_  (.A1(u_multiplier_STAGE1_Full_adder_pp_11__05_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_11__07_ ),
    .B1(u_multiplier_pp_12 [0]),
    .B2(u_multiplier_STAGE1_Full_adder_pp_11__06_ ),
    .ZN(u_multiplier_pp_11 [3]));
 INV_X1 u_multiplier_STAGE1_Full_adder_pp_9__12_  (.A(u_multiplier_STAGE1_pp_8_c4 ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_9__05_ ));
 NAND3_X1 u_multiplier_STAGE1_Full_adder_pp_9__13_  (.A1(u_multiplier_STAGE1__048_ ),
    .A2(u_multiplier_STAGE1__047_ ),
    .A3(u_multiplier_STAGE1_pp_8_c4 ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_9__06_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_9__14_  (.A1(u_multiplier_STAGE1__048_ ),
    .A2(u_multiplier_STAGE1__047_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_9__07_ ));
 AOI21_X1 u_multiplier_STAGE1_Full_adder_pp_9__15_  (.A(u_multiplier_STAGE1_pp_8_c4 ),
    .B1(u_multiplier_STAGE1__047_ ),
    .B2(u_multiplier_STAGE1__048_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_9__08_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_9__16_  (.A1(u_multiplier_STAGE1_Full_adder_pp_9__07_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_9__08_ ),
    .ZN(u_multiplier_pp_10 [0]));
 AOI22_X2 u_multiplier_STAGE1_Full_adder_pp_9__17_  (.A1(u_multiplier_STAGE1_Full_adder_pp_9__05_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_9__07_ ),
    .B1(u_multiplier_pp_10 [0]),
    .B2(u_multiplier_STAGE1_Full_adder_pp_9__06_ ),
    .ZN(u_multiplier_pp_9 [1]));
 AND2_X1 u_multiplier_STAGE1_Half_adder_pp_4__4_  (.A1(u_multiplier_STAGE1__017_ ),
    .A2(u_multiplier_STAGE1__016_ ),
    .ZN(u_multiplier_pp_5 [3]));
 XOR2_X2 u_multiplier_STAGE1_Half_adder_pp_4__5_  (.A(u_multiplier_STAGE1__017_ ),
    .B(u_multiplier_STAGE1__016_ ),
    .Z(u_multiplier_pp_4 [0]));
 AND2_X1 u_multiplier_STAGE1_Half_adder_pp_6__4_  (.A1(u_multiplier_STAGE1__027_ ),
    .A2(u_multiplier_STAGE1__026_ ),
    .ZN(u_multiplier_pp_7 [3]));
 XOR2_X2 u_multiplier_STAGE1_Half_adder_pp_6__5_  (.A(u_multiplier_STAGE1__027_ ),
    .B(u_multiplier_STAGE1__026_ ),
    .Z(u_multiplier_pp_6 [1]));
 AND2_X1 u_multiplier_STAGE1__119_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[0]),
    .ZN(u_multiplier_pp_0 ));
 AND2_X1 u_multiplier_STAGE1__120_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[1]),
    .ZN(u_multiplier_pp_1 [0]));
 AND2_X1 u_multiplier_STAGE1__121_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[1]),
    .ZN(u_multiplier_pp_1 [1]));
 AND2_X1 u_multiplier_STAGE1__122_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[2]),
    .ZN(u_multiplier_pp_2 [0]));
 AND2_X1 u_multiplier_STAGE1__123_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[1]),
    .ZN(u_multiplier_pp_2 [1]));
 AND2_X1 u_multiplier_STAGE1__124_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[2]),
    .ZN(u_multiplier_pp_2 [2]));
 AND2_X1 u_multiplier_STAGE1__125_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[3]),
    .ZN(u_multiplier_pp_3 [0]));
 AND2_X1 u_multiplier_STAGE1__126_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[2]),
    .ZN(u_multiplier_pp_3 [1]));
 AND2_X1 u_multiplier_STAGE1__127_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[2]),
    .ZN(u_multiplier_pp_3 [2]));
 AND2_X1 u_multiplier_STAGE1__128_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[3]),
    .ZN(u_multiplier_pp_3 [3]));
 AND2_X1 u_multiplier_STAGE1__129_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[2]),
    .ZN(u_multiplier_pp_4 [1]));
 AND2_X1 u_multiplier_STAGE1__130_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[3]),
    .ZN(u_multiplier_pp_4 [2]));
 AND2_X1 u_multiplier_STAGE1__131_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[4]),
    .ZN(u_multiplier_pp_4 [3]));
 AND2_X1 u_multiplier_STAGE1__132_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[4]),
    .ZN(u_multiplier_pp_5 [1]));
 AND2_X1 u_multiplier_STAGE1__133_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[5]),
    .ZN(u_multiplier_pp_5 [2]));
 AND2_X1 u_multiplier_STAGE1__134_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[6]),
    .ZN(u_multiplier_pp_6 [2]));
 AND2_X1 u_multiplier_STAGE1__135_  (.A1(data_in_reg[3]),
    .A2(net30),
    .ZN(u_multiplier_pp_10 [2]));
 AND2_X1 u_multiplier_STAGE1__136_  (.A1(net31),
    .A2(data_in_reg[4]),
    .ZN(u_multiplier_pp_11 [1]));
 AND2_X1 u_multiplier_STAGE1__137_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[5]),
    .ZN(u_multiplier_pp_11 [2]));
 AND2_X1 u_multiplier_STAGE1__138_  (.A1(net32),
    .A2(data_in_reg[5]),
    .ZN(u_multiplier_pp_12 [1]));
 AND2_X1 u_multiplier_STAGE1__139_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[6]),
    .ZN(u_multiplier_pp_12 [2]));
 AND2_X1 u_multiplier_STAGE1__140_  (.A1(sram_rdata_reg[5]),
    .A2(net33),
    .ZN(u_multiplier_pp_12 [3]));
 AND2_X1 u_multiplier_STAGE1__141_  (.A1(net34),
    .A2(data_in_reg[6]),
    .ZN(u_multiplier_pp_13 [0]));
 AND2_X1 u_multiplier_STAGE1__142_  (.A1(sram_rdata_reg[6]),
    .A2(net35),
    .ZN(u_multiplier_pp_13 [1]));
 AND2_X1 u_multiplier_STAGE1__143_  (.A1(net36),
    .A2(net37),
    .ZN(u_multiplier_pp_14 ));
 AND2_X1 u_multiplier_STAGE1__144_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[4]),
    .ZN(u_multiplier_STAGE1__016_ ));
 AND2_X1 u_multiplier_STAGE1__145_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[3]),
    .ZN(u_multiplier_STAGE1__017_ ));
 AND2_X1 u_multiplier_STAGE1__146_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[5]),
    .ZN(u_multiplier_STAGE1__018_ ));
 AND2_X1 u_multiplier_STAGE1__147_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[4]),
    .ZN(u_multiplier_STAGE1__019_ ));
 AND2_X1 u_multiplier_STAGE1__148_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[3]),
    .ZN(u_multiplier_STAGE1__020_ ));
 AND2_X1 u_multiplier_STAGE1__149_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[3]),
    .ZN(u_multiplier_STAGE1__021_ ));
 AND2_X1 u_multiplier_STAGE1__150_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[6]),
    .ZN(u_multiplier_STAGE1__022_ ));
 AND2_X1 u_multiplier_STAGE1__151_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[5]),
    .ZN(u_multiplier_STAGE1__023_ ));
 AND2_X1 u_multiplier_STAGE1__152_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[4]),
    .ZN(u_multiplier_STAGE1__024_ ));
 AND2_X1 u_multiplier_STAGE1__153_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[3]),
    .ZN(u_multiplier_STAGE1__025_ ));
 AND2_X1 u_multiplier_STAGE1__154_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[4]),
    .ZN(u_multiplier_STAGE1__026_ ));
 AND2_X1 u_multiplier_STAGE1__155_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[5]),
    .ZN(u_multiplier_STAGE1__027_ ));
 AND2_X1 u_multiplier_STAGE1__156_  (.A1(sram_rdata_reg[0]),
    .A2(net38),
    .ZN(u_multiplier_STAGE1__028_ ));
 AND2_X1 u_multiplier_STAGE1__157_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[6]),
    .ZN(u_multiplier_STAGE1__029_ ));
 AND2_X1 u_multiplier_STAGE1__158_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[5]),
    .ZN(u_multiplier_STAGE1__030_ ));
 AND2_X1 u_multiplier_STAGE1__159_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[4]),
    .ZN(u_multiplier_STAGE1__031_ ));
 AND2_X1 u_multiplier_STAGE1__160_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[4]),
    .ZN(u_multiplier_STAGE1__032_ ));
 AND2_X1 u_multiplier_STAGE1__161_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[5]),
    .ZN(u_multiplier_STAGE1__033_ ));
 AND2_X1 u_multiplier_STAGE1__162_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[6]),
    .ZN(u_multiplier_STAGE1__034_ ));
 AND2_X1 u_multiplier_STAGE1__163_  (.A1(data_in_reg[0]),
    .A2(net39),
    .ZN(u_multiplier_STAGE1__035_ ));
 AND2_X1 u_multiplier_STAGE1__164_  (.A1(sram_rdata_reg[1]),
    .A2(net40),
    .ZN(u_multiplier_STAGE1__036_ ));
 AND2_X1 u_multiplier_STAGE1__165_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[6]),
    .ZN(u_multiplier_STAGE1__037_ ));
 AND2_X1 u_multiplier_STAGE1__166_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[5]),
    .ZN(u_multiplier_STAGE1__038_ ));
 AND2_X1 u_multiplier_STAGE1__167_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[4]),
    .ZN(u_multiplier_STAGE1__039_ ));
 AND2_X1 u_multiplier_STAGE1__168_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[5]),
    .ZN(u_multiplier_STAGE1__040_ ));
 AND2_X1 u_multiplier_STAGE1__169_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[6]),
    .ZN(u_multiplier_STAGE1__041_ ));
 AND2_X1 u_multiplier_STAGE1__170_  (.A1(data_in_reg[1]),
    .A2(net41),
    .ZN(u_multiplier_STAGE1__042_ ));
 AND2_X1 u_multiplier_STAGE1__171_  (.A1(sram_rdata_reg[2]),
    .A2(net42),
    .ZN(u_multiplier_STAGE1__043_ ));
 AND2_X1 u_multiplier_STAGE1__172_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[6]),
    .ZN(u_multiplier_STAGE1__044_ ));
 AND2_X1 u_multiplier_STAGE1__173_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[5]),
    .ZN(u_multiplier_STAGE1__045_ ));
 AND2_X1 u_multiplier_STAGE1__174_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[4]),
    .ZN(u_multiplier_STAGE1__046_ ));
 AND2_X1 u_multiplier_STAGE1__175_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[6]),
    .ZN(u_multiplier_STAGE1__047_ ));
 AND2_X1 u_multiplier_STAGE1__176_  (.A1(data_in_reg[2]),
    .A2(net43),
    .ZN(u_multiplier_STAGE1__048_ ));
 AND2_X1 u_multiplier_STAGE1__177_  (.A1(sram_rdata_reg[3]),
    .A2(net44),
    .ZN(u_multiplier_STAGE1__049_ ));
 AND2_X1 u_multiplier_STAGE1__178_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[6]),
    .ZN(u_multiplier_STAGE1__050_ ));
 AND2_X1 u_multiplier_STAGE1__179_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[5]),
    .ZN(u_multiplier_STAGE1__051_ ));
 AND2_X1 u_multiplier_STAGE1__180_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[4]),
    .ZN(u_multiplier_STAGE1__052_ ));
 AND2_X1 u_multiplier_STAGE1__181_  (.A1(sram_rdata_reg[4]),
    .A2(net45),
    .ZN(u_multiplier_STAGE1__053_ ));
 AND2_X1 u_multiplier_STAGE1__182_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[6]),
    .ZN(u_multiplier_STAGE1__054_ ));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp_10__18_  (.A(u_multiplier_STAGE2_pp_9_c2 ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_10__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_10__19_  (.A1(u_multiplier_pp_10 [1]),
    .A2(u_multiplier_pp_10 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_10__08_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp_10__20_  (.A(u_multiplier_pp_10 [1]),
    .B(u_multiplier_pp_10 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp_10__09_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_10__21_  (.A1(u_multiplier_pp_10 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp_10__09_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_10__10_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp_10__22_  (.A(u_multiplier_pp_10 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp_10__09_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp_10__11_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_10__23_  (.A1(u_multiplier_pp_10 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp_10__11_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_10__12_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp_10__24_  (.A(u_multiplier_pp_10 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp_10__11_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_10__13_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp_10__25_  (.A(u_multiplier_STAGE2_pp_9_c2 ),
    .B(u_multiplier_STAGE2_E_4_2_pp_10__13_ ),
    .ZN(u_multiplier_STAGE2_pp_10_s ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_10__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp_10__08_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp_10__10_ ),
    .ZN(u_multiplier_STAGE2_pp_10_c2 ));
 OAI21_X1 u_multiplier_STAGE2_E_4_2_pp_10__27_  (.A(u_multiplier_STAGE2_E_4_2_pp_10__12_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp_10__13_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp_10__14_ ),
    .ZN(u_multiplier_STAGE2_pp_10_c1 ));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp_11__18_  (.A(u_multiplier_STAGE2_pp_10_c2 ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_11__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_11__19_  (.A1(u_multiplier_pp_11 [1]),
    .A2(u_multiplier_pp_11 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_11__08_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp_11__20_  (.A(u_multiplier_pp_11 [1]),
    .B(u_multiplier_pp_11 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp_11__09_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_11__21_  (.A1(u_multiplier_pp_11 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp_11__09_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_11__10_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp_11__22_  (.A(u_multiplier_pp_11 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp_11__09_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp_11__11_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_11__23_  (.A1(u_multiplier_pp_11 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp_11__11_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_11__12_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp_11__24_  (.A(u_multiplier_pp_11 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp_11__11_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_11__13_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp_11__25_  (.A(u_multiplier_STAGE2_pp_10_c2 ),
    .B(u_multiplier_STAGE2_E_4_2_pp_11__13_ ),
    .ZN(u_multiplier_STAGE2_pp_11_s ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_11__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp_11__08_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp_11__10_ ),
    .ZN(u_multiplier_STAGE2_pp_11_c2 ));
 OAI21_X1 u_multiplier_STAGE2_E_4_2_pp_11__27_  (.A(u_multiplier_STAGE2_E_4_2_pp_11__12_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp_11__13_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp_11__14_ ),
    .ZN(u_multiplier_STAGE2_pp_11_c1 ));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp_12__18_  (.A(u_multiplier_STAGE2_pp_11_c2 ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_12__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_12__19_  (.A1(u_multiplier_pp_12 [1]),
    .A2(u_multiplier_pp_12 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_12__08_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp_12__20_  (.A(u_multiplier_pp_12 [1]),
    .B(u_multiplier_pp_12 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp_12__09_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_12__21_  (.A1(u_multiplier_pp_12 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp_12__09_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_12__10_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp_12__22_  (.A(u_multiplier_pp_12 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp_12__09_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp_12__11_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_12__23_  (.A1(u_multiplier_pp_12 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp_12__11_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_12__12_ ));
 XNOR2_X1 u_multiplier_STAGE2_E_4_2_pp_12__24_  (.A(u_multiplier_pp_12 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp_12__11_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_12__13_ ));
 XNOR2_X1 u_multiplier_STAGE2_E_4_2_pp_12__25_  (.A(u_multiplier_STAGE2_pp_11_c2 ),
    .B(u_multiplier_STAGE2_E_4_2_pp_12__13_ ),
    .ZN(u_multiplier_STAGE2_pp_12_s ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_12__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp_12__08_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp_12__10_ ),
    .ZN(u_multiplier_STAGE2_pp_12_c2 ));
 OAI21_X1 u_multiplier_STAGE2_E_4_2_pp_12__27_  (.A(u_multiplier_STAGE2_E_4_2_pp_12__12_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp_12__13_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp_12__14_ ),
    .ZN(u_multiplier_STAGE2_pp_12_c1 ));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp_3__18_  (.A(net52),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_3__19_  (.A1(u_multiplier_pp_3 [1]),
    .A2(u_multiplier_pp_3 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_3__08_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp_3__20_  (.A(u_multiplier_pp_3 [1]),
    .B(u_multiplier_pp_3 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp_3__09_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_3__21_  (.A1(u_multiplier_pp_3 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp_3__09_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_3__10_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp_3__22_  (.A(u_multiplier_pp_3 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp_3__09_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp_3__11_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_3__23_  (.A1(u_multiplier_pp_3 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp_3__11_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_3__12_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp_3__24_  (.A(u_multiplier_pp_3 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp_3__11_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_3__13_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp_3__25_  (.A(net53),
    .B(u_multiplier_STAGE2_E_4_2_pp_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp_3_s ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp_3__08_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp_3__10_ ),
    .ZN(u_multiplier_STAGE2_pp_3_c2 ));
 OAI21_X1 u_multiplier_STAGE2_E_4_2_pp_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp_3__12_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp_3__13_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp_3__14_ ),
    .ZN(u_multiplier_STAGE2_pp_3_c1 ));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp_4__18_  (.A(u_multiplier_STAGE2_pp_3_c2 ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_4__19_  (.A1(u_multiplier_pp_4 [1]),
    .A2(u_multiplier_pp_4 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_4__08_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp_4__20_  (.A(u_multiplier_pp_4 [1]),
    .B(u_multiplier_pp_4 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp_4__09_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_4__21_  (.A1(u_multiplier_pp_4 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp_4__09_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_4__10_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp_4__22_  (.A(u_multiplier_pp_4 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp_4__09_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp_4__11_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_4__23_  (.A1(u_multiplier_pp_4 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp_4__11_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_4__12_ ));
 XNOR2_X1 u_multiplier_STAGE2_E_4_2_pp_4__24_  (.A(u_multiplier_pp_4 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp_4__11_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_4__13_ ));
 XNOR2_X1 u_multiplier_STAGE2_E_4_2_pp_4__25_  (.A(u_multiplier_STAGE2_pp_3_c2 ),
    .B(u_multiplier_STAGE2_E_4_2_pp_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp_4_s ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp_4__08_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp_4__10_ ),
    .ZN(u_multiplier_STAGE2_pp_4_c2 ));
 OAI21_X1 u_multiplier_STAGE2_E_4_2_pp_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp_4__12_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp_4__13_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp_4__14_ ),
    .ZN(u_multiplier_STAGE2_pp_4_c1 ));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp_5__18_  (.A(u_multiplier_STAGE2_pp_4_c2 ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_5__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_5__19_  (.A1(u_multiplier_pp_5 [1]),
    .A2(u_multiplier_pp_5 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_5__08_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp_5__20_  (.A(u_multiplier_pp_5 [1]),
    .B(u_multiplier_pp_5 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp_5__09_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_5__21_  (.A1(u_multiplier_pp_5 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp_5__09_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_5__10_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp_5__22_  (.A(u_multiplier_pp_5 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp_5__09_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp_5__11_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_5__23_  (.A1(u_multiplier_pp_5 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp_5__11_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_5__12_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp_5__24_  (.A(u_multiplier_pp_5 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp_5__11_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_5__13_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp_5__25_  (.A(u_multiplier_STAGE2_pp_4_c2 ),
    .B(u_multiplier_STAGE2_E_4_2_pp_5__13_ ),
    .ZN(u_multiplier_STAGE2_pp_5_s ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_5__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp_5__08_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp_5__10_ ),
    .ZN(u_multiplier_STAGE2_pp_5_c2 ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp_5__27_  (.A(u_multiplier_STAGE2_E_4_2_pp_5__12_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp_5__13_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp_5__14_ ),
    .ZN(u_multiplier_STAGE2_pp_5_c1 ));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp_6__18_  (.A(u_multiplier_STAGE2_pp_5_c2 ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_6__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_6__19_  (.A1(u_multiplier_pp_6 [1]),
    .A2(u_multiplier_pp_6 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_6__08_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp_6__20_  (.A(u_multiplier_pp_6 [1]),
    .B(u_multiplier_pp_6 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp_6__09_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_6__21_  (.A1(u_multiplier_pp_6 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp_6__09_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_6__10_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp_6__22_  (.A(u_multiplier_pp_6 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp_6__09_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp_6__11_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_6__23_  (.A1(u_multiplier_pp_6 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp_6__11_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_6__12_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp_6__24_  (.A(u_multiplier_pp_6 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp_6__11_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_6__13_ ));
 XNOR2_X1 u_multiplier_STAGE2_E_4_2_pp_6__25_  (.A(u_multiplier_STAGE2_pp_5_c2 ),
    .B(u_multiplier_STAGE2_E_4_2_pp_6__13_ ),
    .ZN(u_multiplier_STAGE2_pp_6_s ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_6__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp_6__08_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp_6__10_ ),
    .ZN(u_multiplier_STAGE2_pp_6_c2 ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp_6__27_  (.A(u_multiplier_STAGE2_E_4_2_pp_6__12_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp_6__13_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp_6__14_ ),
    .ZN(u_multiplier_STAGE2_pp_6_c1 ));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp_7__18_  (.A(u_multiplier_STAGE2_pp_6_c2 ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_7__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_7__19_  (.A1(u_multiplier_pp_7 [1]),
    .A2(u_multiplier_pp_7 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_7__08_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp_7__20_  (.A(u_multiplier_pp_7 [1]),
    .B(u_multiplier_pp_7 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp_7__09_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_7__21_  (.A1(u_multiplier_pp_7 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp_7__09_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_7__10_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp_7__22_  (.A(u_multiplier_pp_7 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp_7__09_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp_7__11_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_7__23_  (.A1(u_multiplier_pp_7 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp_7__11_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_7__12_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp_7__24_  (.A(u_multiplier_pp_7 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp_7__11_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_7__13_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp_7__25_  (.A(u_multiplier_STAGE2_pp_6_c2 ),
    .B(u_multiplier_STAGE2_E_4_2_pp_7__13_ ),
    .ZN(u_multiplier_STAGE2_pp_7_s ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_7__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp_7__08_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp_7__10_ ),
    .ZN(u_multiplier_STAGE2_pp_7_c2 ));
 OAI21_X1 u_multiplier_STAGE2_E_4_2_pp_7__27_  (.A(u_multiplier_STAGE2_E_4_2_pp_7__12_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp_7__13_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp_7__14_ ),
    .ZN(u_multiplier_STAGE2_pp_7_c1 ));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp_8__18_  (.A(u_multiplier_STAGE2_pp_7_c2 ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_8__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_8__19_  (.A1(u_multiplier_pp_8 [1]),
    .A2(u_multiplier_pp_8 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_8__08_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp_8__20_  (.A(u_multiplier_pp_8 [1]),
    .B(u_multiplier_pp_8 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp_8__09_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_8__21_  (.A1(u_multiplier_pp_8 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp_8__09_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_8__10_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp_8__22_  (.A(u_multiplier_pp_8 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp_8__09_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp_8__11_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_8__23_  (.A1(u_multiplier_pp_8 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp_8__11_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_8__12_ ));
 XNOR2_X1 u_multiplier_STAGE2_E_4_2_pp_8__24_  (.A(u_multiplier_pp_8 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp_8__11_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_8__13_ ));
 XNOR2_X1 u_multiplier_STAGE2_E_4_2_pp_8__25_  (.A(u_multiplier_STAGE2_pp_7_c2 ),
    .B(u_multiplier_STAGE2_E_4_2_pp_8__13_ ),
    .ZN(u_multiplier_STAGE2_pp_8_s ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_8__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp_8__08_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp_8__10_ ),
    .ZN(u_multiplier_STAGE2_pp_8_c2 ));
 OAI21_X1 u_multiplier_STAGE2_E_4_2_pp_8__27_  (.A(u_multiplier_STAGE2_E_4_2_pp_8__12_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp_8__13_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp_8__14_ ),
    .ZN(u_multiplier_STAGE2_pp_8_c1 ));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp_9__18_  (.A(u_multiplier_STAGE2_pp_8_c2 ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_9__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_9__19_  (.A1(u_multiplier_pp_9 [1]),
    .A2(u_multiplier_pp_9 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_9__08_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp_9__20_  (.A(u_multiplier_pp_9 [1]),
    .B(u_multiplier_pp_9 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp_9__09_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_9__21_  (.A1(u_multiplier_pp_9 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp_9__09_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_9__10_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp_9__22_  (.A(u_multiplier_pp_9 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp_9__09_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp_9__11_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_9__23_  (.A1(u_multiplier_pp_9 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp_9__11_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_9__12_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp_9__24_  (.A(u_multiplier_pp_9 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp_9__11_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp_9__13_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp_9__25_  (.A(u_multiplier_STAGE2_pp_8_c2 ),
    .B(u_multiplier_STAGE2_E_4_2_pp_9__13_ ),
    .ZN(u_multiplier_STAGE2_pp_9_s ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp_9__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp_9__08_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp_9__10_ ),
    .ZN(u_multiplier_STAGE2_pp_9_c2 ));
 OAI21_X1 u_multiplier_STAGE2_E_4_2_pp_9__27_  (.A(u_multiplier_STAGE2_E_4_2_pp_9__12_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp_9__13_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp_9__14_ ),
    .ZN(u_multiplier_STAGE2_pp_9_c1 ));
 NAND2_X1 u_multiplier_STAGE2_Final_add_cla1__40_  (.A1(u_multiplier_STAGE2_pp_2_c ),
    .A2(u_multiplier_STAGE2_pp_3_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla1__14_ ));
 AND2_X1 u_multiplier_STAGE2_Final_add_cla1__41_  (.A1(u_multiplier_pp_2 [2]),
    .A2(u_multiplier_STAGE2_pp_2_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla1__15_ ));
 NAND2_X1 u_multiplier_STAGE2_Final_add_cla1__42_  (.A1(u_multiplier_pp_1 [0]),
    .A2(u_multiplier_pp_1 [1]),
    .ZN(u_multiplier_STAGE2_Final_add_cla1__16_ ));
 AND2_X1 u_multiplier_STAGE2_Final_add_cla1__43_  (.A1(net54),
    .A2(u_multiplier_pp_0 ),
    .ZN(u_multiplier_STAGE2_Final_add_cla1__17_ ));
 OR2_X1 u_multiplier_STAGE2_Final_add_cla1__44_  (.A1(net55),
    .A2(u_multiplier_pp_0 ),
    .ZN(u_multiplier_STAGE2_Final_add_cla1__18_ ));
 XNOR2_X1 u_multiplier_STAGE2_Final_add_cla1__45_  (.A(net56),
    .B(u_multiplier_pp_0 ),
    .ZN(u_multiplier_STAGE2_Final_add_cla1__19_ ));
 AOI21_X1 u_multiplier_STAGE2_Final_add_cla1__46_  (.A(u_multiplier_STAGE2_Final_add_cla1__17_ ),
    .B1(u_multiplier_STAGE2_Final_add_cla1__18_ ),
    .B2(net57),
    .ZN(u_multiplier_STAGE2_Final_add_cla1__20_ ));
 NOR2_X1 u_multiplier_STAGE2_Final_add_cla1__47_  (.A1(u_multiplier_pp_1 [0]),
    .A2(u_multiplier_pp_1 [1]),
    .ZN(u_multiplier_STAGE2_Final_add_cla1__21_ ));
 XOR2_X1 u_multiplier_STAGE2_Final_add_cla1__48_  (.A(u_multiplier_pp_1 [0]),
    .B(u_multiplier_pp_1 [1]),
    .Z(u_multiplier_STAGE2_Final_add_cla1__22_ ));
 OAI21_X2 u_multiplier_STAGE2_Final_add_cla1__49_  (.A(u_multiplier_STAGE2_Final_add_cla1__16_ ),
    .B1(u_multiplier_STAGE2_Final_add_cla1__20_ ),
    .B2(u_multiplier_STAGE2_Final_add_cla1__21_ ),
    .ZN(u_multiplier_STAGE2_Final_add_cla1__23_ ));
 OR2_X1 u_multiplier_STAGE2_Final_add_cla1__50_  (.A1(u_multiplier_pp_2 [2]),
    .A2(u_multiplier_STAGE2_pp_2_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla1__24_ ));
 XNOR2_X1 u_multiplier_STAGE2_Final_add_cla1__51_  (.A(u_multiplier_pp_2 [2]),
    .B(u_multiplier_STAGE2_pp_2_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla1__25_ ));
 AOI21_X2 u_multiplier_STAGE2_Final_add_cla1__52_  (.A(u_multiplier_STAGE2_Final_add_cla1__15_ ),
    .B1(u_multiplier_STAGE2_Final_add_cla1__23_ ),
    .B2(u_multiplier_STAGE2_Final_add_cla1__24_ ),
    .ZN(u_multiplier_STAGE2_Final_add_cla1__26_ ));
 NOR2_X1 u_multiplier_STAGE2_Final_add_cla1__53_  (.A1(u_multiplier_STAGE2_pp_2_c ),
    .A2(u_multiplier_STAGE2_pp_3_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla1__27_ ));
 XOR2_X1 u_multiplier_STAGE2_Final_add_cla1__54_  (.A(u_multiplier_STAGE2_pp_2_c ),
    .B(u_multiplier_STAGE2_pp_3_s ),
    .Z(u_multiplier_STAGE2_Final_add_cla1__28_ ));
 OAI21_X2 u_multiplier_STAGE2_Final_add_cla1__55_  (.A(u_multiplier_STAGE2_Final_add_cla1__14_ ),
    .B1(u_multiplier_STAGE2_Final_add_cla1__26_ ),
    .B2(u_multiplier_STAGE2_Final_add_cla1__27_ ),
    .ZN(u_multiplier_STAGE2_Final_add_c1 ));
 XNOR2_X1 u_multiplier_STAGE2_Final_add_cla1__56_  (.A(net58),
    .B(u_multiplier_STAGE2_Final_add_cla1__19_ ),
    .ZN(product[0]));
 XNOR2_X1 u_multiplier_STAGE2_Final_add_cla1__57_  (.A(u_multiplier_STAGE2_Final_add_cla1__20_ ),
    .B(u_multiplier_STAGE2_Final_add_cla1__22_ ),
    .ZN(product[1]));
 XNOR2_X1 u_multiplier_STAGE2_Final_add_cla1__58_  (.A(u_multiplier_STAGE2_Final_add_cla1__23_ ),
    .B(u_multiplier_STAGE2_Final_add_cla1__25_ ),
    .ZN(product[2]));
 XNOR2_X1 u_multiplier_STAGE2_Final_add_cla1__59_  (.A(u_multiplier_STAGE2_Final_add_cla1__26_ ),
    .B(u_multiplier_STAGE2_Final_add_cla1__28_ ),
    .ZN(product[3]));
 NAND2_X1 u_multiplier_STAGE2_Final_add_cla2__40_  (.A1(u_multiplier_STAGE2_pp_6_c1 ),
    .A2(u_multiplier_STAGE2_pp_7_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla2__14_ ));
 AND2_X1 u_multiplier_STAGE2_Final_add_cla2__41_  (.A1(u_multiplier_STAGE2_pp_5_c1 ),
    .A2(u_multiplier_STAGE2_pp_6_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla2__15_ ));
 NAND2_X1 u_multiplier_STAGE2_Final_add_cla2__42_  (.A1(u_multiplier_STAGE2_pp_4_c1 ),
    .A2(u_multiplier_STAGE2_pp_5_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla2__16_ ));
 AND2_X1 u_multiplier_STAGE2_Final_add_cla2__43_  (.A1(u_multiplier_STAGE2_pp_3_c1 ),
    .A2(u_multiplier_STAGE2_pp_4_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla2__17_ ));
 OR2_X1 u_multiplier_STAGE2_Final_add_cla2__44_  (.A1(u_multiplier_STAGE2_pp_3_c1 ),
    .A2(u_multiplier_STAGE2_pp_4_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla2__18_ ));
 XNOR2_X1 u_multiplier_STAGE2_Final_add_cla2__45_  (.A(u_multiplier_STAGE2_pp_3_c1 ),
    .B(u_multiplier_STAGE2_pp_4_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla2__19_ ));
 AOI21_X2 u_multiplier_STAGE2_Final_add_cla2__46_  (.A(u_multiplier_STAGE2_Final_add_cla2__17_ ),
    .B1(u_multiplier_STAGE2_Final_add_cla2__18_ ),
    .B2(u_multiplier_STAGE2_Final_add_c1 ),
    .ZN(u_multiplier_STAGE2_Final_add_cla2__20_ ));
 NOR2_X1 u_multiplier_STAGE2_Final_add_cla2__47_  (.A1(u_multiplier_STAGE2_pp_4_c1 ),
    .A2(u_multiplier_STAGE2_pp_5_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla2__21_ ));
 XOR2_X1 u_multiplier_STAGE2_Final_add_cla2__48_  (.A(u_multiplier_STAGE2_pp_4_c1 ),
    .B(u_multiplier_STAGE2_pp_5_s ),
    .Z(u_multiplier_STAGE2_Final_add_cla2__22_ ));
 OAI21_X2 u_multiplier_STAGE2_Final_add_cla2__49_  (.A(u_multiplier_STAGE2_Final_add_cla2__16_ ),
    .B1(u_multiplier_STAGE2_Final_add_cla2__20_ ),
    .B2(u_multiplier_STAGE2_Final_add_cla2__21_ ),
    .ZN(u_multiplier_STAGE2_Final_add_cla2__23_ ));
 OR2_X1 u_multiplier_STAGE2_Final_add_cla2__50_  (.A1(u_multiplier_STAGE2_pp_5_c1 ),
    .A2(u_multiplier_STAGE2_pp_6_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla2__24_ ));
 XNOR2_X1 u_multiplier_STAGE2_Final_add_cla2__51_  (.A(u_multiplier_STAGE2_pp_5_c1 ),
    .B(u_multiplier_STAGE2_pp_6_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla2__25_ ));
 AOI21_X2 u_multiplier_STAGE2_Final_add_cla2__52_  (.A(u_multiplier_STAGE2_Final_add_cla2__15_ ),
    .B1(u_multiplier_STAGE2_Final_add_cla2__23_ ),
    .B2(u_multiplier_STAGE2_Final_add_cla2__24_ ),
    .ZN(u_multiplier_STAGE2_Final_add_cla2__26_ ));
 NOR2_X1 u_multiplier_STAGE2_Final_add_cla2__53_  (.A1(u_multiplier_STAGE2_pp_6_c1 ),
    .A2(u_multiplier_STAGE2_pp_7_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla2__27_ ));
 XOR2_X1 u_multiplier_STAGE2_Final_add_cla2__54_  (.A(u_multiplier_STAGE2_pp_6_c1 ),
    .B(u_multiplier_STAGE2_pp_7_s ),
    .Z(u_multiplier_STAGE2_Final_add_cla2__28_ ));
 OAI21_X2 u_multiplier_STAGE2_Final_add_cla2__55_  (.A(u_multiplier_STAGE2_Final_add_cla2__14_ ),
    .B1(u_multiplier_STAGE2_Final_add_cla2__26_ ),
    .B2(u_multiplier_STAGE2_Final_add_cla2__27_ ),
    .ZN(u_multiplier_STAGE2_Final_add_c2 ));
 XNOR2_X1 u_multiplier_STAGE2_Final_add_cla2__56_  (.A(u_multiplier_STAGE2_Final_add_c1 ),
    .B(u_multiplier_STAGE2_Final_add_cla2__19_ ),
    .ZN(product[4]));
 XNOR2_X1 u_multiplier_STAGE2_Final_add_cla2__57_  (.A(u_multiplier_STAGE2_Final_add_cla2__20_ ),
    .B(u_multiplier_STAGE2_Final_add_cla2__22_ ),
    .ZN(product[5]));
 XNOR2_X1 u_multiplier_STAGE2_Final_add_cla2__58_  (.A(u_multiplier_STAGE2_Final_add_cla2__23_ ),
    .B(u_multiplier_STAGE2_Final_add_cla2__25_ ),
    .ZN(product[6]));
 XNOR2_X1 u_multiplier_STAGE2_Final_add_cla2__59_  (.A(u_multiplier_STAGE2_Final_add_cla2__26_ ),
    .B(u_multiplier_STAGE2_Final_add_cla2__28_ ),
    .ZN(product[7]));
 NAND2_X1 u_multiplier_STAGE2_Final_add_cla3__40_  (.A1(u_multiplier_STAGE2_pp_10_c1 ),
    .A2(u_multiplier_STAGE2_pp_11_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla3__14_ ));
 AND2_X1 u_multiplier_STAGE2_Final_add_cla3__41_  (.A1(u_multiplier_STAGE2_pp_9_c1 ),
    .A2(u_multiplier_STAGE2_pp_10_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla3__15_ ));
 NAND2_X1 u_multiplier_STAGE2_Final_add_cla3__42_  (.A1(u_multiplier_STAGE2_pp_8_c1 ),
    .A2(u_multiplier_STAGE2_pp_9_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla3__16_ ));
 AND2_X1 u_multiplier_STAGE2_Final_add_cla3__43_  (.A1(u_multiplier_STAGE2_pp_7_c1 ),
    .A2(u_multiplier_STAGE2_pp_8_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla3__17_ ));
 OR2_X1 u_multiplier_STAGE2_Final_add_cla3__44_  (.A1(u_multiplier_STAGE2_pp_7_c1 ),
    .A2(u_multiplier_STAGE2_pp_8_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla3__18_ ));
 XNOR2_X1 u_multiplier_STAGE2_Final_add_cla3__45_  (.A(u_multiplier_STAGE2_pp_7_c1 ),
    .B(u_multiplier_STAGE2_pp_8_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla3__19_ ));
 AOI21_X2 u_multiplier_STAGE2_Final_add_cla3__46_  (.A(u_multiplier_STAGE2_Final_add_cla3__17_ ),
    .B1(u_multiplier_STAGE2_Final_add_cla3__18_ ),
    .B2(u_multiplier_STAGE2_Final_add_c2 ),
    .ZN(u_multiplier_STAGE2_Final_add_cla3__20_ ));
 NOR2_X1 u_multiplier_STAGE2_Final_add_cla3__47_  (.A1(u_multiplier_STAGE2_pp_8_c1 ),
    .A2(u_multiplier_STAGE2_pp_9_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla3__21_ ));
 XOR2_X1 u_multiplier_STAGE2_Final_add_cla3__48_  (.A(u_multiplier_STAGE2_pp_8_c1 ),
    .B(u_multiplier_STAGE2_pp_9_s ),
    .Z(u_multiplier_STAGE2_Final_add_cla3__22_ ));
 OAI21_X2 u_multiplier_STAGE2_Final_add_cla3__49_  (.A(u_multiplier_STAGE2_Final_add_cla3__16_ ),
    .B1(u_multiplier_STAGE2_Final_add_cla3__20_ ),
    .B2(u_multiplier_STAGE2_Final_add_cla3__21_ ),
    .ZN(u_multiplier_STAGE2_Final_add_cla3__23_ ));
 OR2_X1 u_multiplier_STAGE2_Final_add_cla3__50_  (.A1(u_multiplier_STAGE2_pp_9_c1 ),
    .A2(u_multiplier_STAGE2_pp_10_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla3__24_ ));
 XNOR2_X1 u_multiplier_STAGE2_Final_add_cla3__51_  (.A(u_multiplier_STAGE2_pp_9_c1 ),
    .B(u_multiplier_STAGE2_pp_10_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla3__25_ ));
 AOI21_X2 u_multiplier_STAGE2_Final_add_cla3__52_  (.A(u_multiplier_STAGE2_Final_add_cla3__15_ ),
    .B1(u_multiplier_STAGE2_Final_add_cla3__23_ ),
    .B2(u_multiplier_STAGE2_Final_add_cla3__24_ ),
    .ZN(u_multiplier_STAGE2_Final_add_cla3__26_ ));
 NOR2_X1 u_multiplier_STAGE2_Final_add_cla3__53_  (.A1(u_multiplier_STAGE2_pp_10_c1 ),
    .A2(u_multiplier_STAGE2_pp_11_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla3__27_ ));
 XOR2_X1 u_multiplier_STAGE2_Final_add_cla3__54_  (.A(u_multiplier_STAGE2_pp_10_c1 ),
    .B(u_multiplier_STAGE2_pp_11_s ),
    .Z(u_multiplier_STAGE2_Final_add_cla3__28_ ));
 OAI21_X2 u_multiplier_STAGE2_Final_add_cla3__55_  (.A(u_multiplier_STAGE2_Final_add_cla3__14_ ),
    .B1(u_multiplier_STAGE2_Final_add_cla3__26_ ),
    .B2(u_multiplier_STAGE2_Final_add_cla3__27_ ),
    .ZN(u_multiplier_STAGE2_Final_add_c3 ));
 XNOR2_X2 u_multiplier_STAGE2_Final_add_cla3__56_  (.A(u_multiplier_STAGE2_Final_add_c2 ),
    .B(u_multiplier_STAGE2_Final_add_cla3__19_ ),
    .ZN(product[8]));
 XNOR2_X1 u_multiplier_STAGE2_Final_add_cla3__57_  (.A(u_multiplier_STAGE2_Final_add_cla3__20_ ),
    .B(u_multiplier_STAGE2_Final_add_cla3__22_ ),
    .ZN(product[9]));
 XNOR2_X1 u_multiplier_STAGE2_Final_add_cla3__58_  (.A(u_multiplier_STAGE2_Final_add_cla3__23_ ),
    .B(u_multiplier_STAGE2_Final_add_cla3__25_ ),
    .ZN(product[10]));
 XNOR2_X1 u_multiplier_STAGE2_Final_add_cla3__59_  (.A(u_multiplier_STAGE2_Final_add_cla3__26_ ),
    .B(u_multiplier_STAGE2_Final_add_cla3__28_ ),
    .ZN(product[11]));
 NAND2_X1 u_multiplier_STAGE2_Final_add_cla4__40_  (.A1(net59),
    .A2(net60),
    .ZN(u_multiplier_STAGE2_Final_add_cla4__14_ ));
 AND2_X1 u_multiplier_STAGE2_Final_add_cla4__41_  (.A1(u_multiplier_STAGE2_pp_13_c ),
    .A2(u_multiplier_pp_14 ),
    .ZN(u_multiplier_STAGE2_Final_add_cla4__15_ ));
 NAND2_X1 u_multiplier_STAGE2_Final_add_cla4__42_  (.A1(u_multiplier_STAGE2_pp_12_c1 ),
    .A2(u_multiplier_STAGE2_pp_13_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla4__16_ ));
 AND2_X1 u_multiplier_STAGE2_Final_add_cla4__43_  (.A1(u_multiplier_STAGE2_pp_11_c1 ),
    .A2(u_multiplier_STAGE2_pp_12_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla4__17_ ));
 OR2_X1 u_multiplier_STAGE2_Final_add_cla4__44_  (.A1(u_multiplier_STAGE2_pp_11_c1 ),
    .A2(u_multiplier_STAGE2_pp_12_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla4__18_ ));
 XNOR2_X1 u_multiplier_STAGE2_Final_add_cla4__45_  (.A(u_multiplier_STAGE2_pp_11_c1 ),
    .B(u_multiplier_STAGE2_pp_12_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla4__19_ ));
 AOI21_X2 u_multiplier_STAGE2_Final_add_cla4__46_  (.A(u_multiplier_STAGE2_Final_add_cla4__17_ ),
    .B1(u_multiplier_STAGE2_Final_add_cla4__18_ ),
    .B2(u_multiplier_STAGE2_Final_add_c3 ),
    .ZN(u_multiplier_STAGE2_Final_add_cla4__20_ ));
 NOR2_X1 u_multiplier_STAGE2_Final_add_cla4__47_  (.A1(u_multiplier_STAGE2_pp_12_c1 ),
    .A2(u_multiplier_STAGE2_pp_13_s ),
    .ZN(u_multiplier_STAGE2_Final_add_cla4__21_ ));
 XOR2_X1 u_multiplier_STAGE2_Final_add_cla4__48_  (.A(u_multiplier_STAGE2_pp_12_c1 ),
    .B(u_multiplier_STAGE2_pp_13_s ),
    .Z(u_multiplier_STAGE2_Final_add_cla4__22_ ));
 OAI21_X2 u_multiplier_STAGE2_Final_add_cla4__49_  (.A(u_multiplier_STAGE2_Final_add_cla4__16_ ),
    .B1(u_multiplier_STAGE2_Final_add_cla4__20_ ),
    .B2(u_multiplier_STAGE2_Final_add_cla4__21_ ),
    .ZN(u_multiplier_STAGE2_Final_add_cla4__23_ ));
 OR2_X1 u_multiplier_STAGE2_Final_add_cla4__50_  (.A1(u_multiplier_STAGE2_pp_13_c ),
    .A2(u_multiplier_pp_14 ),
    .ZN(u_multiplier_STAGE2_Final_add_cla4__24_ ));
 XNOR2_X1 u_multiplier_STAGE2_Final_add_cla4__51_  (.A(u_multiplier_STAGE2_pp_13_c ),
    .B(u_multiplier_pp_14 ),
    .ZN(u_multiplier_STAGE2_Final_add_cla4__25_ ));
 AOI21_X1 u_multiplier_STAGE2_Final_add_cla4__52_  (.A(u_multiplier_STAGE2_Final_add_cla4__15_ ),
    .B1(u_multiplier_STAGE2_Final_add_cla4__23_ ),
    .B2(u_multiplier_STAGE2_Final_add_cla4__24_ ),
    .ZN(u_multiplier_STAGE2_Final_add_cla4__26_ ));
 NOR2_X1 u_multiplier_STAGE2_Final_add_cla4__53_  (.A1(net61),
    .A2(net62),
    .ZN(u_multiplier_STAGE2_Final_add_cla4__27_ ));
 XOR2_X1 u_multiplier_STAGE2_Final_add_cla4__54_  (.A(net63),
    .B(net64),
    .Z(u_multiplier_STAGE2_Final_add_cla4__28_ ));
 OAI21_X1 u_multiplier_STAGE2_Final_add_cla4__55_  (.A(u_multiplier_STAGE2_Final_add_cla4__14_ ),
    .B1(u_multiplier_STAGE2_Final_add_cla4__26_ ),
    .B2(u_multiplier_STAGE2_Final_add_cla4__27_ ),
    .ZN(u_multiplier_STAGE2_Final_add_Cout ));
 XNOR2_X1 u_multiplier_STAGE2_Final_add_cla4__56_  (.A(u_multiplier_STAGE2_Final_add_c3 ),
    .B(u_multiplier_STAGE2_Final_add_cla4__19_ ),
    .ZN(product[12]));
 XNOR2_X1 u_multiplier_STAGE2_Final_add_cla4__57_  (.A(u_multiplier_STAGE2_Final_add_cla4__20_ ),
    .B(u_multiplier_STAGE2_Final_add_cla4__22_ ),
    .ZN(product[13]));
 XNOR2_X2 u_multiplier_STAGE2_Final_add_cla4__58_  (.A(u_multiplier_STAGE2_Final_add_cla4__23_ ),
    .B(u_multiplier_STAGE2_Final_add_cla4__25_ ),
    .ZN(product[14]));
 XNOR2_X1 u_multiplier_STAGE2_Final_add_cla4__59_  (.A(u_multiplier_STAGE2_Final_add_cla4__26_ ),
    .B(u_multiplier_STAGE2_Final_add_cla4__28_ ),
    .ZN(u_multiplier_approx [15]));
 INV_X1 u_multiplier_STAGE2_Full_adder_pp_13__12_  (.A(u_multiplier_STAGE2_pp_12_c2 ),
    .ZN(u_multiplier_STAGE2_Full_adder_pp_13__05_ ));
 NAND3_X1 u_multiplier_STAGE2_Full_adder_pp_13__13_  (.A1(u_multiplier_pp_13 [1]),
    .A2(u_multiplier_pp_13 [0]),
    .A3(u_multiplier_STAGE2_pp_12_c2 ),
    .ZN(u_multiplier_STAGE2_Full_adder_pp_13__06_ ));
 NOR2_X1 u_multiplier_STAGE2_Full_adder_pp_13__14_  (.A1(u_multiplier_pp_13 [1]),
    .A2(u_multiplier_pp_13 [0]),
    .ZN(u_multiplier_STAGE2_Full_adder_pp_13__07_ ));
 AOI21_X1 u_multiplier_STAGE2_Full_adder_pp_13__15_  (.A(u_multiplier_STAGE2_pp_12_c2 ),
    .B1(u_multiplier_pp_13 [0]),
    .B2(u_multiplier_pp_13 [1]),
    .ZN(u_multiplier_STAGE2_Full_adder_pp_13__08_ ));
 NOR2_X1 u_multiplier_STAGE2_Full_adder_pp_13__16_  (.A1(u_multiplier_STAGE2_Full_adder_pp_13__07_ ),
    .A2(u_multiplier_STAGE2_Full_adder_pp_13__08_ ),
    .ZN(u_multiplier_STAGE2_pp_13_c ));
 AOI22_X2 u_multiplier_STAGE2_Full_adder_pp_13__17_  (.A1(u_multiplier_STAGE2_Full_adder_pp_13__05_ ),
    .A2(u_multiplier_STAGE2_Full_adder_pp_13__07_ ),
    .B1(u_multiplier_STAGE2_pp_13_c ),
    .B2(u_multiplier_STAGE2_Full_adder_pp_13__06_ ),
    .ZN(u_multiplier_STAGE2_pp_13_s ));
 AND2_X1 u_multiplier_STAGE2_Half_adder_pp_2__4_  (.A1(u_multiplier_pp_2 [1]),
    .A2(u_multiplier_pp_2 [0]),
    .ZN(u_multiplier_STAGE2_pp_2_c ));
 XOR2_X2 u_multiplier_STAGE2_Half_adder_pp_2__5_  (.A(u_multiplier_pp_2 [1]),
    .B(u_multiplier_pp_2 [0]),
    .Z(u_multiplier_STAGE2_pp_2_s ));
 XOR2_X1 u_multiplier__3_  (.A(net119),
    .B(data_in_reg[7]),
    .Z(product[15]));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_2_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_2_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_2_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_2_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_2_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_2_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_2_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_2_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_2_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_2_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_2_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_2_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_2_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_2_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_2_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_2_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_2_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_2_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_2_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_2_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_2_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_2_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_2_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_2_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_2_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_2_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_2_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_2_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_2_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_2_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_2_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_2_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_2_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_2_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_2_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_2_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_2_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_2_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_2_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_2_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_2_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_2_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_2_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_2_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_2_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_2_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_2_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_2_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_2_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_2_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_2_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_2_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_2_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_2_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_2_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_2_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_2_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_2_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_2_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_2_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_2_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_2_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_2_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_2_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_2_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_2_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_2_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_2_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_2_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_2_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_2_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_2_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_2_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_2_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_1_Left_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_1_Left_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_1_Left_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_1_Left_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_1_Left_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_1_Left_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_1_Left_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_1_Left_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_1_Left_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_1_Left_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_1_Left_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_1_Left_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_1_Left_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_1_Left_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_1_Left_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_1_Left_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_1_Left_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_1_Left_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_1_Left_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_1_Left_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_1_Left_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_1_Left_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_1_Left_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_1_Left_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_1_Left_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_1_Left_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_1_Left_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_1_Left_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_1_Left_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_1_Left_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_1_Left_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_1_Left_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_1_Left_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_1_Left_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_1_Left_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_1_Left_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_1_Left_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_1_Left_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_1_Left_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_1_Left_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_1_Left_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_1_Left_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_1_Left_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_1_Left_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_1_Left_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_1_Left_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_1_Left_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_1_Left_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_1_Left_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_1_Left_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_1_Left_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_1_Left_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_1_Left_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_1_Left_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_1_Left_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_1_Left_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_1_Left_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_1_Left_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_1_Left_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_1_Left_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_1_Left_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_1_Left_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_1_Left_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_1_Left_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_1_Left_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_1_Left_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_1_Left_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_1_Left_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_1_Left_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_1_Left_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_1_Left_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_1_Left_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_1_Left_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Left_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Left_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Left_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Left_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Left_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Left_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Left_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Left_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Left_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_1_Left_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_2_Left_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_2_Left_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_2_Left_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_2_Left_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_2_Left_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_2_Left_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_2_Left_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_2_Left_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_2_Left_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_2_Left_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_2_Left_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_2_Left_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_2_Left_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_2_Left_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_2_Left_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_2_Left_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_2_Left_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_2_Left_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_2_Left_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_2_Left_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_2_Left_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_2_Left_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_2_Left_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_2_Left_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_2_Left_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_2_Left_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_2_Left_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_2_Left_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_2_Left_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_2_Left_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_2_Left_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_2_Left_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_2_Left_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_2_Left_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_2_Left_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_2_Left_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_2_Left_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_2_Left_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_2_Left_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_2_Left_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_2_Left_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_2_Left_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_2_Left_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_2_Left_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_2_Left_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_2_Left_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_2_Left_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_2_Left_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_2_Left_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_2_Left_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_2_Left_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_2_Left_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_2_Left_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_2_Left_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_2_Left_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_2_Left_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_2_Left_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_2_Left_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_2_Left_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_2_Left_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_2_Left_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_2_Left_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_2_Left_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_2_Left_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_2_Left_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_2_Left_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_2_Left_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_2_Left_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_2_Left_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_2_Left_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_2_Left_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_2_Left_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_2_Left_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_2_Left_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_1_Right_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_1_Right_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_1_Right_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_1_Right_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_1_Right_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_1_Right_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_1_Right_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_1_Right_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_1_Right_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_1_Right_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_1_Right_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_1_Right_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_1_Right_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_1_Right_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_1_Right_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_1_Right_265 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_1_Right_266 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_1_Right_267 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_1_Right_268 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_1_Right_269 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_1_Right_270 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_1_Right_271 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_1_Right_272 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_1_Right_273 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_1_Right_274 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_1_Right_275 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_1_Right_276 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_1_Right_277 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_1_Right_278 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_1_Right_279 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_1_Right_280 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_1_Right_281 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_1_Right_282 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_1_Right_283 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_1_Right_284 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_1_Right_285 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_1_Right_286 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_1_Right_287 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_1_Right_288 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_1_Right_289 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_1_Right_290 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_1_Right_291 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_1_Right_292 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_1_Right_293 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_1_Right_294 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_1_Right_295 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_1_Right_296 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_1_Right_297 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_1_Right_298 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_1_Right_299 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_1_Right_300 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_1_Right_301 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_1_Right_302 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_1_Right_303 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_1_Right_304 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_1_Right_305 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_1_Right_306 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_1_Right_307 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_1_Right_308 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_1_Right_309 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_1_Right_310 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_1_Right_311 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_1_Right_312 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_1_Right_313 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_1_Right_314 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_1_Right_315 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_1_Right_316 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_1_Right_317 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_1_Right_318 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_1_Right_319 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_1_Right_320 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_1_Right_321 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_1_Right_322 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_1_Right_323 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_324 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_325 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_326 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_79_327 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_328 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_329 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_330 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_331 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_87_332 ();
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_5__18__46  (.Z(net46));
 LOGIC0_X1 u_multiplier_STAGE2_E_4_2_pp_3__18__52  (.Z(net52));
 CLKBUF_X1 hold65 (.A(net120),
    .Z(net65));
 BUF_X2 input1 (.A(data_in[0]),
    .Z(net1));
 BUF_X1 input2 (.A(data_in[1]),
    .Z(net2));
 BUF_X1 input3 (.A(data_in[2]),
    .Z(net3));
 BUF_X1 input4 (.A(data_in[3]),
    .Z(net4));
 BUF_X1 input5 (.A(data_in[4]),
    .Z(net5));
 BUF_X1 input6 (.A(data_in[5]),
    .Z(net6));
 BUF_X2 input7 (.A(data_in[6]),
    .Z(net7));
 BUF_X1 input8 (.A(data_in[7]),
    .Z(net8));
 BUF_X2 input9 (.A(init_enable),
    .Z(net9));
 BUF_X2 input10 (.A(pe_ce),
    .Z(net10));
 BUF_X8 input11 (.A(rst_n),
    .Z(net11));
 BUF_X1 output12 (.A(net12),
    .Z(curr_state[1]));
 BUF_X1 output13 (.A(net13),
    .Z(data_out[0]));
 BUF_X1 output14 (.A(net14),
    .Z(data_out[10]));
 BUF_X1 output15 (.A(net15),
    .Z(data_out[11]));
 BUF_X1 output16 (.A(net16),
    .Z(data_out[12]));
 BUF_X1 output17 (.A(net17),
    .Z(data_out[13]));
 BUF_X1 output18 (.A(net18),
    .Z(data_out[14]));
 BUF_X1 output19 (.A(net19),
    .Z(data_out[15]));
 BUF_X1 output20 (.A(net20),
    .Z(data_out[1]));
 BUF_X1 output21 (.A(net21),
    .Z(data_out[2]));
 BUF_X1 output22 (.A(net22),
    .Z(data_out[3]));
 BUF_X1 output23 (.A(net23),
    .Z(data_out[4]));
 BUF_X1 output24 (.A(net24),
    .Z(data_out[5]));
 BUF_X1 output25 (.A(net25),
    .Z(data_out[6]));
 BUF_X1 output26 (.A(net26),
    .Z(data_out[7]));
 BUF_X1 output27 (.A(net27),
    .Z(data_out[8]));
 BUF_X1 output28 (.A(net28),
    .Z(data_out[9]));
 BUF_X1 output29 (.A(net29),
    .Z(valid_reg_out));
 LOGIC0_X1 u_multiplier_STAGE1__135__30  (.Z(net30));
 LOGIC0_X1 u_multiplier_STAGE1__136__31  (.Z(net31));
 LOGIC0_X1 u_multiplier_STAGE1__138__32  (.Z(net32));
 LOGIC0_X1 u_multiplier_STAGE1__140__33  (.Z(net33));
 LOGIC0_X1 u_multiplier_STAGE1__141__34  (.Z(net34));
 LOGIC0_X1 u_multiplier_STAGE1__142__35  (.Z(net35));
 LOGIC0_X1 u_multiplier_STAGE1__143__36  (.Z(net36));
 LOGIC0_X1 u_multiplier_STAGE1__143__37  (.Z(net37));
 LOGIC0_X1 u_multiplier_STAGE1__156__38  (.Z(net38));
 LOGIC0_X1 u_multiplier_STAGE1__163__39  (.Z(net39));
 LOGIC0_X1 u_multiplier_STAGE1__164__40  (.Z(net40));
 LOGIC0_X1 u_multiplier_STAGE1__170__41  (.Z(net41));
 LOGIC0_X1 u_multiplier_STAGE1__171__42  (.Z(net42));
 LOGIC0_X1 u_multiplier_STAGE1__176__43  (.Z(net43));
 LOGIC0_X1 u_multiplier_STAGE1__177__44  (.Z(net44));
 LOGIC0_X1 u_multiplier_STAGE1__181__45  (.Z(net45));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_5__25__47  (.Z(net47));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_7_2__18__48  (.Z(net48));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_7_2__25__49  (.Z(net49));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_8_2__18__50  (.Z(net50));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_8_2__25__51  (.Z(net51));
 LOGIC0_X1 u_multiplier_STAGE2_E_4_2_pp_3__25__53  (.Z(net53));
 LOGIC0_X1 u_multiplier_STAGE2_Final_add_cla1__43__54  (.Z(net54));
 LOGIC0_X1 u_multiplier_STAGE2_Final_add_cla1__44__55  (.Z(net55));
 LOGIC0_X1 u_multiplier_STAGE2_Final_add_cla1__45__56  (.Z(net56));
 LOGIC0_X1 u_multiplier_STAGE2_Final_add_cla1__46__57  (.Z(net57));
 LOGIC0_X1 u_multiplier_STAGE2_Final_add_cla1__56__58  (.Z(net58));
 LOGIC0_X1 u_multiplier_STAGE2_Final_add_cla4__40__59  (.Z(net59));
 LOGIC0_X1 u_multiplier_STAGE2_Final_add_cla4__40__60  (.Z(net60));
 LOGIC0_X1 u_multiplier_STAGE2_Final_add_cla4__53__61  (.Z(net61));
 LOGIC0_X1 u_multiplier_STAGE2_Final_add_cla4__53__62  (.Z(net62));
 LOGIC0_X1 u_multiplier_STAGE2_Final_add_cla4__54__63  (.Z(net63));
 LOGIC0_X1 u_multiplier_STAGE2_Final_add_cla4__54__64  (.Z(net64));
 CLKBUF_X1 hold66 (.A(_008_),
    .Z(net66));
 CLKBUF_X1 hold67 (.A(net118),
    .Z(net67));
 CLKBUF_X1 hold68 (.A(_007_),
    .Z(net68));
 CLKBUF_X1 hold69 (.A(net122),
    .Z(net69));
 CLKBUF_X1 hold70 (.A(_047_),
    .Z(net70));
 CLKBUF_X1 hold71 (.A(net95),
    .Z(net71));
 CLKBUF_X1 hold72 (.A(net92),
    .Z(net72));
 CLKBUF_X1 hold73 (.A(net98),
    .Z(net73));
 CLKBUF_X1 hold74 (.A(net101),
    .Z(net74));
 CLKBUF_X1 hold75 (.A(net104),
    .Z(net75));
 CLKBUF_X1 hold76 (.A(net112),
    .Z(net76));
 CLKBUF_X1 hold77 (.A(net110),
    .Z(net77));
 CLKBUF_X1 hold78 (.A(net114),
    .Z(net78));
 CLKBUF_X1 hold79 (.A(net88),
    .Z(net79));
 CLKBUF_X1 hold80 (.A(net115),
    .Z(net80));
 CLKBUF_X1 hold81 (.A(net121),
    .Z(net81));
 CLKBUF_X1 hold82 (.A(net125),
    .Z(net82));
 CLKBUF_X1 hold83 (.A(net127),
    .Z(net83));
 CLKBUF_X1 hold84 (.A(net126),
    .Z(net84));
 CLKBUF_X1 hold85 (.A(net123),
    .Z(net85));
 CLKBUF_X1 hold86 (.A(net124),
    .Z(net86));
 CLKBUF_X1 hold87 (.A(net128),
    .Z(net87));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 CLKBUF_X3 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 CLKBUF_X3 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 CLKBUF_X3 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 INV_X4 clkload0 (.A(clknet_2_0__leaf_clk));
 INV_X2 clkload1 (.A(clknet_2_1__leaf_clk));
 INV_X2 clkload2 (.A(clknet_2_3__leaf_clk));
 CLKBUF_X1 hold1 (.A(_262_),
    .Z(net88));
 CLKBUF_X1 hold2 (.A(_115_),
    .Z(net89));
 CLKBUF_X1 hold3 (.A(_006_),
    .Z(net90));
 CLKBUF_X1 hold4 (.A(net129),
    .Z(net91));
 CLKBUF_X1 hold5 (.A(_269_),
    .Z(net92));
 CLKBUF_X1 hold6 (.A(net72),
    .Z(net93));
 CLKBUF_X1 hold7 (.A(_037_),
    .Z(net94));
 CLKBUF_X1 hold8 (.A(_268_),
    .Z(net95));
 CLKBUF_X1 hold9 (.A(net71),
    .Z(net96));
 CLKBUF_X1 hold10 (.A(_036_),
    .Z(net97));
 CLKBUF_X1 hold11 (.A(_266_),
    .Z(net98));
 CLKBUF_X1 hold12 (.A(net73),
    .Z(net99));
 CLKBUF_X1 hold13 (.A(_034_),
    .Z(net100));
 CLKBUF_X1 hold14 (.A(_265_),
    .Z(net101));
 CLKBUF_X1 hold15 (.A(net74),
    .Z(net102));
 CLKBUF_X1 hold16 (.A(_009_),
    .Z(net103));
 CLKBUF_X1 hold17 (.A(_267_),
    .Z(net104));
 CLKBUF_X1 hold18 (.A(net75),
    .Z(net105));
 CLKBUF_X1 hold19 (.A(_035_),
    .Z(net106));
 CLKBUF_X1 hold20 (.A(curr_state[0]),
    .Z(net107));
 CLKBUF_X1 hold21 (.A(_102_),
    .Z(net108));
 CLKBUF_X1 hold22 (.A(_049_),
    .Z(net109));
 CLKBUF_X1 hold23 (.A(addr_ptr[1]),
    .Z(net110));
 CLKBUF_X1 hold24 (.A(net77),
    .Z(net111));
 CLKBUF_X1 hold25 (.A(addr_ptr[3]),
    .Z(net112));
 CLKBUF_X1 hold26 (.A(net76),
    .Z(net113));
 CLKBUF_X1 hold27 (.A(addr_ptr[2]),
    .Z(net114));
 CLKBUF_X1 hold28 (.A(addr_ptr[0]),
    .Z(net115));
 CLKBUF_X1 hold29 (.A(curr_state[2]),
    .Z(net116));
 CLKBUF_X1 hold30 (.A(_048_),
    .Z(net117));
 CLKBUF_X1 hold31 (.A(_263_),
    .Z(net118));
 CLKBUF_X1 hold32 (.A(sram_rdata_reg[7]),
    .Z(net119));
 CLKBUF_X1 hold33 (.A(_264_),
    .Z(net120));
 CLKBUF_X1 hold34 (.A(data_in_reg[7]),
    .Z(net121));
 CLKBUF_X1 hold35 (.A(_226_),
    .Z(net122));
 CLKBUF_X1 hold36 (.A(data_in_reg[0]),
    .Z(net123));
 CLKBUF_X1 hold37 (.A(data_in_reg[1]),
    .Z(net124));
 CLKBUF_X1 hold38 (.A(data_in_reg[6]),
    .Z(net125));
 CLKBUF_X1 hold39 (.A(data_in_reg[4]),
    .Z(net126));
 CLKBUF_X1 hold40 (.A(data_in_reg[5]),
    .Z(net127));
 CLKBUF_X1 hold41 (.A(data_in_reg[2]),
    .Z(net128));
 CLKBUF_X1 hold42 (.A(data_in_reg[3]),
    .Z(net129));
 FILLCELL_X4 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_8 ();
 FILLCELL_X16 FILLER_0_40 ();
 FILLCELL_X8 FILLER_0_56 ();
 FILLCELL_X4 FILLER_0_64 ();
 FILLCELL_X32 FILLER_0_71 ();
 FILLCELL_X32 FILLER_0_103 ();
 FILLCELL_X16 FILLER_0_135 ();
 FILLCELL_X8 FILLER_0_151 ();
 FILLCELL_X2 FILLER_0_159 ();
 FILLCELL_X1 FILLER_0_161 ();
 FILLCELL_X32 FILLER_0_165 ();
 FILLCELL_X32 FILLER_0_197 ();
 FILLCELL_X16 FILLER_0_229 ();
 FILLCELL_X8 FILLER_0_245 ();
 FILLCELL_X2 FILLER_0_253 ();
 FILLCELL_X1 FILLER_0_255 ();
 FILLCELL_X4 FILLER_0_259 ();
 FILLCELL_X1 FILLER_0_263 ();
 FILLCELL_X32 FILLER_0_268 ();
 FILLCELL_X16 FILLER_0_300 ();
 FILLCELL_X8 FILLER_0_316 ();
 FILLCELL_X4 FILLER_0_324 ();
 FILLCELL_X2 FILLER_0_328 ();
 FILLCELL_X8 FILLER_0_333 ();
 FILLCELL_X4 FILLER_0_341 ();
 FILLCELL_X32 FILLER_0_349 ();
 FILLCELL_X32 FILLER_0_381 ();
 FILLCELL_X16 FILLER_0_413 ();
 FILLCELL_X8 FILLER_0_429 ();
 FILLCELL_X2 FILLER_0_437 ();
 FILLCELL_X32 FILLER_0_442 ();
 FILLCELL_X32 FILLER_0_474 ();
 FILLCELL_X16 FILLER_0_506 ();
 FILLCELL_X8 FILLER_0_522 ();
 FILLCELL_X4 FILLER_0_530 ();
 FILLCELL_X32 FILLER_0_537 ();
 FILLCELL_X32 FILLER_0_569 ();
 FILLCELL_X16 FILLER_0_601 ();
 FILLCELL_X8 FILLER_0_617 ();
 FILLCELL_X4 FILLER_0_625 ();
 FILLCELL_X2 FILLER_0_629 ();
 FILLCELL_X4 FILLER_0_632 ();
 FILLCELL_X8 FILLER_0_639 ();
 FILLCELL_X4 FILLER_0_647 ();
 FILLCELL_X1 FILLER_0_651 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X16 FILLER_1_225 ();
 FILLCELL_X8 FILLER_1_241 ();
 FILLCELL_X4 FILLER_1_249 ();
 FILLCELL_X1 FILLER_1_253 ();
 FILLCELL_X4 FILLER_1_258 ();
 FILLCELL_X32 FILLER_1_281 ();
 FILLCELL_X1 FILLER_1_313 ();
 FILLCELL_X4 FILLER_1_318 ();
 FILLCELL_X32 FILLER_1_341 ();
 FILLCELL_X32 FILLER_1_373 ();
 FILLCELL_X32 FILLER_1_405 ();
 FILLCELL_X32 FILLER_1_437 ();
 FILLCELL_X32 FILLER_1_469 ();
 FILLCELL_X4 FILLER_1_501 ();
 FILLCELL_X2 FILLER_1_505 ();
 FILLCELL_X1 FILLER_1_507 ();
 FILLCELL_X32 FILLER_1_512 ();
 FILLCELL_X32 FILLER_1_544 ();
 FILLCELL_X32 FILLER_1_576 ();
 FILLCELL_X32 FILLER_1_608 ();
 FILLCELL_X8 FILLER_1_640 ();
 FILLCELL_X4 FILLER_1_648 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X16 FILLER_2_193 ();
 FILLCELL_X8 FILLER_2_209 ();
 FILLCELL_X4 FILLER_2_217 ();
 FILLCELL_X2 FILLER_2_221 ();
 FILLCELL_X4 FILLER_2_242 ();
 FILLCELL_X4 FILLER_2_265 ();
 FILLCELL_X8 FILLER_2_288 ();
 FILLCELL_X4 FILLER_2_296 ();
 FILLCELL_X2 FILLER_2_300 ();
 FILLCELL_X1 FILLER_2_302 ();
 FILLCELL_X8 FILLER_2_307 ();
 FILLCELL_X4 FILLER_2_315 ();
 FILLCELL_X8 FILLER_2_338 ();
 FILLCELL_X2 FILLER_2_346 ();
 FILLCELL_X32 FILLER_2_351 ();
 FILLCELL_X32 FILLER_2_383 ();
 FILLCELL_X4 FILLER_2_415 ();
 FILLCELL_X1 FILLER_2_419 ();
 FILLCELL_X8 FILLER_2_439 ();
 FILLCELL_X4 FILLER_2_447 ();
 FILLCELL_X2 FILLER_2_451 ();
 FILLCELL_X1 FILLER_2_453 ();
 FILLCELL_X16 FILLER_2_471 ();
 FILLCELL_X8 FILLER_2_487 ();
 FILLCELL_X2 FILLER_2_495 ();
 FILLCELL_X4 FILLER_2_503 ();
 FILLCELL_X4 FILLER_2_513 ();
 FILLCELL_X4 FILLER_2_523 ();
 FILLCELL_X8 FILLER_2_531 ();
 FILLCELL_X2 FILLER_2_539 ();
 FILLCELL_X32 FILLER_2_545 ();
 FILLCELL_X32 FILLER_2_577 ();
 FILLCELL_X16 FILLER_2_609 ();
 FILLCELL_X4 FILLER_2_625 ();
 FILLCELL_X2 FILLER_2_629 ();
 FILLCELL_X8 FILLER_2_632 ();
 FILLCELL_X4 FILLER_2_640 ();
 FILLCELL_X1 FILLER_2_644 ();
 FILLCELL_X4 FILLER_2_648 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X16 FILLER_3_225 ();
 FILLCELL_X2 FILLER_3_241 ();
 FILLCELL_X1 FILLER_3_243 ();
 FILLCELL_X4 FILLER_3_248 ();
 FILLCELL_X2 FILLER_3_252 ();
 FILLCELL_X4 FILLER_3_273 ();
 FILLCELL_X8 FILLER_3_281 ();
 FILLCELL_X4 FILLER_3_293 ();
 FILLCELL_X2 FILLER_3_297 ();
 FILLCELL_X4 FILLER_3_318 ();
 FILLCELL_X1 FILLER_3_322 ();
 FILLCELL_X4 FILLER_3_342 ();
 FILLCELL_X4 FILLER_3_350 ();
 FILLCELL_X1 FILLER_3_354 ();
 FILLCELL_X8 FILLER_3_358 ();
 FILLCELL_X4 FILLER_3_366 ();
 FILLCELL_X2 FILLER_3_370 ();
 FILLCELL_X1 FILLER_3_372 ();
 FILLCELL_X32 FILLER_3_376 ();
 FILLCELL_X16 FILLER_3_408 ();
 FILLCELL_X2 FILLER_3_424 ();
 FILLCELL_X1 FILLER_3_426 ();
 FILLCELL_X4 FILLER_3_431 ();
 FILLCELL_X32 FILLER_3_439 ();
 FILLCELL_X16 FILLER_3_475 ();
 FILLCELL_X4 FILLER_3_491 ();
 FILLCELL_X4 FILLER_3_499 ();
 FILLCELL_X4 FILLER_3_510 ();
 FILLCELL_X4 FILLER_3_523 ();
 FILLCELL_X8 FILLER_3_531 ();
 FILLCELL_X2 FILLER_3_539 ();
 FILLCELL_X1 FILLER_3_541 ();
 FILLCELL_X32 FILLER_3_561 ();
 FILLCELL_X32 FILLER_3_593 ();
 FILLCELL_X16 FILLER_3_625 ();
 FILLCELL_X8 FILLER_3_641 ();
 FILLCELL_X2 FILLER_3_649 ();
 FILLCELL_X1 FILLER_3_651 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X1 FILLER_4_225 ();
 FILLCELL_X8 FILLER_4_229 ();
 FILLCELL_X4 FILLER_4_237 ();
 FILLCELL_X4 FILLER_4_244 ();
 FILLCELL_X4 FILLER_4_251 ();
 FILLCELL_X4 FILLER_4_258 ();
 FILLCELL_X4 FILLER_4_265 ();
 FILLCELL_X8 FILLER_4_273 ();
 FILLCELL_X1 FILLER_4_281 ();
 FILLCELL_X8 FILLER_4_301 ();
 FILLCELL_X1 FILLER_4_309 ();
 FILLCELL_X4 FILLER_4_314 ();
 FILLCELL_X4 FILLER_4_322 ();
 FILLCELL_X4 FILLER_4_330 ();
 FILLCELL_X4 FILLER_4_353 ();
 FILLCELL_X4 FILLER_4_376 ();
 FILLCELL_X16 FILLER_4_383 ();
 FILLCELL_X8 FILLER_4_399 ();
 FILLCELL_X4 FILLER_4_407 ();
 FILLCELL_X1 FILLER_4_411 ();
 FILLCELL_X8 FILLER_4_415 ();
 FILLCELL_X2 FILLER_4_423 ();
 FILLCELL_X32 FILLER_4_444 ();
 FILLCELL_X16 FILLER_4_476 ();
 FILLCELL_X2 FILLER_4_492 ();
 FILLCELL_X1 FILLER_4_494 ();
 FILLCELL_X8 FILLER_4_498 ();
 FILLCELL_X4 FILLER_4_506 ();
 FILLCELL_X2 FILLER_4_510 ();
 FILLCELL_X1 FILLER_4_512 ();
 FILLCELL_X4 FILLER_4_519 ();
 FILLCELL_X4 FILLER_4_527 ();
 FILLCELL_X4 FILLER_4_535 ();
 FILLCELL_X4 FILLER_4_542 ();
 FILLCELL_X32 FILLER_4_548 ();
 FILLCELL_X32 FILLER_4_580 ();
 FILLCELL_X16 FILLER_4_612 ();
 FILLCELL_X2 FILLER_4_628 ();
 FILLCELL_X1 FILLER_4_630 ();
 FILLCELL_X16 FILLER_4_632 ();
 FILLCELL_X4 FILLER_4_648 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X16 FILLER_5_97 ();
 FILLCELL_X4 FILLER_5_113 ();
 FILLCELL_X1 FILLER_5_117 ();
 FILLCELL_X4 FILLER_5_516 ();
 FILLCELL_X4 FILLER_5_527 ();
 FILLCELL_X4 FILLER_5_534 ();
 FILLCELL_X2 FILLER_5_538 ();
 FILLCELL_X4 FILLER_5_544 ();
 FILLCELL_X32 FILLER_5_565 ();
 FILLCELL_X32 FILLER_5_597 ();
 FILLCELL_X16 FILLER_5_629 ();
 FILLCELL_X4 FILLER_5_645 ();
 FILLCELL_X2 FILLER_5_649 ();
 FILLCELL_X1 FILLER_5_651 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X16 FILLER_6_97 ();
 FILLCELL_X4 FILLER_6_113 ();
 FILLCELL_X1 FILLER_6_117 ();
 FILLCELL_X4 FILLER_6_516 ();
 FILLCELL_X8 FILLER_6_523 ();
 FILLCELL_X4 FILLER_6_537 ();
 FILLCELL_X2 FILLER_6_541 ();
 FILLCELL_X4 FILLER_6_547 ();
 FILLCELL_X16 FILLER_6_555 ();
 FILLCELL_X8 FILLER_6_571 ();
 FILLCELL_X2 FILLER_6_579 ();
 FILLCELL_X4 FILLER_6_584 ();
 FILLCELL_X2 FILLER_6_588 ();
 FILLCELL_X1 FILLER_6_590 ();
 FILLCELL_X8 FILLER_6_595 ();
 FILLCELL_X2 FILLER_6_603 ();
 FILLCELL_X1 FILLER_6_605 ();
 FILLCELL_X32 FILLER_6_610 ();
 FILLCELL_X8 FILLER_6_642 ();
 FILLCELL_X2 FILLER_6_650 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X16 FILLER_7_97 ();
 FILLCELL_X4 FILLER_7_113 ();
 FILLCELL_X1 FILLER_7_117 ();
 FILLCELL_X4 FILLER_7_516 ();
 FILLCELL_X4 FILLER_7_523 ();
 FILLCELL_X4 FILLER_7_537 ();
 FILLCELL_X4 FILLER_7_551 ();
 FILLCELL_X4 FILLER_7_564 ();
 FILLCELL_X4 FILLER_7_572 ();
 FILLCELL_X2 FILLER_7_576 ();
 FILLCELL_X4 FILLER_7_582 ();
 FILLCELL_X4 FILLER_7_590 ();
 FILLCELL_X2 FILLER_7_594 ();
 FILLCELL_X1 FILLER_7_596 ();
 FILLCELL_X4 FILLER_7_614 ();
 FILLCELL_X16 FILLER_7_623 ();
 FILLCELL_X8 FILLER_7_639 ();
 FILLCELL_X4 FILLER_7_647 ();
 FILLCELL_X1 FILLER_7_651 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X16 FILLER_8_97 ();
 FILLCELL_X4 FILLER_8_113 ();
 FILLCELL_X1 FILLER_8_117 ();
 FILLCELL_X8 FILLER_8_516 ();
 FILLCELL_X4 FILLER_8_528 ();
 FILLCELL_X4 FILLER_8_536 ();
 FILLCELL_X4 FILLER_8_542 ();
 FILLCELL_X1 FILLER_8_546 ();
 FILLCELL_X4 FILLER_8_556 ();
 FILLCELL_X4 FILLER_8_563 ();
 FILLCELL_X2 FILLER_8_567 ();
 FILLCELL_X1 FILLER_8_569 ();
 FILLCELL_X4 FILLER_8_574 ();
 FILLCELL_X4 FILLER_8_587 ();
 FILLCELL_X1 FILLER_8_591 ();
 FILLCELL_X4 FILLER_8_596 ();
 FILLCELL_X4 FILLER_8_604 ();
 FILLCELL_X4 FILLER_8_613 ();
 FILLCELL_X4 FILLER_8_626 ();
 FILLCELL_X16 FILLER_8_632 ();
 FILLCELL_X4 FILLER_8_648 ();
 FILLCELL_X4 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_8 ();
 FILLCELL_X32 FILLER_9_40 ();
 FILLCELL_X32 FILLER_9_72 ();
 FILLCELL_X8 FILLER_9_104 ();
 FILLCELL_X4 FILLER_9_112 ();
 FILLCELL_X2 FILLER_9_116 ();
 FILLCELL_X4 FILLER_9_516 ();
 FILLCELL_X8 FILLER_9_522 ();
 FILLCELL_X4 FILLER_9_536 ();
 FILLCELL_X4 FILLER_9_544 ();
 FILLCELL_X4 FILLER_9_552 ();
 FILLCELL_X8 FILLER_9_559 ();
 FILLCELL_X4 FILLER_9_569 ();
 FILLCELL_X1 FILLER_9_573 ();
 FILLCELL_X4 FILLER_9_577 ();
 FILLCELL_X4 FILLER_9_590 ();
 FILLCELL_X4 FILLER_9_598 ();
 FILLCELL_X1 FILLER_9_602 ();
 FILLCELL_X8 FILLER_9_607 ();
 FILLCELL_X1 FILLER_9_615 ();
 FILLCELL_X4 FILLER_9_633 ();
 FILLCELL_X8 FILLER_9_640 ();
 FILLCELL_X4 FILLER_9_648 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X16 FILLER_10_97 ();
 FILLCELL_X4 FILLER_10_113 ();
 FILLCELL_X1 FILLER_10_117 ();
 FILLCELL_X4 FILLER_10_516 ();
 FILLCELL_X8 FILLER_10_523 ();
 FILLCELL_X2 FILLER_10_531 ();
 FILLCELL_X1 FILLER_10_533 ();
 FILLCELL_X4 FILLER_10_541 ();
 FILLCELL_X2 FILLER_10_545 ();
 FILLCELL_X1 FILLER_10_547 ();
 FILLCELL_X4 FILLER_10_551 ();
 FILLCELL_X4 FILLER_10_558 ();
 FILLCELL_X4 FILLER_10_564 ();
 FILLCELL_X4 FILLER_10_570 ();
 FILLCELL_X2 FILLER_10_574 ();
 FILLCELL_X1 FILLER_10_576 ();
 FILLCELL_X16 FILLER_10_579 ();
 FILLCELL_X2 FILLER_10_595 ();
 FILLCELL_X1 FILLER_10_597 ();
 FILLCELL_X8 FILLER_10_601 ();
 FILLCELL_X4 FILLER_10_613 ();
 FILLCELL_X4 FILLER_10_620 ();
 FILLCELL_X1 FILLER_10_624 ();
 FILLCELL_X4 FILLER_10_628 ();
 FILLCELL_X16 FILLER_10_635 ();
 FILLCELL_X1 FILLER_10_651 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X16 FILLER_11_97 ();
 FILLCELL_X4 FILLER_11_113 ();
 FILLCELL_X1 FILLER_11_117 ();
 FILLCELL_X16 FILLER_11_516 ();
 FILLCELL_X2 FILLER_11_532 ();
 FILLCELL_X1 FILLER_11_534 ();
 FILLCELL_X4 FILLER_11_541 ();
 FILLCELL_X2 FILLER_11_545 ();
 FILLCELL_X1 FILLER_11_547 ();
 FILLCELL_X4 FILLER_11_551 ();
 FILLCELL_X4 FILLER_11_561 ();
 FILLCELL_X4 FILLER_11_568 ();
 FILLCELL_X2 FILLER_11_572 ();
 FILLCELL_X4 FILLER_11_584 ();
 FILLCELL_X4 FILLER_11_592 ();
 FILLCELL_X8 FILLER_11_598 ();
 FILLCELL_X4 FILLER_11_606 ();
 FILLCELL_X2 FILLER_11_610 ();
 FILLCELL_X1 FILLER_11_612 ();
 FILLCELL_X4 FILLER_11_615 ();
 FILLCELL_X2 FILLER_11_619 ();
 FILLCELL_X1 FILLER_11_621 ();
 FILLCELL_X8 FILLER_11_631 ();
 FILLCELL_X2 FILLER_11_639 ();
 FILLCELL_X1 FILLER_11_641 ();
 FILLCELL_X4 FILLER_11_646 ();
 FILLCELL_X2 FILLER_11_650 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X16 FILLER_12_97 ();
 FILLCELL_X4 FILLER_12_113 ();
 FILLCELL_X1 FILLER_12_117 ();
 FILLCELL_X4 FILLER_12_516 ();
 FILLCELL_X4 FILLER_12_525 ();
 FILLCELL_X2 FILLER_12_529 ();
 FILLCELL_X4 FILLER_12_535 ();
 FILLCELL_X4 FILLER_12_541 ();
 FILLCELL_X2 FILLER_12_545 ();
 FILLCELL_X4 FILLER_12_551 ();
 FILLCELL_X4 FILLER_12_561 ();
 FILLCELL_X8 FILLER_12_571 ();
 FILLCELL_X4 FILLER_12_585 ();
 FILLCELL_X4 FILLER_12_593 ();
 FILLCELL_X1 FILLER_12_597 ();
 FILLCELL_X4 FILLER_12_602 ();
 FILLCELL_X4 FILLER_12_610 ();
 FILLCELL_X4 FILLER_12_618 ();
 FILLCELL_X4 FILLER_12_625 ();
 FILLCELL_X1 FILLER_12_629 ();
 FILLCELL_X4 FILLER_12_647 ();
 FILLCELL_X1 FILLER_12_651 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X16 FILLER_13_97 ();
 FILLCELL_X4 FILLER_13_113 ();
 FILLCELL_X1 FILLER_13_117 ();
 FILLCELL_X4 FILLER_13_516 ();
 FILLCELL_X4 FILLER_13_526 ();
 FILLCELL_X4 FILLER_13_532 ();
 FILLCELL_X1 FILLER_13_536 ();
 FILLCELL_X4 FILLER_13_543 ();
 FILLCELL_X4 FILLER_13_553 ();
 FILLCELL_X4 FILLER_13_559 ();
 FILLCELL_X4 FILLER_13_582 ();
 FILLCELL_X4 FILLER_13_590 ();
 FILLCELL_X1 FILLER_13_594 ();
 FILLCELL_X4 FILLER_13_599 ();
 FILLCELL_X4 FILLER_13_606 ();
 FILLCELL_X4 FILLER_13_619 ();
 FILLCELL_X2 FILLER_13_623 ();
 FILLCELL_X4 FILLER_13_632 ();
 FILLCELL_X8 FILLER_13_642 ();
 FILLCELL_X2 FILLER_13_650 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X8 FILLER_14_97 ();
 FILLCELL_X4 FILLER_14_105 ();
 FILLCELL_X2 FILLER_14_109 ();
 FILLCELL_X4 FILLER_14_114 ();
 FILLCELL_X4 FILLER_14_516 ();
 FILLCELL_X4 FILLER_14_537 ();
 FILLCELL_X4 FILLER_14_548 ();
 FILLCELL_X4 FILLER_14_556 ();
 FILLCELL_X4 FILLER_14_564 ();
 FILLCELL_X1 FILLER_14_568 ();
 FILLCELL_X8 FILLER_14_571 ();
 FILLCELL_X1 FILLER_14_579 ();
 FILLCELL_X4 FILLER_14_584 ();
 FILLCELL_X4 FILLER_14_590 ();
 FILLCELL_X4 FILLER_14_596 ();
 FILLCELL_X4 FILLER_14_602 ();
 FILLCELL_X1 FILLER_14_606 ();
 FILLCELL_X4 FILLER_14_611 ();
 FILLCELL_X8 FILLER_14_618 ();
 FILLCELL_X1 FILLER_14_626 ();
 FILLCELL_X4 FILLER_14_633 ();
 FILLCELL_X8 FILLER_14_643 ();
 FILLCELL_X1 FILLER_14_651 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X8 FILLER_15_97 ();
 FILLCELL_X4 FILLER_15_105 ();
 FILLCELL_X1 FILLER_15_109 ();
 FILLCELL_X4 FILLER_15_114 ();
 FILLCELL_X4 FILLER_15_516 ();
 FILLCELL_X8 FILLER_15_524 ();
 FILLCELL_X1 FILLER_15_532 ();
 FILLCELL_X4 FILLER_15_535 ();
 FILLCELL_X2 FILLER_15_539 ();
 FILLCELL_X1 FILLER_15_541 ();
 FILLCELL_X4 FILLER_15_545 ();
 FILLCELL_X4 FILLER_15_552 ();
 FILLCELL_X4 FILLER_15_559 ();
 FILLCELL_X8 FILLER_15_565 ();
 FILLCELL_X16 FILLER_15_575 ();
 FILLCELL_X2 FILLER_15_591 ();
 FILLCELL_X16 FILLER_15_596 ();
 FILLCELL_X8 FILLER_15_612 ();
 FILLCELL_X2 FILLER_15_620 ();
 FILLCELL_X4 FILLER_15_625 ();
 FILLCELL_X2 FILLER_15_629 ();
 FILLCELL_X1 FILLER_15_631 ();
 FILLCELL_X4 FILLER_15_636 ();
 FILLCELL_X2 FILLER_15_640 ();
 FILLCELL_X1 FILLER_15_642 ();
 FILLCELL_X4 FILLER_15_647 ();
 FILLCELL_X1 FILLER_15_651 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X16 FILLER_16_65 ();
 FILLCELL_X8 FILLER_16_81 ();
 FILLCELL_X4 FILLER_16_89 ();
 FILLCELL_X2 FILLER_16_93 ();
 FILLCELL_X4 FILLER_16_114 ();
 FILLCELL_X8 FILLER_16_516 ();
 FILLCELL_X4 FILLER_16_524 ();
 FILLCELL_X2 FILLER_16_528 ();
 FILLCELL_X1 FILLER_16_530 ();
 FILLCELL_X4 FILLER_16_534 ();
 FILLCELL_X16 FILLER_16_547 ();
 FILLCELL_X8 FILLER_16_563 ();
 FILLCELL_X4 FILLER_16_571 ();
 FILLCELL_X1 FILLER_16_575 ();
 FILLCELL_X4 FILLER_16_579 ();
 FILLCELL_X4 FILLER_16_587 ();
 FILLCELL_X8 FILLER_16_601 ();
 FILLCELL_X4 FILLER_16_612 ();
 FILLCELL_X4 FILLER_16_619 ();
 FILLCELL_X1 FILLER_16_623 ();
 FILLCELL_X4 FILLER_16_626 ();
 FILLCELL_X8 FILLER_16_636 ();
 FILLCELL_X4 FILLER_16_648 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X16 FILLER_17_97 ();
 FILLCELL_X4 FILLER_17_113 ();
 FILLCELL_X1 FILLER_17_117 ();
 FILLCELL_X8 FILLER_17_516 ();
 FILLCELL_X4 FILLER_17_524 ();
 FILLCELL_X2 FILLER_17_528 ();
 FILLCELL_X1 FILLER_17_530 ();
 FILLCELL_X4 FILLER_17_534 ();
 FILLCELL_X4 FILLER_17_542 ();
 FILLCELL_X4 FILLER_17_550 ();
 FILLCELL_X8 FILLER_17_556 ();
 FILLCELL_X4 FILLER_17_564 ();
 FILLCELL_X4 FILLER_17_572 ();
 FILLCELL_X4 FILLER_17_580 ();
 FILLCELL_X8 FILLER_17_587 ();
 FILLCELL_X1 FILLER_17_595 ();
 FILLCELL_X4 FILLER_17_600 ();
 FILLCELL_X4 FILLER_17_608 ();
 FILLCELL_X2 FILLER_17_612 ();
 FILLCELL_X4 FILLER_17_623 ();
 FILLCELL_X4 FILLER_17_630 ();
 FILLCELL_X1 FILLER_17_634 ();
 FILLCELL_X4 FILLER_17_641 ();
 FILLCELL_X4 FILLER_17_648 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X16 FILLER_18_97 ();
 FILLCELL_X4 FILLER_18_113 ();
 FILLCELL_X1 FILLER_18_117 ();
 FILLCELL_X16 FILLER_18_516 ();
 FILLCELL_X2 FILLER_18_532 ();
 FILLCELL_X1 FILLER_18_534 ();
 FILLCELL_X4 FILLER_18_545 ();
 FILLCELL_X4 FILLER_18_558 ();
 FILLCELL_X2 FILLER_18_562 ();
 FILLCELL_X4 FILLER_18_566 ();
 FILLCELL_X4 FILLER_18_579 ();
 FILLCELL_X8 FILLER_18_587 ();
 FILLCELL_X1 FILLER_18_595 ();
 FILLCELL_X4 FILLER_18_603 ();
 FILLCELL_X4 FILLER_18_616 ();
 FILLCELL_X2 FILLER_18_620 ();
 FILLCELL_X1 FILLER_18_622 ();
 FILLCELL_X4 FILLER_18_633 ();
 FILLCELL_X8 FILLER_18_644 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X16 FILLER_19_97 ();
 FILLCELL_X4 FILLER_19_113 ();
 FILLCELL_X1 FILLER_19_117 ();
 FILLCELL_X4 FILLER_19_516 ();
 FILLCELL_X2 FILLER_19_520 ();
 FILLCELL_X4 FILLER_19_524 ();
 FILLCELL_X4 FILLER_19_532 ();
 FILLCELL_X4 FILLER_19_545 ();
 FILLCELL_X4 FILLER_19_553 ();
 FILLCELL_X4 FILLER_19_561 ();
 FILLCELL_X4 FILLER_19_568 ();
 FILLCELL_X4 FILLER_19_575 ();
 FILLCELL_X4 FILLER_19_588 ();
 FILLCELL_X8 FILLER_19_594 ();
 FILLCELL_X2 FILLER_19_602 ();
 FILLCELL_X4 FILLER_19_614 ();
 FILLCELL_X2 FILLER_19_618 ();
 FILLCELL_X4 FILLER_19_623 ();
 FILLCELL_X4 FILLER_19_631 ();
 FILLCELL_X8 FILLER_19_641 ();
 FILLCELL_X2 FILLER_19_649 ();
 FILLCELL_X1 FILLER_19_651 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X16 FILLER_20_97 ();
 FILLCELL_X4 FILLER_20_113 ();
 FILLCELL_X1 FILLER_20_117 ();
 FILLCELL_X8 FILLER_20_516 ();
 FILLCELL_X4 FILLER_20_524 ();
 FILLCELL_X4 FILLER_20_531 ();
 FILLCELL_X4 FILLER_20_545 ();
 FILLCELL_X8 FILLER_20_556 ();
 FILLCELL_X2 FILLER_20_564 ();
 FILLCELL_X1 FILLER_20_566 ();
 FILLCELL_X4 FILLER_20_571 ();
 FILLCELL_X4 FILLER_20_579 ();
 FILLCELL_X2 FILLER_20_583 ();
 FILLCELL_X4 FILLER_20_588 ();
 FILLCELL_X4 FILLER_20_595 ();
 FILLCELL_X16 FILLER_20_602 ();
 FILLCELL_X8 FILLER_20_618 ();
 FILLCELL_X4 FILLER_20_626 ();
 FILLCELL_X4 FILLER_20_647 ();
 FILLCELL_X1 FILLER_20_651 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X16 FILLER_21_97 ();
 FILLCELL_X4 FILLER_21_113 ();
 FILLCELL_X1 FILLER_21_117 ();
 FILLCELL_X8 FILLER_21_516 ();
 FILLCELL_X4 FILLER_21_524 ();
 FILLCELL_X2 FILLER_21_528 ();
 FILLCELL_X4 FILLER_21_533 ();
 FILLCELL_X1 FILLER_21_537 ();
 FILLCELL_X4 FILLER_21_540 ();
 FILLCELL_X16 FILLER_21_546 ();
 FILLCELL_X8 FILLER_21_562 ();
 FILLCELL_X4 FILLER_21_570 ();
 FILLCELL_X4 FILLER_21_583 ();
 FILLCELL_X2 FILLER_21_587 ();
 FILLCELL_X4 FILLER_21_593 ();
 FILLCELL_X4 FILLER_21_607 ();
 FILLCELL_X8 FILLER_21_613 ();
 FILLCELL_X2 FILLER_21_621 ();
 FILLCELL_X1 FILLER_21_623 ();
 FILLCELL_X8 FILLER_21_626 ();
 FILLCELL_X8 FILLER_21_638 ();
 FILLCELL_X4 FILLER_21_646 ();
 FILLCELL_X2 FILLER_21_650 ();
 FILLCELL_X4 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_8 ();
 FILLCELL_X32 FILLER_22_40 ();
 FILLCELL_X16 FILLER_22_72 ();
 FILLCELL_X8 FILLER_22_88 ();
 FILLCELL_X4 FILLER_22_96 ();
 FILLCELL_X4 FILLER_22_105 ();
 FILLCELL_X4 FILLER_22_114 ();
 FILLCELL_X4 FILLER_22_516 ();
 FILLCELL_X4 FILLER_22_523 ();
 FILLCELL_X1 FILLER_22_527 ();
 FILLCELL_X4 FILLER_22_532 ();
 FILLCELL_X2 FILLER_22_536 ();
 FILLCELL_X1 FILLER_22_538 ();
 FILLCELL_X4 FILLER_22_542 ();
 FILLCELL_X4 FILLER_22_548 ();
 FILLCELL_X2 FILLER_22_552 ();
 FILLCELL_X4 FILLER_22_558 ();
 FILLCELL_X4 FILLER_22_566 ();
 FILLCELL_X8 FILLER_22_574 ();
 FILLCELL_X2 FILLER_22_582 ();
 FILLCELL_X4 FILLER_22_593 ();
 FILLCELL_X4 FILLER_22_600 ();
 FILLCELL_X2 FILLER_22_604 ();
 FILLCELL_X16 FILLER_22_613 ();
 FILLCELL_X8 FILLER_22_639 ();
 FILLCELL_X4 FILLER_22_647 ();
 FILLCELL_X1 FILLER_22_651 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X16 FILLER_23_97 ();
 FILLCELL_X4 FILLER_23_113 ();
 FILLCELL_X1 FILLER_23_117 ();
 FILLCELL_X8 FILLER_23_516 ();
 FILLCELL_X4 FILLER_23_531 ();
 FILLCELL_X4 FILLER_23_539 ();
 FILLCELL_X4 FILLER_23_545 ();
 FILLCELL_X4 FILLER_23_553 ();
 FILLCELL_X4 FILLER_23_561 ();
 FILLCELL_X2 FILLER_23_565 ();
 FILLCELL_X1 FILLER_23_567 ();
 FILLCELL_X4 FILLER_23_577 ();
 FILLCELL_X4 FILLER_23_585 ();
 FILLCELL_X4 FILLER_23_592 ();
 FILLCELL_X8 FILLER_23_598 ();
 FILLCELL_X4 FILLER_23_616 ();
 FILLCELL_X4 FILLER_23_623 ();
 FILLCELL_X4 FILLER_23_630 ();
 FILLCELL_X8 FILLER_23_637 ();
 FILLCELL_X4 FILLER_23_645 ();
 FILLCELL_X2 FILLER_23_649 ();
 FILLCELL_X1 FILLER_23_651 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X16 FILLER_24_97 ();
 FILLCELL_X4 FILLER_24_113 ();
 FILLCELL_X1 FILLER_24_117 ();
 FILLCELL_X4 FILLER_24_516 ();
 FILLCELL_X4 FILLER_24_522 ();
 FILLCELL_X1 FILLER_24_526 ();
 FILLCELL_X4 FILLER_24_533 ();
 FILLCELL_X4 FILLER_24_541 ();
 FILLCELL_X4 FILLER_24_549 ();
 FILLCELL_X4 FILLER_24_556 ();
 FILLCELL_X4 FILLER_24_569 ();
 FILLCELL_X4 FILLER_24_577 ();
 FILLCELL_X4 FILLER_24_584 ();
 FILLCELL_X4 FILLER_24_591 ();
 FILLCELL_X2 FILLER_24_595 ();
 FILLCELL_X4 FILLER_24_600 ();
 FILLCELL_X8 FILLER_24_608 ();
 FILLCELL_X4 FILLER_24_625 ();
 FILLCELL_X4 FILLER_24_638 ();
 FILLCELL_X2 FILLER_24_642 ();
 FILLCELL_X1 FILLER_24_644 ();
 FILLCELL_X4 FILLER_24_648 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X16 FILLER_25_97 ();
 FILLCELL_X4 FILLER_25_113 ();
 FILLCELL_X1 FILLER_25_117 ();
 FILLCELL_X4 FILLER_25_516 ();
 FILLCELL_X4 FILLER_25_537 ();
 FILLCELL_X4 FILLER_25_545 ();
 FILLCELL_X4 FILLER_25_553 ();
 FILLCELL_X2 FILLER_25_557 ();
 FILLCELL_X1 FILLER_25_559 ();
 FILLCELL_X8 FILLER_25_564 ();
 FILLCELL_X2 FILLER_25_572 ();
 FILLCELL_X4 FILLER_25_583 ();
 FILLCELL_X4 FILLER_25_591 ();
 FILLCELL_X16 FILLER_25_605 ();
 FILLCELL_X1 FILLER_25_621 ();
 FILLCELL_X4 FILLER_25_625 ();
 FILLCELL_X4 FILLER_25_639 ();
 FILLCELL_X1 FILLER_25_643 ();
 FILLCELL_X4 FILLER_25_648 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X16 FILLER_26_97 ();
 FILLCELL_X4 FILLER_26_113 ();
 FILLCELL_X1 FILLER_26_117 ();
 FILLCELL_X4 FILLER_26_516 ();
 FILLCELL_X4 FILLER_26_522 ();
 FILLCELL_X4 FILLER_26_532 ();
 FILLCELL_X4 FILLER_26_540 ();
 FILLCELL_X4 FILLER_26_548 ();
 FILLCELL_X4 FILLER_26_555 ();
 FILLCELL_X8 FILLER_26_562 ();
 FILLCELL_X4 FILLER_26_570 ();
 FILLCELL_X1 FILLER_26_574 ();
 FILLCELL_X16 FILLER_26_578 ();
 FILLCELL_X4 FILLER_26_594 ();
 FILLCELL_X1 FILLER_26_598 ();
 FILLCELL_X4 FILLER_26_601 ();
 FILLCELL_X16 FILLER_26_612 ();
 FILLCELL_X2 FILLER_26_628 ();
 FILLCELL_X4 FILLER_26_633 ();
 FILLCELL_X8 FILLER_26_644 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X16 FILLER_27_97 ();
 FILLCELL_X4 FILLER_27_113 ();
 FILLCELL_X1 FILLER_27_117 ();
 FILLCELL_X4 FILLER_27_516 ();
 FILLCELL_X8 FILLER_27_525 ();
 FILLCELL_X1 FILLER_27_533 ();
 FILLCELL_X4 FILLER_27_540 ();
 FILLCELL_X4 FILLER_27_547 ();
 FILLCELL_X4 FILLER_27_560 ();
 FILLCELL_X4 FILLER_27_573 ();
 FILLCELL_X8 FILLER_27_581 ();
 FILLCELL_X4 FILLER_27_589 ();
 FILLCELL_X2 FILLER_27_593 ();
 FILLCELL_X4 FILLER_27_599 ();
 FILLCELL_X4 FILLER_27_613 ();
 FILLCELL_X4 FILLER_27_621 ();
 FILLCELL_X8 FILLER_27_628 ();
 FILLCELL_X4 FILLER_27_642 ();
 FILLCELL_X4 FILLER_27_648 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X16 FILLER_28_97 ();
 FILLCELL_X4 FILLER_28_113 ();
 FILLCELL_X1 FILLER_28_117 ();
 FILLCELL_X4 FILLER_28_516 ();
 FILLCELL_X4 FILLER_28_523 ();
 FILLCELL_X4 FILLER_28_529 ();
 FILLCELL_X1 FILLER_28_533 ();
 FILLCELL_X4 FILLER_28_540 ();
 FILLCELL_X1 FILLER_28_544 ();
 FILLCELL_X16 FILLER_28_549 ();
 FILLCELL_X4 FILLER_28_565 ();
 FILLCELL_X1 FILLER_28_569 ();
 FILLCELL_X4 FILLER_28_573 ();
 FILLCELL_X4 FILLER_28_587 ();
 FILLCELL_X2 FILLER_28_591 ();
 FILLCELL_X8 FILLER_28_597 ();
 FILLCELL_X1 FILLER_28_605 ();
 FILLCELL_X4 FILLER_28_611 ();
 FILLCELL_X4 FILLER_28_624 ();
 FILLCELL_X4 FILLER_28_637 ();
 FILLCELL_X4 FILLER_28_647 ();
 FILLCELL_X1 FILLER_28_651 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X16 FILLER_29_97 ();
 FILLCELL_X4 FILLER_29_113 ();
 FILLCELL_X1 FILLER_29_117 ();
 FILLCELL_X4 FILLER_29_516 ();
 FILLCELL_X16 FILLER_29_525 ();
 FILLCELL_X4 FILLER_29_541 ();
 FILLCELL_X2 FILLER_29_545 ();
 FILLCELL_X4 FILLER_29_556 ();
 FILLCELL_X4 FILLER_29_564 ();
 FILLCELL_X4 FILLER_29_571 ();
 FILLCELL_X4 FILLER_29_577 ();
 FILLCELL_X16 FILLER_29_583 ();
 FILLCELL_X4 FILLER_29_599 ();
 FILLCELL_X4 FILLER_29_607 ();
 FILLCELL_X4 FILLER_29_616 ();
 FILLCELL_X1 FILLER_29_620 ();
 FILLCELL_X4 FILLER_29_624 ();
 FILLCELL_X4 FILLER_29_631 ();
 FILLCELL_X4 FILLER_29_645 ();
 FILLCELL_X2 FILLER_29_649 ();
 FILLCELL_X1 FILLER_29_651 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X16 FILLER_30_97 ();
 FILLCELL_X4 FILLER_30_113 ();
 FILLCELL_X1 FILLER_30_117 ();
 FILLCELL_X8 FILLER_30_516 ();
 FILLCELL_X8 FILLER_30_528 ();
 FILLCELL_X4 FILLER_30_536 ();
 FILLCELL_X8 FILLER_30_544 ();
 FILLCELL_X1 FILLER_30_552 ();
 FILLCELL_X4 FILLER_30_556 ();
 FILLCELL_X8 FILLER_30_570 ();
 FILLCELL_X4 FILLER_30_588 ();
 FILLCELL_X4 FILLER_30_599 ();
 FILLCELL_X4 FILLER_30_607 ();
 FILLCELL_X4 FILLER_30_614 ();
 FILLCELL_X8 FILLER_30_620 ();
 FILLCELL_X1 FILLER_30_628 ();
 FILLCELL_X4 FILLER_30_638 ();
 FILLCELL_X2 FILLER_30_642 ();
 FILLCELL_X1 FILLER_30_644 ();
 FILLCELL_X4 FILLER_30_648 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X16 FILLER_31_97 ();
 FILLCELL_X4 FILLER_31_113 ();
 FILLCELL_X1 FILLER_31_117 ();
 FILLCELL_X16 FILLER_31_516 ();
 FILLCELL_X8 FILLER_31_532 ();
 FILLCELL_X4 FILLER_31_540 ();
 FILLCELL_X1 FILLER_31_544 ();
 FILLCELL_X4 FILLER_31_547 ();
 FILLCELL_X4 FILLER_31_554 ();
 FILLCELL_X8 FILLER_31_560 ();
 FILLCELL_X4 FILLER_31_572 ();
 FILLCELL_X4 FILLER_31_578 ();
 FILLCELL_X1 FILLER_31_582 ();
 FILLCELL_X4 FILLER_31_587 ();
 FILLCELL_X4 FILLER_31_595 ();
 FILLCELL_X1 FILLER_31_599 ();
 FILLCELL_X4 FILLER_31_609 ();
 FILLCELL_X4 FILLER_31_616 ();
 FILLCELL_X8 FILLER_31_623 ();
 FILLCELL_X4 FILLER_31_631 ();
 FILLCELL_X1 FILLER_31_635 ();
 FILLCELL_X8 FILLER_31_640 ();
 FILLCELL_X4 FILLER_31_648 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X16 FILLER_32_97 ();
 FILLCELL_X4 FILLER_32_113 ();
 FILLCELL_X1 FILLER_32_117 ();
 FILLCELL_X4 FILLER_32_516 ();
 FILLCELL_X4 FILLER_32_524 ();
 FILLCELL_X4 FILLER_32_537 ();
 FILLCELL_X4 FILLER_32_551 ();
 FILLCELL_X1 FILLER_32_555 ();
 FILLCELL_X4 FILLER_32_566 ();
 FILLCELL_X8 FILLER_32_577 ();
 FILLCELL_X2 FILLER_32_585 ();
 FILLCELL_X4 FILLER_32_591 ();
 FILLCELL_X8 FILLER_32_599 ();
 FILLCELL_X1 FILLER_32_607 ();
 FILLCELL_X4 FILLER_32_617 ();
 FILLCELL_X2 FILLER_32_621 ();
 FILLCELL_X4 FILLER_32_625 ();
 FILLCELL_X4 FILLER_32_648 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X16 FILLER_33_97 ();
 FILLCELL_X4 FILLER_33_113 ();
 FILLCELL_X1 FILLER_33_117 ();
 FILLCELL_X4 FILLER_33_516 ();
 FILLCELL_X4 FILLER_33_539 ();
 FILLCELL_X4 FILLER_33_547 ();
 FILLCELL_X8 FILLER_33_555 ();
 FILLCELL_X4 FILLER_33_567 ();
 FILLCELL_X4 FILLER_33_575 ();
 FILLCELL_X2 FILLER_33_579 ();
 FILLCELL_X1 FILLER_33_581 ();
 FILLCELL_X4 FILLER_33_586 ();
 FILLCELL_X2 FILLER_33_590 ();
 FILLCELL_X4 FILLER_33_595 ();
 FILLCELL_X8 FILLER_33_602 ();
 FILLCELL_X4 FILLER_33_610 ();
 FILLCELL_X2 FILLER_33_614 ();
 FILLCELL_X4 FILLER_33_619 ();
 FILLCELL_X4 FILLER_33_626 ();
 FILLCELL_X1 FILLER_33_630 ();
 FILLCELL_X8 FILLER_33_634 ();
 FILLCELL_X2 FILLER_33_642 ();
 FILLCELL_X4 FILLER_33_648 ();
 FILLCELL_X4 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_8 ();
 FILLCELL_X32 FILLER_34_40 ();
 FILLCELL_X32 FILLER_34_72 ();
 FILLCELL_X8 FILLER_34_104 ();
 FILLCELL_X4 FILLER_34_112 ();
 FILLCELL_X2 FILLER_34_116 ();
 FILLCELL_X4 FILLER_34_516 ();
 FILLCELL_X2 FILLER_34_520 ();
 FILLCELL_X1 FILLER_34_522 ();
 FILLCELL_X8 FILLER_34_526 ();
 FILLCELL_X1 FILLER_34_534 ();
 FILLCELL_X4 FILLER_34_544 ();
 FILLCELL_X4 FILLER_34_550 ();
 FILLCELL_X4 FILLER_34_557 ();
 FILLCELL_X16 FILLER_34_563 ();
 FILLCELL_X4 FILLER_34_579 ();
 FILLCELL_X2 FILLER_34_583 ();
 FILLCELL_X1 FILLER_34_585 ();
 FILLCELL_X4 FILLER_34_588 ();
 FILLCELL_X8 FILLER_34_601 ();
 FILLCELL_X1 FILLER_34_609 ();
 FILLCELL_X4 FILLER_34_613 ();
 FILLCELL_X1 FILLER_34_617 ();
 FILLCELL_X8 FILLER_34_628 ();
 FILLCELL_X4 FILLER_34_640 ();
 FILLCELL_X4 FILLER_34_648 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X8 FILLER_35_97 ();
 FILLCELL_X4 FILLER_35_105 ();
 FILLCELL_X2 FILLER_35_109 ();
 FILLCELL_X4 FILLER_35_114 ();
 FILLCELL_X8 FILLER_35_516 ();
 FILLCELL_X4 FILLER_35_524 ();
 FILLCELL_X4 FILLER_35_531 ();
 FILLCELL_X4 FILLER_35_538 ();
 FILLCELL_X8 FILLER_35_552 ();
 FILLCELL_X2 FILLER_35_560 ();
 FILLCELL_X8 FILLER_35_571 ();
 FILLCELL_X4 FILLER_35_579 ();
 FILLCELL_X4 FILLER_35_585 ();
 FILLCELL_X4 FILLER_35_598 ();
 FILLCELL_X2 FILLER_35_602 ();
 FILLCELL_X1 FILLER_35_604 ();
 FILLCELL_X4 FILLER_35_614 ();
 FILLCELL_X4 FILLER_35_628 ();
 FILLCELL_X1 FILLER_35_632 ();
 FILLCELL_X8 FILLER_35_643 ();
 FILLCELL_X1 FILLER_35_651 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X8 FILLER_36_97 ();
 FILLCELL_X4 FILLER_36_105 ();
 FILLCELL_X4 FILLER_36_114 ();
 FILLCELL_X4 FILLER_36_516 ();
 FILLCELL_X1 FILLER_36_520 ();
 FILLCELL_X8 FILLER_36_523 ();
 FILLCELL_X4 FILLER_36_531 ();
 FILLCELL_X1 FILLER_36_535 ();
 FILLCELL_X4 FILLER_36_540 ();
 FILLCELL_X4 FILLER_36_551 ();
 FILLCELL_X4 FILLER_36_564 ();
 FILLCELL_X4 FILLER_36_572 ();
 FILLCELL_X2 FILLER_36_576 ();
 FILLCELL_X4 FILLER_36_581 ();
 FILLCELL_X4 FILLER_36_595 ();
 FILLCELL_X2 FILLER_36_599 ();
 FILLCELL_X1 FILLER_36_601 ();
 FILLCELL_X4 FILLER_36_605 ();
 FILLCELL_X8 FILLER_36_618 ();
 FILLCELL_X4 FILLER_36_630 ();
 FILLCELL_X2 FILLER_36_634 ();
 FILLCELL_X1 FILLER_36_636 ();
 FILLCELL_X8 FILLER_36_644 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X16 FILLER_37_97 ();
 FILLCELL_X4 FILLER_37_113 ();
 FILLCELL_X1 FILLER_37_117 ();
 FILLCELL_X16 FILLER_37_516 ();
 FILLCELL_X4 FILLER_37_532 ();
 FILLCELL_X1 FILLER_37_536 ();
 FILLCELL_X4 FILLER_37_540 ();
 FILLCELL_X8 FILLER_37_553 ();
 FILLCELL_X4 FILLER_37_561 ();
 FILLCELL_X2 FILLER_37_565 ();
 FILLCELL_X4 FILLER_37_569 ();
 FILLCELL_X1 FILLER_37_573 ();
 FILLCELL_X4 FILLER_37_583 ();
 FILLCELL_X4 FILLER_37_597 ();
 FILLCELL_X8 FILLER_37_605 ();
 FILLCELL_X2 FILLER_37_613 ();
 FILLCELL_X4 FILLER_37_617 ();
 FILLCELL_X4 FILLER_37_624 ();
 FILLCELL_X4 FILLER_37_638 ();
 FILLCELL_X4 FILLER_37_648 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X16 FILLER_38_97 ();
 FILLCELL_X4 FILLER_38_113 ();
 FILLCELL_X1 FILLER_38_117 ();
 FILLCELL_X8 FILLER_38_516 ();
 FILLCELL_X1 FILLER_38_524 ();
 FILLCELL_X4 FILLER_38_527 ();
 FILLCELL_X4 FILLER_38_534 ();
 FILLCELL_X16 FILLER_38_548 ();
 FILLCELL_X1 FILLER_38_564 ();
 FILLCELL_X8 FILLER_38_568 ();
 FILLCELL_X1 FILLER_38_576 ();
 FILLCELL_X4 FILLER_38_586 ();
 FILLCELL_X4 FILLER_38_593 ();
 FILLCELL_X4 FILLER_38_600 ();
 FILLCELL_X4 FILLER_38_607 ();
 FILLCELL_X4 FILLER_38_613 ();
 FILLCELL_X2 FILLER_38_617 ();
 FILLCELL_X1 FILLER_38_619 ();
 FILLCELL_X4 FILLER_38_622 ();
 FILLCELL_X4 FILLER_38_629 ();
 FILLCELL_X1 FILLER_38_633 ();
 FILLCELL_X8 FILLER_38_640 ();
 FILLCELL_X4 FILLER_38_648 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X16 FILLER_39_97 ();
 FILLCELL_X4 FILLER_39_113 ();
 FILLCELL_X1 FILLER_39_117 ();
 FILLCELL_X8 FILLER_39_516 ();
 FILLCELL_X4 FILLER_39_530 ();
 FILLCELL_X4 FILLER_39_551 ();
 FILLCELL_X4 FILLER_39_562 ();
 FILLCELL_X4 FILLER_39_569 ();
 FILLCELL_X4 FILLER_39_583 ();
 FILLCELL_X2 FILLER_39_587 ();
 FILLCELL_X4 FILLER_39_593 ();
 FILLCELL_X4 FILLER_39_599 ();
 FILLCELL_X4 FILLER_39_609 ();
 FILLCELL_X4 FILLER_39_616 ();
 FILLCELL_X1 FILLER_39_620 ();
 FILLCELL_X8 FILLER_39_624 ();
 FILLCELL_X2 FILLER_39_632 ();
 FILLCELL_X8 FILLER_39_638 ();
 FILLCELL_X4 FILLER_39_646 ();
 FILLCELL_X2 FILLER_39_650 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X16 FILLER_40_97 ();
 FILLCELL_X4 FILLER_40_113 ();
 FILLCELL_X1 FILLER_40_117 ();
 FILLCELL_X8 FILLER_40_516 ();
 FILLCELL_X1 FILLER_40_524 ();
 FILLCELL_X4 FILLER_40_529 ();
 FILLCELL_X4 FILLER_40_539 ();
 FILLCELL_X8 FILLER_40_547 ();
 FILLCELL_X4 FILLER_40_555 ();
 FILLCELL_X4 FILLER_40_561 ();
 FILLCELL_X4 FILLER_40_575 ();
 FILLCELL_X2 FILLER_40_579 ();
 FILLCELL_X8 FILLER_40_585 ();
 FILLCELL_X2 FILLER_40_593 ();
 FILLCELL_X1 FILLER_40_595 ();
 FILLCELL_X8 FILLER_40_602 ();
 FILLCELL_X1 FILLER_40_610 ();
 FILLCELL_X4 FILLER_40_615 ();
 FILLCELL_X4 FILLER_40_626 ();
 FILLCELL_X4 FILLER_40_647 ();
 FILLCELL_X1 FILLER_40_651 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X4 FILLER_41_97 ();
 FILLCELL_X2 FILLER_41_101 ();
 FILLCELL_X1 FILLER_41_103 ();
 FILLCELL_X4 FILLER_41_106 ();
 FILLCELL_X4 FILLER_41_114 ();
 FILLCELL_X8 FILLER_41_516 ();
 FILLCELL_X1 FILLER_41_524 ();
 FILLCELL_X8 FILLER_41_531 ();
 FILLCELL_X2 FILLER_41_539 ();
 FILLCELL_X4 FILLER_41_548 ();
 FILLCELL_X2 FILLER_41_552 ();
 FILLCELL_X4 FILLER_41_560 ();
 FILLCELL_X4 FILLER_41_567 ();
 FILLCELL_X8 FILLER_41_574 ();
 FILLCELL_X2 FILLER_41_582 ();
 FILLCELL_X4 FILLER_41_588 ();
 FILLCELL_X16 FILLER_41_599 ();
 FILLCELL_X1 FILLER_41_615 ();
 FILLCELL_X4 FILLER_41_622 ();
 FILLCELL_X8 FILLER_41_632 ();
 FILLCELL_X4 FILLER_41_640 ();
 FILLCELL_X1 FILLER_41_644 ();
 FILLCELL_X4 FILLER_41_648 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X16 FILLER_42_65 ();
 FILLCELL_X4 FILLER_42_81 ();
 FILLCELL_X2 FILLER_42_85 ();
 FILLCELL_X1 FILLER_42_87 ();
 FILLCELL_X4 FILLER_42_93 ();
 FILLCELL_X4 FILLER_42_114 ();
 FILLCELL_X32 FILLER_42_516 ();
 FILLCELL_X2 FILLER_42_548 ();
 FILLCELL_X1 FILLER_42_550 ();
 FILLCELL_X4 FILLER_42_557 ();
 FILLCELL_X4 FILLER_42_568 ();
 FILLCELL_X4 FILLER_42_582 ();
 FILLCELL_X16 FILLER_42_592 ();
 FILLCELL_X8 FILLER_42_608 ();
 FILLCELL_X4 FILLER_42_616 ();
 FILLCELL_X2 FILLER_42_620 ();
 FILLCELL_X16 FILLER_42_626 ();
 FILLCELL_X8 FILLER_42_642 ();
 FILLCELL_X2 FILLER_42_650 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X8 FILLER_43_65 ();
 FILLCELL_X4 FILLER_43_73 ();
 FILLCELL_X2 FILLER_43_77 ();
 FILLCELL_X4 FILLER_43_96 ();
 FILLCELL_X2 FILLER_43_100 ();
 FILLCELL_X4 FILLER_43_105 ();
 FILLCELL_X4 FILLER_43_112 ();
 FILLCELL_X2 FILLER_43_116 ();
 FILLCELL_X16 FILLER_43_516 ();
 FILLCELL_X1 FILLER_43_532 ();
 FILLCELL_X32 FILLER_43_537 ();
 FILLCELL_X32 FILLER_43_569 ();
 FILLCELL_X16 FILLER_43_601 ();
 FILLCELL_X4 FILLER_43_617 ();
 FILLCELL_X1 FILLER_43_621 ();
 FILLCELL_X8 FILLER_43_641 ();
 FILLCELL_X2 FILLER_43_649 ();
 FILLCELL_X1 FILLER_43_651 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X16 FILLER_44_33 ();
 FILLCELL_X8 FILLER_44_49 ();
 FILLCELL_X4 FILLER_44_57 ();
 FILLCELL_X4 FILLER_44_64 ();
 FILLCELL_X1 FILLER_44_68 ();
 FILLCELL_X4 FILLER_44_72 ();
 FILLCELL_X4 FILLER_44_79 ();
 FILLCELL_X4 FILLER_44_102 ();
 FILLCELL_X8 FILLER_44_110 ();
 FILLCELL_X8 FILLER_44_516 ();
 FILLCELL_X4 FILLER_44_524 ();
 FILLCELL_X2 FILLER_44_528 ();
 FILLCELL_X1 FILLER_44_530 ();
 FILLCELL_X4 FILLER_44_548 ();
 FILLCELL_X2 FILLER_44_552 ();
 FILLCELL_X1 FILLER_44_554 ();
 FILLCELL_X32 FILLER_44_559 ();
 FILLCELL_X32 FILLER_44_591 ();
 FILLCELL_X16 FILLER_44_623 ();
 FILLCELL_X8 FILLER_44_639 ();
 FILLCELL_X4 FILLER_44_647 ();
 FILLCELL_X1 FILLER_44_651 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X16 FILLER_45_33 ();
 FILLCELL_X8 FILLER_45_49 ();
 FILLCELL_X2 FILLER_45_57 ();
 FILLCELL_X4 FILLER_45_63 ();
 FILLCELL_X8 FILLER_45_72 ();
 FILLCELL_X4 FILLER_45_83 ();
 FILLCELL_X4 FILLER_45_90 ();
 FILLCELL_X4 FILLER_45_99 ();
 FILLCELL_X4 FILLER_45_106 ();
 FILLCELL_X4 FILLER_45_113 ();
 FILLCELL_X1 FILLER_45_117 ();
 FILLCELL_X32 FILLER_45_516 ();
 FILLCELL_X4 FILLER_45_548 ();
 FILLCELL_X2 FILLER_45_552 ();
 FILLCELL_X32 FILLER_45_571 ();
 FILLCELL_X32 FILLER_45_603 ();
 FILLCELL_X16 FILLER_45_635 ();
 FILLCELL_X1 FILLER_45_651 ();
 FILLCELL_X4 FILLER_46_1 ();
 FILLCELL_X32 FILLER_46_9 ();
 FILLCELL_X4 FILLER_46_44 ();
 FILLCELL_X4 FILLER_46_65 ();
 FILLCELL_X4 FILLER_46_74 ();
 FILLCELL_X2 FILLER_46_78 ();
 FILLCELL_X4 FILLER_46_83 ();
 FILLCELL_X4 FILLER_46_106 ();
 FILLCELL_X4 FILLER_46_113 ();
 FILLCELL_X1 FILLER_46_117 ();
 FILLCELL_X16 FILLER_46_516 ();
 FILLCELL_X8 FILLER_46_532 ();
 FILLCELL_X4 FILLER_46_540 ();
 FILLCELL_X2 FILLER_46_544 ();
 FILLCELL_X1 FILLER_46_546 ();
 FILLCELL_X32 FILLER_46_564 ();
 FILLCELL_X32 FILLER_46_596 ();
 FILLCELL_X16 FILLER_46_628 ();
 FILLCELL_X8 FILLER_46_644 ();
 FILLCELL_X16 FILLER_47_1 ();
 FILLCELL_X8 FILLER_47_17 ();
 FILLCELL_X4 FILLER_47_25 ();
 FILLCELL_X4 FILLER_47_31 ();
 FILLCELL_X4 FILLER_47_38 ();
 FILLCELL_X4 FILLER_47_45 ();
 FILLCELL_X8 FILLER_47_66 ();
 FILLCELL_X1 FILLER_47_74 ();
 FILLCELL_X8 FILLER_47_80 ();
 FILLCELL_X1 FILLER_47_88 ();
 FILLCELL_X8 FILLER_47_93 ();
 FILLCELL_X8 FILLER_47_110 ();
 FILLCELL_X32 FILLER_47_516 ();
 FILLCELL_X32 FILLER_47_548 ();
 FILLCELL_X32 FILLER_47_580 ();
 FILLCELL_X32 FILLER_47_612 ();
 FILLCELL_X8 FILLER_47_644 ();
 FILLCELL_X32 FILLER_48_1 ();
 FILLCELL_X8 FILLER_48_33 ();
 FILLCELL_X1 FILLER_48_41 ();
 FILLCELL_X4 FILLER_48_45 ();
 FILLCELL_X4 FILLER_48_53 ();
 FILLCELL_X4 FILLER_48_62 ();
 FILLCELL_X4 FILLER_48_71 ();
 FILLCELL_X4 FILLER_48_78 ();
 FILLCELL_X4 FILLER_48_86 ();
 FILLCELL_X4 FILLER_48_95 ();
 FILLCELL_X4 FILLER_48_104 ();
 FILLCELL_X4 FILLER_48_111 ();
 FILLCELL_X2 FILLER_48_115 ();
 FILLCELL_X1 FILLER_48_117 ();
 FILLCELL_X32 FILLER_48_516 ();
 FILLCELL_X32 FILLER_48_548 ();
 FILLCELL_X32 FILLER_48_580 ();
 FILLCELL_X32 FILLER_48_612 ();
 FILLCELL_X8 FILLER_48_644 ();
 FILLCELL_X32 FILLER_49_1 ();
 FILLCELL_X8 FILLER_49_33 ();
 FILLCELL_X4 FILLER_49_41 ();
 FILLCELL_X1 FILLER_49_45 ();
 FILLCELL_X4 FILLER_49_49 ();
 FILLCELL_X4 FILLER_49_56 ();
 FILLCELL_X8 FILLER_49_65 ();
 FILLCELL_X4 FILLER_49_77 ();
 FILLCELL_X4 FILLER_49_84 ();
 FILLCELL_X4 FILLER_49_91 ();
 FILLCELL_X2 FILLER_49_95 ();
 FILLCELL_X4 FILLER_49_100 ();
 FILLCELL_X2 FILLER_49_104 ();
 FILLCELL_X4 FILLER_49_108 ();
 FILLCELL_X4 FILLER_49_114 ();
 FILLCELL_X32 FILLER_49_516 ();
 FILLCELL_X32 FILLER_49_548 ();
 FILLCELL_X32 FILLER_49_580 ();
 FILLCELL_X32 FILLER_49_612 ();
 FILLCELL_X8 FILLER_49_644 ();
 FILLCELL_X32 FILLER_50_1 ();
 FILLCELL_X8 FILLER_50_33 ();
 FILLCELL_X2 FILLER_50_41 ();
 FILLCELL_X1 FILLER_50_43 ();
 FILLCELL_X4 FILLER_50_48 ();
 FILLCELL_X4 FILLER_50_56 ();
 FILLCELL_X4 FILLER_50_65 ();
 FILLCELL_X8 FILLER_50_74 ();
 FILLCELL_X2 FILLER_50_82 ();
 FILLCELL_X4 FILLER_50_87 ();
 FILLCELL_X8 FILLER_50_94 ();
 FILLCELL_X1 FILLER_50_102 ();
 FILLCELL_X4 FILLER_50_107 ();
 FILLCELL_X4 FILLER_50_114 ();
 FILLCELL_X32 FILLER_50_516 ();
 FILLCELL_X32 FILLER_50_548 ();
 FILLCELL_X32 FILLER_50_580 ();
 FILLCELL_X32 FILLER_50_612 ();
 FILLCELL_X8 FILLER_50_644 ();
 FILLCELL_X32 FILLER_51_1 ();
 FILLCELL_X8 FILLER_51_33 ();
 FILLCELL_X2 FILLER_51_41 ();
 FILLCELL_X1 FILLER_51_43 ();
 FILLCELL_X4 FILLER_51_48 ();
 FILLCELL_X4 FILLER_51_71 ();
 FILLCELL_X8 FILLER_51_80 ();
 FILLCELL_X1 FILLER_51_88 ();
 FILLCELL_X4 FILLER_51_93 ();
 FILLCELL_X4 FILLER_51_101 ();
 FILLCELL_X2 FILLER_51_105 ();
 FILLCELL_X1 FILLER_51_107 ();
 FILLCELL_X4 FILLER_51_112 ();
 FILLCELL_X2 FILLER_51_116 ();
 FILLCELL_X32 FILLER_51_516 ();
 FILLCELL_X32 FILLER_51_548 ();
 FILLCELL_X32 FILLER_51_580 ();
 FILLCELL_X32 FILLER_51_612 ();
 FILLCELL_X8 FILLER_51_644 ();
 FILLCELL_X32 FILLER_52_1 ();
 FILLCELL_X16 FILLER_52_33 ();
 FILLCELL_X1 FILLER_52_49 ();
 FILLCELL_X8 FILLER_52_69 ();
 FILLCELL_X4 FILLER_52_82 ();
 FILLCELL_X4 FILLER_52_92 ();
 FILLCELL_X4 FILLER_52_113 ();
 FILLCELL_X1 FILLER_52_117 ();
 FILLCELL_X32 FILLER_52_516 ();
 FILLCELL_X32 FILLER_52_548 ();
 FILLCELL_X32 FILLER_52_580 ();
 FILLCELL_X32 FILLER_52_612 ();
 FILLCELL_X8 FILLER_52_644 ();
 FILLCELL_X32 FILLER_53_1 ();
 FILLCELL_X8 FILLER_53_33 ();
 FILLCELL_X2 FILLER_53_41 ();
 FILLCELL_X1 FILLER_53_43 ();
 FILLCELL_X4 FILLER_53_46 ();
 FILLCELL_X4 FILLER_53_53 ();
 FILLCELL_X4 FILLER_53_60 ();
 FILLCELL_X4 FILLER_53_67 ();
 FILLCELL_X4 FILLER_53_76 ();
 FILLCELL_X2 FILLER_53_80 ();
 FILLCELL_X1 FILLER_53_82 ();
 FILLCELL_X4 FILLER_53_102 ();
 FILLCELL_X2 FILLER_53_106 ();
 FILLCELL_X1 FILLER_53_108 ();
 FILLCELL_X4 FILLER_53_112 ();
 FILLCELL_X2 FILLER_53_116 ();
 FILLCELL_X32 FILLER_53_516 ();
 FILLCELL_X32 FILLER_53_548 ();
 FILLCELL_X32 FILLER_53_580 ();
 FILLCELL_X32 FILLER_53_612 ();
 FILLCELL_X8 FILLER_53_644 ();
 FILLCELL_X32 FILLER_54_1 ();
 FILLCELL_X16 FILLER_54_33 ();
 FILLCELL_X4 FILLER_54_49 ();
 FILLCELL_X2 FILLER_54_53 ();
 FILLCELL_X4 FILLER_54_58 ();
 FILLCELL_X4 FILLER_54_65 ();
 FILLCELL_X4 FILLER_54_72 ();
 FILLCELL_X4 FILLER_54_79 ();
 FILLCELL_X4 FILLER_54_86 ();
 FILLCELL_X4 FILLER_54_95 ();
 FILLCELL_X2 FILLER_54_99 ();
 FILLCELL_X4 FILLER_54_107 ();
 FILLCELL_X4 FILLER_54_114 ();
 FILLCELL_X32 FILLER_54_516 ();
 FILLCELL_X32 FILLER_54_548 ();
 FILLCELL_X32 FILLER_54_580 ();
 FILLCELL_X32 FILLER_54_612 ();
 FILLCELL_X8 FILLER_54_644 ();
 FILLCELL_X32 FILLER_55_1 ();
 FILLCELL_X16 FILLER_55_33 ();
 FILLCELL_X4 FILLER_55_49 ();
 FILLCELL_X2 FILLER_55_53 ();
 FILLCELL_X1 FILLER_55_55 ();
 FILLCELL_X4 FILLER_55_59 ();
 FILLCELL_X4 FILLER_55_66 ();
 FILLCELL_X4 FILLER_55_73 ();
 FILLCELL_X4 FILLER_55_80 ();
 FILLCELL_X8 FILLER_55_101 ();
 FILLCELL_X4 FILLER_55_114 ();
 FILLCELL_X32 FILLER_55_516 ();
 FILLCELL_X32 FILLER_55_548 ();
 FILLCELL_X32 FILLER_55_580 ();
 FILLCELL_X32 FILLER_55_612 ();
 FILLCELL_X8 FILLER_55_644 ();
 FILLCELL_X32 FILLER_56_1 ();
 FILLCELL_X32 FILLER_56_33 ();
 FILLCELL_X1 FILLER_56_65 ();
 FILLCELL_X4 FILLER_56_69 ();
 FILLCELL_X2 FILLER_56_73 ();
 FILLCELL_X1 FILLER_56_75 ();
 FILLCELL_X4 FILLER_56_79 ();
 FILLCELL_X4 FILLER_56_100 ();
 FILLCELL_X8 FILLER_56_110 ();
 FILLCELL_X32 FILLER_56_516 ();
 FILLCELL_X32 FILLER_56_548 ();
 FILLCELL_X32 FILLER_56_580 ();
 FILLCELL_X32 FILLER_56_612 ();
 FILLCELL_X8 FILLER_56_644 ();
 FILLCELL_X32 FILLER_57_1 ();
 FILLCELL_X32 FILLER_57_33 ();
 FILLCELL_X16 FILLER_57_65 ();
 FILLCELL_X1 FILLER_57_81 ();
 FILLCELL_X4 FILLER_57_85 ();
 FILLCELL_X4 FILLER_57_92 ();
 FILLCELL_X8 FILLER_57_102 ();
 FILLCELL_X1 FILLER_57_110 ();
 FILLCELL_X4 FILLER_57_114 ();
 FILLCELL_X32 FILLER_57_516 ();
 FILLCELL_X32 FILLER_57_548 ();
 FILLCELL_X32 FILLER_57_580 ();
 FILLCELL_X32 FILLER_57_612 ();
 FILLCELL_X8 FILLER_57_644 ();
 FILLCELL_X32 FILLER_58_1 ();
 FILLCELL_X32 FILLER_58_33 ();
 FILLCELL_X16 FILLER_58_65 ();
 FILLCELL_X2 FILLER_58_81 ();
 FILLCELL_X1 FILLER_58_83 ();
 FILLCELL_X4 FILLER_58_86 ();
 FILLCELL_X2 FILLER_58_90 ();
 FILLCELL_X4 FILLER_58_95 ();
 FILLCELL_X4 FILLER_58_102 ();
 FILLCELL_X8 FILLER_58_109 ();
 FILLCELL_X1 FILLER_58_117 ();
 FILLCELL_X32 FILLER_58_516 ();
 FILLCELL_X32 FILLER_58_548 ();
 FILLCELL_X32 FILLER_58_580 ();
 FILLCELL_X32 FILLER_58_612 ();
 FILLCELL_X8 FILLER_58_644 ();
 FILLCELL_X4 FILLER_59_1 ();
 FILLCELL_X32 FILLER_59_8 ();
 FILLCELL_X32 FILLER_59_40 ();
 FILLCELL_X16 FILLER_59_72 ();
 FILLCELL_X4 FILLER_59_88 ();
 FILLCELL_X2 FILLER_59_92 ();
 FILLCELL_X4 FILLER_59_97 ();
 FILLCELL_X4 FILLER_59_104 ();
 FILLCELL_X1 FILLER_59_108 ();
 FILLCELL_X4 FILLER_59_112 ();
 FILLCELL_X2 FILLER_59_116 ();
 FILLCELL_X32 FILLER_59_516 ();
 FILLCELL_X32 FILLER_59_548 ();
 FILLCELL_X32 FILLER_59_580 ();
 FILLCELL_X32 FILLER_59_612 ();
 FILLCELL_X8 FILLER_59_644 ();
 FILLCELL_X32 FILLER_60_1 ();
 FILLCELL_X32 FILLER_60_33 ();
 FILLCELL_X32 FILLER_60_65 ();
 FILLCELL_X4 FILLER_60_97 ();
 FILLCELL_X2 FILLER_60_101 ();
 FILLCELL_X1 FILLER_60_103 ();
 FILLCELL_X4 FILLER_60_107 ();
 FILLCELL_X4 FILLER_60_114 ();
 FILLCELL_X32 FILLER_60_516 ();
 FILLCELL_X32 FILLER_60_548 ();
 FILLCELL_X32 FILLER_60_580 ();
 FILLCELL_X32 FILLER_60_612 ();
 FILLCELL_X8 FILLER_60_644 ();
 FILLCELL_X32 FILLER_61_1 ();
 FILLCELL_X32 FILLER_61_33 ();
 FILLCELL_X32 FILLER_61_65 ();
 FILLCELL_X8 FILLER_61_97 ();
 FILLCELL_X4 FILLER_61_105 ();
 FILLCELL_X2 FILLER_61_109 ();
 FILLCELL_X4 FILLER_61_114 ();
 FILLCELL_X32 FILLER_61_516 ();
 FILLCELL_X32 FILLER_61_548 ();
 FILLCELL_X32 FILLER_61_580 ();
 FILLCELL_X32 FILLER_61_612 ();
 FILLCELL_X8 FILLER_61_644 ();
 FILLCELL_X32 FILLER_62_1 ();
 FILLCELL_X32 FILLER_62_33 ();
 FILLCELL_X32 FILLER_62_65 ();
 FILLCELL_X8 FILLER_62_97 ();
 FILLCELL_X1 FILLER_62_105 ();
 FILLCELL_X8 FILLER_62_109 ();
 FILLCELL_X1 FILLER_62_117 ();
 FILLCELL_X32 FILLER_62_516 ();
 FILLCELL_X32 FILLER_62_548 ();
 FILLCELL_X32 FILLER_62_580 ();
 FILLCELL_X32 FILLER_62_612 ();
 FILLCELL_X8 FILLER_62_644 ();
 FILLCELL_X32 FILLER_63_1 ();
 FILLCELL_X32 FILLER_63_33 ();
 FILLCELL_X32 FILLER_63_65 ();
 FILLCELL_X16 FILLER_63_97 ();
 FILLCELL_X4 FILLER_63_113 ();
 FILLCELL_X1 FILLER_63_117 ();
 FILLCELL_X32 FILLER_63_516 ();
 FILLCELL_X32 FILLER_63_548 ();
 FILLCELL_X32 FILLER_63_580 ();
 FILLCELL_X32 FILLER_63_612 ();
 FILLCELL_X8 FILLER_63_644 ();
 FILLCELL_X32 FILLER_64_1 ();
 FILLCELL_X32 FILLER_64_33 ();
 FILLCELL_X32 FILLER_64_65 ();
 FILLCELL_X8 FILLER_64_97 ();
 FILLCELL_X4 FILLER_64_105 ();
 FILLCELL_X2 FILLER_64_109 ();
 FILLCELL_X4 FILLER_64_114 ();
 FILLCELL_X32 FILLER_64_516 ();
 FILLCELL_X32 FILLER_64_548 ();
 FILLCELL_X32 FILLER_64_580 ();
 FILLCELL_X32 FILLER_64_612 ();
 FILLCELL_X8 FILLER_64_644 ();
 FILLCELL_X32 FILLER_65_1 ();
 FILLCELL_X32 FILLER_65_33 ();
 FILLCELL_X32 FILLER_65_65 ();
 FILLCELL_X8 FILLER_65_97 ();
 FILLCELL_X4 FILLER_65_105 ();
 FILLCELL_X2 FILLER_65_109 ();
 FILLCELL_X4 FILLER_65_114 ();
 FILLCELL_X32 FILLER_65_516 ();
 FILLCELL_X32 FILLER_65_548 ();
 FILLCELL_X32 FILLER_65_580 ();
 FILLCELL_X32 FILLER_65_612 ();
 FILLCELL_X8 FILLER_65_644 ();
 FILLCELL_X32 FILLER_66_1 ();
 FILLCELL_X32 FILLER_66_33 ();
 FILLCELL_X32 FILLER_66_65 ();
 FILLCELL_X16 FILLER_66_97 ();
 FILLCELL_X4 FILLER_66_113 ();
 FILLCELL_X1 FILLER_66_117 ();
 FILLCELL_X32 FILLER_66_516 ();
 FILLCELL_X32 FILLER_66_548 ();
 FILLCELL_X32 FILLER_66_580 ();
 FILLCELL_X32 FILLER_66_612 ();
 FILLCELL_X1 FILLER_66_644 ();
 FILLCELL_X4 FILLER_66_648 ();
 FILLCELL_X32 FILLER_67_1 ();
 FILLCELL_X32 FILLER_67_33 ();
 FILLCELL_X32 FILLER_67_65 ();
 FILLCELL_X8 FILLER_67_97 ();
 FILLCELL_X4 FILLER_67_105 ();
 FILLCELL_X2 FILLER_67_109 ();
 FILLCELL_X4 FILLER_67_114 ();
 FILLCELL_X32 FILLER_67_516 ();
 FILLCELL_X32 FILLER_67_548 ();
 FILLCELL_X32 FILLER_67_580 ();
 FILLCELL_X32 FILLER_67_612 ();
 FILLCELL_X8 FILLER_67_644 ();
 FILLCELL_X32 FILLER_68_1 ();
 FILLCELL_X32 FILLER_68_33 ();
 FILLCELL_X32 FILLER_68_65 ();
 FILLCELL_X16 FILLER_68_97 ();
 FILLCELL_X4 FILLER_68_113 ();
 FILLCELL_X1 FILLER_68_117 ();
 FILLCELL_X32 FILLER_68_516 ();
 FILLCELL_X32 FILLER_68_548 ();
 FILLCELL_X32 FILLER_68_580 ();
 FILLCELL_X32 FILLER_68_612 ();
 FILLCELL_X8 FILLER_68_644 ();
 FILLCELL_X32 FILLER_69_1 ();
 FILLCELL_X32 FILLER_69_33 ();
 FILLCELL_X32 FILLER_69_65 ();
 FILLCELL_X16 FILLER_69_97 ();
 FILLCELL_X4 FILLER_69_113 ();
 FILLCELL_X1 FILLER_69_117 ();
 FILLCELL_X32 FILLER_69_516 ();
 FILLCELL_X32 FILLER_69_548 ();
 FILLCELL_X32 FILLER_69_580 ();
 FILLCELL_X32 FILLER_69_612 ();
 FILLCELL_X8 FILLER_69_644 ();
 FILLCELL_X32 FILLER_70_1 ();
 FILLCELL_X32 FILLER_70_33 ();
 FILLCELL_X32 FILLER_70_65 ();
 FILLCELL_X16 FILLER_70_97 ();
 FILLCELL_X4 FILLER_70_113 ();
 FILLCELL_X1 FILLER_70_117 ();
 FILLCELL_X32 FILLER_70_516 ();
 FILLCELL_X32 FILLER_70_548 ();
 FILLCELL_X32 FILLER_70_580 ();
 FILLCELL_X32 FILLER_70_612 ();
 FILLCELL_X8 FILLER_70_644 ();
 FILLCELL_X32 FILLER_71_1 ();
 FILLCELL_X32 FILLER_71_33 ();
 FILLCELL_X32 FILLER_71_65 ();
 FILLCELL_X8 FILLER_71_97 ();
 FILLCELL_X4 FILLER_71_105 ();
 FILLCELL_X2 FILLER_71_109 ();
 FILLCELL_X4 FILLER_71_114 ();
 FILLCELL_X32 FILLER_71_516 ();
 FILLCELL_X32 FILLER_71_548 ();
 FILLCELL_X32 FILLER_71_580 ();
 FILLCELL_X32 FILLER_71_612 ();
 FILLCELL_X8 FILLER_71_644 ();
 FILLCELL_X4 FILLER_72_1 ();
 FILLCELL_X32 FILLER_72_9 ();
 FILLCELL_X32 FILLER_72_41 ();
 FILLCELL_X32 FILLER_72_73 ();
 FILLCELL_X8 FILLER_72_105 ();
 FILLCELL_X4 FILLER_72_113 ();
 FILLCELL_X1 FILLER_72_117 ();
 FILLCELL_X32 FILLER_72_516 ();
 FILLCELL_X32 FILLER_72_548 ();
 FILLCELL_X32 FILLER_72_580 ();
 FILLCELL_X32 FILLER_72_612 ();
 FILLCELL_X8 FILLER_72_644 ();
 FILLCELL_X32 FILLER_73_1 ();
 FILLCELL_X32 FILLER_73_33 ();
 FILLCELL_X32 FILLER_73_65 ();
 FILLCELL_X16 FILLER_73_97 ();
 FILLCELL_X4 FILLER_73_113 ();
 FILLCELL_X1 FILLER_73_117 ();
 FILLCELL_X32 FILLER_73_516 ();
 FILLCELL_X32 FILLER_73_548 ();
 FILLCELL_X32 FILLER_73_580 ();
 FILLCELL_X32 FILLER_73_612 ();
 FILLCELL_X8 FILLER_73_644 ();
 FILLCELL_X32 FILLER_74_1 ();
 FILLCELL_X32 FILLER_74_33 ();
 FILLCELL_X32 FILLER_74_65 ();
 FILLCELL_X16 FILLER_74_97 ();
 FILLCELL_X4 FILLER_74_113 ();
 FILLCELL_X1 FILLER_74_117 ();
 FILLCELL_X32 FILLER_74_516 ();
 FILLCELL_X32 FILLER_74_548 ();
 FILLCELL_X32 FILLER_74_580 ();
 FILLCELL_X32 FILLER_74_612 ();
 FILLCELL_X8 FILLER_74_644 ();
 FILLCELL_X32 FILLER_75_1 ();
 FILLCELL_X32 FILLER_75_33 ();
 FILLCELL_X32 FILLER_75_65 ();
 FILLCELL_X16 FILLER_75_97 ();
 FILLCELL_X4 FILLER_75_113 ();
 FILLCELL_X1 FILLER_75_117 ();
 FILLCELL_X32 FILLER_75_516 ();
 FILLCELL_X32 FILLER_75_548 ();
 FILLCELL_X32 FILLER_75_580 ();
 FILLCELL_X32 FILLER_75_612 ();
 FILLCELL_X8 FILLER_75_644 ();
 FILLCELL_X32 FILLER_76_1 ();
 FILLCELL_X32 FILLER_76_33 ();
 FILLCELL_X32 FILLER_76_65 ();
 FILLCELL_X16 FILLER_76_97 ();
 FILLCELL_X4 FILLER_76_113 ();
 FILLCELL_X1 FILLER_76_117 ();
 FILLCELL_X32 FILLER_76_516 ();
 FILLCELL_X32 FILLER_76_548 ();
 FILLCELL_X32 FILLER_76_580 ();
 FILLCELL_X32 FILLER_76_612 ();
 FILLCELL_X8 FILLER_76_644 ();
 FILLCELL_X32 FILLER_77_1 ();
 FILLCELL_X32 FILLER_77_33 ();
 FILLCELL_X32 FILLER_77_65 ();
 FILLCELL_X16 FILLER_77_97 ();
 FILLCELL_X4 FILLER_77_113 ();
 FILLCELL_X1 FILLER_77_117 ();
 FILLCELL_X32 FILLER_77_516 ();
 FILLCELL_X32 FILLER_77_548 ();
 FILLCELL_X32 FILLER_77_580 ();
 FILLCELL_X32 FILLER_77_612 ();
 FILLCELL_X8 FILLER_77_644 ();
 FILLCELL_X32 FILLER_78_1 ();
 FILLCELL_X32 FILLER_78_33 ();
 FILLCELL_X32 FILLER_78_65 ();
 FILLCELL_X16 FILLER_78_97 ();
 FILLCELL_X4 FILLER_78_113 ();
 FILLCELL_X1 FILLER_78_117 ();
 FILLCELL_X32 FILLER_78_516 ();
 FILLCELL_X32 FILLER_78_548 ();
 FILLCELL_X32 FILLER_78_580 ();
 FILLCELL_X32 FILLER_78_612 ();
 FILLCELL_X1 FILLER_78_644 ();
 FILLCELL_X4 FILLER_78_648 ();
 FILLCELL_X32 FILLER_79_1 ();
 FILLCELL_X32 FILLER_79_33 ();
 FILLCELL_X32 FILLER_79_65 ();
 FILLCELL_X32 FILLER_79_97 ();
 FILLCELL_X32 FILLER_79_129 ();
 FILLCELL_X32 FILLER_79_161 ();
 FILLCELL_X32 FILLER_79_193 ();
 FILLCELL_X32 FILLER_79_225 ();
 FILLCELL_X32 FILLER_79_257 ();
 FILLCELL_X32 FILLER_79_289 ();
 FILLCELL_X32 FILLER_79_321 ();
 FILLCELL_X32 FILLER_79_353 ();
 FILLCELL_X32 FILLER_79_385 ();
 FILLCELL_X32 FILLER_79_417 ();
 FILLCELL_X32 FILLER_79_449 ();
 FILLCELL_X32 FILLER_79_481 ();
 FILLCELL_X32 FILLER_79_513 ();
 FILLCELL_X32 FILLER_79_545 ();
 FILLCELL_X32 FILLER_79_577 ();
 FILLCELL_X16 FILLER_79_609 ();
 FILLCELL_X4 FILLER_79_625 ();
 FILLCELL_X2 FILLER_79_629 ();
 FILLCELL_X16 FILLER_79_632 ();
 FILLCELL_X4 FILLER_79_648 ();
 FILLCELL_X32 FILLER_80_1 ();
 FILLCELL_X32 FILLER_80_33 ();
 FILLCELL_X32 FILLER_80_65 ();
 FILLCELL_X32 FILLER_80_97 ();
 FILLCELL_X32 FILLER_80_129 ();
 FILLCELL_X32 FILLER_80_161 ();
 FILLCELL_X32 FILLER_80_193 ();
 FILLCELL_X32 FILLER_80_225 ();
 FILLCELL_X32 FILLER_80_257 ();
 FILLCELL_X32 FILLER_80_289 ();
 FILLCELL_X32 FILLER_80_321 ();
 FILLCELL_X32 FILLER_80_353 ();
 FILLCELL_X32 FILLER_80_385 ();
 FILLCELL_X32 FILLER_80_417 ();
 FILLCELL_X32 FILLER_80_449 ();
 FILLCELL_X32 FILLER_80_481 ();
 FILLCELL_X32 FILLER_80_513 ();
 FILLCELL_X32 FILLER_80_545 ();
 FILLCELL_X32 FILLER_80_577 ();
 FILLCELL_X16 FILLER_80_609 ();
 FILLCELL_X4 FILLER_80_625 ();
 FILLCELL_X2 FILLER_80_629 ();
 FILLCELL_X16 FILLER_80_632 ();
 FILLCELL_X4 FILLER_80_648 ();
 FILLCELL_X32 FILLER_81_1 ();
 FILLCELL_X32 FILLER_81_33 ();
 FILLCELL_X32 FILLER_81_65 ();
 FILLCELL_X32 FILLER_81_97 ();
 FILLCELL_X32 FILLER_81_129 ();
 FILLCELL_X32 FILLER_81_161 ();
 FILLCELL_X32 FILLER_81_193 ();
 FILLCELL_X32 FILLER_81_225 ();
 FILLCELL_X32 FILLER_81_257 ();
 FILLCELL_X32 FILLER_81_289 ();
 FILLCELL_X32 FILLER_81_321 ();
 FILLCELL_X32 FILLER_81_353 ();
 FILLCELL_X32 FILLER_81_385 ();
 FILLCELL_X32 FILLER_81_417 ();
 FILLCELL_X32 FILLER_81_449 ();
 FILLCELL_X32 FILLER_81_481 ();
 FILLCELL_X32 FILLER_81_513 ();
 FILLCELL_X32 FILLER_81_545 ();
 FILLCELL_X32 FILLER_81_577 ();
 FILLCELL_X32 FILLER_81_609 ();
 FILLCELL_X8 FILLER_81_641 ();
 FILLCELL_X2 FILLER_81_649 ();
 FILLCELL_X1 FILLER_81_651 ();
 FILLCELL_X32 FILLER_82_1 ();
 FILLCELL_X32 FILLER_82_33 ();
 FILLCELL_X32 FILLER_82_65 ();
 FILLCELL_X32 FILLER_82_97 ();
 FILLCELL_X32 FILLER_82_129 ();
 FILLCELL_X32 FILLER_82_161 ();
 FILLCELL_X32 FILLER_82_193 ();
 FILLCELL_X32 FILLER_82_225 ();
 FILLCELL_X32 FILLER_82_257 ();
 FILLCELL_X32 FILLER_82_289 ();
 FILLCELL_X32 FILLER_82_321 ();
 FILLCELL_X32 FILLER_82_353 ();
 FILLCELL_X32 FILLER_82_385 ();
 FILLCELL_X32 FILLER_82_417 ();
 FILLCELL_X32 FILLER_82_449 ();
 FILLCELL_X32 FILLER_82_481 ();
 FILLCELL_X32 FILLER_82_513 ();
 FILLCELL_X32 FILLER_82_545 ();
 FILLCELL_X32 FILLER_82_577 ();
 FILLCELL_X16 FILLER_82_609 ();
 FILLCELL_X4 FILLER_82_625 ();
 FILLCELL_X2 FILLER_82_629 ();
 FILLCELL_X16 FILLER_82_632 ();
 FILLCELL_X4 FILLER_82_648 ();
 FILLCELL_X32 FILLER_83_1 ();
 FILLCELL_X32 FILLER_83_33 ();
 FILLCELL_X32 FILLER_83_65 ();
 FILLCELL_X32 FILLER_83_97 ();
 FILLCELL_X32 FILLER_83_129 ();
 FILLCELL_X32 FILLER_83_161 ();
 FILLCELL_X32 FILLER_83_193 ();
 FILLCELL_X32 FILLER_83_225 ();
 FILLCELL_X32 FILLER_83_257 ();
 FILLCELL_X32 FILLER_83_289 ();
 FILLCELL_X32 FILLER_83_321 ();
 FILLCELL_X32 FILLER_83_353 ();
 FILLCELL_X32 FILLER_83_385 ();
 FILLCELL_X32 FILLER_83_417 ();
 FILLCELL_X32 FILLER_83_449 ();
 FILLCELL_X32 FILLER_83_481 ();
 FILLCELL_X32 FILLER_83_513 ();
 FILLCELL_X32 FILLER_83_545 ();
 FILLCELL_X32 FILLER_83_577 ();
 FILLCELL_X32 FILLER_83_609 ();
 FILLCELL_X8 FILLER_83_641 ();
 FILLCELL_X2 FILLER_83_649 ();
 FILLCELL_X1 FILLER_83_651 ();
 FILLCELL_X32 FILLER_84_1 ();
 FILLCELL_X32 FILLER_84_33 ();
 FILLCELL_X32 FILLER_84_65 ();
 FILLCELL_X32 FILLER_84_97 ();
 FILLCELL_X32 FILLER_84_129 ();
 FILLCELL_X32 FILLER_84_161 ();
 FILLCELL_X32 FILLER_84_193 ();
 FILLCELL_X32 FILLER_84_225 ();
 FILLCELL_X32 FILLER_84_257 ();
 FILLCELL_X32 FILLER_84_289 ();
 FILLCELL_X32 FILLER_84_321 ();
 FILLCELL_X32 FILLER_84_353 ();
 FILLCELL_X32 FILLER_84_385 ();
 FILLCELL_X32 FILLER_84_417 ();
 FILLCELL_X32 FILLER_84_449 ();
 FILLCELL_X32 FILLER_84_481 ();
 FILLCELL_X32 FILLER_84_513 ();
 FILLCELL_X32 FILLER_84_545 ();
 FILLCELL_X32 FILLER_84_577 ();
 FILLCELL_X16 FILLER_84_609 ();
 FILLCELL_X4 FILLER_84_625 ();
 FILLCELL_X2 FILLER_84_629 ();
 FILLCELL_X16 FILLER_84_632 ();
 FILLCELL_X4 FILLER_84_648 ();
 FILLCELL_X4 FILLER_85_1 ();
 FILLCELL_X32 FILLER_85_18 ();
 FILLCELL_X32 FILLER_85_50 ();
 FILLCELL_X32 FILLER_85_82 ();
 FILLCELL_X32 FILLER_85_114 ();
 FILLCELL_X32 FILLER_85_146 ();
 FILLCELL_X32 FILLER_85_178 ();
 FILLCELL_X32 FILLER_85_210 ();
 FILLCELL_X32 FILLER_85_242 ();
 FILLCELL_X32 FILLER_85_274 ();
 FILLCELL_X32 FILLER_85_306 ();
 FILLCELL_X32 FILLER_85_338 ();
 FILLCELL_X32 FILLER_85_370 ();
 FILLCELL_X32 FILLER_85_402 ();
 FILLCELL_X32 FILLER_85_434 ();
 FILLCELL_X32 FILLER_85_466 ();
 FILLCELL_X32 FILLER_85_498 ();
 FILLCELL_X32 FILLER_85_530 ();
 FILLCELL_X32 FILLER_85_562 ();
 FILLCELL_X32 FILLER_85_594 ();
 FILLCELL_X16 FILLER_85_626 ();
 FILLCELL_X8 FILLER_85_642 ();
 FILLCELL_X2 FILLER_85_650 ();
 FILLCELL_X32 FILLER_86_1 ();
 FILLCELL_X32 FILLER_86_33 ();
 FILLCELL_X32 FILLER_86_65 ();
 FILLCELL_X32 FILLER_86_97 ();
 FILLCELL_X32 FILLER_86_129 ();
 FILLCELL_X32 FILLER_86_161 ();
 FILLCELL_X32 FILLER_86_193 ();
 FILLCELL_X32 FILLER_86_225 ();
 FILLCELL_X32 FILLER_86_257 ();
 FILLCELL_X32 FILLER_86_289 ();
 FILLCELL_X32 FILLER_86_321 ();
 FILLCELL_X32 FILLER_86_353 ();
 FILLCELL_X32 FILLER_86_385 ();
 FILLCELL_X32 FILLER_86_417 ();
 FILLCELL_X32 FILLER_86_449 ();
 FILLCELL_X32 FILLER_86_481 ();
 FILLCELL_X32 FILLER_86_513 ();
 FILLCELL_X32 FILLER_86_545 ();
 FILLCELL_X32 FILLER_86_577 ();
 FILLCELL_X16 FILLER_86_609 ();
 FILLCELL_X4 FILLER_86_625 ();
 FILLCELL_X2 FILLER_86_629 ();
 FILLCELL_X16 FILLER_86_632 ();
 FILLCELL_X4 FILLER_86_648 ();
 FILLCELL_X16 FILLER_87_1 ();
 FILLCELL_X4 FILLER_87_17 ();
 FILLCELL_X32 FILLER_87_24 ();
 FILLCELL_X32 FILLER_87_56 ();
 FILLCELL_X16 FILLER_87_88 ();
 FILLCELL_X8 FILLER_87_104 ();
 FILLCELL_X2 FILLER_87_112 ();
 FILLCELL_X1 FILLER_87_114 ();
 FILLCELL_X32 FILLER_87_118 ();
 FILLCELL_X32 FILLER_87_150 ();
 FILLCELL_X16 FILLER_87_182 ();
 FILLCELL_X8 FILLER_87_198 ();
 FILLCELL_X2 FILLER_87_206 ();
 FILLCELL_X1 FILLER_87_208 ();
 FILLCELL_X32 FILLER_87_213 ();
 FILLCELL_X32 FILLER_87_245 ();
 FILLCELL_X16 FILLER_87_277 ();
 FILLCELL_X8 FILLER_87_293 ();
 FILLCELL_X2 FILLER_87_301 ();
 FILLCELL_X1 FILLER_87_303 ();
 FILLCELL_X32 FILLER_87_307 ();
 FILLCELL_X32 FILLER_87_339 ();
 FILLCELL_X16 FILLER_87_371 ();
 FILLCELL_X4 FILLER_87_387 ();
 FILLCELL_X1 FILLER_87_391 ();
 FILLCELL_X32 FILLER_87_395 ();
 FILLCELL_X32 FILLER_87_427 ();
 FILLCELL_X16 FILLER_87_459 ();
 FILLCELL_X8 FILLER_87_475 ();
 FILLCELL_X2 FILLER_87_483 ();
 FILLCELL_X1 FILLER_87_485 ();
 FILLCELL_X32 FILLER_87_489 ();
 FILLCELL_X32 FILLER_87_521 ();
 FILLCELL_X16 FILLER_87_553 ();
 FILLCELL_X8 FILLER_87_569 ();
 FILLCELL_X4 FILLER_87_577 ();
 FILLCELL_X32 FILLER_87_584 ();
 FILLCELL_X8 FILLER_87_616 ();
 FILLCELL_X4 FILLER_87_624 ();
 FILLCELL_X2 FILLER_87_628 ();
 FILLCELL_X1 FILLER_87_630 ();
 FILLCELL_X8 FILLER_87_632 ();
 FILLCELL_X4 FILLER_87_640 ();
 FILLCELL_X1 FILLER_87_644 ();
 FILLCELL_X4 FILLER_87_648 ();
 assign init_done = curr_state[1];
 assign valid_out = valid_reg_out;
endmodule
