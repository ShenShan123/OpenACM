module sram_multiplier_system (clk,
    init_done,
    init_enable,
    pe_ce,
    rst_n,
    valid_out,
    data_in,
    data_out);
 input clk;
 output init_done;
 input init_enable;
 input pe_ce;
 input rst_n;
 output valid_out;
 input [15:0] data_in;
 output [31:0] data_out;

 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire \u_multiplier/pp_0 ;
 wire \u_multiplier/pp_30 ;
 wire \u_multiplier/s_0 ;
 wire \u_multiplier/s_30 ;
 wire \u_multiplier/STAGE1/_178_ ;
 wire \u_multiplier/STAGE1/_179_ ;
 wire \u_multiplier/STAGE1/_180_ ;
 wire \u_multiplier/STAGE1/_181_ ;
 wire \u_multiplier/STAGE1/_182_ ;
 wire \u_multiplier/STAGE1/_183_ ;
 wire \u_multiplier/STAGE1/_184_ ;
 wire \u_multiplier/STAGE1/_185_ ;
 wire \u_multiplier/STAGE1/_186_ ;
 wire \u_multiplier/STAGE1/_187_ ;
 wire \u_multiplier/STAGE1/_188_ ;
 wire \u_multiplier/STAGE1/_189_ ;
 wire \u_multiplier/STAGE1/_190_ ;
 wire \u_multiplier/STAGE1/_191_ ;
 wire \u_multiplier/STAGE1/_192_ ;
 wire \u_multiplier/STAGE1/_193_ ;
 wire \u_multiplier/STAGE1/_194_ ;
 wire \u_multiplier/STAGE1/_195_ ;
 wire \u_multiplier/STAGE1/_196_ ;
 wire \u_multiplier/STAGE1/_197_ ;
 wire \u_multiplier/STAGE1/_198_ ;
 wire \u_multiplier/STAGE1/_199_ ;
 wire \u_multiplier/STAGE1/_200_ ;
 wire \u_multiplier/STAGE1/_201_ ;
 wire \u_multiplier/STAGE1/_202_ ;
 wire \u_multiplier/STAGE1/_203_ ;
 wire \u_multiplier/STAGE1/_204_ ;
 wire \u_multiplier/STAGE1/_205_ ;
 wire \u_multiplier/STAGE1/_206_ ;
 wire \u_multiplier/STAGE1/_207_ ;
 wire \u_multiplier/STAGE1/_208_ ;
 wire \u_multiplier/STAGE1/_209_ ;
 wire \u_multiplier/STAGE1/_210_ ;
 wire \u_multiplier/STAGE1/_211_ ;
 wire \u_multiplier/STAGE1/_212_ ;
 wire \u_multiplier/STAGE1/_213_ ;
 wire \u_multiplier/STAGE1/_214_ ;
 wire \u_multiplier/STAGE1/_215_ ;
 wire \u_multiplier/STAGE1/_216_ ;
 wire \u_multiplier/STAGE1/_217_ ;
 wire \u_multiplier/STAGE1/_218_ ;
 wire \u_multiplier/STAGE1/_219_ ;
 wire \u_multiplier/STAGE1/_220_ ;
 wire \u_multiplier/STAGE1/_221_ ;
 wire \u_multiplier/STAGE1/_222_ ;
 wire \u_multiplier/STAGE1/_223_ ;
 wire \u_multiplier/STAGE1/_224_ ;
 wire \u_multiplier/STAGE1/_225_ ;
 wire \u_multiplier/STAGE1/_226_ ;
 wire \u_multiplier/STAGE1/_227_ ;
 wire \u_multiplier/STAGE1/_228_ ;
 wire \u_multiplier/STAGE1/_229_ ;
 wire \u_multiplier/STAGE1/_230_ ;
 wire \u_multiplier/STAGE1/_231_ ;
 wire \u_multiplier/STAGE1/_232_ ;
 wire \u_multiplier/STAGE1/_233_ ;
 wire \u_multiplier/STAGE1/_234_ ;
 wire \u_multiplier/STAGE1/_235_ ;
 wire \u_multiplier/STAGE1/_236_ ;
 wire \u_multiplier/STAGE1/_237_ ;
 wire \u_multiplier/STAGE1/_238_ ;
 wire \u_multiplier/STAGE1/_239_ ;
 wire \u_multiplier/STAGE1/_240_ ;
 wire \u_multiplier/STAGE1/_241_ ;
 wire \u_multiplier/STAGE1/_242_ ;
 wire \u_multiplier/STAGE1/_243_ ;
 wire \u_multiplier/STAGE1/_244_ ;
 wire \u_multiplier/STAGE1/_245_ ;
 wire \u_multiplier/STAGE1/_246_ ;
 wire \u_multiplier/STAGE1/_247_ ;
 wire \u_multiplier/STAGE1/_248_ ;
 wire \u_multiplier/STAGE1/_249_ ;
 wire \u_multiplier/STAGE1/_250_ ;
 wire \u_multiplier/STAGE1/_251_ ;
 wire \u_multiplier/STAGE1/_252_ ;
 wire \u_multiplier/STAGE1/_253_ ;
 wire \u_multiplier/STAGE1/_254_ ;
 wire \u_multiplier/STAGE1/_255_ ;
 wire \u_multiplier/STAGE1/_256_ ;
 wire \u_multiplier/STAGE1/_257_ ;
 wire \u_multiplier/STAGE1/_258_ ;
 wire \u_multiplier/STAGE1/_259_ ;
 wire \u_multiplier/STAGE1/_260_ ;
 wire \u_multiplier/STAGE1/_261_ ;
 wire \u_multiplier/STAGE1/_262_ ;
 wire \u_multiplier/STAGE1/_263_ ;
 wire \u_multiplier/STAGE1/_264_ ;
 wire \u_multiplier/STAGE1/_265_ ;
 wire \u_multiplier/STAGE1/_266_ ;
 wire \u_multiplier/STAGE1/_267_ ;
 wire \u_multiplier/STAGE1/_268_ ;
 wire \u_multiplier/STAGE1/_269_ ;
 wire \u_multiplier/STAGE1/_270_ ;
 wire \u_multiplier/STAGE1/_271_ ;
 wire \u_multiplier/STAGE1/_272_ ;
 wire \u_multiplier/STAGE1/_273_ ;
 wire \u_multiplier/STAGE1/_274_ ;
 wire \u_multiplier/STAGE1/_275_ ;
 wire \u_multiplier/STAGE1/_276_ ;
 wire \u_multiplier/STAGE1/_277_ ;
 wire \u_multiplier/STAGE1/_278_ ;
 wire \u_multiplier/STAGE1/_279_ ;
 wire \u_multiplier/STAGE1/_280_ ;
 wire \u_multiplier/STAGE1/_281_ ;
 wire \u_multiplier/STAGE1/_282_ ;
 wire \u_multiplier/STAGE1/_283_ ;
 wire \u_multiplier/STAGE1/_284_ ;
 wire \u_multiplier/STAGE1/_285_ ;
 wire \u_multiplier/STAGE1/_286_ ;
 wire \u_multiplier/STAGE1/_287_ ;
 wire \u_multiplier/STAGE1/_288_ ;
 wire \u_multiplier/STAGE1/_289_ ;
 wire \u_multiplier/STAGE1/_290_ ;
 wire \u_multiplier/STAGE1/_291_ ;
 wire \u_multiplier/STAGE1/_292_ ;
 wire \u_multiplier/STAGE1/_293_ ;
 wire \u_multiplier/STAGE1/_294_ ;
 wire \u_multiplier/STAGE1/_295_ ;
 wire \u_multiplier/STAGE1/_296_ ;
 wire \u_multiplier/STAGE1/_297_ ;
 wire \u_multiplier/STAGE1/_298_ ;
 wire \u_multiplier/STAGE1/_299_ ;
 wire \u_multiplier/STAGE1/_300_ ;
 wire \u_multiplier/STAGE1/_301_ ;
 wire \u_multiplier/STAGE1/_302_ ;
 wire \u_multiplier/STAGE1/_303_ ;
 wire \u_multiplier/STAGE1/_304_ ;
 wire \u_multiplier/STAGE1/_305_ ;
 wire \u_multiplier/STAGE1/_306_ ;
 wire \u_multiplier/STAGE1/_307_ ;
 wire \u_multiplier/STAGE1/_308_ ;
 wire \u_multiplier/STAGE1/_309_ ;
 wire \u_multiplier/STAGE1/_310_ ;
 wire \u_multiplier/STAGE1/_311_ ;
 wire \u_multiplier/STAGE1/_312_ ;
 wire \u_multiplier/STAGE1/_313_ ;
 wire \u_multiplier/STAGE1/_314_ ;
 wire \u_multiplier/STAGE1/_315_ ;
 wire \u_multiplier/STAGE1/_316_ ;
 wire \u_multiplier/STAGE1/_317_ ;
 wire \u_multiplier/STAGE1/_318_ ;
 wire \u_multiplier/STAGE1/_319_ ;
 wire \u_multiplier/STAGE1/_320_ ;
 wire \u_multiplier/STAGE1/_321_ ;
 wire \u_multiplier/STAGE1/_322_ ;
 wire \u_multiplier/STAGE1/_323_ ;
 wire \u_multiplier/STAGE1/pp_10_c2 ;
 wire \u_multiplier/STAGE1/pp_11_c2 ;
 wire \u_multiplier/STAGE1/pp_11_c4 ;
 wire \u_multiplier/STAGE1/pp_12_c2 ;
 wire \u_multiplier/STAGE1/pp_12_c4 ;
 wire \u_multiplier/STAGE1/pp_13_c2 ;
 wire \u_multiplier/STAGE1/pp_13_c4 ;
 wire \u_multiplier/STAGE1/pp_13_c6 ;
 wire \u_multiplier/STAGE1/pp_14_c2 ;
 wire \u_multiplier/STAGE1/pp_14_c4 ;
 wire \u_multiplier/STAGE1/pp_14_c6 ;
 wire \u_multiplier/STAGE1/pp_15_c2 ;
 wire \u_multiplier/STAGE1/pp_15_c4 ;
 wire \u_multiplier/STAGE1/pp_15_c6 ;
 wire \u_multiplier/STAGE1/pp_15_c8 ;
 wire \u_multiplier/STAGE1/pp_16_c2 ;
 wire \u_multiplier/STAGE1/pp_16_c4 ;
 wire \u_multiplier/STAGE1/pp_16_c6 ;
 wire \u_multiplier/STAGE1/pp_16_c8 ;
 wire \u_multiplier/STAGE1/pp_17_c2 ;
 wire \u_multiplier/STAGE1/pp_17_c4 ;
 wire \u_multiplier/STAGE1/pp_17_c6 ;
 wire \u_multiplier/STAGE1/pp_18_c2 ;
 wire \u_multiplier/STAGE1/pp_18_c4 ;
 wire \u_multiplier/STAGE1/pp_19_c2 ;
 wire \u_multiplier/STAGE1/pp_19_c4 ;
 wire \u_multiplier/STAGE1/pp_20_c2 ;
 wire \u_multiplier/STAGE1/pp_21_c2 ;
 wire \u_multiplier/STAGE1/pp_9_c2 ;
 wire net64;
 wire \u_multiplier/STAGE1/E_4_2_pp_10/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_10/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_10/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_10/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_10/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_10/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_10/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_11_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_11_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_11_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_11_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_11_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_11_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_11_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_11_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_11_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_11_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_11_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_11_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_11_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_11_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_12_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_12_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_12_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_12_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_12_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_12_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_12_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_12_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_12_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_12_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_12_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_12_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_12_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_12_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_13_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_13_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_13_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_13_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_13_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_13_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_13_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_13_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_13_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_13_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_13_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_13_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_13_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_13_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_13_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_13_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_13_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_13_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_13_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_13_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_13_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_14_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_14_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_14_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_14_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_14_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_14_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_14_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_14_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_14_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_14_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_14_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_14_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_14_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_14_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_14_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_14_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_14_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_14_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_14_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_14_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_14_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_4/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_4/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_4/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_4/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_4/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_4/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_15_4/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_4/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_4/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_4/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_4/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_4/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_4/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_16_4/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_9/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_9/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_9/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_9/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_9/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_9/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_9/_17_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_17/_08_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_17/_09_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_17/_10_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_17/_11_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_19/_08_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_19/_09_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_19/_10_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_19/_11_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_21/_08_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_21/_09_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_21/_10_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_21/_11_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_23/_08_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_23/_09_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_23/_10_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_23/_11_ ;
 wire \u_multiplier/STAGE2/pp_10_c2 ;
 wire \u_multiplier/STAGE2/pp_10_c4 ;
 wire \u_multiplier/STAGE2/pp_11_c2 ;
 wire \u_multiplier/STAGE2/pp_11_c4 ;
 wire \u_multiplier/STAGE2/pp_12_c2 ;
 wire \u_multiplier/STAGE2/pp_12_c4 ;
 wire \u_multiplier/STAGE2/pp_13_c2 ;
 wire \u_multiplier/STAGE2/pp_13_c4 ;
 wire \u_multiplier/STAGE2/pp_14_c2 ;
 wire \u_multiplier/STAGE2/pp_14_c4 ;
 wire \u_multiplier/STAGE2/pp_15_c2 ;
 wire \u_multiplier/STAGE2/pp_15_c4 ;
 wire \u_multiplier/STAGE2/pp_16_c2 ;
 wire \u_multiplier/STAGE2/pp_16_c4 ;
 wire \u_multiplier/STAGE2/pp_17_c2 ;
 wire \u_multiplier/STAGE2/pp_17_c4 ;
 wire \u_multiplier/STAGE2/pp_18_c2 ;
 wire \u_multiplier/STAGE2/pp_18_c4 ;
 wire \u_multiplier/STAGE2/pp_19_c2 ;
 wire \u_multiplier/STAGE2/pp_19_c4 ;
 wire \u_multiplier/STAGE2/pp_20_c2 ;
 wire \u_multiplier/STAGE2/pp_20_c4 ;
 wire \u_multiplier/STAGE2/pp_21_c2 ;
 wire \u_multiplier/STAGE2/pp_21_c4 ;
 wire \u_multiplier/STAGE2/pp_22_c2 ;
 wire \u_multiplier/STAGE2/pp_22_c4 ;
 wire \u_multiplier/STAGE2/pp_23_c2 ;
 wire \u_multiplier/STAGE2/pp_23_c4 ;
 wire \u_multiplier/STAGE2/pp_24_c2 ;
 wire \u_multiplier/STAGE2/pp_24_c4 ;
 wire \u_multiplier/STAGE2/pp_25_c2 ;
 wire \u_multiplier/STAGE2/pp_5_c2 ;
 wire \u_multiplier/STAGE2/pp_6_c2 ;
 wire \u_multiplier/STAGE2/pp_7_c2 ;
 wire \u_multiplier/STAGE2/pp_7_c4 ;
 wire \u_multiplier/STAGE2/pp_8_c2 ;
 wire \u_multiplier/STAGE2/pp_8_c4 ;
 wire \u_multiplier/STAGE2/pp_9_c2 ;
 wire \u_multiplier/STAGE2/pp_9_c4 ;
 wire net68;
 wire \u_multiplier/STAGE2/E_4_2_pp_10_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_10_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_10_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_10_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_10_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_10_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_10_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_10_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_10_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_10_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_10_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_10_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_10_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_10_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_11_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_11_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_11_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_11_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_11_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_11_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_11_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_11_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_11_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_11_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_11_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_11_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_11_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_11_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_12_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_12_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_12_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_12_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_12_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_12_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_12_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_12_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_12_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_12_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_12_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_12_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_12_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_12_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_13_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_13_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_13_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_13_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_13_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_13_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_13_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_13_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_13_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_13_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_13_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_13_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_13_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_13_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_14_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_14_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_14_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_14_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_14_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_14_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_14_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_14_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_14_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_14_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_14_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_14_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_14_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_14_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_15_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_15_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_15_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_15_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_15_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_15_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_15_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_15_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_15_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_15_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_15_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_15_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_15_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_15_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_16_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_17_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_18_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_19_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_20_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_21_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_22_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_23_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_24_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_25_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_25_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_25_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_25_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_25_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_25_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_25_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_26_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_26_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_26_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_26_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_26_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_26_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_26_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_5/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_5/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_5/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_5/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_5/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_5/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_5/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_6/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_6/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_6/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_6/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_6/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_6/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_6/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_7_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_7_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_7_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_7_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_7_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_7_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_7_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_7_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_7_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_7_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_7_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_7_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_7_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_7_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_8_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_8_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_8_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_8_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_8_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_8_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_8_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_8_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_8_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_8_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_8_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_8_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_8_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_8_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_9_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_9_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_9_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_9_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_9_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_9_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_9_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_9_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_9_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_9_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_9_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_9_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_9_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp_9_2/_17_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp_25/_08_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp_25/_09_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp_25/_10_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp_25/_11_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp_27/_08_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp_27/_09_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp_27/_10_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp_27/_11_ ;
 wire \u_multiplier/STAGE3/pp_10_c1 ;
 wire \u_multiplier/STAGE3/pp_10_c2 ;
 wire \u_multiplier/STAGE3/pp_10_s ;
 wire \u_multiplier/STAGE3/pp_11_c1 ;
 wire \u_multiplier/STAGE3/pp_11_c2 ;
 wire \u_multiplier/STAGE3/pp_11_s ;
 wire \u_multiplier/STAGE3/pp_12_c1 ;
 wire \u_multiplier/STAGE3/pp_12_c2 ;
 wire \u_multiplier/STAGE3/pp_12_s ;
 wire \u_multiplier/STAGE3/pp_13_c1 ;
 wire \u_multiplier/STAGE3/pp_13_c2 ;
 wire \u_multiplier/STAGE3/pp_13_s ;
 wire \u_multiplier/STAGE3/pp_14_c1 ;
 wire \u_multiplier/STAGE3/pp_14_c2 ;
 wire \u_multiplier/STAGE3/pp_14_s ;
 wire \u_multiplier/STAGE3/pp_15_c1 ;
 wire \u_multiplier/STAGE3/pp_15_c2 ;
 wire \u_multiplier/STAGE3/pp_15_s ;
 wire \u_multiplier/STAGE3/pp_16_c1 ;
 wire \u_multiplier/STAGE3/pp_16_c2 ;
 wire \u_multiplier/STAGE3/pp_16_s ;
 wire \u_multiplier/STAGE3/pp_17_c1 ;
 wire \u_multiplier/STAGE3/pp_17_c2 ;
 wire \u_multiplier/STAGE3/pp_17_s ;
 wire \u_multiplier/STAGE3/pp_18_c1 ;
 wire \u_multiplier/STAGE3/pp_18_c2 ;
 wire \u_multiplier/STAGE3/pp_18_s ;
 wire \u_multiplier/STAGE3/pp_19_c1 ;
 wire \u_multiplier/STAGE3/pp_19_c2 ;
 wire \u_multiplier/STAGE3/pp_19_s ;
 wire \u_multiplier/STAGE3/pp_20_c1 ;
 wire \u_multiplier/STAGE3/pp_20_c2 ;
 wire \u_multiplier/STAGE3/pp_20_s ;
 wire \u_multiplier/STAGE3/pp_21_c1 ;
 wire \u_multiplier/STAGE3/pp_21_c2 ;
 wire \u_multiplier/STAGE3/pp_21_s ;
 wire \u_multiplier/STAGE3/pp_22_c1 ;
 wire \u_multiplier/STAGE3/pp_22_c2 ;
 wire \u_multiplier/STAGE3/pp_22_s ;
 wire \u_multiplier/STAGE3/pp_23_c1 ;
 wire \u_multiplier/STAGE3/pp_23_c2 ;
 wire \u_multiplier/STAGE3/pp_23_s ;
 wire \u_multiplier/STAGE3/pp_24_c1 ;
 wire \u_multiplier/STAGE3/pp_24_c2 ;
 wire \u_multiplier/STAGE3/pp_24_s ;
 wire \u_multiplier/STAGE3/pp_25_c1 ;
 wire \u_multiplier/STAGE3/pp_25_c2 ;
 wire \u_multiplier/STAGE3/pp_25_s ;
 wire \u_multiplier/STAGE3/pp_26_c1 ;
 wire \u_multiplier/STAGE3/pp_26_c2 ;
 wire \u_multiplier/STAGE3/pp_26_s ;
 wire \u_multiplier/STAGE3/pp_27_c1 ;
 wire \u_multiplier/STAGE3/pp_27_c2 ;
 wire \u_multiplier/STAGE3/pp_27_s ;
 wire \u_multiplier/STAGE3/pp_28_c1 ;
 wire \u_multiplier/STAGE3/pp_28_c2 ;
 wire \u_multiplier/STAGE3/pp_28_s ;
 wire \u_multiplier/STAGE3/pp_29_c ;
 wire \u_multiplier/STAGE3/pp_29_s ;
 wire \u_multiplier/STAGE3/pp_2_c ;
 wire \u_multiplier/STAGE3/pp_2_s ;
 wire \u_multiplier/STAGE3/pp_3_c1 ;
 wire \u_multiplier/STAGE3/pp_3_c2 ;
 wire \u_multiplier/STAGE3/pp_3_s ;
 wire \u_multiplier/STAGE3/pp_4_c1 ;
 wire \u_multiplier/STAGE3/pp_4_c2 ;
 wire \u_multiplier/STAGE3/pp_4_s ;
 wire \u_multiplier/STAGE3/pp_5_c1 ;
 wire \u_multiplier/STAGE3/pp_5_c2 ;
 wire \u_multiplier/STAGE3/pp_5_s ;
 wire \u_multiplier/STAGE3/pp_6_c1 ;
 wire \u_multiplier/STAGE3/pp_6_c2 ;
 wire \u_multiplier/STAGE3/pp_6_s ;
 wire \u_multiplier/STAGE3/pp_7_c1 ;
 wire \u_multiplier/STAGE3/pp_7_c2 ;
 wire \u_multiplier/STAGE3/pp_7_s ;
 wire \u_multiplier/STAGE3/pp_8_c1 ;
 wire \u_multiplier/STAGE3/pp_8_c2 ;
 wire \u_multiplier/STAGE3/pp_8_s ;
 wire \u_multiplier/STAGE3/pp_9_c1 ;
 wire \u_multiplier/STAGE3/pp_9_c2 ;
 wire \u_multiplier/STAGE3/pp_9_s ;
 wire net81;
 wire \u_multiplier/STAGE3/E_4_2_pp_10_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_10_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_10_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_10_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_10_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_10_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_10_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_11_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_11_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_11_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_11_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_11_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_11_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_11_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_12_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_12_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_12_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_12_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_12_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_12_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_12_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_13_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_13_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_13_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_13_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_13_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_13_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_13_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_14_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_14_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_14_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_14_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_14_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_14_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_14_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_15_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_15_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_15_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_15_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_15_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_15_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_15_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_16_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_16_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_16_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_16_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_16_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_16_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_16_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_17_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_17_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_17_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_17_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_17_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_17_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_17_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_18_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_18_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_18_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_18_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_18_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_18_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_18_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_19_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_19_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_19_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_19_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_19_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_19_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_19_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_20_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_20_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_20_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_20_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_20_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_20_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_20_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_21_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_21_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_21_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_21_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_21_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_21_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_21_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_22_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_22_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_22_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_22_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_22_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_22_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_22_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_23_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_23_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_23_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_23_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_23_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_23_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_23_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_24_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_24_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_24_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_24_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_24_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_24_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_24_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_25_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_25_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_25_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_25_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_25_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_25_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_25_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_26_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_26_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_26_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_26_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_26_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_26_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_26_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_27_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_27_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_27_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_27_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_27_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_27_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_27_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_28_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_28_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_28_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_28_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_28_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_28_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_28_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_3/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_3/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_3/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_3/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_3/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_3/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_3/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_4/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_4/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_4/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_4/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_4/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_4/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_4/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_5/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_5/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_5/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_5/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_5/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_5/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_5/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_6/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_6/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_6/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_6/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_6/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_6/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_6/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_7/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_7/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_7/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_7/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_7/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_7/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_7/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_8/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_8/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_8/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_8/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_8/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_8/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_8/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_9/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_9/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_9/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_9/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_9/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_9/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp_9/_17_ ;
 wire \u_multiplier/STAGE3/Final_add/Cout ;
 wire \u_multiplier/STAGE3/Final_add/c1 ;
 wire \u_multiplier/STAGE3/Final_add/cla1/c1 ;
 wire \u_multiplier/STAGE3/Final_add/cla1/c2 ;
 wire \u_multiplier/STAGE3/Final_add/cla1/c3 ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_25_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_26_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_27_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_28_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_29_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_30_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_31_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_32_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_33_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_34_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_35_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_36_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_37_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_38_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla1/_39_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_25_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_26_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_27_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_28_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_29_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_30_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_31_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_32_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_33_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_34_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_35_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_36_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_37_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_38_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla2/_39_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_25_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_26_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_27_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_28_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_29_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_30_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_31_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_32_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_33_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_34_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_35_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_36_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_37_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_38_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla3/_39_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_25_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_26_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_27_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_28_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_29_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_30_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_31_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_32_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_33_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_34_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_35_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_36_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_37_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_38_ ;
 wire \u_multiplier/STAGE3/Final_add/cla1/cla4/_39_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/c1 ;
 wire \u_multiplier/STAGE3/Final_add/cla2/c2 ;
 wire \u_multiplier/STAGE3/Final_add/cla2/c3 ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_25_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_26_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_27_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_28_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_29_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_30_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_31_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_32_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_33_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_34_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_35_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_36_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_37_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_38_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla1/_39_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_25_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_26_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_27_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_28_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_29_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_30_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_31_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_32_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_33_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_34_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_35_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_36_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_37_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_38_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla2/_39_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_25_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_26_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_27_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_28_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_29_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_30_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_31_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_32_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_33_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_34_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_35_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_36_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_37_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_38_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla3/_39_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_25_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_26_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_27_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_28_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_29_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_30_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_31_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_32_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_33_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_34_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_35_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_36_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_37_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_38_ ;
 wire \u_multiplier/STAGE3/Final_add/cla2/cla4/_39_ ;
 wire \u_multiplier/STAGE3/Full_adder_pp_29/_08_ ;
 wire \u_multiplier/STAGE3/Full_adder_pp_29/_09_ ;
 wire \u_multiplier/STAGE3/Full_adder_pp_29/_10_ ;
 wire \u_multiplier/STAGE3/Full_adder_pp_29/_11_ ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire valid_reg_out;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net65;
 wire net66;
 wire net67;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire clknet_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire [4:0] addr_ptr;
 wire [2:0] curr_state;
 wire [15:0] data_in_reg;
 wire [4:0] init_count;
 wire [31:0] product;
 wire [15:0] sram_rdata;
 wire [15:0] sram_rdata_reg;
 wire [1:0] \u_multiplier/pp_1 ;
 wire [7:0] \u_multiplier/pp_10 ;
 wire [7:0] \u_multiplier/pp_11 ;
 wire [7:0] \u_multiplier/pp_12 ;
 wire [7:0] \u_multiplier/pp_13 ;
 wire [7:0] \u_multiplier/pp_14 ;
 wire [7:0] \u_multiplier/pp_15 ;
 wire [7:0] \u_multiplier/pp_16 ;
 wire [7:0] \u_multiplier/pp_17 ;
 wire [7:0] \u_multiplier/pp_18 ;
 wire [7:0] \u_multiplier/pp_19 ;
 wire [2:0] \u_multiplier/pp_2 ;
 wire [7:0] \u_multiplier/pp_20 ;
 wire [7:0] \u_multiplier/pp_21 ;
 wire [7:0] \u_multiplier/pp_22 ;
 wire [7:0] \u_multiplier/pp_23 ;
 wire [7:0] \u_multiplier/pp_24 ;
 wire [5:0] \u_multiplier/pp_25 ;
 wire [4:0] \u_multiplier/pp_26 ;
 wire [3:0] \u_multiplier/pp_27 ;
 wire [2:0] \u_multiplier/pp_28 ;
 wire [1:0] \u_multiplier/pp_29 ;
 wire [3:0] \u_multiplier/pp_3 ;
 wire [4:0] \u_multiplier/pp_4 ;
 wire [5:0] \u_multiplier/pp_5 ;
 wire [6:0] \u_multiplier/pp_6 ;
 wire [7:0] \u_multiplier/pp_7 ;
 wire [7:0] \u_multiplier/pp_8 ;
 wire [7:0] \u_multiplier/pp_9 ;
 wire [1:0] \u_multiplier/s_1 ;
 wire [3:0] \u_multiplier/s_10 ;
 wire [3:0] \u_multiplier/s_11 ;
 wire [3:0] \u_multiplier/s_12 ;
 wire [3:0] \u_multiplier/s_13 ;
 wire [3:0] \u_multiplier/s_14 ;
 wire [3:0] \u_multiplier/s_15 ;
 wire [3:0] \u_multiplier/s_16 ;
 wire [3:0] \u_multiplier/s_17 ;
 wire [3:0] \u_multiplier/s_18 ;
 wire [3:0] \u_multiplier/s_19 ;
 wire [2:0] \u_multiplier/s_2 ;
 wire [3:0] \u_multiplier/s_20 ;
 wire [3:0] \u_multiplier/s_21 ;
 wire [3:0] \u_multiplier/s_22 ;
 wire [3:0] \u_multiplier/s_23 ;
 wire [3:0] \u_multiplier/s_24 ;
 wire [3:0] \u_multiplier/s_25 ;
 wire [3:0] \u_multiplier/s_26 ;
 wire [3:0] \u_multiplier/s_27 ;
 wire [3:0] \u_multiplier/s_28 ;
 wire [1:0] \u_multiplier/s_29 ;
 wire [3:0] \u_multiplier/s_3 ;
 wire [3:0] \u_multiplier/s_4 ;
 wire [3:0] \u_multiplier/s_5 ;
 wire [3:0] \u_multiplier/s_6 ;
 wire [3:0] \u_multiplier/s_7 ;
 wire [3:0] \u_multiplier/s_8 ;
 wire [3:0] \u_multiplier/s_9 ;

 INV_X1 _420_ (.A(net19),
    .ZN(_238_));
 INV_X2 _421_ (.A(net18),
    .ZN(_195_));
 INV_X1 _422_ (.A(curr_state[2]),
    .ZN(_239_));
 INV_X1 _423_ (.A(_408_),
    .ZN(_240_));
 INV_X1 _424_ (.A(addr_ptr[0]),
    .ZN(_241_));
 INV_X1 _425_ (.A(_401_),
    .ZN(_242_));
 AND2_X4 _426_ (.A1(net19),
    .A2(net20),
    .ZN(_191_));
 INV_X1 _427_ (.A(_191_),
    .ZN(_243_));
 NAND2_X1 _428_ (.A1(net19),
    .A2(net151),
    .ZN(_196_));
 NAND2_X1 _429_ (.A1(init_count[1]),
    .A2(init_count[0]),
    .ZN(_244_));
 AND3_X1 _430_ (.A1(init_count[1]),
    .A2(init_count[0]),
    .A3(init_count[2]),
    .ZN(_245_));
 AND4_X2 _431_ (.A1(init_count[1]),
    .A2(init_count[0]),
    .A3(init_count[3]),
    .A4(init_count[2]),
    .ZN(_246_));
 AND3_X1 _432_ (.A1(net18),
    .A2(init_count[4]),
    .A3(_246_),
    .ZN(_247_));
 NOR2_X1 _433_ (.A1(_191_),
    .A2(_247_),
    .ZN(_248_));
 AOI21_X1 _434_ (.A(_248_),
    .B1(_196_),
    .B2(_243_),
    .ZN(_193_));
 NOR2_X2 _435_ (.A1(_238_),
    .A2(_195_),
    .ZN(_249_));
 NAND2_X2 _436_ (.A1(net19),
    .A2(net18),
    .ZN(_250_));
 NAND3_X1 _437_ (.A1(net17),
    .A2(net114),
    .A3(_249_),
    .ZN(_251_));
 OAI21_X1 _438_ (.A(net115),
    .B1(_247_),
    .B2(_196_),
    .ZN(_194_));
 AOI22_X1 _439_ (.A1(net19),
    .A2(net83),
    .B1(_249_),
    .B2(net17),
    .ZN(_192_));
 AND2_X1 _440_ (.A1(net19),
    .A2(sram_rdata[0]),
    .ZN(_175_));
 AND2_X1 _441_ (.A1(net19),
    .A2(sram_rdata[1]),
    .ZN(_182_));
 AND2_X1 _442_ (.A1(net19),
    .A2(sram_rdata[2]),
    .ZN(_183_));
 AND2_X1 _443_ (.A1(net19),
    .A2(sram_rdata[3]),
    .ZN(_184_));
 AND2_X1 _444_ (.A1(net19),
    .A2(sram_rdata[4]),
    .ZN(_185_));
 AND2_X1 _445_ (.A1(net19),
    .A2(sram_rdata[5]),
    .ZN(_186_));
 AND2_X1 _446_ (.A1(net19),
    .A2(sram_rdata[6]),
    .ZN(_187_));
 AND2_X1 _447_ (.A1(net19),
    .A2(sram_rdata[7]),
    .ZN(_188_));
 AND2_X1 _448_ (.A1(net19),
    .A2(sram_rdata[8]),
    .ZN(_189_));
 AND2_X1 _449_ (.A1(net19),
    .A2(sram_rdata[9]),
    .ZN(_190_));
 AND2_X1 _450_ (.A1(net19),
    .A2(sram_rdata[10]),
    .ZN(_176_));
 AND2_X1 _451_ (.A1(net19),
    .A2(sram_rdata[11]),
    .ZN(_177_));
 AND2_X1 _452_ (.A1(net19),
    .A2(sram_rdata[12]),
    .ZN(_178_));
 AND2_X1 _453_ (.A1(net19),
    .A2(sram_rdata[13]),
    .ZN(_179_));
 AND2_X1 _454_ (.A1(net19),
    .A2(sram_rdata[14]),
    .ZN(_180_));
 AND2_X1 _455_ (.A1(net19),
    .A2(sram_rdata[15]),
    .ZN(_181_));
 AND2_X1 _456_ (.A1(product[0]),
    .A2(_191_),
    .ZN(_138_));
 AND2_X1 _457_ (.A1(product[1]),
    .A2(_191_),
    .ZN(_149_));
 AND2_X1 _458_ (.A1(product[2]),
    .A2(_191_),
    .ZN(_160_));
 AND2_X1 _459_ (.A1(product[3]),
    .A2(_191_),
    .ZN(_163_));
 AND2_X1 _460_ (.A1(product[4]),
    .A2(_191_),
    .ZN(_164_));
 AND2_X1 _461_ (.A1(product[5]),
    .A2(_191_),
    .ZN(_165_));
 AND2_X1 _462_ (.A1(product[6]),
    .A2(_191_),
    .ZN(_166_));
 AND2_X1 _463_ (.A1(product[7]),
    .A2(_191_),
    .ZN(_167_));
 AND2_X1 _464_ (.A1(product[8]),
    .A2(_191_),
    .ZN(_168_));
 AND2_X1 _465_ (.A1(product[9]),
    .A2(_191_),
    .ZN(_169_));
 AND2_X1 _466_ (.A1(product[10]),
    .A2(_191_),
    .ZN(_139_));
 AND2_X1 _467_ (.A1(product[11]),
    .A2(_191_),
    .ZN(_140_));
 AND2_X1 _468_ (.A1(product[12]),
    .A2(_191_),
    .ZN(_141_));
 AND2_X1 _469_ (.A1(product[13]),
    .A2(_191_),
    .ZN(_142_));
 AND2_X1 _470_ (.A1(product[14]),
    .A2(_191_),
    .ZN(_143_));
 AND2_X1 _471_ (.A1(product[15]),
    .A2(_191_),
    .ZN(_144_));
 AND2_X1 _472_ (.A1(product[16]),
    .A2(_191_),
    .ZN(_145_));
 AND2_X1 _473_ (.A1(product[17]),
    .A2(_191_),
    .ZN(_146_));
 AND2_X1 _474_ (.A1(product[18]),
    .A2(_191_),
    .ZN(_147_));
 AND2_X1 _475_ (.A1(product[19]),
    .A2(_191_),
    .ZN(_148_));
 AND2_X1 _476_ (.A1(product[20]),
    .A2(_191_),
    .ZN(_150_));
 AND2_X1 _477_ (.A1(product[21]),
    .A2(_191_),
    .ZN(_151_));
 AND2_X1 _478_ (.A1(product[22]),
    .A2(_191_),
    .ZN(_152_));
 AND2_X1 _479_ (.A1(product[23]),
    .A2(_191_),
    .ZN(_153_));
 AND2_X1 _480_ (.A1(product[24]),
    .A2(_191_),
    .ZN(_154_));
 AND2_X1 _481_ (.A1(product[25]),
    .A2(_191_),
    .ZN(_155_));
 AND2_X1 _482_ (.A1(product[26]),
    .A2(_191_),
    .ZN(_156_));
 AND2_X1 _483_ (.A1(product[27]),
    .A2(_191_),
    .ZN(_157_));
 AND2_X1 _484_ (.A1(product[28]),
    .A2(_191_),
    .ZN(_158_));
 AND2_X1 _485_ (.A1(product[29]),
    .A2(_191_),
    .ZN(_159_));
 AND2_X1 _486_ (.A1(product[30]),
    .A2(_191_),
    .ZN(_161_));
 AND2_X1 _487_ (.A1(product[31]),
    .A2(_191_),
    .ZN(_162_));
 AND2_X1 _488_ (.A1(net19),
    .A2(net1),
    .ZN(_122_));
 AND2_X1 _489_ (.A1(net19),
    .A2(net8),
    .ZN(_129_));
 AND2_X1 _490_ (.A1(net19),
    .A2(net9),
    .ZN(_130_));
 AND2_X1 _491_ (.A1(net19),
    .A2(net10),
    .ZN(_131_));
 AND2_X1 _492_ (.A1(net19),
    .A2(net11),
    .ZN(_132_));
 AND2_X1 _493_ (.A1(net19),
    .A2(net12),
    .ZN(_133_));
 AND2_X1 _494_ (.A1(net19),
    .A2(net13),
    .ZN(_134_));
 AND2_X1 _495_ (.A1(net19),
    .A2(net14),
    .ZN(_135_));
 AND2_X1 _496_ (.A1(net19),
    .A2(net15),
    .ZN(_136_));
 AND2_X1 _497_ (.A1(net19),
    .A2(net16),
    .ZN(_137_));
 AND2_X1 _498_ (.A1(net19),
    .A2(net2),
    .ZN(_123_));
 AND2_X1 _499_ (.A1(net19),
    .A2(net3),
    .ZN(_124_));
 AND2_X1 _500_ (.A1(net19),
    .A2(net4),
    .ZN(_125_));
 AND2_X1 _501_ (.A1(net19),
    .A2(net5),
    .ZN(_126_));
 AND2_X1 _502_ (.A1(net19),
    .A2(net6),
    .ZN(_127_));
 AND2_X1 _503_ (.A1(net19),
    .A2(net7),
    .ZN(_128_));
 NAND2_X2 _504_ (.A1(net19),
    .A2(_195_),
    .ZN(_252_));
 NAND2_X2 _505_ (.A1(_240_),
    .A2(_246_),
    .ZN(_253_));
 XNOR2_X1 _506_ (.A(net117),
    .B(_253_),
    .ZN(_254_));
 AOI22_X1 _507_ (.A1(init_count[0]),
    .A2(net20),
    .B1(_254_),
    .B2(curr_state[2]),
    .ZN(_255_));
 OAI22_X1 _508_ (.A1(net118),
    .A2(_252_),
    .B1(_255_),
    .B2(_250_),
    .ZN(_170_));
 XNOR2_X1 _509_ (.A(init_count[1]),
    .B(init_count[0]),
    .ZN(_256_));
 AOI21_X1 _510_ (.A(_239_),
    .B1(_253_),
    .B2(_256_),
    .ZN(_257_));
 AOI21_X1 _511_ (.A(_257_),
    .B1(net20),
    .B2(init_count[1]),
    .ZN(_258_));
 OAI22_X1 _512_ (.A1(net112),
    .A2(_252_),
    .B1(_258_),
    .B2(_250_),
    .ZN(_171_));
 XNOR2_X1 _513_ (.A(_406_),
    .B(_244_),
    .ZN(_259_));
 AOI21_X1 _514_ (.A(_239_),
    .B1(_253_),
    .B2(_259_),
    .ZN(_260_));
 AOI21_X1 _515_ (.A(_260_),
    .B1(net20),
    .B2(init_count[2]),
    .ZN(_261_));
 OAI22_X1 _516_ (.A1(net109),
    .A2(_252_),
    .B1(_261_),
    .B2(_250_),
    .ZN(_172_));
 OAI21_X1 _517_ (.A(curr_state[2]),
    .B1(_245_),
    .B2(init_count[3]),
    .ZN(_262_));
 AOI21_X1 _518_ (.A(_262_),
    .B1(_246_),
    .B2(_408_),
    .ZN(_263_));
 AOI21_X1 _519_ (.A(_263_),
    .B1(net20),
    .B2(init_count[3]),
    .ZN(_264_));
 OAI22_X1 _520_ (.A1(net81),
    .A2(_252_),
    .B1(_264_),
    .B2(_250_),
    .ZN(_173_));
 AND2_X1 _521_ (.A1(init_count[4]),
    .A2(net20),
    .ZN(_265_));
 OAI221_X1 _522_ (.A(_249_),
    .B1(_265_),
    .B2(curr_state[2]),
    .C1(_246_),
    .C2(init_count[4]),
    .ZN(_266_));
 OAI21_X1 _523_ (.A(_266_),
    .B1(_252_),
    .B2(net131),
    .ZN(_174_));
 AND2_X1 _524_ (.A1(curr_state[2]),
    .A2(net97),
    .ZN(_267_));
 AOI22_X1 _525_ (.A1(net20),
    .A2(_241_),
    .B1(_253_),
    .B2(_267_),
    .ZN(_268_));
 OAI22_X1 _526_ (.A1(net98),
    .A2(_252_),
    .B1(_268_),
    .B2(_250_),
    .ZN(_117_));
 AOI21_X2 _527_ (.A(_239_),
    .B1(_246_),
    .B2(init_count[4]),
    .ZN(_269_));
 AND2_X1 _528_ (.A1(addr_ptr[0]),
    .A2(addr_ptr[1]),
    .ZN(_270_));
 NOR2_X1 _529_ (.A1(_250_),
    .A2(_270_),
    .ZN(_271_));
 OAI221_X1 _530_ (.A(_271_),
    .B1(addr_ptr[1]),
    .B2(addr_ptr[0]),
    .C1(net20),
    .C2(_269_),
    .ZN(_272_));
 OAI21_X1 _531_ (.A(_272_),
    .B1(_252_),
    .B2(net101),
    .ZN(_118_));
 NAND4_X1 _532_ (.A1(addr_ptr[3]),
    .A2(addr_ptr[2]),
    .A3(addr_ptr[4]),
    .A4(_270_),
    .ZN(_273_));
 AOI21_X2 _533_ (.A(_269_),
    .B1(_273_),
    .B2(net20),
    .ZN(_274_));
 XNOR2_X1 _534_ (.A(net120),
    .B(_270_),
    .ZN(_275_));
 NAND2_X1 _535_ (.A1(_249_),
    .A2(_275_),
    .ZN(_276_));
 OAI22_X1 _536_ (.A1(net121),
    .A2(_252_),
    .B1(_274_),
    .B2(_276_),
    .ZN(_119_));
 NAND3_X1 _537_ (.A1(net18),
    .A2(_242_),
    .A3(_270_),
    .ZN(_277_));
 XNOR2_X1 _538_ (.A(net103),
    .B(_277_),
    .ZN(_278_));
 AOI211_X1 _539_ (.A(_238_),
    .B(net104),
    .C1(_274_),
    .C2(net18),
    .ZN(_120_));
 NAND4_X1 _540_ (.A1(net18),
    .A2(addr_ptr[3]),
    .A3(addr_ptr[2]),
    .A4(_270_),
    .ZN(_279_));
 XNOR2_X1 _541_ (.A(net105),
    .B(_279_),
    .ZN(_280_));
 AOI211_X1 _542_ (.A(_238_),
    .B(net106),
    .C1(_274_),
    .C2(net18),
    .ZN(_121_));
 DFF_X1 _543_ (.D(net84),
    .CK(clknet_3_3_0_clk),
    .Q(curr_state[0]),
    .QN(_331_));
 DFF_X2 _544_ (.D(_193_),
    .CK(clknet_3_3_0_clk),
    .Q(net20),
    .QN(_332_));
 DFF_X2 _545_ (.D(net116),
    .CK(clknet_3_3_0_clk),
    .Q(curr_state[2]),
    .QN(_333_));
 DFF_X1 _546_ (.D(_138_),
    .CK(clknet_3_7_0_clk),
    .Q(net21),
    .QN(_334_));
 DFF_X1 _547_ (.D(_149_),
    .CK(clknet_3_6_0_clk),
    .Q(net32),
    .QN(_335_));
 DFF_X1 _548_ (.D(_160_),
    .CK(clknet_3_7_0_clk),
    .Q(net43),
    .QN(_336_));
 DFF_X2 _549_ (.D(_163_),
    .CK(clknet_3_6_0_clk),
    .Q(net46),
    .QN(_337_));
 DFF_X2 _550_ (.D(_164_),
    .CK(clknet_3_4_0_clk),
    .Q(net47),
    .QN(_338_));
 DFF_X2 _551_ (.D(_165_),
    .CK(clknet_3_6_0_clk),
    .Q(net48),
    .QN(_339_));
 DFF_X1 _552_ (.D(_166_),
    .CK(clknet_3_3_0_clk),
    .Q(net49),
    .QN(_340_));
 DFF_X1 _553_ (.D(_167_),
    .CK(clknet_3_6_0_clk),
    .Q(net50),
    .QN(_341_));
 DFF_X2 _554_ (.D(_168_),
    .CK(clknet_3_7_0_clk),
    .Q(net51),
    .QN(_342_));
 DFF_X2 _555_ (.D(_169_),
    .CK(clknet_3_7_0_clk),
    .Q(net52),
    .QN(_343_));
 DFF_X2 _556_ (.D(_139_),
    .CK(clknet_3_6_0_clk),
    .Q(net22),
    .QN(_344_));
 DFF_X2 _557_ (.D(_140_),
    .CK(clknet_3_7_0_clk),
    .Q(net23),
    .QN(_345_));
 DFF_X1 _558_ (.D(_141_),
    .CK(clknet_3_2_0_clk),
    .Q(net24),
    .QN(_346_));
 DFF_X2 _559_ (.D(_142_),
    .CK(clknet_3_6_0_clk),
    .Q(net25),
    .QN(_347_));
 DFF_X2 _560_ (.D(_143_),
    .CK(clknet_3_7_0_clk),
    .Q(net26),
    .QN(_348_));
 DFF_X2 _561_ (.D(_144_),
    .CK(clknet_3_7_0_clk),
    .Q(net27),
    .QN(_349_));
 DFF_X2 _562_ (.D(_145_),
    .CK(clknet_3_2_0_clk),
    .Q(net28),
    .QN(_350_));
 DFF_X2 _563_ (.D(_146_),
    .CK(clknet_3_5_0_clk),
    .Q(net29),
    .QN(_351_));
 DFF_X1 _564_ (.D(_147_),
    .CK(clknet_3_3_0_clk),
    .Q(net30),
    .QN(_352_));
 DFF_X2 _565_ (.D(_148_),
    .CK(clknet_3_5_0_clk),
    .Q(net31),
    .QN(_353_));
 DFF_X2 _566_ (.D(_150_),
    .CK(clknet_3_0_0_clk),
    .Q(net33),
    .QN(_354_));
 DFF_X2 _567_ (.D(_151_),
    .CK(clknet_3_4_0_clk),
    .Q(net34),
    .QN(_355_));
 DFF_X2 _568_ (.D(_152_),
    .CK(clknet_3_4_0_clk),
    .Q(net35),
    .QN(_356_));
 DFF_X2 _569_ (.D(_153_),
    .CK(clknet_3_4_0_clk),
    .Q(net36),
    .QN(_357_));
 DFF_X2 _570_ (.D(_154_),
    .CK(clknet_3_3_0_clk),
    .Q(net37),
    .QN(_358_));
 DFF_X2 _571_ (.D(_155_),
    .CK(clknet_3_5_0_clk),
    .Q(net38),
    .QN(_359_));
 DFF_X2 _572_ (.D(_156_),
    .CK(clknet_3_4_0_clk),
    .Q(net39),
    .QN(_360_));
 DFF_X2 _573_ (.D(_157_),
    .CK(clknet_3_4_0_clk),
    .Q(net40),
    .QN(_361_));
 DFF_X1 _574_ (.D(_158_),
    .CK(clknet_3_5_0_clk),
    .Q(net41),
    .QN(_362_));
 DFF_X2 _575_ (.D(_159_),
    .CK(clknet_3_5_0_clk),
    .Q(net42),
    .QN(_363_));
 DFF_X2 _576_ (.D(_161_),
    .CK(clknet_3_5_0_clk),
    .Q(net44),
    .QN(_364_));
 DFF_X2 _577_ (.D(_162_),
    .CK(clknet_3_5_0_clk),
    .Q(net45),
    .QN(_365_));
 DFF_X2 _578_ (.D(_122_),
    .CK(clknet_3_7_0_clk),
    .Q(data_in_reg[0]),
    .QN(_366_));
 DFF_X2 _579_ (.D(_129_),
    .CK(clknet_3_2_0_clk),
    .Q(data_in_reg[1]),
    .QN(_367_));
 DFF_X2 _580_ (.D(_130_),
    .CK(clknet_3_5_0_clk),
    .Q(data_in_reg[2]),
    .QN(_368_));
 DFF_X2 _581_ (.D(_131_),
    .CK(clknet_3_7_0_clk),
    .Q(data_in_reg[3]),
    .QN(_369_));
 DFF_X2 _582_ (.D(_132_),
    .CK(clknet_3_3_0_clk),
    .Q(data_in_reg[4]),
    .QN(_370_));
 DFF_X2 _583_ (.D(_133_),
    .CK(clknet_3_1_0_clk),
    .Q(data_in_reg[5]),
    .QN(_371_));
 DFF_X2 _584_ (.D(_134_),
    .CK(clknet_3_5_0_clk),
    .Q(data_in_reg[6]),
    .QN(_372_));
 DFF_X2 _585_ (.D(_135_),
    .CK(clknet_3_7_0_clk),
    .Q(data_in_reg[7]),
    .QN(_373_));
 DFF_X2 _586_ (.D(_136_),
    .CK(clknet_3_2_0_clk),
    .Q(data_in_reg[8]),
    .QN(_374_));
 DFF_X2 _587_ (.D(_137_),
    .CK(clknet_3_2_0_clk),
    .Q(data_in_reg[9]),
    .QN(_375_));
 DFF_X2 _588_ (.D(_123_),
    .CK(clknet_3_4_0_clk),
    .Q(data_in_reg[10]),
    .QN(_376_));
 DFF_X2 _589_ (.D(_124_),
    .CK(clknet_3_7_0_clk),
    .Q(data_in_reg[11]),
    .QN(_377_));
 DFF_X2 _590_ (.D(_125_),
    .CK(clknet_3_6_0_clk),
    .Q(data_in_reg[12]),
    .QN(_378_));
 DFF_X2 _591_ (.D(_126_),
    .CK(clknet_3_5_0_clk),
    .Q(data_in_reg[13]),
    .QN(_379_));
 DFF_X2 _592_ (.D(_127_),
    .CK(clknet_3_0_0_clk),
    .Q(data_in_reg[14]),
    .QN(_380_));
 DFF_X2 _593_ (.D(_128_),
    .CK(clknet_3_4_0_clk),
    .Q(data_in_reg[15]),
    .QN(_381_));
 DFF_X2 _594_ (.D(_175_),
    .CK(clknet_3_0_0_clk),
    .Q(sram_rdata_reg[0]),
    .QN(_382_));
 DFF_X2 _595_ (.D(_182_),
    .CK(clknet_3_0_0_clk),
    .Q(sram_rdata_reg[1]),
    .QN(_383_));
 DFF_X2 _596_ (.D(_183_),
    .CK(clknet_3_0_0_clk),
    .Q(sram_rdata_reg[2]),
    .QN(_384_));
 DFF_X2 _597_ (.D(_184_),
    .CK(clknet_3_0_0_clk),
    .Q(sram_rdata_reg[3]),
    .QN(_385_));
 DFF_X2 _598_ (.D(_185_),
    .CK(clknet_3_0_0_clk),
    .Q(sram_rdata_reg[4]),
    .QN(_386_));
 DFF_X2 _599_ (.D(_186_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[5]),
    .QN(_387_));
 DFF_X2 _600_ (.D(_187_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[6]),
    .QN(_388_));
 DFF_X2 _601_ (.D(_188_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[7]),
    .QN(_389_));
 DFF_X2 _602_ (.D(_189_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[8]),
    .QN(_390_));
 DFF_X2 _603_ (.D(_190_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[9]),
    .QN(_391_));
 DFF_X2 _604_ (.D(_176_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[10]),
    .QN(_392_));
 DFF_X2 _605_ (.D(_177_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[11]),
    .QN(_393_));
 DFF_X2 _606_ (.D(_178_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[12]),
    .QN(_394_));
 DFF_X2 _607_ (.D(_179_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[13]),
    .QN(_395_));
 DFF_X2 _608_ (.D(_180_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[14]),
    .QN(_396_));
 DFF_X2 _609_ (.D(_181_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[15]),
    .QN(_397_));
 DFF_X1 _610_ (.D(_191_),
    .CK(clknet_3_6_0_clk),
    .Q(net53),
    .QN(_398_));
 DFF_X1 _611_ (.D(net99),
    .CK(clknet_3_3_0_clk),
    .Q(addr_ptr[0]),
    .QN(_399_));
 DFF_X1 _612_ (.D(net102),
    .CK(clknet_3_2_0_clk),
    .Q(addr_ptr[1]),
    .QN(_400_));
 DFF_X1 _613_ (.D(_119_),
    .CK(clknet_3_2_0_clk),
    .Q(addr_ptr[2]),
    .QN(_401_));
 DFF_X1 _614_ (.D(_120_),
    .CK(clknet_3_2_0_clk),
    .Q(addr_ptr[3]),
    .QN(_402_));
 DFF_X1 _615_ (.D(_121_),
    .CK(clknet_3_2_0_clk),
    .Q(addr_ptr[4]),
    .QN(_403_));
 DFF_X2 _616_ (.D(net119),
    .CK(clknet_3_3_0_clk),
    .Q(init_count[0]),
    .QN(_404_));
 DFF_X2 _617_ (.D(net113),
    .CK(clknet_3_3_0_clk),
    .Q(init_count[1]),
    .QN(_405_));
 DFF_X1 _618_ (.D(net110),
    .CK(clknet_3_3_0_clk),
    .Q(init_count[2]),
    .QN(_406_));
 DFF_X1 _619_ (.D(net82),
    .CK(clknet_3_3_0_clk),
    .Q(init_count[3]),
    .QN(_407_));
 DFF_X1 _620_ (.D(net132),
    .CK(clknet_3_3_0_clk),
    .Q(init_count[4]),
    .QN(_408_));
 SRAM_6T_CORE_32x16_MC_TB sram_inst (.ce_in(_195_),
    .we_in(_196_),
    .clk(clknet_3_0_0_clk),
    .addr_in({net129,
    net136,
    net134,
    net124,
    net95}),
    .rd_out({sram_rdata[15],
    sram_rdata[14],
    sram_rdata[13],
    sram_rdata[12],
    sram_rdata[11],
    sram_rdata[10],
    sram_rdata[9],
    sram_rdata[8],
    sram_rdata[7],
    sram_rdata[6],
    sram_rdata[5],
    sram_rdata[4],
    sram_rdata[3],
    sram_rdata[2],
    sram_rdata[1],
    sram_rdata[0]}),
    .wd_in({net126,
    net127,
    net138,
    net137,
    net139,
    net122,
    net150,
    net149,
    net141,
    net140,
    net107,
    net147,
    net145,
    net144,
    net125,
    net148}));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_10/_18_  (.A(\u_multiplier/STAGE1/pp_9_c2 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_10/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_10/_19_  (.A1(\u_multiplier/STAGE1/_185_ ),
    .A2(\u_multiplier/STAGE1/_184_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_10/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_10/_20_  (.A(\u_multiplier/STAGE1/_185_ ),
    .B(\u_multiplier/STAGE1/_184_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_10/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_10/_21_  (.A1(\u_multiplier/STAGE1/_186_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_10/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_10/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_10/_22_  (.A(\u_multiplier/STAGE1/_186_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_10/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_10/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_10/_23_  (.A1(\u_multiplier/STAGE1/_187_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_10/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_10/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_10/_24_  (.A(\u_multiplier/STAGE1/_187_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_10/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_10/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_10/_25_  (.A(\u_multiplier/STAGE1/pp_9_c2 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_10/_16_ ),
    .ZN(\u_multiplier/pp_10 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_10/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_10/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_10/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_10_c2 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_10/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_10/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_10/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_10/_17_ ),
    .ZN(\u_multiplier/pp_11 [2]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_11_1/_18_  (.A(\u_multiplier/STAGE1/pp_10_c2 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_11_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_11_1/_19_  (.A1(\u_multiplier/STAGE1/_191_ ),
    .A2(\u_multiplier/STAGE1/_190_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_11_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_11_1/_20_  (.A(\u_multiplier/STAGE1/_191_ ),
    .B(\u_multiplier/STAGE1/_190_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_11_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_11_1/_21_  (.A1(\u_multiplier/STAGE1/_192_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_11_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_11_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_11_1/_22_  (.A(\u_multiplier/STAGE1/_192_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_11_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_11_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_11_1/_23_  (.A1(\u_multiplier/STAGE1/_193_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_11_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_11_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_11_1/_24_  (.A(\u_multiplier/STAGE1/_193_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_11_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_11_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_11_1/_25_  (.A(\u_multiplier/STAGE1/pp_10_c2 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_11_1/_16_ ),
    .ZN(\u_multiplier/pp_11 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_11_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_11_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_11_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_11_c2 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_11_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_11_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_11_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_11_1/_17_ ),
    .ZN(\u_multiplier/pp_12 [4]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_11_2/_18_  (.A(net54),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_11_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_11_2/_19_  (.A1(\u_multiplier/STAGE1/_195_ ),
    .A2(\u_multiplier/STAGE1/_194_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_11_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_11_2/_20_  (.A(\u_multiplier/STAGE1/_195_ ),
    .B(\u_multiplier/STAGE1/_194_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_11_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_11_2/_21_  (.A1(\u_multiplier/STAGE1/_196_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_11_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_11_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_11_2/_22_  (.A(\u_multiplier/STAGE1/_196_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_11_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_11_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_11_2/_23_  (.A1(\u_multiplier/STAGE1/_197_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_11_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_11_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_11_2/_24_  (.A(\u_multiplier/STAGE1/_197_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_11_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_11_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_11_2/_25_  (.A(net55),
    .B(\u_multiplier/STAGE1/E_4_2_pp_11_2/_16_ ),
    .ZN(\u_multiplier/pp_11 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_11_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_11_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_11_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_11_c4 ));
 OAI21_X1 \u_multiplier/STAGE1/E_4_2_pp_11_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_11_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_11_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_11_2/_17_ ),
    .ZN(\u_multiplier/pp_12 [3]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_12_1/_18_  (.A(\u_multiplier/STAGE1/pp_11_c2 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_12_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_12_1/_19_  (.A1(\u_multiplier/STAGE1/_199_ ),
    .A2(\u_multiplier/STAGE1/_198_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_12_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_12_1/_20_  (.A(\u_multiplier/STAGE1/_199_ ),
    .B(\u_multiplier/STAGE1/_198_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_12_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_12_1/_21_  (.A1(\u_multiplier/STAGE1/_200_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_12_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_12_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_12_1/_22_  (.A(\u_multiplier/STAGE1/_200_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_12_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_12_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_12_1/_23_  (.A1(\u_multiplier/STAGE1/_201_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_12_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_12_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_12_1/_24_  (.A(\u_multiplier/STAGE1/_201_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_12_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_12_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_12_1/_25_  (.A(\u_multiplier/STAGE1/pp_11_c2 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_12_1/_16_ ),
    .ZN(\u_multiplier/pp_12 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_12_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_12_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_12_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_12_c2 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_12_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_12_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_12_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_12_1/_17_ ),
    .ZN(\u_multiplier/pp_13 [5]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_12_2/_18_  (.A(\u_multiplier/STAGE1/pp_11_c4 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_12_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_12_2/_19_  (.A1(\u_multiplier/STAGE1/_203_ ),
    .A2(\u_multiplier/STAGE1/_202_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_12_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_12_2/_20_  (.A(\u_multiplier/STAGE1/_203_ ),
    .B(\u_multiplier/STAGE1/_202_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_12_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_12_2/_21_  (.A1(\u_multiplier/STAGE1/_204_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_12_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_12_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_12_2/_22_  (.A(\u_multiplier/STAGE1/_204_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_12_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_12_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_12_2/_23_  (.A1(\u_multiplier/STAGE1/_205_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_12_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_12_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_12_2/_24_  (.A(\u_multiplier/STAGE1/_205_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_12_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_12_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_12_2/_25_  (.A(\u_multiplier/STAGE1/pp_11_c4 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_12_2/_16_ ),
    .ZN(\u_multiplier/pp_12 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_12_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_12_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_12_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_12_c4 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_12_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_12_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_12_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_12_2/_17_ ),
    .ZN(\u_multiplier/pp_13 [4]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_13_1/_18_  (.A(\u_multiplier/STAGE1/pp_12_c2 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_13_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_13_1/_19_  (.A1(\u_multiplier/STAGE1/_209_ ),
    .A2(\u_multiplier/STAGE1/_208_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_13_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_13_1/_20_  (.A(\u_multiplier/STAGE1/_209_ ),
    .B(\u_multiplier/STAGE1/_208_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_13_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_13_1/_21_  (.A1(\u_multiplier/STAGE1/_210_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_13_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_13_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_13_1/_22_  (.A(\u_multiplier/STAGE1/_210_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_13_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_13_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_13_1/_23_  (.A1(\u_multiplier/STAGE1/_211_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_13_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_13_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_13_1/_24_  (.A(\u_multiplier/STAGE1/_211_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_13_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_13_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_13_1/_25_  (.A(\u_multiplier/STAGE1/pp_12_c2 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_13_1/_16_ ),
    .ZN(\u_multiplier/pp_13 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_13_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_13_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_13_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_13_c2 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_13_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_13_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_13_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_13_1/_17_ ),
    .ZN(\u_multiplier/pp_14 [6]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_13_2/_18_  (.A(\u_multiplier/STAGE1/pp_12_c4 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_13_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_13_2/_19_  (.A1(\u_multiplier/STAGE1/_213_ ),
    .A2(\u_multiplier/STAGE1/_212_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_13_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_13_2/_20_  (.A(\u_multiplier/STAGE1/_213_ ),
    .B(\u_multiplier/STAGE1/_212_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_13_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_13_2/_21_  (.A1(\u_multiplier/STAGE1/_214_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_13_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_13_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_13_2/_22_  (.A(\u_multiplier/STAGE1/_214_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_13_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_13_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_13_2/_23_  (.A1(\u_multiplier/STAGE1/_215_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_13_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_13_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_13_2/_24_  (.A(\u_multiplier/STAGE1/_215_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_13_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_13_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_13_2/_25_  (.A(\u_multiplier/STAGE1/pp_12_c4 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_13_2/_16_ ),
    .ZN(\u_multiplier/pp_13 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_13_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_13_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_13_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_13_c4 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_13_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_13_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_13_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_13_2/_17_ ),
    .ZN(\u_multiplier/pp_14 [5]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_13_3/_18_  (.A(net56),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_13_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_13_3/_19_  (.A1(\u_multiplier/STAGE1/_217_ ),
    .A2(\u_multiplier/STAGE1/_216_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_13_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_13_3/_20_  (.A(\u_multiplier/STAGE1/_217_ ),
    .B(\u_multiplier/STAGE1/_216_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_13_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_13_3/_21_  (.A1(\u_multiplier/STAGE1/_218_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_13_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_13_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_13_3/_22_  (.A(\u_multiplier/STAGE1/_218_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_13_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_13_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_13_3/_23_  (.A1(\u_multiplier/STAGE1/_219_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_13_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_13_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_13_3/_24_  (.A(\u_multiplier/STAGE1/_219_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_13_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_13_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_13_3/_25_  (.A(net57),
    .B(\u_multiplier/STAGE1/E_4_2_pp_13_3/_16_ ),
    .ZN(\u_multiplier/pp_13 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_13_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_13_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_13_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_13_c6 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_13_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_13_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_13_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_13_3/_17_ ),
    .ZN(\u_multiplier/pp_14 [4]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_14_1/_18_  (.A(\u_multiplier/STAGE1/pp_13_c2 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_14_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_14_1/_19_  (.A1(\u_multiplier/STAGE1/_221_ ),
    .A2(\u_multiplier/STAGE1/_220_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_14_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_14_1/_20_  (.A(\u_multiplier/STAGE1/_221_ ),
    .B(\u_multiplier/STAGE1/_220_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_14_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_14_1/_21_  (.A1(\u_multiplier/STAGE1/_222_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_14_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_14_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_14_1/_22_  (.A(\u_multiplier/STAGE1/_222_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_14_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_14_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_14_1/_23_  (.A1(\u_multiplier/STAGE1/_223_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_14_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_14_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_14_1/_24_  (.A(\u_multiplier/STAGE1/_223_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_14_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_14_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_14_1/_25_  (.A(\u_multiplier/STAGE1/pp_13_c2 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_14_1/_16_ ),
    .ZN(\u_multiplier/pp_14 [3]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_14_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_14_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_14_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_14_c2 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_14_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_14_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_14_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_14_1/_17_ ),
    .ZN(\u_multiplier/pp_15 [7]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_14_2/_18_  (.A(\u_multiplier/STAGE1/pp_13_c4 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_14_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_14_2/_19_  (.A1(\u_multiplier/STAGE1/_225_ ),
    .A2(\u_multiplier/STAGE1/_224_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_14_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_14_2/_20_  (.A(\u_multiplier/STAGE1/_225_ ),
    .B(\u_multiplier/STAGE1/_224_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_14_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_14_2/_21_  (.A1(\u_multiplier/STAGE1/_226_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_14_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_14_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_14_2/_22_  (.A(\u_multiplier/STAGE1/_226_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_14_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_14_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_14_2/_23_  (.A1(\u_multiplier/STAGE1/_227_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_14_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_14_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_14_2/_24_  (.A(\u_multiplier/STAGE1/_227_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_14_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_14_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_14_2/_25_  (.A(\u_multiplier/STAGE1/pp_13_c4 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_14_2/_16_ ),
    .ZN(\u_multiplier/pp_14 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_14_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_14_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_14_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_14_c4 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_14_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_14_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_14_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_14_2/_17_ ),
    .ZN(\u_multiplier/pp_15 [6]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_14_3/_18_  (.A(\u_multiplier/STAGE1/pp_13_c6 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_14_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_14_3/_19_  (.A1(\u_multiplier/STAGE1/_229_ ),
    .A2(\u_multiplier/STAGE1/_228_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_14_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_14_3/_20_  (.A(\u_multiplier/STAGE1/_229_ ),
    .B(\u_multiplier/STAGE1/_228_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_14_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_14_3/_21_  (.A1(\u_multiplier/STAGE1/_230_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_14_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_14_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_14_3/_22_  (.A(\u_multiplier/STAGE1/_230_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_14_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_14_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_14_3/_23_  (.A1(\u_multiplier/STAGE1/_231_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_14_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_14_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_14_3/_24_  (.A(\u_multiplier/STAGE1/_231_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_14_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_14_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_14_3/_25_  (.A(\u_multiplier/STAGE1/pp_13_c6 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_14_3/_16_ ),
    .ZN(\u_multiplier/pp_14 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_14_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_14_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_14_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_14_c6 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_14_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_14_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_14_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_14_3/_17_ ),
    .ZN(\u_multiplier/pp_15 [5]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_15_1/_18_  (.A(\u_multiplier/STAGE1/pp_14_c2 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_15_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_15_1/_19_  (.A1(\u_multiplier/STAGE1/_235_ ),
    .A2(\u_multiplier/STAGE1/_234_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_15_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_15_1/_20_  (.A(\u_multiplier/STAGE1/_235_ ),
    .B(\u_multiplier/STAGE1/_234_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_15_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_15_1/_21_  (.A1(\u_multiplier/STAGE1/_236_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_15_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_15_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_15_1/_22_  (.A(\u_multiplier/STAGE1/_236_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_15_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_15_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_15_1/_23_  (.A1(\u_multiplier/STAGE1/_237_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_15_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_15_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_15_1/_24_  (.A(\u_multiplier/STAGE1/_237_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_15_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_15_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_15_1/_25_  (.A(\u_multiplier/STAGE1/pp_14_c2 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_15_1/_16_ ),
    .ZN(\u_multiplier/pp_15 [3]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_15_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_15_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_15_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_15_c2 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_15_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_15_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_15_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_15_1/_17_ ),
    .ZN(\u_multiplier/pp_16 [7]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_15_2/_18_  (.A(\u_multiplier/STAGE1/pp_14_c4 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_15_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_15_2/_19_  (.A1(\u_multiplier/STAGE1/_239_ ),
    .A2(\u_multiplier/STAGE1/_238_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_15_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_15_2/_20_  (.A(\u_multiplier/STAGE1/_239_ ),
    .B(\u_multiplier/STAGE1/_238_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_15_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_15_2/_21_  (.A1(\u_multiplier/STAGE1/_240_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_15_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_15_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_15_2/_22_  (.A(\u_multiplier/STAGE1/_240_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_15_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_15_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_15_2/_23_  (.A1(\u_multiplier/STAGE1/_241_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_15_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_15_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_15_2/_24_  (.A(\u_multiplier/STAGE1/_241_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_15_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_15_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_15_2/_25_  (.A(\u_multiplier/STAGE1/pp_14_c4 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_15_2/_16_ ),
    .ZN(\u_multiplier/pp_15 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_15_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_15_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_15_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_15_c4 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_15_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_15_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_15_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_15_2/_17_ ),
    .ZN(\u_multiplier/pp_16 [6]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_15_3/_18_  (.A(\u_multiplier/STAGE1/pp_14_c6 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_15_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_15_3/_19_  (.A1(\u_multiplier/STAGE1/_243_ ),
    .A2(\u_multiplier/STAGE1/_242_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_15_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_15_3/_20_  (.A(\u_multiplier/STAGE1/_243_ ),
    .B(\u_multiplier/STAGE1/_242_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_15_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_15_3/_21_  (.A1(\u_multiplier/STAGE1/_244_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_15_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_15_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_15_3/_22_  (.A(\u_multiplier/STAGE1/_244_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_15_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_15_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_15_3/_23_  (.A1(\u_multiplier/STAGE1/_245_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_15_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_15_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_15_3/_24_  (.A(\u_multiplier/STAGE1/_245_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_15_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_15_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_15_3/_25_  (.A(\u_multiplier/STAGE1/pp_14_c6 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_15_3/_16_ ),
    .ZN(\u_multiplier/pp_15 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_15_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_15_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_15_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_15_c6 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_15_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_15_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_15_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_15_3/_17_ ),
    .ZN(\u_multiplier/pp_16 [5]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_15_4/_18_  (.A(net58),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_15_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_15_4/_19_  (.A1(\u_multiplier/STAGE1/_247_ ),
    .A2(\u_multiplier/STAGE1/_246_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_15_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_15_4/_20_  (.A(\u_multiplier/STAGE1/_247_ ),
    .B(\u_multiplier/STAGE1/_246_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_15_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_15_4/_21_  (.A1(\u_multiplier/STAGE1/_248_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_15_4/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_15_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_15_4/_22_  (.A(\u_multiplier/STAGE1/_248_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_15_4/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_15_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_15_4/_23_  (.A1(\u_multiplier/STAGE1/_249_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_15_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_15_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_15_4/_24_  (.A(\u_multiplier/STAGE1/_249_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_15_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_15_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_15_4/_25_  (.A(net59),
    .B(\u_multiplier/STAGE1/E_4_2_pp_15_4/_16_ ),
    .ZN(\u_multiplier/pp_15 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_15_4/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_15_4/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_15_4/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_15_c8 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_15_4/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_15_4/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_15_4/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_15_4/_17_ ),
    .ZN(\u_multiplier/pp_16 [4]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_16_1/_18_  (.A(\u_multiplier/STAGE1/pp_15_c2 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_1/_19_  (.A1(\u_multiplier/STAGE1/_251_ ),
    .A2(\u_multiplier/STAGE1/_250_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_1/_20_  (.A(\u_multiplier/STAGE1/_251_ ),
    .B(\u_multiplier/STAGE1/_250_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_16_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_1/_21_  (.A1(\u_multiplier/STAGE1/_252_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_16_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_1/_22_  (.A(\u_multiplier/STAGE1/_252_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_16_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_16_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_1/_23_  (.A1(\u_multiplier/STAGE1/_253_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_16_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_1/_24_  (.A(\u_multiplier/STAGE1/_253_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_16_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_1/_25_  (.A(\u_multiplier/STAGE1/pp_15_c2 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_16_1/_16_ ),
    .ZN(\u_multiplier/pp_16 [3]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_16_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_16_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_16_c2 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_16_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_16_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_16_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_16_1/_17_ ),
    .ZN(\u_multiplier/pp_17 [7]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_16_2/_18_  (.A(\u_multiplier/STAGE1/pp_15_c4 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_2/_19_  (.A1(\u_multiplier/STAGE1/_255_ ),
    .A2(\u_multiplier/STAGE1/_254_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_2/_20_  (.A(\u_multiplier/STAGE1/_255_ ),
    .B(\u_multiplier/STAGE1/_254_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_16_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_2/_21_  (.A1(\u_multiplier/STAGE1/_256_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_16_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_2/_22_  (.A(\u_multiplier/STAGE1/_256_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_16_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_16_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_2/_23_  (.A1(\u_multiplier/STAGE1/_257_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_16_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_2/_24_  (.A(\u_multiplier/STAGE1/_257_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_16_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_2/_25_  (.A(\u_multiplier/STAGE1/pp_15_c4 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_16_2/_16_ ),
    .ZN(\u_multiplier/pp_16 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_16_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_16_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_16_c4 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_16_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_16_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_16_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_16_2/_17_ ),
    .ZN(\u_multiplier/pp_17 [6]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_16_3/_18_  (.A(\u_multiplier/STAGE1/pp_15_c6 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_3/_19_  (.A1(\u_multiplier/STAGE1/_259_ ),
    .A2(\u_multiplier/STAGE1/_258_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_3/_20_  (.A(\u_multiplier/STAGE1/_259_ ),
    .B(\u_multiplier/STAGE1/_258_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_16_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_3/_21_  (.A1(\u_multiplier/STAGE1/_260_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_16_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_3/_22_  (.A(\u_multiplier/STAGE1/_260_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_16_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_16_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_3/_23_  (.A1(\u_multiplier/STAGE1/_261_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_16_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_3/_24_  (.A(\u_multiplier/STAGE1/_261_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_16_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_3/_25_  (.A(\u_multiplier/STAGE1/pp_15_c6 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_16_3/_16_ ),
    .ZN(\u_multiplier/pp_16 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_16_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_16_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_16_c6 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_16_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_16_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_16_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_16_3/_17_ ),
    .ZN(\u_multiplier/pp_17 [5]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_16_4/_18_  (.A(net60),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_4/_19_  (.A1(\u_multiplier/STAGE1/_263_ ),
    .A2(\u_multiplier/STAGE1/_262_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_4/_20_  (.A(\u_multiplier/STAGE1/_263_ ),
    .B(\u_multiplier/STAGE1/_262_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_16_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_4/_21_  (.A1(\u_multiplier/STAGE1/_264_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_16_4/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_4/_22_  (.A(\u_multiplier/STAGE1/_264_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_16_4/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_16_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_4/_23_  (.A1(\u_multiplier/STAGE1/pp_15_c8 ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_16_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_4/_24_  (.A(\u_multiplier/STAGE1/pp_15_c8 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_16_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_16_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_16_4/_25_  (.A(net61),
    .B(\u_multiplier/STAGE1/E_4_2_pp_16_4/_16_ ),
    .ZN(\u_multiplier/pp_16 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_16_4/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_16_4/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_16_4/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_16_c8 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_16_4/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_16_4/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_16_4/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_16_4/_17_ ),
    .ZN(\u_multiplier/pp_17 [4]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_17_1/_18_  (.A(\u_multiplier/STAGE1/pp_16_c2 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_1/_19_  (.A1(\u_multiplier/STAGE1/_266_ ),
    .A2(\u_multiplier/STAGE1/_265_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_1/_20_  (.A(\u_multiplier/STAGE1/_266_ ),
    .B(\u_multiplier/STAGE1/_265_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_17_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_1/_21_  (.A1(\u_multiplier/STAGE1/_267_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_17_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_1/_22_  (.A(\u_multiplier/STAGE1/_267_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_17_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_17_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_1/_23_  (.A1(\u_multiplier/STAGE1/_268_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_17_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_1/_24_  (.A(\u_multiplier/STAGE1/_268_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_17_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_1/_25_  (.A(\u_multiplier/STAGE1/pp_16_c2 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_17_1/_16_ ),
    .ZN(\u_multiplier/pp_17 [3]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_17_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_17_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_17_c2 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_17_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_17_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_17_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_17_1/_17_ ),
    .ZN(\u_multiplier/pp_18 [6]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_17_2/_18_  (.A(\u_multiplier/STAGE1/pp_16_c4 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_2/_19_  (.A1(\u_multiplier/STAGE1/_270_ ),
    .A2(\u_multiplier/STAGE1/_269_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_2/_20_  (.A(\u_multiplier/STAGE1/_270_ ),
    .B(\u_multiplier/STAGE1/_269_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_17_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_2/_21_  (.A1(\u_multiplier/STAGE1/_271_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_17_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_2/_22_  (.A(\u_multiplier/STAGE1/_271_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_17_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_17_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_2/_23_  (.A1(\u_multiplier/STAGE1/_272_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_17_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_2/_24_  (.A(\u_multiplier/STAGE1/_272_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_17_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_2/_25_  (.A(\u_multiplier/STAGE1/pp_16_c4 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_17_2/_16_ ),
    .ZN(\u_multiplier/pp_17 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_17_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_17_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_17_c4 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_17_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_17_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_17_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_17_2/_17_ ),
    .ZN(\u_multiplier/pp_18 [5]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_17_3/_18_  (.A(\u_multiplier/STAGE1/pp_16_c6 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_3/_19_  (.A1(\u_multiplier/STAGE1/_274_ ),
    .A2(\u_multiplier/STAGE1/_273_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_3/_20_  (.A(\u_multiplier/STAGE1/_274_ ),
    .B(\u_multiplier/STAGE1/_273_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_17_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_3/_21_  (.A1(\u_multiplier/STAGE1/_275_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_17_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_3/_22_  (.A(\u_multiplier/STAGE1/_275_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_17_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_17_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_3/_23_  (.A1(\u_multiplier/STAGE1/_276_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_17_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_3/_24_  (.A(\u_multiplier/STAGE1/_276_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_17_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_3/_25_  (.A(\u_multiplier/STAGE1/pp_16_c6 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_17_3/_16_ ),
    .ZN(\u_multiplier/pp_17 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_17_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_17_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_17_c6 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_17_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_17_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_17_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_17_3/_17_ ),
    .ZN(\u_multiplier/pp_18 [4]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_18_1/_18_  (.A(\u_multiplier/STAGE1/pp_17_c2 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_18_1/_19_  (.A1(\u_multiplier/STAGE1/_280_ ),
    .A2(\u_multiplier/STAGE1/_279_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_1/_20_  (.A(\u_multiplier/STAGE1/_280_ ),
    .B(\u_multiplier/STAGE1/_279_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_18_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_18_1/_21_  (.A1(\u_multiplier/STAGE1/_281_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_18_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_1/_22_  (.A(\u_multiplier/STAGE1/_281_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_18_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_18_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_18_1/_23_  (.A1(\u_multiplier/STAGE1/_282_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_18_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_1/_24_  (.A(\u_multiplier/STAGE1/_282_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_18_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_1/_25_  (.A(\u_multiplier/STAGE1/pp_17_c2 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_18_1/_16_ ),
    .ZN(\u_multiplier/pp_18 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_18_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_18_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_18_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_18_c2 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_18_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_18_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_18_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_18_1/_17_ ),
    .ZN(\u_multiplier/pp_19 [6]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_18_2/_18_  (.A(\u_multiplier/STAGE1/pp_17_c4 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_18_2/_19_  (.A1(\u_multiplier/STAGE1/_284_ ),
    .A2(\u_multiplier/STAGE1/_283_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_2/_20_  (.A(\u_multiplier/STAGE1/_284_ ),
    .B(\u_multiplier/STAGE1/_283_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_18_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_18_2/_21_  (.A1(\u_multiplier/STAGE1/_285_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_18_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_2/_22_  (.A(\u_multiplier/STAGE1/_285_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_18_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_18_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_18_2/_23_  (.A1(\u_multiplier/STAGE1/_286_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_18_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_2/_24_  (.A(\u_multiplier/STAGE1/_286_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_18_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_2/_25_  (.A(\u_multiplier/STAGE1/pp_17_c4 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_18_2/_16_ ),
    .ZN(\u_multiplier/pp_18 [1]));
 NAND2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_18_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_18_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_18_c4 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_18_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_18_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_18_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_18_2/_17_ ),
    .ZN(\u_multiplier/pp_19 [5]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_18_3/_18_  (.A(\u_multiplier/STAGE1/pp_17_c6 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_18_3/_19_  (.A1(\u_multiplier/STAGE1/_288_ ),
    .A2(\u_multiplier/STAGE1/_287_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_3/_20_  (.A(\u_multiplier/STAGE1/_288_ ),
    .B(\u_multiplier/STAGE1/_287_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_18_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_18_3/_21_  (.A1(\u_multiplier/STAGE1/_289_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_18_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_3/_22_  (.A(\u_multiplier/STAGE1/_289_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_18_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_18_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_18_3/_23_  (.A1(\u_multiplier/STAGE1/_290_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_18_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_3/_24_  (.A(\u_multiplier/STAGE1/_290_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_18_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_3/_25_  (.A(\u_multiplier/STAGE1/pp_17_c6 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_18_3/_16_ ),
    .ZN(\u_multiplier/pp_18 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_18_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_18_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_18_3/_13_ ),
    .ZN(\u_multiplier/pp_19 [3]));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_18_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_18_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_18_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_18_3/_17_ ),
    .ZN(\u_multiplier/pp_19 [4]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_19_1/_18_  (.A(\u_multiplier/STAGE1/pp_18_c2 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_19_1/_19_  (.A1(\u_multiplier/STAGE1/_292_ ),
    .A2(\u_multiplier/STAGE1/_291_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_19_1/_20_  (.A(\u_multiplier/STAGE1/_292_ ),
    .B(\u_multiplier/STAGE1/_291_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_19_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_19_1/_21_  (.A1(\u_multiplier/STAGE1/_293_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_19_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_19_1/_22_  (.A(\u_multiplier/STAGE1/_293_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_19_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_19_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_19_1/_23_  (.A1(\u_multiplier/STAGE1/_294_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_19_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_19_1/_24_  (.A(\u_multiplier/STAGE1/_294_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_19_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_19_1/_25_  (.A(\u_multiplier/STAGE1/pp_18_c2 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_19_1/_16_ ),
    .ZN(\u_multiplier/pp_19 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_19_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_19_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_19_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_19_c2 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_19_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_19_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_19_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_19_1/_17_ ),
    .ZN(\u_multiplier/pp_20 [4]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_19_2/_18_  (.A(\u_multiplier/STAGE1/pp_18_c4 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_19_2/_19_  (.A1(\u_multiplier/STAGE1/_296_ ),
    .A2(\u_multiplier/STAGE1/_295_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_19_2/_20_  (.A(\u_multiplier/STAGE1/_296_ ),
    .B(\u_multiplier/STAGE1/_295_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_19_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_19_2/_21_  (.A1(\u_multiplier/STAGE1/_297_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_19_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_19_2/_22_  (.A(\u_multiplier/STAGE1/_297_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_19_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_19_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_19_2/_23_  (.A1(\u_multiplier/STAGE1/_298_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_19_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_19_2/_24_  (.A(\u_multiplier/STAGE1/_298_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_19_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_19_2/_25_  (.A(\u_multiplier/STAGE1/pp_18_c4 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_19_2/_16_ ),
    .ZN(\u_multiplier/pp_19 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_19_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_19_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_19_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_19_c4 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_19_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_19_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_19_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_19_2/_17_ ),
    .ZN(\u_multiplier/pp_20 [3]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_20_1/_18_  (.A(\u_multiplier/STAGE1/pp_19_c2 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_20_1/_19_  (.A1(\u_multiplier/STAGE1/_303_ ),
    .A2(\u_multiplier/STAGE1/_302_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_20_1/_20_  (.A(\u_multiplier/STAGE1/_303_ ),
    .B(\u_multiplier/STAGE1/_302_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_20_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_20_1/_21_  (.A1(\u_multiplier/STAGE1/_304_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_20_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_20_1/_22_  (.A(\u_multiplier/STAGE1/_304_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_20_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_20_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_20_1/_23_  (.A1(\u_multiplier/STAGE1/_305_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_20_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_20_1/_24_  (.A(\u_multiplier/STAGE1/_305_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_20_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_20_1/_25_  (.A(\u_multiplier/STAGE1/pp_19_c2 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_20_1/_16_ ),
    .ZN(\u_multiplier/pp_20 [1]));
 NAND2_X2 \u_multiplier/STAGE1/E_4_2_pp_20_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_20_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_20_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_20_c2 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_20_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_20_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_20_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_20_1/_17_ ),
    .ZN(\u_multiplier/pp_21 [4]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_20_2/_18_  (.A(\u_multiplier/STAGE1/pp_19_c4 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_20_2/_19_  (.A1(\u_multiplier/STAGE1/_307_ ),
    .A2(\u_multiplier/STAGE1/_306_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_20_2/_20_  (.A(\u_multiplier/STAGE1/_307_ ),
    .B(\u_multiplier/STAGE1/_306_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_20_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_20_2/_21_  (.A1(\u_multiplier/STAGE1/_308_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_20_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_20_2/_22_  (.A(\u_multiplier/STAGE1/_308_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_20_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_20_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_20_2/_23_  (.A1(\u_multiplier/STAGE1/_309_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_20_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_20_2/_24_  (.A(\u_multiplier/STAGE1/_309_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_20_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_20_2/_25_  (.A(\u_multiplier/STAGE1/pp_19_c4 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_20_2/_16_ ),
    .ZN(\u_multiplier/pp_20 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_20_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_20_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_20_2/_13_ ),
    .ZN(\u_multiplier/pp_21 [2]));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_20_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_20_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_20_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_20_2/_17_ ),
    .ZN(\u_multiplier/pp_21 [3]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_21_1/_18_  (.A(\u_multiplier/STAGE1/pp_20_c2 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_21_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_21_1/_19_  (.A1(\u_multiplier/STAGE1/_311_ ),
    .A2(\u_multiplier/STAGE1/_310_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_21_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_21_1/_20_  (.A(\u_multiplier/STAGE1/_311_ ),
    .B(\u_multiplier/STAGE1/_310_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_21_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_21_1/_21_  (.A1(\u_multiplier/STAGE1/_312_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_21_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_21_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_21_1/_22_  (.A(\u_multiplier/STAGE1/_312_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_21_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_21_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_21_1/_23_  (.A1(\u_multiplier/STAGE1/_313_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_21_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_21_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_21_1/_24_  (.A(\u_multiplier/STAGE1/_313_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_21_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_21_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_21_1/_25_  (.A(\u_multiplier/STAGE1/pp_20_c2 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_21_1/_16_ ),
    .ZN(\u_multiplier/pp_21 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_21_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_21_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_21_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_21_c2 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_21_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_21_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_21_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_21_1/_17_ ),
    .ZN(\u_multiplier/pp_22 [2]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_22/_18_  (.A(\u_multiplier/STAGE1/pp_21_c2 ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_22/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_22/_19_  (.A1(\u_multiplier/STAGE1/_318_ ),
    .A2(\u_multiplier/STAGE1/_317_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_22/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_22/_20_  (.A(\u_multiplier/STAGE1/_318_ ),
    .B(\u_multiplier/STAGE1/_317_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_22/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_22/_21_  (.A1(\u_multiplier/STAGE1/_319_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_22/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_22/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_22/_22_  (.A(\u_multiplier/STAGE1/_319_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_22/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_22/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_22/_23_  (.A1(\u_multiplier/STAGE1/_320_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_22/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_22/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_22/_24_  (.A(\u_multiplier/STAGE1/_320_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_22/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_22/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_22/_25_  (.A(\u_multiplier/STAGE1/pp_21_c2 ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_22/_16_ ),
    .ZN(\u_multiplier/pp_22 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_22/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_22/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_22/_13_ ),
    .ZN(\u_multiplier/pp_23 [1]));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_22/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_22/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_22/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_22/_17_ ),
    .ZN(\u_multiplier/pp_23 [2]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_9/_18_  (.A(net62),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_9/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_9/_19_  (.A1(\u_multiplier/STAGE1/_181_ ),
    .A2(\u_multiplier/STAGE1/_180_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_9/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_9/_20_  (.A(\u_multiplier/STAGE1/_181_ ),
    .B(\u_multiplier/STAGE1/_180_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_9/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_9/_21_  (.A1(\u_multiplier/STAGE1/_182_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_9/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_9/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_9/_22_  (.A(\u_multiplier/STAGE1/_182_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_9/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_9/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_9/_23_  (.A1(\u_multiplier/STAGE1/_183_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_9/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_9/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_9/_24_  (.A(\u_multiplier/STAGE1/_183_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_9/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_9/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_9/_25_  (.A(net63),
    .B(\u_multiplier/STAGE1/E_4_2_pp_9/_16_ ),
    .ZN(\u_multiplier/pp_9 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_9/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_9/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_9/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp_9_c2 ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_9/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_9/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_9/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_9/_17_ ),
    .ZN(\u_multiplier/pp_10 [2]));
 INV_X1 \u_multiplier/STAGE1/Full_adder_pp_17/_12_  (.A(\u_multiplier/STAGE1/pp_16_c8 ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_17/_08_ ));
 NAND3_X2 \u_multiplier/STAGE1/Full_adder_pp_17/_13_  (.A1(\u_multiplier/STAGE1/_278_ ),
    .A2(\u_multiplier/STAGE1/_277_ ),
    .A3(\u_multiplier/STAGE1/pp_16_c8 ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_17/_09_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_17/_14_  (.A1(\u_multiplier/STAGE1/_278_ ),
    .A2(\u_multiplier/STAGE1/_277_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_17/_10_ ));
 AOI21_X1 \u_multiplier/STAGE1/Full_adder_pp_17/_15_  (.A(\u_multiplier/STAGE1/pp_16_c8 ),
    .B1(\u_multiplier/STAGE1/_277_ ),
    .B2(\u_multiplier/STAGE1/_278_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_17/_11_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_17/_16_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_17/_10_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_17/_11_ ),
    .ZN(\u_multiplier/pp_18 [3]));
 AOI22_X4 \u_multiplier/STAGE1/Full_adder_pp_17/_17_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_17/_08_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_17/_10_ ),
    .B1(\u_multiplier/pp_18 [3]),
    .B2(\u_multiplier/STAGE1/Full_adder_pp_17/_09_ ),
    .ZN(\u_multiplier/pp_17 [0]));
 INV_X1 \u_multiplier/STAGE1/Full_adder_pp_19/_12_  (.A(\u_multiplier/STAGE1/_301_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_19/_08_ ));
 NAND3_X2 \u_multiplier/STAGE1/Full_adder_pp_19/_13_  (.A1(\u_multiplier/STAGE1/_300_ ),
    .A2(\u_multiplier/STAGE1/_299_ ),
    .A3(\u_multiplier/STAGE1/_301_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_19/_09_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_19/_14_  (.A1(\u_multiplier/STAGE1/_300_ ),
    .A2(\u_multiplier/STAGE1/_299_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_19/_10_ ));
 AOI21_X1 \u_multiplier/STAGE1/Full_adder_pp_19/_15_  (.A(\u_multiplier/STAGE1/_301_ ),
    .B1(\u_multiplier/STAGE1/_299_ ),
    .B2(\u_multiplier/STAGE1/_300_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_19/_11_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_19/_16_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_19/_10_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_19/_11_ ),
    .ZN(\u_multiplier/pp_20 [2]));
 AOI22_X4 \u_multiplier/STAGE1/Full_adder_pp_19/_17_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_19/_08_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_19/_10_ ),
    .B1(\u_multiplier/pp_20 [2]),
    .B2(\u_multiplier/STAGE1/Full_adder_pp_19/_09_ ),
    .ZN(\u_multiplier/pp_19 [0]));
 INV_X1 \u_multiplier/STAGE1/Full_adder_pp_21/_12_  (.A(\u_multiplier/STAGE1/_316_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_21/_08_ ));
 NAND3_X2 \u_multiplier/STAGE1/Full_adder_pp_21/_13_  (.A1(\u_multiplier/STAGE1/_315_ ),
    .A2(\u_multiplier/STAGE1/_314_ ),
    .A3(\u_multiplier/STAGE1/_316_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_21/_09_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_21/_14_  (.A1(\u_multiplier/STAGE1/_315_ ),
    .A2(\u_multiplier/STAGE1/_314_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_21/_10_ ));
 AOI21_X1 \u_multiplier/STAGE1/Full_adder_pp_21/_15_  (.A(\u_multiplier/STAGE1/_316_ ),
    .B1(\u_multiplier/STAGE1/_314_ ),
    .B2(\u_multiplier/STAGE1/_315_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_21/_11_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_21/_16_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_21/_10_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_21/_11_ ),
    .ZN(\u_multiplier/pp_22 [1]));
 AOI22_X4 \u_multiplier/STAGE1/Full_adder_pp_21/_17_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_21/_08_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_21/_10_ ),
    .B1(\u_multiplier/pp_22 [1]),
    .B2(\u_multiplier/STAGE1/Full_adder_pp_21/_09_ ),
    .ZN(\u_multiplier/pp_21 [0]));
 INV_X1 \u_multiplier/STAGE1/Full_adder_pp_23/_12_  (.A(\u_multiplier/STAGE1/_323_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_23/_08_ ));
 NAND3_X2 \u_multiplier/STAGE1/Full_adder_pp_23/_13_  (.A1(\u_multiplier/STAGE1/_322_ ),
    .A2(\u_multiplier/STAGE1/_321_ ),
    .A3(\u_multiplier/STAGE1/_323_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_23/_09_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_23/_14_  (.A1(\u_multiplier/STAGE1/_322_ ),
    .A2(\u_multiplier/STAGE1/_321_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_23/_10_ ));
 AOI21_X1 \u_multiplier/STAGE1/Full_adder_pp_23/_15_  (.A(\u_multiplier/STAGE1/_323_ ),
    .B1(\u_multiplier/STAGE1/_321_ ),
    .B2(\u_multiplier/STAGE1/_322_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_23/_11_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_23/_16_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_23/_10_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_23/_11_ ),
    .ZN(\u_multiplier/pp_24 [0]));
 AOI22_X4 \u_multiplier/STAGE1/Full_adder_pp_23/_17_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_23/_08_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_23/_10_ ),
    .B1(\u_multiplier/pp_24 [0]),
    .B2(\u_multiplier/STAGE1/Full_adder_pp_23/_09_ ),
    .ZN(\u_multiplier/pp_23 [0]));
 AND2_X1 \u_multiplier/STAGE1/Half_adder_pp_10/_4_  (.A1(\u_multiplier/STAGE1/_189_ ),
    .A2(\u_multiplier/STAGE1/_188_ ),
    .ZN(\u_multiplier/pp_11 [3]));
 XOR2_X2 \u_multiplier/STAGE1/Half_adder_pp_10/_5_  (.A(\u_multiplier/STAGE1/_189_ ),
    .B(\u_multiplier/STAGE1/_188_ ),
    .Z(\u_multiplier/pp_10 [0]));
 AND2_X1 \u_multiplier/STAGE1/Half_adder_pp_12/_4_  (.A1(\u_multiplier/STAGE1/_207_ ),
    .A2(\u_multiplier/STAGE1/_206_ ),
    .ZN(\u_multiplier/pp_13 [3]));
 XOR2_X2 \u_multiplier/STAGE1/Half_adder_pp_12/_5_  (.A(\u_multiplier/STAGE1/_207_ ),
    .B(\u_multiplier/STAGE1/_206_ ),
    .Z(\u_multiplier/pp_12 [0]));
 AND2_X1 \u_multiplier/STAGE1/Half_adder_pp_14/_4_  (.A1(\u_multiplier/STAGE1/_233_ ),
    .A2(\u_multiplier/STAGE1/_232_ ),
    .ZN(\u_multiplier/pp_15 [4]));
 XOR2_X2 \u_multiplier/STAGE1/Half_adder_pp_14/_5_  (.A(\u_multiplier/STAGE1/_233_ ),
    .B(\u_multiplier/STAGE1/_232_ ),
    .Z(\u_multiplier/pp_14 [0]));
 AND2_X1 \u_multiplier/STAGE1/Half_adder_pp_8/_4_  (.A1(\u_multiplier/STAGE1/_179_ ),
    .A2(\u_multiplier/STAGE1/_178_ ),
    .ZN(\u_multiplier/pp_9 [1]));
 XOR2_X2 \u_multiplier/STAGE1/Half_adder_pp_8/_5_  (.A(\u_multiplier/STAGE1/_179_ ),
    .B(\u_multiplier/STAGE1/_178_ ),
    .Z(\u_multiplier/pp_8 [0]));
 AND2_X1 \u_multiplier/STAGE1/_434_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[0]),
    .ZN(\u_multiplier/s_0 ));
 AND2_X1 \u_multiplier/STAGE1/_435_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[1]),
    .ZN(\u_multiplier/s_1 [0]));
 AND2_X1 \u_multiplier/STAGE1/_436_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[1]),
    .ZN(\u_multiplier/s_1 [1]));
 AND2_X1 \u_multiplier/STAGE1/_437_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[2]),
    .ZN(\u_multiplier/s_2 [0]));
 AND2_X1 \u_multiplier/STAGE1/_438_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[1]),
    .ZN(\u_multiplier/s_2 [1]));
 AND2_X1 \u_multiplier/STAGE1/_439_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[2]),
    .ZN(\u_multiplier/s_2 [2]));
 AND2_X1 \u_multiplier/STAGE1/_440_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[3]),
    .ZN(\u_multiplier/s_3 [0]));
 AND2_X1 \u_multiplier/STAGE1/_441_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[2]),
    .ZN(\u_multiplier/s_3 [1]));
 AND2_X1 \u_multiplier/STAGE1/_442_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[2]),
    .ZN(\u_multiplier/s_3 [2]));
 AND2_X1 \u_multiplier/STAGE1/_443_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[3]),
    .ZN(\u_multiplier/s_3 [3]));
 AND2_X1 \u_multiplier/STAGE1/_444_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[4]),
    .ZN(\u_multiplier/pp_4 [0]));
 AND2_X1 \u_multiplier/STAGE1/_445_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[3]),
    .ZN(\u_multiplier/pp_4 [1]));
 AND2_X1 \u_multiplier/STAGE1/_446_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[2]),
    .ZN(\u_multiplier/s_4 [1]));
 AND2_X1 \u_multiplier/STAGE1/_447_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[3]),
    .ZN(\u_multiplier/s_4 [2]));
 AND2_X1 \u_multiplier/STAGE1/_448_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[4]),
    .ZN(\u_multiplier/s_4 [3]));
 AND2_X1 \u_multiplier/STAGE1/_449_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[5]),
    .ZN(\u_multiplier/pp_5 [0]));
 AND2_X1 \u_multiplier/STAGE1/_450_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[4]),
    .ZN(\u_multiplier/pp_5 [1]));
 AND2_X1 \u_multiplier/STAGE1/_451_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[3]),
    .ZN(\u_multiplier/pp_5 [2]));
 AND2_X1 \u_multiplier/STAGE1/_452_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[3]),
    .ZN(\u_multiplier/pp_5 [3]));
 AND2_X1 \u_multiplier/STAGE1/_453_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[4]),
    .ZN(\u_multiplier/s_5 [2]));
 AND2_X1 \u_multiplier/STAGE1/_454_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[5]),
    .ZN(\u_multiplier/s_5 [3]));
 AND2_X1 \u_multiplier/STAGE1/_455_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[6]),
    .ZN(\u_multiplier/pp_6 [0]));
 AND2_X1 \u_multiplier/STAGE1/_456_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[5]),
    .ZN(\u_multiplier/pp_6 [1]));
 AND2_X1 \u_multiplier/STAGE1/_457_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[4]),
    .ZN(\u_multiplier/pp_6 [2]));
 AND2_X1 \u_multiplier/STAGE1/_458_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[3]),
    .ZN(\u_multiplier/pp_6 [3]));
 AND2_X1 \u_multiplier/STAGE1/_459_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[4]),
    .ZN(\u_multiplier/pp_6 [4]));
 AND2_X1 \u_multiplier/STAGE1/_460_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[5]),
    .ZN(\u_multiplier/pp_6 [5]));
 AND2_X1 \u_multiplier/STAGE1/_461_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[6]),
    .ZN(\u_multiplier/s_6 [3]));
 AND2_X1 \u_multiplier/STAGE1/_462_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[7]),
    .ZN(\u_multiplier/pp_7 [0]));
 AND2_X1 \u_multiplier/STAGE1/_463_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[6]),
    .ZN(\u_multiplier/pp_7 [1]));
 AND2_X1 \u_multiplier/STAGE1/_464_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[5]),
    .ZN(\u_multiplier/pp_7 [2]));
 AND2_X1 \u_multiplier/STAGE1/_465_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[4]),
    .ZN(\u_multiplier/pp_7 [3]));
 AND2_X1 \u_multiplier/STAGE1/_466_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[4]),
    .ZN(\u_multiplier/pp_7 [4]));
 AND2_X1 \u_multiplier/STAGE1/_467_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[5]),
    .ZN(\u_multiplier/pp_7 [5]));
 AND2_X1 \u_multiplier/STAGE1/_468_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[6]),
    .ZN(\u_multiplier/pp_7 [6]));
 AND2_X1 \u_multiplier/STAGE1/_469_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[7]),
    .ZN(\u_multiplier/pp_7 [7]));
 AND2_X1 \u_multiplier/STAGE1/_470_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[6]),
    .ZN(\u_multiplier/pp_8 [1]));
 AND2_X1 \u_multiplier/STAGE1/_471_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[5]),
    .ZN(\u_multiplier/pp_8 [2]));
 AND2_X1 \u_multiplier/STAGE1/_472_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[4]),
    .ZN(\u_multiplier/pp_8 [3]));
 AND2_X1 \u_multiplier/STAGE1/_473_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[5]),
    .ZN(\u_multiplier/pp_8 [4]));
 AND2_X1 \u_multiplier/STAGE1/_474_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[6]),
    .ZN(\u_multiplier/pp_8 [5]));
 AND2_X1 \u_multiplier/STAGE1/_475_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[7]),
    .ZN(\u_multiplier/pp_8 [6]));
 AND2_X1 \u_multiplier/STAGE1/_476_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/pp_8 [7]));
 AND2_X1 \u_multiplier/STAGE1/_477_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[5]),
    .ZN(\u_multiplier/pp_9 [2]));
 AND2_X1 \u_multiplier/STAGE1/_478_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[5]),
    .ZN(\u_multiplier/pp_9 [3]));
 AND2_X1 \u_multiplier/STAGE1/_479_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[6]),
    .ZN(\u_multiplier/pp_9 [4]));
 AND2_X1 \u_multiplier/STAGE1/_480_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[7]),
    .ZN(\u_multiplier/pp_9 [5]));
 AND2_X1 \u_multiplier/STAGE1/_481_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/pp_9 [6]));
 AND2_X1 \u_multiplier/STAGE1/_482_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/pp_9 [7]));
 AND2_X1 \u_multiplier/STAGE1/_483_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[6]),
    .ZN(\u_multiplier/pp_10 [3]));
 AND2_X1 \u_multiplier/STAGE1/_484_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[7]),
    .ZN(\u_multiplier/pp_10 [4]));
 AND2_X1 \u_multiplier/STAGE1/_485_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/pp_10 [5]));
 AND2_X1 \u_multiplier/STAGE1/_486_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/pp_10 [6]));
 AND2_X1 \u_multiplier/STAGE1/_487_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/pp_10 [7]));
 AND2_X1 \u_multiplier/STAGE1/_488_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/pp_11 [4]));
 AND2_X1 \u_multiplier/STAGE1/_489_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/pp_11 [5]));
 AND2_X1 \u_multiplier/STAGE1/_490_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/pp_11 [6]));
 AND2_X1 \u_multiplier/STAGE1/_491_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/pp_11 [7]));
 AND2_X1 \u_multiplier/STAGE1/_492_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/pp_12 [5]));
 AND2_X1 \u_multiplier/STAGE1/_493_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/pp_12 [6]));
 AND2_X1 \u_multiplier/STAGE1/_494_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/pp_12 [7]));
 AND2_X1 \u_multiplier/STAGE1/_495_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/pp_13 [6]));
 AND2_X1 \u_multiplier/STAGE1/_496_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/pp_13 [7]));
 AND2_X1 \u_multiplier/STAGE1/_497_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/pp_14 [7]));
 AND2_X1 \u_multiplier/STAGE1/_498_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/pp_18 [7]));
 AND2_X1 \u_multiplier/STAGE1/_499_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/pp_19 [7]));
 AND2_X1 \u_multiplier/STAGE1/_500_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/pp_20 [5]));
 AND2_X1 \u_multiplier/STAGE1/_501_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/pp_20 [6]));
 AND2_X1 \u_multiplier/STAGE1/_502_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/pp_20 [7]));
 AND2_X1 \u_multiplier/STAGE1/_503_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/pp_21 [5]));
 AND2_X1 \u_multiplier/STAGE1/_504_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/pp_21 [6]));
 AND2_X1 \u_multiplier/STAGE1/_505_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/pp_21 [7]));
 AND2_X1 \u_multiplier/STAGE1/_506_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/pp_22 [3]));
 AND2_X1 \u_multiplier/STAGE1/_507_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/pp_22 [4]));
 AND2_X1 \u_multiplier/STAGE1/_508_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/pp_22 [5]));
 AND2_X1 \u_multiplier/STAGE1/_509_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/pp_22 [6]));
 AND2_X1 \u_multiplier/STAGE1/_510_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/pp_22 [7]));
 AND2_X1 \u_multiplier/STAGE1/_511_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/pp_23 [3]));
 AND2_X1 \u_multiplier/STAGE1/_512_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/pp_23 [4]));
 AND2_X1 \u_multiplier/STAGE1/_513_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/pp_23 [5]));
 AND2_X1 \u_multiplier/STAGE1/_514_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/pp_23 [6]));
 AND2_X1 \u_multiplier/STAGE1/_515_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/pp_23 [7]));
 AND2_X1 \u_multiplier/STAGE1/_516_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/pp_24 [1]));
 AND2_X1 \u_multiplier/STAGE1/_517_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/pp_24 [2]));
 AND2_X1 \u_multiplier/STAGE1/_518_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/pp_24 [3]));
 AND2_X1 \u_multiplier/STAGE1/_519_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/pp_24 [4]));
 AND2_X1 \u_multiplier/STAGE1/_520_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/pp_24 [5]));
 AND2_X1 \u_multiplier/STAGE1/_521_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/pp_24 [6]));
 AND2_X1 \u_multiplier/STAGE1/_522_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/pp_24 [7]));
 AND2_X1 \u_multiplier/STAGE1/_523_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/pp_25 [0]));
 AND2_X1 \u_multiplier/STAGE1/_524_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/pp_25 [1]));
 AND2_X1 \u_multiplier/STAGE1/_525_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/pp_25 [2]));
 AND2_X1 \u_multiplier/STAGE1/_526_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/pp_25 [3]));
 AND2_X1 \u_multiplier/STAGE1/_527_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/pp_25 [4]));
 AND2_X1 \u_multiplier/STAGE1/_528_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/pp_25 [5]));
 AND2_X1 \u_multiplier/STAGE1/_529_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/pp_26 [0]));
 AND2_X1 \u_multiplier/STAGE1/_530_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/pp_26 [1]));
 AND2_X1 \u_multiplier/STAGE1/_531_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/pp_26 [2]));
 AND2_X1 \u_multiplier/STAGE1/_532_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/pp_26 [3]));
 AND2_X1 \u_multiplier/STAGE1/_533_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/s_26 [3]));
 AND2_X1 \u_multiplier/STAGE1/_534_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/pp_27 [0]));
 AND2_X1 \u_multiplier/STAGE1/_535_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/pp_27 [1]));
 AND2_X1 \u_multiplier/STAGE1/_536_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/pp_27 [2]));
 AND2_X1 \u_multiplier/STAGE1/_537_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/s_27 [3]));
 AND2_X1 \u_multiplier/STAGE1/_538_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/s_28 [1]));
 AND2_X1 \u_multiplier/STAGE1/_539_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/s_28 [2]));
 AND2_X1 \u_multiplier/STAGE1/_540_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/s_28 [3]));
 AND2_X1 \u_multiplier/STAGE1/_541_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/s_29 [0]));
 AND2_X1 \u_multiplier/STAGE1/_542_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/s_29 [1]));
 AND2_X1 \u_multiplier/STAGE1/_543_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/s_30 ));
 AND2_X1 \u_multiplier/STAGE1/_544_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/STAGE1/_178_ ));
 AND2_X1 \u_multiplier/STAGE1/_545_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[7]),
    .ZN(\u_multiplier/STAGE1/_179_ ));
 AND2_X1 \u_multiplier/STAGE1/_546_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/STAGE1/_180_ ));
 AND2_X1 \u_multiplier/STAGE1/_547_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/STAGE1/_181_ ));
 AND2_X1 \u_multiplier/STAGE1/_548_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[7]),
    .ZN(\u_multiplier/STAGE1/_182_ ));
 AND2_X1 \u_multiplier/STAGE1/_549_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[6]),
    .ZN(\u_multiplier/STAGE1/_183_ ));
 AND2_X1 \u_multiplier/STAGE1/_550_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/STAGE1/_184_ ));
 AND2_X1 \u_multiplier/STAGE1/_551_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/STAGE1/_185_ ));
 AND2_X1 \u_multiplier/STAGE1/_552_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/STAGE1/_186_ ));
 AND2_X1 \u_multiplier/STAGE1/_553_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[7]),
    .ZN(\u_multiplier/STAGE1/_187_ ));
 AND2_X1 \u_multiplier/STAGE1/_554_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[6]),
    .ZN(\u_multiplier/STAGE1/_188_ ));
 AND2_X1 \u_multiplier/STAGE1/_555_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[5]),
    .ZN(\u_multiplier/STAGE1/_189_ ));
 AND2_X1 \u_multiplier/STAGE1/_556_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/STAGE1/_190_ ));
 AND2_X1 \u_multiplier/STAGE1/_557_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/STAGE1/_191_ ));
 AND2_X1 \u_multiplier/STAGE1/_558_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/STAGE1/_192_ ));
 AND2_X1 \u_multiplier/STAGE1/_559_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/STAGE1/_193_ ));
 AND2_X1 \u_multiplier/STAGE1/_560_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[7]),
    .ZN(\u_multiplier/STAGE1/_194_ ));
 AND2_X1 \u_multiplier/STAGE1/_561_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[6]),
    .ZN(\u_multiplier/STAGE1/_195_ ));
 AND2_X1 \u_multiplier/STAGE1/_562_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[6]),
    .ZN(\u_multiplier/STAGE1/_196_ ));
 AND2_X1 \u_multiplier/STAGE1/_563_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[7]),
    .ZN(\u_multiplier/STAGE1/_197_ ));
 AND2_X1 \u_multiplier/STAGE1/_564_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/STAGE1/_198_ ));
 AND2_X1 \u_multiplier/STAGE1/_565_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/STAGE1/_199_ ));
 AND2_X1 \u_multiplier/STAGE1/_566_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/STAGE1/_200_ ));
 AND2_X1 \u_multiplier/STAGE1/_567_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/STAGE1/_201_ ));
 AND2_X1 \u_multiplier/STAGE1/_568_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/STAGE1/_202_ ));
 AND2_X1 \u_multiplier/STAGE1/_569_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[7]),
    .ZN(\u_multiplier/STAGE1/_203_ ));
 AND2_X1 \u_multiplier/STAGE1/_570_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[6]),
    .ZN(\u_multiplier/STAGE1/_204_ ));
 AND2_X1 \u_multiplier/STAGE1/_571_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[7]),
    .ZN(\u_multiplier/STAGE1/_205_ ));
 AND2_X1 \u_multiplier/STAGE1/_572_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/STAGE1/_206_ ));
 AND2_X1 \u_multiplier/STAGE1/_573_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/STAGE1/_207_ ));
 AND2_X1 \u_multiplier/STAGE1/_574_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/STAGE1/_208_ ));
 AND2_X1 \u_multiplier/STAGE1/_575_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/STAGE1/_209_ ));
 AND2_X1 \u_multiplier/STAGE1/_576_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/STAGE1/_210_ ));
 AND2_X1 \u_multiplier/STAGE1/_577_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/STAGE1/_211_ ));
 AND2_X1 \u_multiplier/STAGE1/_578_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/STAGE1/_212_ ));
 AND2_X1 \u_multiplier/STAGE1/_579_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/STAGE1/_213_ ));
 AND2_X1 \u_multiplier/STAGE1/_580_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[7]),
    .ZN(\u_multiplier/STAGE1/_214_ ));
 AND2_X1 \u_multiplier/STAGE1/_581_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[7]),
    .ZN(\u_multiplier/STAGE1/_215_ ));
 AND2_X1 \u_multiplier/STAGE1/_582_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/STAGE1/_216_ ));
 AND2_X1 \u_multiplier/STAGE1/_583_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/STAGE1/_217_ ));
 AND2_X1 \u_multiplier/STAGE1/_584_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/STAGE1/_218_ ));
 AND2_X1 \u_multiplier/STAGE1/_585_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/STAGE1/_219_ ));
 AND2_X1 \u_multiplier/STAGE1/_586_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/STAGE1/_220_ ));
 AND2_X1 \u_multiplier/STAGE1/_587_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/STAGE1/_221_ ));
 AND2_X1 \u_multiplier/STAGE1/_588_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/STAGE1/_222_ ));
 AND2_X1 \u_multiplier/STAGE1/_589_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/STAGE1/_223_ ));
 AND2_X1 \u_multiplier/STAGE1/_590_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/STAGE1/_224_ ));
 AND2_X1 \u_multiplier/STAGE1/_591_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/STAGE1/_225_ ));
 AND2_X1 \u_multiplier/STAGE1/_592_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/STAGE1/_226_ ));
 AND2_X1 \u_multiplier/STAGE1/_593_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[7]),
    .ZN(\u_multiplier/STAGE1/_227_ ));
 AND2_X1 \u_multiplier/STAGE1/_594_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/STAGE1/_228_ ));
 AND2_X1 \u_multiplier/STAGE1/_595_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/STAGE1/_229_ ));
 AND2_X1 \u_multiplier/STAGE1/_596_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/STAGE1/_230_ ));
 AND2_X1 \u_multiplier/STAGE1/_597_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/STAGE1/_231_ ));
 AND2_X1 \u_multiplier/STAGE1/_598_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/STAGE1/_232_ ));
 AND2_X1 \u_multiplier/STAGE1/_599_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/STAGE1/_233_ ));
 AND2_X1 \u_multiplier/STAGE1/_600_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/STAGE1/_234_ ));
 AND2_X1 \u_multiplier/STAGE1/_601_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/STAGE1/_235_ ));
 AND2_X1 \u_multiplier/STAGE1/_602_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/STAGE1/_236_ ));
 AND2_X1 \u_multiplier/STAGE1/_603_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/STAGE1/_237_ ));
 AND2_X1 \u_multiplier/STAGE1/_604_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/STAGE1/_238_ ));
 AND2_X1 \u_multiplier/STAGE1/_605_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/STAGE1/_239_ ));
 AND2_X1 \u_multiplier/STAGE1/_606_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/STAGE1/_240_ ));
 AND2_X1 \u_multiplier/STAGE1/_607_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/STAGE1/_241_ ));
 AND2_X1 \u_multiplier/STAGE1/_608_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/STAGE1/_242_ ));
 AND2_X1 \u_multiplier/STAGE1/_609_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/STAGE1/_243_ ));
 AND2_X1 \u_multiplier/STAGE1/_610_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/STAGE1/_244_ ));
 AND2_X1 \u_multiplier/STAGE1/_611_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/STAGE1/_245_ ));
 AND2_X1 \u_multiplier/STAGE1/_612_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/STAGE1/_246_ ));
 AND2_X1 \u_multiplier/STAGE1/_613_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/STAGE1/_247_ ));
 AND2_X1 \u_multiplier/STAGE1/_614_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/STAGE1/_248_ ));
 AND2_X1 \u_multiplier/STAGE1/_615_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/STAGE1/_249_ ));
 AND2_X1 \u_multiplier/STAGE1/_616_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/STAGE1/_250_ ));
 AND2_X1 \u_multiplier/STAGE1/_617_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/STAGE1/_251_ ));
 AND2_X1 \u_multiplier/STAGE1/_618_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/STAGE1/_252_ ));
 AND2_X1 \u_multiplier/STAGE1/_619_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/STAGE1/_253_ ));
 AND2_X1 \u_multiplier/STAGE1/_620_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/STAGE1/_254_ ));
 AND2_X1 \u_multiplier/STAGE1/_621_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/STAGE1/_255_ ));
 AND2_X1 \u_multiplier/STAGE1/_622_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/STAGE1/_256_ ));
 AND2_X1 \u_multiplier/STAGE1/_623_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/STAGE1/_257_ ));
 AND2_X1 \u_multiplier/STAGE1/_624_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/STAGE1/_258_ ));
 AND2_X1 \u_multiplier/STAGE1/_625_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/STAGE1/_259_ ));
 AND2_X1 \u_multiplier/STAGE1/_626_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/STAGE1/_260_ ));
 AND2_X1 \u_multiplier/STAGE1/_627_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/STAGE1/_261_ ));
 AND2_X1 \u_multiplier/STAGE1/_628_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/STAGE1/_262_ ));
 AND2_X1 \u_multiplier/STAGE1/_629_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/STAGE1/_263_ ));
 AND2_X1 \u_multiplier/STAGE1/_630_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/STAGE1/_264_ ));
 AND2_X1 \u_multiplier/STAGE1/_631_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/STAGE1/_265_ ));
 AND2_X1 \u_multiplier/STAGE1/_632_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/STAGE1/_266_ ));
 AND2_X1 \u_multiplier/STAGE1/_633_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/STAGE1/_267_ ));
 AND2_X1 \u_multiplier/STAGE1/_634_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/STAGE1/_268_ ));
 AND2_X1 \u_multiplier/STAGE1/_635_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/STAGE1/_269_ ));
 AND2_X1 \u_multiplier/STAGE1/_636_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/STAGE1/_270_ ));
 AND2_X1 \u_multiplier/STAGE1/_637_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/STAGE1/_271_ ));
 AND2_X1 \u_multiplier/STAGE1/_638_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/STAGE1/_272_ ));
 AND2_X1 \u_multiplier/STAGE1/_639_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/STAGE1/_273_ ));
 AND2_X1 \u_multiplier/STAGE1/_640_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/STAGE1/_274_ ));
 AND2_X1 \u_multiplier/STAGE1/_641_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/STAGE1/_275_ ));
 AND2_X1 \u_multiplier/STAGE1/_642_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/STAGE1/_276_ ));
 AND2_X1 \u_multiplier/STAGE1/_643_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/STAGE1/_277_ ));
 AND2_X1 \u_multiplier/STAGE1/_644_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/STAGE1/_278_ ));
 AND2_X1 \u_multiplier/STAGE1/_645_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/STAGE1/_279_ ));
 AND2_X1 \u_multiplier/STAGE1/_646_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/STAGE1/_280_ ));
 AND2_X1 \u_multiplier/STAGE1/_647_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/STAGE1/_281_ ));
 AND2_X1 \u_multiplier/STAGE1/_648_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/STAGE1/_282_ ));
 AND2_X1 \u_multiplier/STAGE1/_649_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/STAGE1/_283_ ));
 AND2_X1 \u_multiplier/STAGE1/_650_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/STAGE1/_284_ ));
 AND2_X1 \u_multiplier/STAGE1/_651_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/STAGE1/_285_ ));
 AND2_X1 \u_multiplier/STAGE1/_652_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/STAGE1/_286_ ));
 AND2_X1 \u_multiplier/STAGE1/_653_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/STAGE1/_287_ ));
 AND2_X1 \u_multiplier/STAGE1/_654_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/STAGE1/_288_ ));
 AND2_X1 \u_multiplier/STAGE1/_655_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/STAGE1/_289_ ));
 AND2_X1 \u_multiplier/STAGE1/_656_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/STAGE1/_290_ ));
 AND2_X1 \u_multiplier/STAGE1/_657_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/STAGE1/_291_ ));
 AND2_X1 \u_multiplier/STAGE1/_658_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/STAGE1/_292_ ));
 AND2_X1 \u_multiplier/STAGE1/_659_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/STAGE1/_293_ ));
 AND2_X1 \u_multiplier/STAGE1/_660_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/STAGE1/_294_ ));
 AND2_X1 \u_multiplier/STAGE1/_661_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/STAGE1/_295_ ));
 AND2_X1 \u_multiplier/STAGE1/_662_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/STAGE1/_296_ ));
 AND2_X1 \u_multiplier/STAGE1/_663_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/STAGE1/_297_ ));
 AND2_X1 \u_multiplier/STAGE1/_664_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/STAGE1/_298_ ));
 AND2_X1 \u_multiplier/STAGE1/_665_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/STAGE1/_299_ ));
 AND2_X1 \u_multiplier/STAGE1/_666_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/STAGE1/_300_ ));
 AND2_X1 \u_multiplier/STAGE1/_667_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/STAGE1/_301_ ));
 AND2_X1 \u_multiplier/STAGE1/_668_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/STAGE1/_302_ ));
 AND2_X1 \u_multiplier/STAGE1/_669_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/STAGE1/_303_ ));
 AND2_X1 \u_multiplier/STAGE1/_670_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/STAGE1/_304_ ));
 AND2_X1 \u_multiplier/STAGE1/_671_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/STAGE1/_305_ ));
 AND2_X1 \u_multiplier/STAGE1/_672_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/STAGE1/_306_ ));
 AND2_X1 \u_multiplier/STAGE1/_673_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/STAGE1/_307_ ));
 AND2_X1 \u_multiplier/STAGE1/_674_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/STAGE1/_308_ ));
 AND2_X1 \u_multiplier/STAGE1/_675_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/STAGE1/_309_ ));
 AND2_X1 \u_multiplier/STAGE1/_676_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/STAGE1/_310_ ));
 AND2_X1 \u_multiplier/STAGE1/_677_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/STAGE1/_311_ ));
 AND2_X1 \u_multiplier/STAGE1/_678_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/STAGE1/_312_ ));
 AND2_X1 \u_multiplier/STAGE1/_679_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/STAGE1/_313_ ));
 AND2_X1 \u_multiplier/STAGE1/_680_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/STAGE1/_314_ ));
 AND2_X1 \u_multiplier/STAGE1/_681_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/STAGE1/_315_ ));
 AND2_X1 \u_multiplier/STAGE1/_682_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/STAGE1/_316_ ));
 AND2_X1 \u_multiplier/STAGE1/_683_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/STAGE1/_317_ ));
 AND2_X1 \u_multiplier/STAGE1/_684_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/STAGE1/_318_ ));
 AND2_X1 \u_multiplier/STAGE1/_685_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/STAGE1/_319_ ));
 AND2_X1 \u_multiplier/STAGE1/_686_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/STAGE1/_320_ ));
 AND2_X1 \u_multiplier/STAGE1/_687_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/STAGE1/_321_ ));
 AND2_X1 \u_multiplier/STAGE1/_688_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/STAGE1/_322_ ));
 AND2_X1 \u_multiplier/STAGE1/_689_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/STAGE1/_323_ ));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_10_1/_18_  (.A(\u_multiplier/STAGE2/pp_9_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_10_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_10_1/_19_  (.A1(\u_multiplier/pp_10 [1]),
    .A2(\u_multiplier/pp_10 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_10_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_10_1/_20_  (.A(\u_multiplier/pp_10 [1]),
    .B(\u_multiplier/pp_10 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_10_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_10_1/_21_  (.A1(\u_multiplier/pp_10 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_10_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_10_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_10_1/_22_  (.A(\u_multiplier/pp_10 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_10_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_10_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_10_1/_23_  (.A1(\u_multiplier/pp_10 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_10_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_10_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_10_1/_24_  (.A(\u_multiplier/pp_10 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_10_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_10_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_10_1/_25_  (.A(\u_multiplier/STAGE2/pp_9_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_10_1/_16_ ),
    .ZN(\u_multiplier/s_10 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_10_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_10_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_10_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_10_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_10_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_10_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_10_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_10_1/_17_ ),
    .ZN(\u_multiplier/s_11 [1]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_10_2/_18_  (.A(\u_multiplier/STAGE2/pp_9_c4 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_10_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_10_2/_19_  (.A1(\u_multiplier/pp_10 [5]),
    .A2(\u_multiplier/pp_10 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_10_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_10_2/_20_  (.A(\u_multiplier/pp_10 [5]),
    .B(\u_multiplier/pp_10 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_10_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_10_2/_21_  (.A1(\u_multiplier/pp_10 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_10_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_10_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_10_2/_22_  (.A(\u_multiplier/pp_10 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_10_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_10_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_10_2/_23_  (.A1(\u_multiplier/pp_10 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_10_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_10_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_10_2/_24_  (.A(\u_multiplier/pp_10 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_10_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_10_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_10_2/_25_  (.A(\u_multiplier/STAGE2/pp_9_c4 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_10_2/_16_ ),
    .ZN(\u_multiplier/s_10 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_10_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_10_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_10_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_10_c4 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_10_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_10_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_10_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_10_2/_17_ ),
    .ZN(\u_multiplier/s_11 [0]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_11_1/_18_  (.A(\u_multiplier/STAGE2/pp_10_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_11_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_11_1/_19_  (.A1(\u_multiplier/pp_11 [1]),
    .A2(\u_multiplier/pp_11 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_11_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_11_1/_20_  (.A(\u_multiplier/pp_11 [1]),
    .B(\u_multiplier/pp_11 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_11_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_11_1/_21_  (.A1(\u_multiplier/pp_11 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_11_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_11_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_11_1/_22_  (.A(\u_multiplier/pp_11 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_11_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_11_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_11_1/_23_  (.A1(\u_multiplier/pp_11 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_11_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_11_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_11_1/_24_  (.A(\u_multiplier/pp_11 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_11_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_11_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_11_1/_25_  (.A(\u_multiplier/STAGE2/pp_10_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_11_1/_16_ ),
    .ZN(\u_multiplier/s_11 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_11_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_11_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_11_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_11_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_11_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_11_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_11_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_11_1/_17_ ),
    .ZN(\u_multiplier/s_12 [1]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_11_2/_18_  (.A(\u_multiplier/STAGE2/pp_10_c4 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_11_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_11_2/_19_  (.A1(\u_multiplier/pp_11 [5]),
    .A2(\u_multiplier/pp_11 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_11_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_11_2/_20_  (.A(\u_multiplier/pp_11 [5]),
    .B(\u_multiplier/pp_11 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_11_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_11_2/_21_  (.A1(\u_multiplier/pp_11 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_11_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_11_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_11_2/_22_  (.A(\u_multiplier/pp_11 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_11_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_11_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_11_2/_23_  (.A1(\u_multiplier/pp_11 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_11_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_11_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_11_2/_24_  (.A(\u_multiplier/pp_11 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_11_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_11_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_11_2/_25_  (.A(\u_multiplier/STAGE2/pp_10_c4 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_11_2/_16_ ),
    .ZN(\u_multiplier/s_11 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_11_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_11_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_11_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_11_c4 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_11_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_11_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_11_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_11_2/_17_ ),
    .ZN(\u_multiplier/s_12 [0]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_12_1/_18_  (.A(\u_multiplier/STAGE2/pp_11_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_12_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_12_1/_19_  (.A1(\u_multiplier/pp_12 [1]),
    .A2(\u_multiplier/pp_12 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_12_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_12_1/_20_  (.A(\u_multiplier/pp_12 [1]),
    .B(\u_multiplier/pp_12 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_12_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_12_1/_21_  (.A1(\u_multiplier/pp_12 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_12_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_12_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_12_1/_22_  (.A(\u_multiplier/pp_12 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_12_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_12_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_12_1/_23_  (.A1(\u_multiplier/pp_12 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_12_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_12_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_12_1/_24_  (.A(\u_multiplier/pp_12 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_12_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_12_1/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE2/E_4_2_pp_12_1/_25_  (.A(\u_multiplier/STAGE2/pp_11_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_12_1/_16_ ),
    .ZN(\u_multiplier/s_12 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_12_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_12_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_12_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_12_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_12_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_12_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_12_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_12_1/_17_ ),
    .ZN(\u_multiplier/s_13 [1]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_12_2/_18_  (.A(\u_multiplier/STAGE2/pp_11_c4 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_12_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_12_2/_19_  (.A1(\u_multiplier/pp_12 [5]),
    .A2(\u_multiplier/pp_12 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_12_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_12_2/_20_  (.A(\u_multiplier/pp_12 [5]),
    .B(\u_multiplier/pp_12 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_12_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_12_2/_21_  (.A1(\u_multiplier/pp_12 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_12_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_12_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_12_2/_22_  (.A(\u_multiplier/pp_12 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_12_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_12_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_12_2/_23_  (.A1(\u_multiplier/pp_12 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_12_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_12_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_12_2/_24_  (.A(\u_multiplier/pp_12 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_12_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_12_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_12_2/_25_  (.A(\u_multiplier/STAGE2/pp_11_c4 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_12_2/_16_ ),
    .ZN(\u_multiplier/s_12 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_12_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_12_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_12_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_12_c4 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_12_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_12_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_12_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_12_2/_17_ ),
    .ZN(\u_multiplier/s_13 [0]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_13_1/_18_  (.A(\u_multiplier/STAGE2/pp_12_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_13_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_13_1/_19_  (.A1(\u_multiplier/pp_13 [1]),
    .A2(\u_multiplier/pp_13 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_13_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_13_1/_20_  (.A(\u_multiplier/pp_13 [1]),
    .B(\u_multiplier/pp_13 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_13_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_13_1/_21_  (.A1(\u_multiplier/pp_13 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_13_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_13_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_13_1/_22_  (.A(\u_multiplier/pp_13 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_13_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_13_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_13_1/_23_  (.A1(\u_multiplier/pp_13 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_13_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_13_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_13_1/_24_  (.A(\u_multiplier/pp_13 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_13_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_13_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_13_1/_25_  (.A(\u_multiplier/STAGE2/pp_12_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_13_1/_16_ ),
    .ZN(\u_multiplier/s_13 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_13_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_13_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_13_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_13_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_13_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_13_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_13_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_13_1/_17_ ),
    .ZN(\u_multiplier/s_14 [1]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_13_2/_18_  (.A(\u_multiplier/STAGE2/pp_12_c4 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_13_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_13_2/_19_  (.A1(\u_multiplier/pp_13 [5]),
    .A2(\u_multiplier/pp_13 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_13_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_13_2/_20_  (.A(\u_multiplier/pp_13 [5]),
    .B(\u_multiplier/pp_13 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_13_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_13_2/_21_  (.A1(\u_multiplier/pp_13 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_13_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_13_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_13_2/_22_  (.A(\u_multiplier/pp_13 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_13_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_13_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_13_2/_23_  (.A1(\u_multiplier/pp_13 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_13_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_13_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_13_2/_24_  (.A(\u_multiplier/pp_13 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_13_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_13_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_13_2/_25_  (.A(\u_multiplier/STAGE2/pp_12_c4 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_13_2/_16_ ),
    .ZN(\u_multiplier/s_13 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_13_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_13_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_13_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_13_c4 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_13_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_13_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_13_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_13_2/_17_ ),
    .ZN(\u_multiplier/s_14 [0]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_14_1/_18_  (.A(\u_multiplier/STAGE2/pp_13_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_14_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_14_1/_19_  (.A1(\u_multiplier/pp_14 [1]),
    .A2(\u_multiplier/pp_14 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_14_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_14_1/_20_  (.A(\u_multiplier/pp_14 [1]),
    .B(\u_multiplier/pp_14 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_14_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_14_1/_21_  (.A1(\u_multiplier/pp_14 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_14_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_14_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_14_1/_22_  (.A(\u_multiplier/pp_14 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_14_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_14_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_14_1/_23_  (.A1(\u_multiplier/pp_14 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_14_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_14_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_14_1/_24_  (.A(\u_multiplier/pp_14 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_14_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_14_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_14_1/_25_  (.A(\u_multiplier/STAGE2/pp_13_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_14_1/_16_ ),
    .ZN(\u_multiplier/s_14 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_14_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_14_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_14_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_14_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_14_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_14_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_14_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_14_1/_17_ ),
    .ZN(\u_multiplier/s_15 [1]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_14_2/_18_  (.A(\u_multiplier/STAGE2/pp_13_c4 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_14_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_14_2/_19_  (.A1(\u_multiplier/pp_14 [5]),
    .A2(\u_multiplier/pp_14 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_14_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_14_2/_20_  (.A(\u_multiplier/pp_14 [5]),
    .B(\u_multiplier/pp_14 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_14_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_14_2/_21_  (.A1(\u_multiplier/pp_14 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_14_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_14_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_14_2/_22_  (.A(\u_multiplier/pp_14 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_14_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_14_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_14_2/_23_  (.A1(\u_multiplier/pp_14 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_14_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_14_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_14_2/_24_  (.A(\u_multiplier/pp_14 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_14_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_14_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_14_2/_25_  (.A(\u_multiplier/STAGE2/pp_13_c4 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_14_2/_16_ ),
    .ZN(\u_multiplier/s_14 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_14_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_14_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_14_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_14_c4 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_14_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_14_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_14_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_14_2/_17_ ),
    .ZN(\u_multiplier/s_15 [0]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_15_1/_18_  (.A(\u_multiplier/STAGE2/pp_14_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_15_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_15_1/_19_  (.A1(\u_multiplier/pp_15 [1]),
    .A2(\u_multiplier/pp_15 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_15_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_15_1/_20_  (.A(\u_multiplier/pp_15 [1]),
    .B(\u_multiplier/pp_15 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_15_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_15_1/_21_  (.A1(\u_multiplier/pp_15 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_15_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_15_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_15_1/_22_  (.A(\u_multiplier/pp_15 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_15_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_15_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_15_1/_23_  (.A1(\u_multiplier/pp_15 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_15_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_15_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_15_1/_24_  (.A(\u_multiplier/pp_15 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_15_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_15_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_15_1/_25_  (.A(\u_multiplier/STAGE2/pp_14_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_15_1/_16_ ),
    .ZN(\u_multiplier/s_15 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_15_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_15_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_15_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_15_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_15_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_15_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_15_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_15_1/_17_ ),
    .ZN(\u_multiplier/s_16 [1]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_15_2/_18_  (.A(\u_multiplier/STAGE2/pp_14_c4 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_15_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_15_2/_19_  (.A1(\u_multiplier/pp_15 [5]),
    .A2(\u_multiplier/pp_15 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_15_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_15_2/_20_  (.A(\u_multiplier/pp_15 [5]),
    .B(\u_multiplier/pp_15 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_15_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_15_2/_21_  (.A1(\u_multiplier/pp_15 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_15_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_15_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_15_2/_22_  (.A(\u_multiplier/pp_15 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_15_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_15_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_15_2/_23_  (.A1(\u_multiplier/pp_15 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_15_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_15_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_15_2/_24_  (.A(\u_multiplier/pp_15 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_15_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_15_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_15_2/_25_  (.A(\u_multiplier/STAGE2/pp_14_c4 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_15_2/_16_ ),
    .ZN(\u_multiplier/s_15 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_15_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_15_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_15_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_15_c4 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_15_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_15_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_15_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_15_2/_17_ ),
    .ZN(\u_multiplier/s_16 [0]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_16_1/_18_  (.A(\u_multiplier/STAGE2/pp_15_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_16_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_16_1/_19_  (.A1(\u_multiplier/pp_16 [1]),
    .A2(\u_multiplier/pp_16 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_16_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_16_1/_20_  (.A(\u_multiplier/pp_16 [1]),
    .B(\u_multiplier/pp_16 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_16_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_16_1/_21_  (.A1(\u_multiplier/pp_16 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_16_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_16_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_16_1/_22_  (.A(\u_multiplier/pp_16 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_16_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_16_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_16_1/_23_  (.A1(\u_multiplier/pp_16 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_16_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_16_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_16_1/_24_  (.A(\u_multiplier/pp_16 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_16_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_16_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_16_1/_25_  (.A(\u_multiplier/STAGE2/pp_15_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_16_1/_16_ ),
    .ZN(\u_multiplier/s_16 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_16_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_16_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_16_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_16_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_16_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_16_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_16_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_16_1/_17_ ),
    .ZN(\u_multiplier/s_17 [1]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_16_2/_18_  (.A(\u_multiplier/STAGE2/pp_15_c4 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_16_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_16_2/_19_  (.A1(\u_multiplier/pp_16 [5]),
    .A2(\u_multiplier/pp_16 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_16_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_16_2/_20_  (.A(\u_multiplier/pp_16 [5]),
    .B(\u_multiplier/pp_16 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_16_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_16_2/_21_  (.A1(\u_multiplier/pp_16 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_16_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_16_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_16_2/_22_  (.A(\u_multiplier/pp_16 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_16_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_16_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_16_2/_23_  (.A1(\u_multiplier/pp_16 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_16_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_16_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_16_2/_24_  (.A(\u_multiplier/pp_16 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_16_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_16_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_16_2/_25_  (.A(\u_multiplier/STAGE2/pp_15_c4 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_16_2/_16_ ),
    .ZN(\u_multiplier/s_16 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_16_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_16_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_16_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_16_c4 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_16_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_16_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_16_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_16_2/_17_ ),
    .ZN(\u_multiplier/s_17 [0]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_17_1/_18_  (.A(\u_multiplier/STAGE2/pp_16_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_17_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_17_1/_19_  (.A1(\u_multiplier/pp_17 [1]),
    .A2(\u_multiplier/pp_17 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_17_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_17_1/_20_  (.A(\u_multiplier/pp_17 [1]),
    .B(\u_multiplier/pp_17 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_17_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_17_1/_21_  (.A1(\u_multiplier/pp_17 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_17_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_17_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_17_1/_22_  (.A(\u_multiplier/pp_17 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_17_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_17_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_17_1/_23_  (.A1(\u_multiplier/pp_17 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_17_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_17_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_17_1/_24_  (.A(\u_multiplier/pp_17 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_17_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_17_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_17_1/_25_  (.A(\u_multiplier/STAGE2/pp_16_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_17_1/_16_ ),
    .ZN(\u_multiplier/s_17 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_17_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_17_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_17_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_17_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_17_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_17_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_17_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_17_1/_17_ ),
    .ZN(\u_multiplier/s_18 [1]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_17_2/_18_  (.A(\u_multiplier/STAGE2/pp_16_c4 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_17_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_17_2/_19_  (.A1(\u_multiplier/pp_17 [5]),
    .A2(\u_multiplier/pp_17 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_17_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_17_2/_20_  (.A(\u_multiplier/pp_17 [5]),
    .B(\u_multiplier/pp_17 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_17_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_17_2/_21_  (.A1(\u_multiplier/pp_17 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_17_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_17_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_17_2/_22_  (.A(\u_multiplier/pp_17 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_17_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_17_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_17_2/_23_  (.A1(\u_multiplier/pp_17 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_17_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_17_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_17_2/_24_  (.A(\u_multiplier/pp_17 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_17_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_17_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_17_2/_25_  (.A(\u_multiplier/STAGE2/pp_16_c4 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_17_2/_16_ ),
    .ZN(\u_multiplier/s_17 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_17_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_17_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_17_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_17_c4 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_17_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_17_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_17_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_17_2/_17_ ),
    .ZN(\u_multiplier/s_18 [0]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_18_1/_18_  (.A(\u_multiplier/STAGE2/pp_17_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_18_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_18_1/_19_  (.A1(\u_multiplier/pp_18 [1]),
    .A2(\u_multiplier/pp_18 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_18_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_18_1/_20_  (.A(\u_multiplier/pp_18 [1]),
    .B(\u_multiplier/pp_18 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_18_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_18_1/_21_  (.A1(\u_multiplier/pp_18 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_18_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_18_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_18_1/_22_  (.A(\u_multiplier/pp_18 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_18_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_18_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_18_1/_23_  (.A1(\u_multiplier/pp_18 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_18_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_18_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_18_1/_24_  (.A(\u_multiplier/pp_18 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_18_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_18_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_18_1/_25_  (.A(\u_multiplier/STAGE2/pp_17_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_18_1/_16_ ),
    .ZN(\u_multiplier/s_18 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_18_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_18_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_18_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_18_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_18_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_18_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_18_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_18_1/_17_ ),
    .ZN(\u_multiplier/s_19 [1]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_18_2/_18_  (.A(\u_multiplier/STAGE2/pp_17_c4 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_18_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_18_2/_19_  (.A1(\u_multiplier/pp_18 [5]),
    .A2(\u_multiplier/pp_18 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_18_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_18_2/_20_  (.A(\u_multiplier/pp_18 [5]),
    .B(\u_multiplier/pp_18 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_18_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_18_2/_21_  (.A1(\u_multiplier/pp_18 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_18_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_18_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_18_2/_22_  (.A(\u_multiplier/pp_18 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_18_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_18_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_18_2/_23_  (.A1(\u_multiplier/pp_18 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_18_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_18_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_18_2/_24_  (.A(\u_multiplier/pp_18 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_18_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_18_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_18_2/_25_  (.A(\u_multiplier/STAGE2/pp_17_c4 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_18_2/_16_ ),
    .ZN(\u_multiplier/s_18 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_18_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_18_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_18_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_18_c4 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_18_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_18_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_18_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_18_2/_17_ ),
    .ZN(\u_multiplier/s_19 [0]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_19_1/_18_  (.A(\u_multiplier/STAGE2/pp_18_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_19_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_19_1/_19_  (.A1(\u_multiplier/pp_19 [1]),
    .A2(\u_multiplier/pp_19 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_19_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_19_1/_20_  (.A(\u_multiplier/pp_19 [1]),
    .B(\u_multiplier/pp_19 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_19_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_19_1/_21_  (.A1(\u_multiplier/pp_19 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_19_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_19_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_19_1/_22_  (.A(\u_multiplier/pp_19 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_19_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_19_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_19_1/_23_  (.A1(\u_multiplier/pp_19 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_19_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_19_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_19_1/_24_  (.A(\u_multiplier/pp_19 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_19_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_19_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_19_1/_25_  (.A(\u_multiplier/STAGE2/pp_18_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_19_1/_16_ ),
    .ZN(\u_multiplier/s_19 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_19_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_19_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_19_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_19_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_19_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_19_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_19_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_19_1/_17_ ),
    .ZN(\u_multiplier/s_20 [1]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_19_2/_18_  (.A(\u_multiplier/STAGE2/pp_18_c4 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_19_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_19_2/_19_  (.A1(\u_multiplier/pp_19 [5]),
    .A2(\u_multiplier/pp_19 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_19_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_19_2/_20_  (.A(\u_multiplier/pp_19 [5]),
    .B(\u_multiplier/pp_19 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_19_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_19_2/_21_  (.A1(\u_multiplier/pp_19 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_19_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_19_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_19_2/_22_  (.A(\u_multiplier/pp_19 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_19_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_19_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_19_2/_23_  (.A1(\u_multiplier/pp_19 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_19_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_19_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_19_2/_24_  (.A(\u_multiplier/pp_19 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_19_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_19_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_19_2/_25_  (.A(\u_multiplier/STAGE2/pp_18_c4 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_19_2/_16_ ),
    .ZN(\u_multiplier/s_19 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_19_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_19_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_19_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_19_c4 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_19_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_19_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_19_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_19_2/_17_ ),
    .ZN(\u_multiplier/s_20 [0]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_20_1/_18_  (.A(\u_multiplier/STAGE2/pp_19_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_20_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_20_1/_19_  (.A1(\u_multiplier/pp_20 [1]),
    .A2(\u_multiplier/pp_20 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_20_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_20_1/_20_  (.A(\u_multiplier/pp_20 [1]),
    .B(\u_multiplier/pp_20 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_20_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_20_1/_21_  (.A1(\u_multiplier/pp_20 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_20_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_20_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_20_1/_22_  (.A(\u_multiplier/pp_20 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_20_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_20_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_20_1/_23_  (.A1(\u_multiplier/pp_20 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_20_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_20_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_20_1/_24_  (.A(\u_multiplier/pp_20 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_20_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_20_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_20_1/_25_  (.A(\u_multiplier/STAGE2/pp_19_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_20_1/_16_ ),
    .ZN(\u_multiplier/s_20 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_20_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_20_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_20_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_20_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_20_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_20_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_20_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_20_1/_17_ ),
    .ZN(\u_multiplier/s_21 [1]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_20_2/_18_  (.A(\u_multiplier/STAGE2/pp_19_c4 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_20_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_20_2/_19_  (.A1(\u_multiplier/pp_20 [5]),
    .A2(\u_multiplier/pp_20 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_20_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_20_2/_20_  (.A(\u_multiplier/pp_20 [5]),
    .B(\u_multiplier/pp_20 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_20_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_20_2/_21_  (.A1(\u_multiplier/pp_20 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_20_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_20_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_20_2/_22_  (.A(\u_multiplier/pp_20 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_20_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_20_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_20_2/_23_  (.A1(\u_multiplier/pp_20 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_20_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_20_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_20_2/_24_  (.A(\u_multiplier/pp_20 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_20_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_20_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_20_2/_25_  (.A(\u_multiplier/STAGE2/pp_19_c4 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_20_2/_16_ ),
    .ZN(\u_multiplier/s_20 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_20_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_20_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_20_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_20_c4 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_20_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_20_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_20_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_20_2/_17_ ),
    .ZN(\u_multiplier/s_21 [0]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_21_1/_18_  (.A(\u_multiplier/STAGE2/pp_20_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_21_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_21_1/_19_  (.A1(\u_multiplier/pp_21 [1]),
    .A2(\u_multiplier/pp_21 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_21_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_21_1/_20_  (.A(\u_multiplier/pp_21 [1]),
    .B(\u_multiplier/pp_21 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_21_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_21_1/_21_  (.A1(\u_multiplier/pp_21 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_21_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_21_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_21_1/_22_  (.A(\u_multiplier/pp_21 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_21_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_21_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_21_1/_23_  (.A1(\u_multiplier/pp_21 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_21_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_21_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_21_1/_24_  (.A(\u_multiplier/pp_21 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_21_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_21_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_21_1/_25_  (.A(\u_multiplier/STAGE2/pp_20_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_21_1/_16_ ),
    .ZN(\u_multiplier/s_21 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_21_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_21_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_21_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_21_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_21_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_21_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_21_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_21_1/_17_ ),
    .ZN(\u_multiplier/s_22 [1]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_21_2/_18_  (.A(\u_multiplier/STAGE2/pp_20_c4 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_21_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_21_2/_19_  (.A1(\u_multiplier/pp_21 [5]),
    .A2(\u_multiplier/pp_21 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_21_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_21_2/_20_  (.A(\u_multiplier/pp_21 [5]),
    .B(\u_multiplier/pp_21 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_21_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_21_2/_21_  (.A1(\u_multiplier/pp_21 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_21_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_21_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_21_2/_22_  (.A(\u_multiplier/pp_21 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_21_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_21_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_21_2/_23_  (.A1(\u_multiplier/pp_21 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_21_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_21_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_21_2/_24_  (.A(\u_multiplier/pp_21 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_21_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_21_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_21_2/_25_  (.A(\u_multiplier/STAGE2/pp_20_c4 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_21_2/_16_ ),
    .ZN(\u_multiplier/s_21 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_21_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_21_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_21_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_21_c4 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_21_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_21_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_21_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_21_2/_17_ ),
    .ZN(\u_multiplier/s_22 [0]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_22_1/_18_  (.A(\u_multiplier/STAGE2/pp_21_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_22_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_22_1/_19_  (.A1(\u_multiplier/pp_22 [1]),
    .A2(\u_multiplier/pp_22 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_22_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_22_1/_20_  (.A(\u_multiplier/pp_22 [1]),
    .B(\u_multiplier/pp_22 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_22_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_22_1/_21_  (.A1(\u_multiplier/pp_22 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_22_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_22_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_22_1/_22_  (.A(\u_multiplier/pp_22 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_22_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_22_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_22_1/_23_  (.A1(\u_multiplier/pp_22 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_22_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_22_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_22_1/_24_  (.A(\u_multiplier/pp_22 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_22_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_22_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_22_1/_25_  (.A(\u_multiplier/STAGE2/pp_21_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_22_1/_16_ ),
    .ZN(\u_multiplier/s_22 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_22_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_22_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_22_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_22_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_22_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_22_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_22_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_22_1/_17_ ),
    .ZN(\u_multiplier/s_23 [1]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_22_2/_18_  (.A(\u_multiplier/STAGE2/pp_21_c4 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_22_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_22_2/_19_  (.A1(\u_multiplier/pp_22 [5]),
    .A2(\u_multiplier/pp_22 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_22_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_22_2/_20_  (.A(\u_multiplier/pp_22 [5]),
    .B(\u_multiplier/pp_22 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_22_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_22_2/_21_  (.A1(\u_multiplier/pp_22 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_22_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_22_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_22_2/_22_  (.A(\u_multiplier/pp_22 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_22_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_22_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_22_2/_23_  (.A1(\u_multiplier/pp_22 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_22_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_22_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_22_2/_24_  (.A(\u_multiplier/pp_22 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_22_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_22_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_22_2/_25_  (.A(\u_multiplier/STAGE2/pp_21_c4 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_22_2/_16_ ),
    .ZN(\u_multiplier/s_22 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_22_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_22_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_22_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_22_c4 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_22_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_22_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_22_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_22_2/_17_ ),
    .ZN(\u_multiplier/s_23 [0]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_23_1/_18_  (.A(\u_multiplier/STAGE2/pp_22_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_23_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_23_1/_19_  (.A1(\u_multiplier/pp_23 [1]),
    .A2(\u_multiplier/pp_23 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_23_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_23_1/_20_  (.A(\u_multiplier/pp_23 [1]),
    .B(\u_multiplier/pp_23 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_23_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_23_1/_21_  (.A1(\u_multiplier/pp_23 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_23_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_23_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_23_1/_22_  (.A(\u_multiplier/pp_23 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_23_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_23_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_23_1/_23_  (.A1(\u_multiplier/pp_23 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_23_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_23_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_23_1/_24_  (.A(\u_multiplier/pp_23 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_23_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_23_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_23_1/_25_  (.A(\u_multiplier/STAGE2/pp_22_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_23_1/_16_ ),
    .ZN(\u_multiplier/s_23 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_23_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_23_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_23_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_23_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_23_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_23_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_23_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_23_1/_17_ ),
    .ZN(\u_multiplier/s_24 [1]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_23_2/_18_  (.A(\u_multiplier/STAGE2/pp_22_c4 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_23_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_23_2/_19_  (.A1(\u_multiplier/pp_23 [5]),
    .A2(\u_multiplier/pp_23 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_23_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_23_2/_20_  (.A(\u_multiplier/pp_23 [5]),
    .B(\u_multiplier/pp_23 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_23_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_23_2/_21_  (.A1(\u_multiplier/pp_23 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_23_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_23_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_23_2/_22_  (.A(\u_multiplier/pp_23 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_23_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_23_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_23_2/_23_  (.A1(\u_multiplier/pp_23 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_23_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_23_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_23_2/_24_  (.A(\u_multiplier/pp_23 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_23_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_23_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_23_2/_25_  (.A(\u_multiplier/STAGE2/pp_22_c4 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_23_2/_16_ ),
    .ZN(\u_multiplier/s_23 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_23_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_23_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_23_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_23_c4 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_23_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_23_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_23_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_23_2/_17_ ),
    .ZN(\u_multiplier/s_24 [0]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_24_1/_18_  (.A(\u_multiplier/STAGE2/pp_23_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_24_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_24_1/_19_  (.A1(\u_multiplier/pp_24 [1]),
    .A2(\u_multiplier/pp_24 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_24_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_24_1/_20_  (.A(\u_multiplier/pp_24 [1]),
    .B(\u_multiplier/pp_24 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_24_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_24_1/_21_  (.A1(\u_multiplier/pp_24 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_24_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_24_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_24_1/_22_  (.A(\u_multiplier/pp_24 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_24_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_24_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_24_1/_23_  (.A1(\u_multiplier/pp_24 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_24_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_24_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_24_1/_24_  (.A(\u_multiplier/pp_24 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_24_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_24_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_24_1/_25_  (.A(\u_multiplier/STAGE2/pp_23_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_24_1/_16_ ),
    .ZN(\u_multiplier/s_24 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_24_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_24_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_24_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_24_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_24_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_24_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_24_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_24_1/_17_ ),
    .ZN(\u_multiplier/s_25 [1]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_24_2/_18_  (.A(\u_multiplier/STAGE2/pp_23_c4 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_24_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_24_2/_19_  (.A1(\u_multiplier/pp_24 [5]),
    .A2(\u_multiplier/pp_24 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_24_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_24_2/_20_  (.A(\u_multiplier/pp_24 [5]),
    .B(\u_multiplier/pp_24 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_24_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_24_2/_21_  (.A1(\u_multiplier/pp_24 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_24_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_24_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_24_2/_22_  (.A(\u_multiplier/pp_24 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_24_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_24_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_24_2/_23_  (.A1(\u_multiplier/pp_24 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_24_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_24_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_24_2/_24_  (.A(\u_multiplier/pp_24 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_24_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_24_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_24_2/_25_  (.A(\u_multiplier/STAGE2/pp_23_c4 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_24_2/_16_ ),
    .ZN(\u_multiplier/s_24 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_24_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_24_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_24_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_24_c4 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_24_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_24_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_24_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_24_2/_17_ ),
    .ZN(\u_multiplier/s_25 [0]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_25_1/_18_  (.A(\u_multiplier/STAGE2/pp_24_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_25_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_25_1/_19_  (.A1(\u_multiplier/pp_25 [1]),
    .A2(\u_multiplier/pp_25 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_25_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_25_1/_20_  (.A(\u_multiplier/pp_25 [1]),
    .B(\u_multiplier/pp_25 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_25_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_25_1/_21_  (.A1(\u_multiplier/pp_25 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_25_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_25_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_25_1/_22_  (.A(\u_multiplier/pp_25 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_25_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_25_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_25_1/_23_  (.A1(\u_multiplier/pp_25 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_25_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_25_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_25_1/_24_  (.A(\u_multiplier/pp_25 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_25_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_25_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_25_1/_25_  (.A(\u_multiplier/STAGE2/pp_24_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_25_1/_16_ ),
    .ZN(\u_multiplier/s_25 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_25_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_25_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_25_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_25_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_25_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_25_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_25_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_25_1/_17_ ),
    .ZN(\u_multiplier/s_26 [1]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_26_1/_18_  (.A(\u_multiplier/STAGE2/pp_25_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_26_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_26_1/_19_  (.A1(\u_multiplier/pp_26 [1]),
    .A2(\u_multiplier/pp_26 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_26_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_26_1/_20_  (.A(\u_multiplier/pp_26 [1]),
    .B(\u_multiplier/pp_26 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_26_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_26_1/_21_  (.A1(\u_multiplier/pp_26 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_26_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_26_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_26_1/_22_  (.A(\u_multiplier/pp_26 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_26_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_26_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_26_1/_23_  (.A1(\u_multiplier/pp_26 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_26_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_26_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_26_1/_24_  (.A(\u_multiplier/pp_26 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_26_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_26_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_26_1/_25_  (.A(\u_multiplier/STAGE2/pp_25_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_26_1/_16_ ),
    .ZN(\u_multiplier/s_26 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_26_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_26_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_26_1/_13_ ),
    .ZN(\u_multiplier/s_27 [0]));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_26_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_26_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_26_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_26_1/_17_ ),
    .ZN(\u_multiplier/s_27 [1]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_5/_18_  (.A(net64),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_5/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_5/_19_  (.A1(\u_multiplier/pp_5 [1]),
    .A2(\u_multiplier/pp_5 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_5/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_5/_20_  (.A(\u_multiplier/pp_5 [1]),
    .B(\u_multiplier/pp_5 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_5/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_5/_21_  (.A1(\u_multiplier/pp_5 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_5/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_5/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_5/_22_  (.A(\u_multiplier/pp_5 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_5/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_5/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_5/_23_  (.A1(\u_multiplier/pp_5 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_5/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_5/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_5/_24_  (.A(\u_multiplier/pp_5 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_5/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_5/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_5/_25_  (.A(net65),
    .B(\u_multiplier/STAGE2/E_4_2_pp_5/_16_ ),
    .ZN(\u_multiplier/s_5 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_5/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_5/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_5/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_5_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_5/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_5/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_5/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_5/_17_ ),
    .ZN(\u_multiplier/s_6 [2]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_6/_18_  (.A(\u_multiplier/STAGE2/pp_5_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_6/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_6/_19_  (.A1(\u_multiplier/pp_6 [1]),
    .A2(\u_multiplier/pp_6 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_6/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_6/_20_  (.A(\u_multiplier/pp_6 [1]),
    .B(\u_multiplier/pp_6 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_6/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_6/_21_  (.A1(\u_multiplier/pp_6 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_6/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_6/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_6/_22_  (.A(\u_multiplier/pp_6 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_6/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_6/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_6/_23_  (.A1(\u_multiplier/pp_6 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_6/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_6/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_6/_24_  (.A(\u_multiplier/pp_6 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_6/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_6/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_6/_25_  (.A(\u_multiplier/STAGE2/pp_5_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_6/_16_ ),
    .ZN(\u_multiplier/s_6 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_6/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_6/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_6/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_6_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_6/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_6/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_6/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_6/_17_ ),
    .ZN(\u_multiplier/s_7 [1]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_7_1/_18_  (.A(\u_multiplier/STAGE2/pp_6_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_7_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_7_1/_19_  (.A1(\u_multiplier/pp_7 [1]),
    .A2(\u_multiplier/pp_7 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_7_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_7_1/_20_  (.A(\u_multiplier/pp_7 [1]),
    .B(\u_multiplier/pp_7 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_7_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_7_1/_21_  (.A1(\u_multiplier/pp_7 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_7_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_7_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_7_1/_22_  (.A(\u_multiplier/pp_7 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_7_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_7_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_7_1/_23_  (.A1(\u_multiplier/pp_7 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_7_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_7_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_7_1/_24_  (.A(\u_multiplier/pp_7 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_7_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_7_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_7_1/_25_  (.A(\u_multiplier/STAGE2/pp_6_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_7_1/_16_ ),
    .ZN(\u_multiplier/s_7 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_7_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_7_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_7_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_7_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_7_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_7_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_7_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_7_1/_17_ ),
    .ZN(\u_multiplier/s_8 [1]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_7_2/_18_  (.A(net66),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_7_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_7_2/_19_  (.A1(\u_multiplier/pp_7 [5]),
    .A2(\u_multiplier/pp_7 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_7_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_7_2/_20_  (.A(\u_multiplier/pp_7 [5]),
    .B(\u_multiplier/pp_7 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_7_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_7_2/_21_  (.A1(\u_multiplier/pp_7 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_7_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_7_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_7_2/_22_  (.A(\u_multiplier/pp_7 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_7_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_7_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_7_2/_23_  (.A1(\u_multiplier/pp_7 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_7_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_7_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_7_2/_24_  (.A(\u_multiplier/pp_7 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_7_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_7_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_7_2/_25_  (.A(net67),
    .B(\u_multiplier/STAGE2/E_4_2_pp_7_2/_16_ ),
    .ZN(\u_multiplier/s_7 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_7_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_7_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_7_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_7_c4 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_7_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_7_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_7_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_7_2/_17_ ),
    .ZN(\u_multiplier/s_8 [0]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_8_1/_18_  (.A(\u_multiplier/STAGE2/pp_7_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_8_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_8_1/_19_  (.A1(\u_multiplier/pp_8 [1]),
    .A2(\u_multiplier/pp_8 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_8_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_8_1/_20_  (.A(\u_multiplier/pp_8 [1]),
    .B(\u_multiplier/pp_8 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_8_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_8_1/_21_  (.A1(\u_multiplier/pp_8 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_8_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_8_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_8_1/_22_  (.A(\u_multiplier/pp_8 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_8_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_8_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_8_1/_23_  (.A1(\u_multiplier/pp_8 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_8_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_8_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_8_1/_24_  (.A(\u_multiplier/pp_8 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_8_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_8_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_8_1/_25_  (.A(\u_multiplier/STAGE2/pp_7_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_8_1/_16_ ),
    .ZN(\u_multiplier/s_8 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_8_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_8_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_8_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_8_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_8_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_8_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_8_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_8_1/_17_ ),
    .ZN(\u_multiplier/s_9 [1]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_8_2/_18_  (.A(\u_multiplier/STAGE2/pp_7_c4 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_8_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_8_2/_19_  (.A1(\u_multiplier/pp_8 [5]),
    .A2(\u_multiplier/pp_8 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_8_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_8_2/_20_  (.A(\u_multiplier/pp_8 [5]),
    .B(\u_multiplier/pp_8 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_8_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_8_2/_21_  (.A1(\u_multiplier/pp_8 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_8_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_8_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_8_2/_22_  (.A(\u_multiplier/pp_8 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_8_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_8_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_8_2/_23_  (.A1(\u_multiplier/pp_8 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_8_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_8_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_8_2/_24_  (.A(\u_multiplier/pp_8 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_8_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_8_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_8_2/_25_  (.A(\u_multiplier/STAGE2/pp_7_c4 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_8_2/_16_ ),
    .ZN(\u_multiplier/s_8 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_8_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_8_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_8_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_8_c4 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_8_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_8_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_8_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_8_2/_17_ ),
    .ZN(\u_multiplier/s_9 [0]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_9_1/_18_  (.A(\u_multiplier/STAGE2/pp_8_c2 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_9_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_9_1/_19_  (.A1(\u_multiplier/pp_9 [1]),
    .A2(\u_multiplier/pp_9 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_9_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_9_1/_20_  (.A(\u_multiplier/pp_9 [1]),
    .B(\u_multiplier/pp_9 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_9_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_9_1/_21_  (.A1(\u_multiplier/pp_9 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_9_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_9_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_9_1/_22_  (.A(\u_multiplier/pp_9 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_9_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_9_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_9_1/_23_  (.A1(\u_multiplier/pp_9 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_9_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_9_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_9_1/_24_  (.A(\u_multiplier/pp_9 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_9_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_9_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_9_1/_25_  (.A(\u_multiplier/STAGE2/pp_8_c2 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_9_1/_16_ ),
    .ZN(\u_multiplier/s_9 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_9_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_9_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_9_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_9_c2 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_9_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_9_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_9_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_9_1/_17_ ),
    .ZN(\u_multiplier/s_10 [1]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp_9_2/_18_  (.A(\u_multiplier/STAGE2/pp_8_c4 ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_9_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_9_2/_19_  (.A1(\u_multiplier/pp_9 [5]),
    .A2(\u_multiplier/pp_9 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_9_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_9_2/_20_  (.A(\u_multiplier/pp_9 [5]),
    .B(\u_multiplier/pp_9 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_9_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_9_2/_21_  (.A1(\u_multiplier/pp_9 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_9_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_9_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_9_2/_22_  (.A(\u_multiplier/pp_9 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_9_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp_9_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_9_2/_23_  (.A1(\u_multiplier/pp_9 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_9_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_9_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_9_2/_24_  (.A(\u_multiplier/pp_9 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp_9_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp_9_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp_9_2/_25_  (.A(\u_multiplier/STAGE2/pp_8_c4 ),
    .B(\u_multiplier/STAGE2/E_4_2_pp_9_2/_16_ ),
    .ZN(\u_multiplier/s_9 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp_9_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp_9_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp_9_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp_9_c4 ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp_9_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp_9_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp_9_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp_9_2/_17_ ),
    .ZN(\u_multiplier/s_10 [0]));
 INV_X1 \u_multiplier/STAGE2/Full_adder_pp_25/_12_  (.A(\u_multiplier/STAGE2/pp_24_c4 ),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp_25/_08_ ));
 NAND3_X2 \u_multiplier/STAGE2/Full_adder_pp_25/_13_  (.A1(\u_multiplier/pp_25 [5]),
    .A2(\u_multiplier/pp_25 [4]),
    .A3(\u_multiplier/STAGE2/pp_24_c4 ),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp_25/_09_ ));
 NOR2_X2 \u_multiplier/STAGE2/Full_adder_pp_25/_14_  (.A1(\u_multiplier/pp_25 [5]),
    .A2(\u_multiplier/pp_25 [4]),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp_25/_10_ ));
 AOI21_X1 \u_multiplier/STAGE2/Full_adder_pp_25/_15_  (.A(\u_multiplier/STAGE2/pp_24_c4 ),
    .B1(\u_multiplier/pp_25 [4]),
    .B2(\u_multiplier/pp_25 [5]),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp_25/_11_ ));
 NOR2_X2 \u_multiplier/STAGE2/Full_adder_pp_25/_16_  (.A1(\u_multiplier/STAGE2/Full_adder_pp_25/_10_ ),
    .A2(\u_multiplier/STAGE2/Full_adder_pp_25/_11_ ),
    .ZN(\u_multiplier/s_26 [0]));
 AOI22_X4 \u_multiplier/STAGE2/Full_adder_pp_25/_17_  (.A1(\u_multiplier/STAGE2/Full_adder_pp_25/_08_ ),
    .A2(\u_multiplier/STAGE2/Full_adder_pp_25/_10_ ),
    .B1(\u_multiplier/s_26 [0]),
    .B2(\u_multiplier/STAGE2/Full_adder_pp_25/_09_ ),
    .ZN(\u_multiplier/s_25 [2]));
 INV_X1 \u_multiplier/STAGE2/Full_adder_pp_27/_12_  (.A(\u_multiplier/pp_27 [2]),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp_27/_08_ ));
 NAND3_X1 \u_multiplier/STAGE2/Full_adder_pp_27/_13_  (.A1(\u_multiplier/pp_27 [1]),
    .A2(\u_multiplier/pp_27 [0]),
    .A3(\u_multiplier/pp_27 [2]),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp_27/_09_ ));
 NOR2_X2 \u_multiplier/STAGE2/Full_adder_pp_27/_14_  (.A1(\u_multiplier/pp_27 [1]),
    .A2(\u_multiplier/pp_27 [0]),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp_27/_10_ ));
 AOI21_X1 \u_multiplier/STAGE2/Full_adder_pp_27/_15_  (.A(\u_multiplier/pp_27 [2]),
    .B1(\u_multiplier/pp_27 [0]),
    .B2(\u_multiplier/pp_27 [1]),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp_27/_11_ ));
 NOR2_X2 \u_multiplier/STAGE2/Full_adder_pp_27/_16_  (.A1(\u_multiplier/STAGE2/Full_adder_pp_27/_10_ ),
    .A2(\u_multiplier/STAGE2/Full_adder_pp_27/_11_ ),
    .ZN(\u_multiplier/s_28 [0]));
 AOI22_X2 \u_multiplier/STAGE2/Full_adder_pp_27/_17_  (.A1(\u_multiplier/STAGE2/Full_adder_pp_27/_08_ ),
    .A2(\u_multiplier/STAGE2/Full_adder_pp_27/_10_ ),
    .B1(\u_multiplier/s_28 [0]),
    .B2(\u_multiplier/STAGE2/Full_adder_pp_27/_09_ ),
    .ZN(\u_multiplier/s_27 [2]));
 AND2_X1 \u_multiplier/STAGE2/Half_adder_pp_4/_4_  (.A1(\u_multiplier/pp_4 [1]),
    .A2(\u_multiplier/pp_4 [0]),
    .ZN(\u_multiplier/s_5 [1]));
 XOR2_X2 \u_multiplier/STAGE2/Half_adder_pp_4/_5_  (.A(\u_multiplier/pp_4 [1]),
    .B(\u_multiplier/pp_4 [0]),
    .Z(\u_multiplier/s_4 [0]));
 AND2_X1 \u_multiplier/STAGE2/Half_adder_pp_6/_4_  (.A1(\u_multiplier/pp_6 [5]),
    .A2(\u_multiplier/pp_6 [4]),
    .ZN(\u_multiplier/s_7 [0]));
 XOR2_X2 \u_multiplier/STAGE2/Half_adder_pp_6/_5_  (.A(\u_multiplier/pp_6 [5]),
    .B(\u_multiplier/pp_6 [4]),
    .Z(\u_multiplier/s_6 [0]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_10_1/_18_  (.A(\u_multiplier/STAGE3/pp_9_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_10_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_10_1/_19_  (.A1(\u_multiplier/s_10 [1]),
    .A2(\u_multiplier/s_10 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_10_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_10_1/_20_  (.A(\u_multiplier/s_10 [1]),
    .B(\u_multiplier/s_10 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_10_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_10_1/_21_  (.A1(\u_multiplier/s_10 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_10_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_10_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_10_1/_22_  (.A(\u_multiplier/s_10 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_10_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_10_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_10_1/_23_  (.A1(\u_multiplier/s_10 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_10_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_10_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_10_1/_24_  (.A(\u_multiplier/s_10 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_10_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_10_1/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE3/E_4_2_pp_10_1/_25_  (.A(\u_multiplier/STAGE3/pp_9_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_10_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_10_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_10_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_10_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_10_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_10_c2 ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp_10_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_10_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_10_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_10_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_10_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_11_1/_18_  (.A(\u_multiplier/STAGE3/pp_10_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_11_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_11_1/_19_  (.A1(\u_multiplier/s_11 [1]),
    .A2(\u_multiplier/s_11 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_11_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_11_1/_20_  (.A(\u_multiplier/s_11 [1]),
    .B(\u_multiplier/s_11 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_11_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_11_1/_21_  (.A1(\u_multiplier/s_11 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_11_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_11_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_11_1/_22_  (.A(\u_multiplier/s_11 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_11_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_11_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_11_1/_23_  (.A1(\u_multiplier/s_11 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_11_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_11_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_11_1/_24_  (.A(\u_multiplier/s_11 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_11_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_11_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_11_1/_25_  (.A(\u_multiplier/STAGE3/pp_10_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_11_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_11_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_11_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_11_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_11_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_11_c2 ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp_11_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_11_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_11_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_11_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_11_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_12_1/_18_  (.A(\u_multiplier/STAGE3/pp_11_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_12_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_12_1/_19_  (.A1(\u_multiplier/s_12 [1]),
    .A2(\u_multiplier/s_12 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_12_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_12_1/_20_  (.A(\u_multiplier/s_12 [1]),
    .B(\u_multiplier/s_12 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_12_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_12_1/_21_  (.A1(\u_multiplier/s_12 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_12_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_12_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_12_1/_22_  (.A(\u_multiplier/s_12 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_12_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_12_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_12_1/_23_  (.A1(\u_multiplier/s_12 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_12_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_12_1/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE3/E_4_2_pp_12_1/_24_  (.A(\u_multiplier/s_12 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_12_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_12_1/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE3/E_4_2_pp_12_1/_25_  (.A(\u_multiplier/STAGE3/pp_11_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_12_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_12_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_12_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_12_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_12_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_12_c2 ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp_12_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_12_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_12_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_12_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_12_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_13_1/_18_  (.A(\u_multiplier/STAGE3/pp_12_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_13_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_13_1/_19_  (.A1(\u_multiplier/s_13 [1]),
    .A2(\u_multiplier/s_13 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_13_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_13_1/_20_  (.A(\u_multiplier/s_13 [1]),
    .B(\u_multiplier/s_13 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_13_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_13_1/_21_  (.A1(\u_multiplier/s_13 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_13_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_13_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_13_1/_22_  (.A(\u_multiplier/s_13 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_13_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_13_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_13_1/_23_  (.A1(\u_multiplier/s_13 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_13_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_13_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_13_1/_24_  (.A(\u_multiplier/s_13 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_13_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_13_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_13_1/_25_  (.A(\u_multiplier/STAGE3/pp_12_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_13_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_13_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_13_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_13_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_13_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_13_c2 ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp_13_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_13_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_13_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_13_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_13_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_14_1/_18_  (.A(\u_multiplier/STAGE3/pp_13_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_14_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_14_1/_19_  (.A1(\u_multiplier/s_14 [1]),
    .A2(\u_multiplier/s_14 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_14_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_14_1/_20_  (.A(\u_multiplier/s_14 [1]),
    .B(\u_multiplier/s_14 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_14_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_14_1/_21_  (.A1(\u_multiplier/s_14 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_14_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_14_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_14_1/_22_  (.A(\u_multiplier/s_14 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_14_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_14_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_14_1/_23_  (.A1(\u_multiplier/s_14 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_14_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_14_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_14_1/_24_  (.A(\u_multiplier/s_14 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_14_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_14_1/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE3/E_4_2_pp_14_1/_25_  (.A(\u_multiplier/STAGE3/pp_13_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_14_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_14_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_14_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_14_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_14_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_14_c2 ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp_14_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_14_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_14_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_14_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_14_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_15_1/_18_  (.A(\u_multiplier/STAGE3/pp_14_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_15_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_15_1/_19_  (.A1(\u_multiplier/s_15 [1]),
    .A2(\u_multiplier/s_15 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_15_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_15_1/_20_  (.A(\u_multiplier/s_15 [1]),
    .B(\u_multiplier/s_15 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_15_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_15_1/_21_  (.A1(\u_multiplier/s_15 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_15_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_15_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_15_1/_22_  (.A(\u_multiplier/s_15 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_15_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_15_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_15_1/_23_  (.A1(\u_multiplier/s_15 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_15_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_15_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_15_1/_24_  (.A(\u_multiplier/s_15 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_15_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_15_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_15_1/_25_  (.A(\u_multiplier/STAGE3/pp_14_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_15_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_15_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_15_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_15_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_15_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_15_c2 ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp_15_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_15_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_15_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_15_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_15_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_16_1/_18_  (.A(\u_multiplier/STAGE3/pp_15_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_16_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_16_1/_19_  (.A1(\u_multiplier/s_16 [1]),
    .A2(\u_multiplier/s_16 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_16_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_16_1/_20_  (.A(\u_multiplier/s_16 [1]),
    .B(\u_multiplier/s_16 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_16_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_16_1/_21_  (.A1(\u_multiplier/s_16 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_16_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_16_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_16_1/_22_  (.A(\u_multiplier/s_16 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_16_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_16_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_16_1/_23_  (.A1(\u_multiplier/s_16 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_16_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_16_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_16_1/_24_  (.A(\u_multiplier/s_16 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_16_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_16_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_16_1/_25_  (.A(\u_multiplier/STAGE3/pp_15_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_16_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_16_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_16_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_16_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_16_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_16_c2 ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp_16_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_16_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_16_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_16_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_16_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_17_1/_18_  (.A(\u_multiplier/STAGE3/pp_16_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_17_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_17_1/_19_  (.A1(\u_multiplier/s_17 [1]),
    .A2(\u_multiplier/s_17 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_17_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_17_1/_20_  (.A(\u_multiplier/s_17 [1]),
    .B(\u_multiplier/s_17 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_17_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_17_1/_21_  (.A1(\u_multiplier/s_17 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_17_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_17_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_17_1/_22_  (.A(\u_multiplier/s_17 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_17_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_17_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_17_1/_23_  (.A1(\u_multiplier/s_17 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_17_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_17_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_17_1/_24_  (.A(\u_multiplier/s_17 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_17_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_17_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_17_1/_25_  (.A(\u_multiplier/STAGE3/pp_16_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_17_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_17_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_17_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_17_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_17_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_17_c2 ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp_17_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_17_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_17_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_17_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_17_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_18_1/_18_  (.A(\u_multiplier/STAGE3/pp_17_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_18_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_18_1/_19_  (.A1(\u_multiplier/s_18 [1]),
    .A2(\u_multiplier/s_18 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_18_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_18_1/_20_  (.A(\u_multiplier/s_18 [1]),
    .B(\u_multiplier/s_18 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_18_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_18_1/_21_  (.A1(\u_multiplier/s_18 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_18_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_18_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_18_1/_22_  (.A(\u_multiplier/s_18 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_18_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_18_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_18_1/_23_  (.A1(\u_multiplier/s_18 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_18_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_18_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_18_1/_24_  (.A(\u_multiplier/s_18 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_18_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_18_1/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE3/E_4_2_pp_18_1/_25_  (.A(\u_multiplier/STAGE3/pp_17_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_18_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_18_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_18_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_18_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_18_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_18_c2 ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp_18_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_18_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_18_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_18_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_18_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_19_1/_18_  (.A(\u_multiplier/STAGE3/pp_18_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_19_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_19_1/_19_  (.A1(\u_multiplier/s_19 [1]),
    .A2(\u_multiplier/s_19 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_19_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_19_1/_20_  (.A(\u_multiplier/s_19 [1]),
    .B(\u_multiplier/s_19 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_19_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_19_1/_21_  (.A1(\u_multiplier/s_19 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_19_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_19_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_19_1/_22_  (.A(\u_multiplier/s_19 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_19_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_19_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_19_1/_23_  (.A1(\u_multiplier/s_19 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_19_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_19_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_19_1/_24_  (.A(\u_multiplier/s_19 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_19_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_19_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_19_1/_25_  (.A(\u_multiplier/STAGE3/pp_18_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_19_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_19_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_19_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_19_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_19_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_19_c2 ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp_19_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_19_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_19_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_19_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_19_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_20_1/_18_  (.A(\u_multiplier/STAGE3/pp_19_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_20_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_20_1/_19_  (.A1(\u_multiplier/s_20 [1]),
    .A2(\u_multiplier/s_20 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_20_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_20_1/_20_  (.A(\u_multiplier/s_20 [1]),
    .B(\u_multiplier/s_20 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_20_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_20_1/_21_  (.A1(\u_multiplier/s_20 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_20_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_20_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_20_1/_22_  (.A(\u_multiplier/s_20 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_20_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_20_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_20_1/_23_  (.A1(\u_multiplier/s_20 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_20_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_20_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_20_1/_24_  (.A(\u_multiplier/s_20 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_20_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_20_1/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE3/E_4_2_pp_20_1/_25_  (.A(\u_multiplier/STAGE3/pp_19_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_20_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_20_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_20_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_20_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_20_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_20_c2 ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp_20_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_20_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_20_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_20_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_20_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_21_1/_18_  (.A(\u_multiplier/STAGE3/pp_20_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_21_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_21_1/_19_  (.A1(\u_multiplier/s_21 [1]),
    .A2(\u_multiplier/s_21 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_21_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_21_1/_20_  (.A(\u_multiplier/s_21 [1]),
    .B(\u_multiplier/s_21 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_21_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_21_1/_21_  (.A1(\u_multiplier/s_21 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_21_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_21_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_21_1/_22_  (.A(\u_multiplier/s_21 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_21_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_21_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_21_1/_23_  (.A1(\u_multiplier/s_21 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_21_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_21_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_21_1/_24_  (.A(\u_multiplier/s_21 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_21_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_21_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_21_1/_25_  (.A(\u_multiplier/STAGE3/pp_20_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_21_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_21_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_21_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_21_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_21_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_21_c2 ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp_21_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_21_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_21_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_21_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_21_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_22_1/_18_  (.A(\u_multiplier/STAGE3/pp_21_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_22_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_22_1/_19_  (.A1(\u_multiplier/s_22 [1]),
    .A2(\u_multiplier/s_22 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_22_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_22_1/_20_  (.A(\u_multiplier/s_22 [1]),
    .B(\u_multiplier/s_22 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_22_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_22_1/_21_  (.A1(\u_multiplier/s_22 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_22_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_22_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_22_1/_22_  (.A(\u_multiplier/s_22 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_22_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_22_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_22_1/_23_  (.A1(\u_multiplier/s_22 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_22_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_22_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_22_1/_24_  (.A(\u_multiplier/s_22 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_22_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_22_1/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE3/E_4_2_pp_22_1/_25_  (.A(\u_multiplier/STAGE3/pp_21_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_22_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_22_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_22_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_22_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_22_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_22_c2 ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp_22_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_22_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_22_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_22_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_22_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_23_1/_18_  (.A(\u_multiplier/STAGE3/pp_22_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_23_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_23_1/_19_  (.A1(\u_multiplier/s_23 [1]),
    .A2(\u_multiplier/s_23 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_23_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_23_1/_20_  (.A(\u_multiplier/s_23 [1]),
    .B(\u_multiplier/s_23 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_23_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_23_1/_21_  (.A1(\u_multiplier/s_23 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_23_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_23_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_23_1/_22_  (.A(\u_multiplier/s_23 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_23_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_23_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_23_1/_23_  (.A1(\u_multiplier/s_23 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_23_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_23_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_23_1/_24_  (.A(\u_multiplier/s_23 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_23_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_23_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_23_1/_25_  (.A(\u_multiplier/STAGE3/pp_22_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_23_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_23_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_23_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_23_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_23_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_23_c2 ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp_23_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_23_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_23_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_23_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_23_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_24_1/_18_  (.A(\u_multiplier/STAGE3/pp_23_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_24_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_24_1/_19_  (.A1(\u_multiplier/s_24 [1]),
    .A2(\u_multiplier/s_24 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_24_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_24_1/_20_  (.A(\u_multiplier/s_24 [1]),
    .B(\u_multiplier/s_24 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_24_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_24_1/_21_  (.A1(\u_multiplier/s_24 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_24_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_24_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_24_1/_22_  (.A(\u_multiplier/s_24 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_24_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_24_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_24_1/_23_  (.A1(\u_multiplier/s_24 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_24_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_24_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_24_1/_24_  (.A(\u_multiplier/s_24 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_24_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_24_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_24_1/_25_  (.A(\u_multiplier/STAGE3/pp_23_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_24_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_24_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_24_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_24_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_24_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_24_c2 ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp_24_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_24_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_24_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_24_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_24_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_25_1/_18_  (.A(\u_multiplier/STAGE3/pp_24_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_25_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_25_1/_19_  (.A1(\u_multiplier/s_25 [1]),
    .A2(\u_multiplier/s_25 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_25_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_25_1/_20_  (.A(\u_multiplier/s_25 [1]),
    .B(\u_multiplier/s_25 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_25_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_25_1/_21_  (.A1(\u_multiplier/s_25 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_25_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_25_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_25_1/_22_  (.A(\u_multiplier/s_25 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_25_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_25_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_25_1/_23_  (.A1(\u_multiplier/s_25 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_25_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_25_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_25_1/_24_  (.A(\u_multiplier/s_25 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_25_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_25_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_25_1/_25_  (.A(\u_multiplier/STAGE3/pp_24_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_25_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_25_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_25_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_25_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_25_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_25_c2 ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp_25_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_25_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_25_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_25_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_25_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_26_1/_18_  (.A(\u_multiplier/STAGE3/pp_25_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_26_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_26_1/_19_  (.A1(\u_multiplier/s_26 [1]),
    .A2(\u_multiplier/s_26 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_26_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_26_1/_20_  (.A(\u_multiplier/s_26 [1]),
    .B(\u_multiplier/s_26 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_26_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_26_1/_21_  (.A1(\u_multiplier/s_26 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_26_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_26_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_26_1/_22_  (.A(\u_multiplier/s_26 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_26_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_26_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_26_1/_23_  (.A1(\u_multiplier/s_26 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_26_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_26_1/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE3/E_4_2_pp_26_1/_24_  (.A(\u_multiplier/s_26 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_26_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_26_1/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE3/E_4_2_pp_26_1/_25_  (.A(\u_multiplier/STAGE3/pp_25_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_26_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_26_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_26_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_26_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_26_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_26_c2 ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp_26_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_26_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_26_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_26_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_26_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_27_1/_18_  (.A(\u_multiplier/STAGE3/pp_26_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_27_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_27_1/_19_  (.A1(\u_multiplier/s_27 [1]),
    .A2(\u_multiplier/s_27 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_27_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_27_1/_20_  (.A(\u_multiplier/s_27 [1]),
    .B(\u_multiplier/s_27 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_27_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_27_1/_21_  (.A1(\u_multiplier/s_27 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_27_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_27_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_27_1/_22_  (.A(\u_multiplier/s_27 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_27_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_27_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_27_1/_23_  (.A1(\u_multiplier/s_27 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_27_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_27_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_27_1/_24_  (.A(\u_multiplier/s_27 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_27_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_27_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_27_1/_25_  (.A(\u_multiplier/STAGE3/pp_26_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_27_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_27_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_27_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_27_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_27_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_27_c2 ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp_27_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_27_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_27_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_27_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_27_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_28_1/_18_  (.A(\u_multiplier/STAGE3/pp_27_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_28_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_28_1/_19_  (.A1(\u_multiplier/s_28 [1]),
    .A2(\u_multiplier/s_28 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_28_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_28_1/_20_  (.A(\u_multiplier/s_28 [1]),
    .B(\u_multiplier/s_28 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_28_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_28_1/_21_  (.A1(\u_multiplier/s_28 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_28_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_28_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_28_1/_22_  (.A(\u_multiplier/s_28 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_28_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_28_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_28_1/_23_  (.A1(\u_multiplier/s_28 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_28_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_28_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_28_1/_24_  (.A(\u_multiplier/s_28 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_28_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_28_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_28_1/_25_  (.A(\u_multiplier/STAGE3/pp_27_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_28_1/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_28_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_28_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_28_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_28_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_28_c2 ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp_28_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_28_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_28_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_28_1/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_28_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_3/_18_  (.A(net68),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_3/_19_  (.A1(\u_multiplier/s_3 [1]),
    .A2(\u_multiplier/s_3 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_3/_20_  (.A(\u_multiplier/s_3 [1]),
    .B(\u_multiplier/s_3 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_3/_21_  (.A1(\u_multiplier/s_3 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_3/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_3/_22_  (.A(\u_multiplier/s_3 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_3/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_3/_23_  (.A1(\u_multiplier/s_3 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_3/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_3/_24_  (.A(\u_multiplier/s_3 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_3/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_3/_25_  (.A(net69),
    .B(\u_multiplier/STAGE3/E_4_2_pp_3/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_3_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_3/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_3/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_3/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_3_c2 ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp_3/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_3/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_3/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_3/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_3_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_4/_18_  (.A(\u_multiplier/STAGE3/pp_3_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_4/_19_  (.A1(\u_multiplier/s_4 [1]),
    .A2(\u_multiplier/s_4 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_4/_20_  (.A(\u_multiplier/s_4 [1]),
    .B(\u_multiplier/s_4 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_4/_21_  (.A1(\u_multiplier/s_4 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_4/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_4/_22_  (.A(\u_multiplier/s_4 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_4/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_4/_23_  (.A1(\u_multiplier/s_4 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_4/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_4/_24_  (.A(\u_multiplier/s_4 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_4/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_4/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE3/E_4_2_pp_4/_25_  (.A(\u_multiplier/STAGE3/pp_3_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_4/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_4_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_4/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_4/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_4/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_4_c2 ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp_4/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_4/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_4/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_4/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_4_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_5/_18_  (.A(\u_multiplier/STAGE3/pp_4_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_5/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_5/_19_  (.A1(\u_multiplier/s_5 [1]),
    .A2(\u_multiplier/s_5 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_5/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_5/_20_  (.A(\u_multiplier/s_5 [1]),
    .B(\u_multiplier/s_5 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_5/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_5/_21_  (.A1(\u_multiplier/s_5 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_5/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_5/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_5/_22_  (.A(\u_multiplier/s_5 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_5/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_5/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_5/_23_  (.A1(\u_multiplier/s_5 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_5/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_5/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_5/_24_  (.A(\u_multiplier/s_5 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_5/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_5/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_5/_25_  (.A(\u_multiplier/STAGE3/pp_4_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_5/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_5_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_5/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_5/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_5/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_5_c2 ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp_5/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_5/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_5/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_5/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_5_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_6/_18_  (.A(\u_multiplier/STAGE3/pp_5_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_6/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_6/_19_  (.A1(\u_multiplier/s_6 [1]),
    .A2(\u_multiplier/s_6 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_6/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_6/_20_  (.A(\u_multiplier/s_6 [1]),
    .B(\u_multiplier/s_6 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_6/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_6/_21_  (.A1(\u_multiplier/s_6 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_6/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_6/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_6/_22_  (.A(\u_multiplier/s_6 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_6/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_6/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_6/_23_  (.A1(\u_multiplier/s_6 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_6/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_6/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_6/_24_  (.A(\u_multiplier/s_6 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_6/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_6/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE3/E_4_2_pp_6/_25_  (.A(\u_multiplier/STAGE3/pp_5_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_6/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_6_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_6/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_6/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_6/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_6_c2 ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp_6/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_6/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_6/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_6/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_6_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_7/_18_  (.A(\u_multiplier/STAGE3/pp_6_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_7/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_7/_19_  (.A1(\u_multiplier/s_7 [1]),
    .A2(\u_multiplier/s_7 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_7/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_7/_20_  (.A(\u_multiplier/s_7 [1]),
    .B(\u_multiplier/s_7 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_7/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_7/_21_  (.A1(\u_multiplier/s_7 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_7/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_7/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_7/_22_  (.A(\u_multiplier/s_7 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_7/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_7/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_7/_23_  (.A1(\u_multiplier/s_7 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_7/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_7/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_7/_24_  (.A(\u_multiplier/s_7 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_7/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_7/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_7/_25_  (.A(\u_multiplier/STAGE3/pp_6_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_7/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_7_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_7/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_7/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_7/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_7_c2 ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp_7/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_7/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_7/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_7/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_7_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_8/_18_  (.A(\u_multiplier/STAGE3/pp_7_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_8/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_8/_19_  (.A1(\u_multiplier/s_8 [1]),
    .A2(\u_multiplier/s_8 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_8/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_8/_20_  (.A(\u_multiplier/s_8 [1]),
    .B(\u_multiplier/s_8 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_8/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_8/_21_  (.A1(\u_multiplier/s_8 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_8/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_8/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_8/_22_  (.A(\u_multiplier/s_8 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_8/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_8/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_8/_23_  (.A1(\u_multiplier/s_8 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_8/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_8/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_8/_24_  (.A(\u_multiplier/s_8 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_8/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_8/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE3/E_4_2_pp_8/_25_  (.A(\u_multiplier/STAGE3/pp_7_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_8/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_8_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_8/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_8/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_8/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_8_c2 ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp_8/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_8/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_8/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_8/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_8_c1 ));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp_9/_18_  (.A(\u_multiplier/STAGE3/pp_8_c2 ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_9/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_9/_19_  (.A1(\u_multiplier/s_9 [1]),
    .A2(\u_multiplier/s_9 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_9/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_9/_20_  (.A(\u_multiplier/s_9 [1]),
    .B(\u_multiplier/s_9 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_9/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_9/_21_  (.A1(\u_multiplier/s_9 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_9/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_9/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_9/_22_  (.A(\u_multiplier/s_9 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_9/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp_9/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_9/_23_  (.A1(\u_multiplier/s_9 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_9/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_9/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_9/_24_  (.A(\u_multiplier/s_9 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp_9/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp_9/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp_9/_25_  (.A(\u_multiplier/STAGE3/pp_8_c2 ),
    .B(\u_multiplier/STAGE3/E_4_2_pp_9/_16_ ),
    .ZN(\u_multiplier/STAGE3/pp_9_s ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp_9/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp_9/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp_9/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp_9_c2 ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp_9/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp_9/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp_9/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp_9/_17_ ),
    .ZN(\u_multiplier/STAGE3/pp_9_c1 ));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_40_  (.A1(\u_multiplier/STAGE3/pp_2_c ),
    .A2(\u_multiplier/STAGE3/pp_3_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla1/_25_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_41_  (.A1(\u_multiplier/s_2 [2]),
    .A2(\u_multiplier/STAGE3/pp_2_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla1/_26_ ));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_42_  (.A1(\u_multiplier/s_1 [0]),
    .A2(\u_multiplier/s_1 [1]),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla1/_27_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_43_  (.A1(net70),
    .A2(\u_multiplier/s_0 ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla1/_28_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_44_  (.A1(net71),
    .A2(\u_multiplier/s_0 ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla1/_29_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_45_  (.A(net72),
    .B(\u_multiplier/s_0 ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla1/_30_ ));
 AOI21_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_46_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla1/_28_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla1/_29_ ),
    .B2(net73),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla1/_31_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_47_  (.A1(\u_multiplier/s_1 [0]),
    .A2(\u_multiplier/s_1 [1]),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla1/_32_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_48_  (.A(\u_multiplier/s_1 [0]),
    .B(\u_multiplier/s_1 [1]),
    .Z(\u_multiplier/STAGE3/Final_add/cla1/cla1/_33_ ));
 OAI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla1/_49_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla1/_27_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla1/_31_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/cla1/_32_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla1/_34_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_50_  (.A1(\u_multiplier/s_2 [2]),
    .A2(\u_multiplier/STAGE3/pp_2_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla1/_35_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_51_  (.A(\u_multiplier/s_2 [2]),
    .B(\u_multiplier/STAGE3/pp_2_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla1/_36_ ));
 AOI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla1/_52_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla1/_26_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla1/_34_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/cla1/_35_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla1/_37_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_53_  (.A1(\u_multiplier/STAGE3/pp_2_c ),
    .A2(\u_multiplier/STAGE3/pp_3_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla1/_38_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_54_  (.A(\u_multiplier/STAGE3/pp_2_c ),
    .B(\u_multiplier/STAGE3/pp_3_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla1/cla1/_39_ ));
 OAI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla1/_55_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla1/_25_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla1/_37_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/cla1/_38_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/c1 ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_56_  (.A(net74),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla1/_30_ ),
    .ZN(product[0]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_57_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla1/_31_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla1/_33_ ),
    .ZN(product[1]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_58_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla1/_34_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla1/_36_ ),
    .ZN(product[2]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_59_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla1/_37_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla1/_39_ ),
    .ZN(product[3]));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_40_  (.A1(\u_multiplier/STAGE3/pp_6_c1 ),
    .A2(\u_multiplier/STAGE3/pp_7_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla2/_25_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_41_  (.A1(\u_multiplier/STAGE3/pp_5_c1 ),
    .A2(\u_multiplier/STAGE3/pp_6_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla2/_26_ ));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_42_  (.A1(\u_multiplier/STAGE3/pp_4_c1 ),
    .A2(\u_multiplier/STAGE3/pp_5_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla2/_27_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_43_  (.A1(\u_multiplier/STAGE3/pp_3_c1 ),
    .A2(\u_multiplier/STAGE3/pp_4_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla2/_28_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_44_  (.A1(\u_multiplier/STAGE3/pp_3_c1 ),
    .A2(\u_multiplier/STAGE3/pp_4_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla2/_29_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_45_  (.A(\u_multiplier/STAGE3/pp_3_c1 ),
    .B(\u_multiplier/STAGE3/pp_4_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla2/_30_ ));
 AOI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla2/_46_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla2/_28_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla2/_29_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/c1 ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla2/_31_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_47_  (.A1(\u_multiplier/STAGE3/pp_4_c1 ),
    .A2(\u_multiplier/STAGE3/pp_5_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla2/_32_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_48_  (.A(\u_multiplier/STAGE3/pp_4_c1 ),
    .B(\u_multiplier/STAGE3/pp_5_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla1/cla2/_33_ ));
 OAI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla2/_49_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla2/_27_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla2/_31_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/cla2/_32_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla2/_34_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_50_  (.A1(\u_multiplier/STAGE3/pp_5_c1 ),
    .A2(\u_multiplier/STAGE3/pp_6_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla2/_35_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_51_  (.A(\u_multiplier/STAGE3/pp_5_c1 ),
    .B(\u_multiplier/STAGE3/pp_6_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla2/_36_ ));
 AOI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla2/_52_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla2/_26_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla2/_34_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/cla2/_35_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla2/_37_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_53_  (.A1(\u_multiplier/STAGE3/pp_6_c1 ),
    .A2(\u_multiplier/STAGE3/pp_7_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla2/_38_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_54_  (.A(\u_multiplier/STAGE3/pp_6_c1 ),
    .B(\u_multiplier/STAGE3/pp_7_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla1/cla2/_39_ ));
 OAI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla2/_55_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla2/_25_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla2/_37_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/cla2/_38_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/c2 ));
 XNOR2_X2 \u_multiplier/STAGE3/Final_add/cla1/cla2/_56_  (.A(\u_multiplier/STAGE3/Final_add/cla1/c1 ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla2/_30_ ),
    .ZN(product[4]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_57_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla2/_31_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla2/_33_ ),
    .ZN(product[5]));
 XNOR2_X2 \u_multiplier/STAGE3/Final_add/cla1/cla2/_58_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla2/_34_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla2/_36_ ),
    .ZN(product[6]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla2/_59_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla2/_37_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla2/_39_ ),
    .ZN(product[7]));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_40_  (.A1(\u_multiplier/STAGE3/pp_10_c1 ),
    .A2(\u_multiplier/STAGE3/pp_11_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla3/_25_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_41_  (.A1(\u_multiplier/STAGE3/pp_9_c1 ),
    .A2(\u_multiplier/STAGE3/pp_10_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla3/_26_ ));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_42_  (.A1(\u_multiplier/STAGE3/pp_8_c1 ),
    .A2(\u_multiplier/STAGE3/pp_9_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla3/_27_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_43_  (.A1(\u_multiplier/STAGE3/pp_7_c1 ),
    .A2(\u_multiplier/STAGE3/pp_8_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla3/_28_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_44_  (.A1(\u_multiplier/STAGE3/pp_7_c1 ),
    .A2(\u_multiplier/STAGE3/pp_8_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla3/_29_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_45_  (.A(\u_multiplier/STAGE3/pp_7_c1 ),
    .B(\u_multiplier/STAGE3/pp_8_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla3/_30_ ));
 AOI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla3/_46_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla3/_28_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla3/_29_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/c2 ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla3/_31_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_47_  (.A1(\u_multiplier/STAGE3/pp_8_c1 ),
    .A2(\u_multiplier/STAGE3/pp_9_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla3/_32_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_48_  (.A(\u_multiplier/STAGE3/pp_8_c1 ),
    .B(\u_multiplier/STAGE3/pp_9_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla1/cla3/_33_ ));
 OAI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla3/_49_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla3/_27_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla3/_31_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/cla3/_32_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla3/_34_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_50_  (.A1(\u_multiplier/STAGE3/pp_9_c1 ),
    .A2(\u_multiplier/STAGE3/pp_10_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla3/_35_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_51_  (.A(\u_multiplier/STAGE3/pp_9_c1 ),
    .B(\u_multiplier/STAGE3/pp_10_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla3/_36_ ));
 AOI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla3/_52_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla3/_26_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla3/_34_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/cla3/_35_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla3/_37_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_53_  (.A1(\u_multiplier/STAGE3/pp_10_c1 ),
    .A2(\u_multiplier/STAGE3/pp_11_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla3/_38_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_54_  (.A(\u_multiplier/STAGE3/pp_10_c1 ),
    .B(\u_multiplier/STAGE3/pp_11_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla1/cla3/_39_ ));
 OAI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla3/_55_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla3/_25_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla3/_37_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/cla3/_38_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/c3 ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_56_  (.A(\u_multiplier/STAGE3/Final_add/cla1/c2 ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla3/_30_ ),
    .ZN(product[8]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_57_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla3/_31_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla3/_33_ ),
    .ZN(product[9]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_58_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla3/_34_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla3/_36_ ),
    .ZN(product[10]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla3/_59_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla3/_37_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla3/_39_ ),
    .ZN(product[11]));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_40_  (.A1(\u_multiplier/STAGE3/pp_14_c1 ),
    .A2(\u_multiplier/STAGE3/pp_15_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla4/_25_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_41_  (.A1(\u_multiplier/STAGE3/pp_13_c1 ),
    .A2(\u_multiplier/STAGE3/pp_14_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla4/_26_ ));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_42_  (.A1(\u_multiplier/STAGE3/pp_12_c1 ),
    .A2(\u_multiplier/STAGE3/pp_13_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla4/_27_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_43_  (.A1(\u_multiplier/STAGE3/pp_11_c1 ),
    .A2(\u_multiplier/STAGE3/pp_12_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla4/_28_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_44_  (.A1(\u_multiplier/STAGE3/pp_11_c1 ),
    .A2(\u_multiplier/STAGE3/pp_12_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla4/_29_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_45_  (.A(\u_multiplier/STAGE3/pp_11_c1 ),
    .B(\u_multiplier/STAGE3/pp_12_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla4/_30_ ));
 AOI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla4/_46_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla4/_28_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla4/_29_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/c3 ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla4/_31_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_47_  (.A1(\u_multiplier/STAGE3/pp_12_c1 ),
    .A2(\u_multiplier/STAGE3/pp_13_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla4/_32_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_48_  (.A(\u_multiplier/STAGE3/pp_12_c1 ),
    .B(\u_multiplier/STAGE3/pp_13_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla1/cla4/_33_ ));
 OAI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla4/_49_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla4/_27_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla4/_31_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/cla4/_32_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla4/_34_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_50_  (.A1(\u_multiplier/STAGE3/pp_13_c1 ),
    .A2(\u_multiplier/STAGE3/pp_14_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla4/_35_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_51_  (.A(\u_multiplier/STAGE3/pp_13_c1 ),
    .B(\u_multiplier/STAGE3/pp_14_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla4/_36_ ));
 AOI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla4/_52_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla4/_26_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla4/_34_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/cla4/_35_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla4/_37_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_53_  (.A1(\u_multiplier/STAGE3/pp_14_c1 ),
    .A2(\u_multiplier/STAGE3/pp_15_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla1/cla4/_38_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_54_  (.A(\u_multiplier/STAGE3/pp_14_c1 ),
    .B(\u_multiplier/STAGE3/pp_15_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla1/cla4/_39_ ));
 OAI21_X2 \u_multiplier/STAGE3/Final_add/cla1/cla4/_55_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla4/_25_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla1/cla4/_37_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla1/cla4/_38_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/c1 ));
 XNOR2_X2 \u_multiplier/STAGE3/Final_add/cla1/cla4/_56_  (.A(\u_multiplier/STAGE3/Final_add/cla1/c3 ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla4/_30_ ),
    .ZN(product[12]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_57_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla4/_31_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla4/_33_ ),
    .ZN(product[13]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_58_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla4/_34_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla4/_36_ ),
    .ZN(product[14]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla1/cla4/_59_  (.A(\u_multiplier/STAGE3/Final_add/cla1/cla4/_37_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla1/cla4/_39_ ),
    .ZN(product[15]));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_40_  (.A1(\u_multiplier/STAGE3/pp_18_c1 ),
    .A2(\u_multiplier/STAGE3/pp_19_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla1/_25_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_41_  (.A1(\u_multiplier/STAGE3/pp_17_c1 ),
    .A2(\u_multiplier/STAGE3/pp_18_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla1/_26_ ));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_42_  (.A1(\u_multiplier/STAGE3/pp_16_c1 ),
    .A2(\u_multiplier/STAGE3/pp_17_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla1/_27_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_43_  (.A1(\u_multiplier/STAGE3/pp_15_c1 ),
    .A2(\u_multiplier/STAGE3/pp_16_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla1/_28_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_44_  (.A1(\u_multiplier/STAGE3/pp_15_c1 ),
    .A2(\u_multiplier/STAGE3/pp_16_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla1/_29_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_45_  (.A(\u_multiplier/STAGE3/pp_15_c1 ),
    .B(\u_multiplier/STAGE3/pp_16_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla1/_30_ ));
 AOI21_X2 \u_multiplier/STAGE3/Final_add/cla2/cla1/_46_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla1/_28_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla1/_29_ ),
    .B2(\u_multiplier/STAGE3/Final_add/c1 ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla1/_31_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_47_  (.A1(\u_multiplier/STAGE3/pp_16_c1 ),
    .A2(\u_multiplier/STAGE3/pp_17_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla1/_32_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_48_  (.A(\u_multiplier/STAGE3/pp_16_c1 ),
    .B(\u_multiplier/STAGE3/pp_17_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla2/cla1/_33_ ));
 OAI21_X2 \u_multiplier/STAGE3/Final_add/cla2/cla1/_49_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla1/_27_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla1/_31_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/cla1/_32_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla1/_34_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_50_  (.A1(\u_multiplier/STAGE3/pp_17_c1 ),
    .A2(\u_multiplier/STAGE3/pp_18_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla1/_35_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_51_  (.A(\u_multiplier/STAGE3/pp_17_c1 ),
    .B(\u_multiplier/STAGE3/pp_18_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla1/_36_ ));
 AOI21_X2 \u_multiplier/STAGE3/Final_add/cla2/cla1/_52_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla1/_26_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla1/_34_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/cla1/_35_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla1/_37_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_53_  (.A1(\u_multiplier/STAGE3/pp_18_c1 ),
    .A2(\u_multiplier/STAGE3/pp_19_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla1/_38_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_54_  (.A(\u_multiplier/STAGE3/pp_18_c1 ),
    .B(\u_multiplier/STAGE3/pp_19_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla2/cla1/_39_ ));
 OAI21_X2 \u_multiplier/STAGE3/Final_add/cla2/cla1/_55_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla1/_25_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla1/_37_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/cla1/_38_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/c1 ));
 XNOR2_X2 \u_multiplier/STAGE3/Final_add/cla2/cla1/_56_  (.A(\u_multiplier/STAGE3/Final_add/c1 ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla1/_30_ ),
    .ZN(product[16]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_57_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla1/_31_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla1/_33_ ),
    .ZN(product[17]));
 XNOR2_X2 \u_multiplier/STAGE3/Final_add/cla2/cla1/_58_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla1/_34_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla1/_36_ ),
    .ZN(product[18]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla1/_59_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla1/_37_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla1/_39_ ),
    .ZN(product[19]));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_40_  (.A1(\u_multiplier/STAGE3/pp_22_c1 ),
    .A2(\u_multiplier/STAGE3/pp_23_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla2/_25_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_41_  (.A1(\u_multiplier/STAGE3/pp_21_c1 ),
    .A2(\u_multiplier/STAGE3/pp_22_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla2/_26_ ));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_42_  (.A1(\u_multiplier/STAGE3/pp_20_c1 ),
    .A2(\u_multiplier/STAGE3/pp_21_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla2/_27_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_43_  (.A1(\u_multiplier/STAGE3/pp_19_c1 ),
    .A2(\u_multiplier/STAGE3/pp_20_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla2/_28_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_44_  (.A1(\u_multiplier/STAGE3/pp_19_c1 ),
    .A2(\u_multiplier/STAGE3/pp_20_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla2/_29_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_45_  (.A(\u_multiplier/STAGE3/pp_19_c1 ),
    .B(\u_multiplier/STAGE3/pp_20_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla2/_30_ ));
 AOI21_X2 \u_multiplier/STAGE3/Final_add/cla2/cla2/_46_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla2/_28_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla2/_29_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/c1 ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla2/_31_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_47_  (.A1(\u_multiplier/STAGE3/pp_20_c1 ),
    .A2(\u_multiplier/STAGE3/pp_21_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla2/_32_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_48_  (.A(\u_multiplier/STAGE3/pp_20_c1 ),
    .B(\u_multiplier/STAGE3/pp_21_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla2/cla2/_33_ ));
 OAI21_X2 \u_multiplier/STAGE3/Final_add/cla2/cla2/_49_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla2/_27_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla2/_31_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/cla2/_32_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla2/_34_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_50_  (.A1(\u_multiplier/STAGE3/pp_21_c1 ),
    .A2(\u_multiplier/STAGE3/pp_22_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla2/_35_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_51_  (.A(\u_multiplier/STAGE3/pp_21_c1 ),
    .B(\u_multiplier/STAGE3/pp_22_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla2/_36_ ));
 AOI21_X2 \u_multiplier/STAGE3/Final_add/cla2/cla2/_52_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla2/_26_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla2/_34_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/cla2/_35_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla2/_37_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_53_  (.A1(\u_multiplier/STAGE3/pp_22_c1 ),
    .A2(\u_multiplier/STAGE3/pp_23_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla2/_38_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_54_  (.A(\u_multiplier/STAGE3/pp_22_c1 ),
    .B(\u_multiplier/STAGE3/pp_23_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla2/cla2/_39_ ));
 OAI21_X2 \u_multiplier/STAGE3/Final_add/cla2/cla2/_55_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla2/_25_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla2/_37_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/cla2/_38_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/c2 ));
 XNOR2_X2 \u_multiplier/STAGE3/Final_add/cla2/cla2/_56_  (.A(\u_multiplier/STAGE3/Final_add/cla2/c1 ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla2/_30_ ),
    .ZN(product[20]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_57_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla2/_31_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla2/_33_ ),
    .ZN(product[21]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_58_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla2/_34_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla2/_36_ ),
    .ZN(product[22]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla2/_59_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla2/_37_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla2/_39_ ),
    .ZN(product[23]));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_40_  (.A1(\u_multiplier/STAGE3/pp_26_c1 ),
    .A2(\u_multiplier/STAGE3/pp_27_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla3/_25_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_41_  (.A1(\u_multiplier/STAGE3/pp_25_c1 ),
    .A2(\u_multiplier/STAGE3/pp_26_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla3/_26_ ));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_42_  (.A1(\u_multiplier/STAGE3/pp_24_c1 ),
    .A2(\u_multiplier/STAGE3/pp_25_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla3/_27_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_43_  (.A1(\u_multiplier/STAGE3/pp_23_c1 ),
    .A2(\u_multiplier/STAGE3/pp_24_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla3/_28_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_44_  (.A1(\u_multiplier/STAGE3/pp_23_c1 ),
    .A2(\u_multiplier/STAGE3/pp_24_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla3/_29_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_45_  (.A(\u_multiplier/STAGE3/pp_23_c1 ),
    .B(\u_multiplier/STAGE3/pp_24_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla3/_30_ ));
 AOI21_X2 \u_multiplier/STAGE3/Final_add/cla2/cla3/_46_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla3/_28_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla3/_29_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/c2 ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla3/_31_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_47_  (.A1(\u_multiplier/STAGE3/pp_24_c1 ),
    .A2(\u_multiplier/STAGE3/pp_25_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla3/_32_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_48_  (.A(\u_multiplier/STAGE3/pp_24_c1 ),
    .B(\u_multiplier/STAGE3/pp_25_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla2/cla3/_33_ ));
 OAI21_X2 \u_multiplier/STAGE3/Final_add/cla2/cla3/_49_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla3/_27_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla3/_31_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/cla3/_32_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla3/_34_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_50_  (.A1(\u_multiplier/STAGE3/pp_25_c1 ),
    .A2(\u_multiplier/STAGE3/pp_26_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla3/_35_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_51_  (.A(\u_multiplier/STAGE3/pp_25_c1 ),
    .B(\u_multiplier/STAGE3/pp_26_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla3/_36_ ));
 AOI21_X2 \u_multiplier/STAGE3/Final_add/cla2/cla3/_52_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla3/_26_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla3/_34_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/cla3/_35_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla3/_37_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_53_  (.A1(\u_multiplier/STAGE3/pp_26_c1 ),
    .A2(\u_multiplier/STAGE3/pp_27_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla3/_38_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_54_  (.A(\u_multiplier/STAGE3/pp_26_c1 ),
    .B(\u_multiplier/STAGE3/pp_27_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla2/cla3/_39_ ));
 OAI21_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_55_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla3/_25_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla3/_37_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/cla3/_38_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/c3 ));
 XNOR2_X2 \u_multiplier/STAGE3/Final_add/cla2/cla3/_56_  (.A(\u_multiplier/STAGE3/Final_add/cla2/c2 ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla3/_30_ ),
    .ZN(product[24]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_57_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla3/_31_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla3/_33_ ),
    .ZN(product[25]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_58_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla3/_34_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla3/_36_ ),
    .ZN(product[26]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla3/_59_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla3/_37_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla3/_39_ ),
    .ZN(product[27]));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_40_  (.A1(net75),
    .A2(net76),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla4/_25_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_41_  (.A1(\u_multiplier/STAGE3/pp_29_c ),
    .A2(\u_multiplier/s_30 ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla4/_26_ ));
 NAND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_42_  (.A1(\u_multiplier/STAGE3/pp_28_c1 ),
    .A2(\u_multiplier/STAGE3/pp_29_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla4/_27_ ));
 AND2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_43_  (.A1(\u_multiplier/STAGE3/pp_27_c1 ),
    .A2(\u_multiplier/STAGE3/pp_28_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla4/_28_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_44_  (.A1(\u_multiplier/STAGE3/pp_27_c1 ),
    .A2(\u_multiplier/STAGE3/pp_28_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla4/_29_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_45_  (.A(\u_multiplier/STAGE3/pp_27_c1 ),
    .B(\u_multiplier/STAGE3/pp_28_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla4/_30_ ));
 AOI21_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_46_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla4/_28_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla4/_29_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/c3 ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla4/_31_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_47_  (.A1(\u_multiplier/STAGE3/pp_28_c1 ),
    .A2(\u_multiplier/STAGE3/pp_29_s ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla4/_32_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_48_  (.A(\u_multiplier/STAGE3/pp_28_c1 ),
    .B(\u_multiplier/STAGE3/pp_29_s ),
    .Z(\u_multiplier/STAGE3/Final_add/cla2/cla4/_33_ ));
 OAI21_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_49_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla4/_27_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla4/_31_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/cla4/_32_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla4/_34_ ));
 OR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_50_  (.A1(\u_multiplier/STAGE3/pp_29_c ),
    .A2(\u_multiplier/s_30 ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla4/_35_ ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_51_  (.A(\u_multiplier/STAGE3/pp_29_c ),
    .B(\u_multiplier/s_30 ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla4/_36_ ));
 AOI21_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_52_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla4/_26_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla4/_34_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/cla4/_35_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla4/_37_ ));
 NOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_53_  (.A1(net77),
    .A2(net78),
    .ZN(\u_multiplier/STAGE3/Final_add/cla2/cla4/_38_ ));
 XOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_54_  (.A(net79),
    .B(net80),
    .Z(\u_multiplier/STAGE3/Final_add/cla2/cla4/_39_ ));
 OAI21_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_55_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla4/_25_ ),
    .B1(\u_multiplier/STAGE3/Final_add/cla2/cla4/_37_ ),
    .B2(\u_multiplier/STAGE3/Final_add/cla2/cla4/_38_ ),
    .ZN(\u_multiplier/STAGE3/Final_add/Cout ));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_56_  (.A(\u_multiplier/STAGE3/Final_add/cla2/c3 ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla4/_30_ ),
    .ZN(product[28]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_57_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla4/_31_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla4/_33_ ),
    .ZN(product[29]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_58_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla4/_34_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla4/_36_ ),
    .ZN(product[30]));
 XNOR2_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_59_  (.A(\u_multiplier/STAGE3/Final_add/cla2/cla4/_37_ ),
    .B(\u_multiplier/STAGE3/Final_add/cla2/cla4/_39_ ),
    .ZN(product[31]));
 INV_X1 \u_multiplier/STAGE3/Full_adder_pp_29/_12_  (.A(\u_multiplier/STAGE3/pp_28_c2 ),
    .ZN(\u_multiplier/STAGE3/Full_adder_pp_29/_08_ ));
 NAND3_X1 \u_multiplier/STAGE3/Full_adder_pp_29/_13_  (.A1(\u_multiplier/s_29 [1]),
    .A2(\u_multiplier/s_29 [0]),
    .A3(\u_multiplier/STAGE3/pp_28_c2 ),
    .ZN(\u_multiplier/STAGE3/Full_adder_pp_29/_09_ ));
 NOR2_X2 \u_multiplier/STAGE3/Full_adder_pp_29/_14_  (.A1(\u_multiplier/s_29 [1]),
    .A2(\u_multiplier/s_29 [0]),
    .ZN(\u_multiplier/STAGE3/Full_adder_pp_29/_10_ ));
 AOI21_X1 \u_multiplier/STAGE3/Full_adder_pp_29/_15_  (.A(\u_multiplier/STAGE3/pp_28_c2 ),
    .B1(\u_multiplier/s_29 [0]),
    .B2(\u_multiplier/s_29 [1]),
    .ZN(\u_multiplier/STAGE3/Full_adder_pp_29/_11_ ));
 NOR2_X2 \u_multiplier/STAGE3/Full_adder_pp_29/_16_  (.A1(\u_multiplier/STAGE3/Full_adder_pp_29/_10_ ),
    .A2(\u_multiplier/STAGE3/Full_adder_pp_29/_11_ ),
    .ZN(\u_multiplier/STAGE3/pp_29_c ));
 AOI22_X2 \u_multiplier/STAGE3/Full_adder_pp_29/_17_  (.A1(\u_multiplier/STAGE3/Full_adder_pp_29/_08_ ),
    .A2(\u_multiplier/STAGE3/Full_adder_pp_29/_10_ ),
    .B1(\u_multiplier/STAGE3/pp_29_c ),
    .B2(\u_multiplier/STAGE3/Full_adder_pp_29/_09_ ),
    .ZN(\u_multiplier/STAGE3/pp_29_s ));
 AND2_X1 \u_multiplier/STAGE3/Half_adder_pp_2/_4_  (.A1(\u_multiplier/s_2 [1]),
    .A2(\u_multiplier/s_2 [0]),
    .ZN(\u_multiplier/STAGE3/pp_2_c ));
 XOR2_X2 \u_multiplier/STAGE3/Half_adder_pp_2/_5_  (.A(\u_multiplier/s_2 [1]),
    .B(\u_multiplier/s_2 [0]),
    .Z(\u_multiplier/STAGE3/pp_2_s ));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_2_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_2_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_2_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_2_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_2_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_2_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_2_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_2_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_2_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_2_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_2_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_2_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_2_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_2_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_2_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_2_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_2_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_2_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_2_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_2_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_2_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_2_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_2_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_2_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_2_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_2_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_2_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_2_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_2_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_2_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_2_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_2_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_2_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_2_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_2_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_2_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_2_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_2_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_2_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_2_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_2_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_2_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_2_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_2_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_2_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_2_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_2_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_2_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_2_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_2_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_2_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_2_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_2_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_2_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_2_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_2_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_2_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_2_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_2_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_2_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_2_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_2_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_2_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_2_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_2_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_2_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_2_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_2_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_2_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_2_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_2_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_2_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_2_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_2_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_2_Right_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_2_Right_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_2_Right_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_2_Right_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_2_Right_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_2_Right_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_2_Right_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_2_Right_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_2_Right_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_2_Right_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_2_Right_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_2_Right_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_2_Right_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_2_Right_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_2_Right_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_2_Right_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_2_Right_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_2_Right_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_2_Right_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_2_Right_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_2_Right_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_2_Right_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_2_Right_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_2_Right_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_2_Right_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_2_Right_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_2_Right_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_2_Right_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_2_Right_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_2_Right_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_2_Right_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_1_Left_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_1_Left_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_1_Left_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_1_Left_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_1_Left_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_1_Left_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_1_Left_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_1_Left_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_1_Left_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_1_Left_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_1_Left_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_1_Left_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_1_Left_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_1_Left_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_1_Left_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_1_Left_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_1_Left_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_1_Left_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_1_Left_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_1_Left_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_1_Left_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_1_Left_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_1_Left_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_1_Left_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_1_Left_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_1_Left_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_1_Left_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_1_Left_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_1_Left_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_1_Left_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_1_Left_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_1_Left_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_1_Left_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_1_Left_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_1_Left_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_1_Left_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_1_Left_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_1_Left_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_1_Left_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_1_Left_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_1_Left_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_1_Left_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_1_Left_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_1_Left_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_1_Left_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_1_Left_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_1_Left_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_1_Left_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_1_Left_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_1_Left_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_1_Left_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_1_Left_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_1_Left_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_1_Left_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_1_Left_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_1_Left_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_1_Left_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_1_Left_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_1_Left_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_1_Left_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_1_Left_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_1_Left_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_1_Left_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_1_Left_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_1_Left_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_1_Left_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_1_Left_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_1_Left_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_1_Left_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_1_Left_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_1_Left_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_1_Left_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_1_Left_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_1_Left_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_1_Left_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_1_Left_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_1_Left_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_1_Left_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_1_Left_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_1_Left_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_1_Left_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_1_Left_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_1_Left_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_1_Left_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_1_Left_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_1_Left_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_1_Left_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_1_Left_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_1_Left_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_1_Left_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_1_Left_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_1_Left_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_1_Left_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_1_Left_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_1_Left_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_1_Left_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_1_Left_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_1_Left_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_1_Left_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_1_Left_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_1_Left_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_1_Left_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_1_Left_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_1_Left_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Left_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Left_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Left_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Left_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Left_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Left_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Left_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Left_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Left_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Left_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Left_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Left_265 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Left_266 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Left_267 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Left_268 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Left_269 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Left_270 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Left_271 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Left_272 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Left_273 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Left_274 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_1_Left_275 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_2_Left_276 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_2_Left_277 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_2_Left_278 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_2_Left_279 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_2_Left_280 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_2_Left_281 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_2_Left_282 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_2_Left_283 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_2_Left_284 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_2_Left_285 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_2_Left_286 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_2_Left_287 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_2_Left_288 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_2_Left_289 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_2_Left_290 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_2_Left_291 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_2_Left_292 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_2_Left_293 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_2_Left_294 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_2_Left_295 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_2_Left_296 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_2_Left_297 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_2_Left_298 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_2_Left_299 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_2_Left_300 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_2_Left_301 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_2_Left_302 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_2_Left_303 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_2_Left_304 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_2_Left_305 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_2_Left_306 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_2_Left_307 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_2_Left_308 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_2_Left_309 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_2_Left_310 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_2_Left_311 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_2_Left_312 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_2_Left_313 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_2_Left_314 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_2_Left_315 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_2_Left_316 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_2_Left_317 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_2_Left_318 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_2_Left_319 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_2_Left_320 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_2_Left_321 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_2_Left_322 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_2_Left_323 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_2_Left_324 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_2_Left_325 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_2_Left_326 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_2_Left_327 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_2_Left_328 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_2_Left_329 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_2_Left_330 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_2_Left_331 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_2_Left_332 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_2_Left_333 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_2_Left_334 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_2_Left_335 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_2_Left_336 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_2_Left_337 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_2_Left_338 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_2_Left_339 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_2_Left_340 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_2_Left_341 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_2_Left_342 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_2_Left_343 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_2_Left_344 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_2_Left_345 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_2_Left_346 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_2_Left_347 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_2_Left_348 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_2_Left_349 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_2_Left_350 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_2_Left_351 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_2_Left_352 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_2_Left_353 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_2_Left_354 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_2_Left_355 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_2_Left_356 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_2_Left_357 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_2_Left_358 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_2_Left_359 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_2_Left_360 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_2_Left_361 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_2_Left_362 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_2_Left_363 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_2_Left_364 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_2_Left_365 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_2_Left_366 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_2_Left_367 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_2_Left_368 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_2_Left_369 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_2_Left_370 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_2_Left_371 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_2_Left_372 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_2_Left_373 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_2_Left_374 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_2_Left_375 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_2_Left_376 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_2_Left_377 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_2_Left_378 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_2_Left_379 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_2_Left_380 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_1_Right_381 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_1_Right_382 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_1_Right_383 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_1_Right_384 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_1_Right_385 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_1_Right_386 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_1_Right_387 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_1_Right_388 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_1_Right_389 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_1_Right_390 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_1_Right_391 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_1_Right_392 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_1_Right_393 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_1_Right_394 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_1_Right_395 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_1_Right_396 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_1_Right_397 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_1_Right_398 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_1_Right_399 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_1_Right_400 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_1_Right_401 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_1_Right_402 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_1_Right_403 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_1_Right_404 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_1_Right_405 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_1_Right_406 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_1_Right_407 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_1_Right_408 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_1_Right_409 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_1_Right_410 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_1_Right_411 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_1_Right_412 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_1_Right_413 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_1_Right_414 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_1_Right_415 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_1_Right_416 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_1_Right_417 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_1_Right_418 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_1_Right_419 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_1_Right_420 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_1_Right_421 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_1_Right_422 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_1_Right_423 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_1_Right_424 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_1_Right_425 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_1_Right_426 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_1_Right_427 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_1_Right_428 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_1_Right_429 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_1_Right_430 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_1_Right_431 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_1_Right_432 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_1_Right_433 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_1_Right_434 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_1_Right_435 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_1_Right_436 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_1_Right_437 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_1_Right_438 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_1_Right_439 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_1_Right_440 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_1_Right_441 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_1_Right_442 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_1_Right_443 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_1_Right_444 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_1_Right_445 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_1_Right_446 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_1_Right_447 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_1_Right_448 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_1_Right_449 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_1_Right_450 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_1_Right_451 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_1_Right_452 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_1_Right_453 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_1_Right_454 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_1_Right_455 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_1_Right_456 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_1_Right_457 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_1_Right_458 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_1_Right_459 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_1_Right_460 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_1_Right_461 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_1_Right_462 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_1_Right_463 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_1_Right_464 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_1_Right_465 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_1_Right_466 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_1_Right_467 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_1_Right_468 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_1_Right_469 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_1_Right_470 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_1_Right_471 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_1_Right_472 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_1_Right_473 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_1_Right_474 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_1_Right_475 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_1_Right_476 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_1_Right_477 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_1_Right_478 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_1_Right_479 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_1_Right_480 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_1_Right_481 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_1_Right_482 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_1_Right_483 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_1_Right_484 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_1_Right_485 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_486 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_487 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_488 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_489 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_490 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_491 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_492 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_117_493 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_494 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_495 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_496 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_497 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_498 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_499 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_500 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_501 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_502 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_503 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_137_504 ();
 LOGIC0_X1 \u_multiplier/STAGE2/E_4_2_pp_5/_18__64  (.Z(net64));
 LOGIC0_X1 \u_multiplier/STAGE3/E_4_2_pp_3/_18__68  (.Z(net68));
 CLKBUF_X1 hold81 (.A(net143),
    .Z(net81));
 BUF_X1 input1 (.A(data_in[0]),
    .Z(net1));
 BUF_X1 input2 (.A(data_in[10]),
    .Z(net2));
 BUF_X1 input3 (.A(data_in[11]),
    .Z(net3));
 CLKBUF_X2 input4 (.A(data_in[12]),
    .Z(net4));
 BUF_X1 input5 (.A(data_in[13]),
    .Z(net5));
 BUF_X1 input6 (.A(data_in[14]),
    .Z(net6));
 BUF_X2 input7 (.A(data_in[15]),
    .Z(net7));
 CLKBUF_X2 input8 (.A(data_in[1]),
    .Z(net8));
 BUF_X1 input9 (.A(data_in[2]),
    .Z(net9));
 BUF_X2 input10 (.A(data_in[3]),
    .Z(net10));
 BUF_X1 input11 (.A(data_in[4]),
    .Z(net11));
 BUF_X1 input12 (.A(data_in[5]),
    .Z(net12));
 BUF_X1 input13 (.A(data_in[6]),
    .Z(net13));
 BUF_X1 input14 (.A(data_in[7]),
    .Z(net14));
 CLKBUF_X2 input15 (.A(data_in[8]),
    .Z(net15));
 BUF_X1 input16 (.A(data_in[9]),
    .Z(net16));
 CLKBUF_X3 input17 (.A(init_enable),
    .Z(net17));
 BUF_X2 input18 (.A(pe_ce),
    .Z(net18));
 BUF_X8 input19 (.A(rst_n),
    .Z(net19));
 BUF_X1 output20 (.A(net20),
    .Z(curr_state[1]));
 BUF_X1 output21 (.A(net21),
    .Z(data_out[0]));
 BUF_X1 output22 (.A(net22),
    .Z(data_out[10]));
 BUF_X1 output23 (.A(net23),
    .Z(data_out[11]));
 BUF_X1 output24 (.A(net24),
    .Z(data_out[12]));
 BUF_X1 output25 (.A(net25),
    .Z(data_out[13]));
 BUF_X1 output26 (.A(net26),
    .Z(data_out[14]));
 BUF_X1 output27 (.A(net27),
    .Z(data_out[15]));
 BUF_X1 output28 (.A(net28),
    .Z(data_out[16]));
 BUF_X1 output29 (.A(net29),
    .Z(data_out[17]));
 BUF_X1 output30 (.A(net30),
    .Z(data_out[18]));
 BUF_X1 output31 (.A(net31),
    .Z(data_out[19]));
 BUF_X1 output32 (.A(net32),
    .Z(data_out[1]));
 BUF_X1 output33 (.A(net33),
    .Z(data_out[20]));
 BUF_X1 output34 (.A(net34),
    .Z(data_out[21]));
 BUF_X1 output35 (.A(net35),
    .Z(data_out[22]));
 BUF_X1 output36 (.A(net36),
    .Z(data_out[23]));
 BUF_X1 output37 (.A(net37),
    .Z(data_out[24]));
 BUF_X1 output38 (.A(net38),
    .Z(data_out[25]));
 BUF_X1 output39 (.A(net39),
    .Z(data_out[26]));
 BUF_X1 output40 (.A(net40),
    .Z(data_out[27]));
 BUF_X1 output41 (.A(net41),
    .Z(data_out[28]));
 BUF_X1 output42 (.A(net42),
    .Z(data_out[29]));
 BUF_X1 output43 (.A(net43),
    .Z(data_out[2]));
 BUF_X1 output44 (.A(net44),
    .Z(data_out[30]));
 BUF_X1 output45 (.A(net45),
    .Z(data_out[31]));
 BUF_X1 output46 (.A(net46),
    .Z(data_out[3]));
 BUF_X1 output47 (.A(net47),
    .Z(data_out[4]));
 BUF_X1 output48 (.A(net48),
    .Z(data_out[5]));
 BUF_X1 output49 (.A(net49),
    .Z(data_out[6]));
 BUF_X1 output50 (.A(net50),
    .Z(data_out[7]));
 BUF_X1 output51 (.A(net51),
    .Z(data_out[8]));
 BUF_X1 output52 (.A(net52),
    .Z(data_out[9]));
 BUF_X1 output53 (.A(net53),
    .Z(valid_reg_out));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_11_2/_18__54  (.Z(net54));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_11_2/_25__55  (.Z(net55));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_13_3/_18__56  (.Z(net56));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_13_3/_25__57  (.Z(net57));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_15_4/_18__58  (.Z(net58));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_15_4/_25__59  (.Z(net59));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_16_4/_18__60  (.Z(net60));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_16_4/_25__61  (.Z(net61));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_9/_18__62  (.Z(net62));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_9/_25__63  (.Z(net63));
 LOGIC0_X1 \u_multiplier/STAGE2/E_4_2_pp_5/_25__65  (.Z(net65));
 LOGIC0_X1 \u_multiplier/STAGE2/E_4_2_pp_7_2/_18__66  (.Z(net66));
 LOGIC0_X1 \u_multiplier/STAGE2/E_4_2_pp_7_2/_25__67  (.Z(net67));
 LOGIC0_X1 \u_multiplier/STAGE3/E_4_2_pp_3/_25__69  (.Z(net69));
 LOGIC0_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_43__70  (.Z(net70));
 LOGIC0_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_44__71  (.Z(net71));
 LOGIC0_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_45__72  (.Z(net72));
 LOGIC0_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_46__73  (.Z(net73));
 LOGIC0_X1 \u_multiplier/STAGE3/Final_add/cla1/cla1/_56__74  (.Z(net74));
 LOGIC0_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_40__75  (.Z(net75));
 LOGIC0_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_40__76  (.Z(net76));
 LOGIC0_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_53__77  (.Z(net77));
 LOGIC0_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_53__78  (.Z(net78));
 LOGIC0_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_54__79  (.Z(net79));
 LOGIC0_X1 \u_multiplier/STAGE3/Final_add/cla2/cla4/_54__80  (.Z(net80));
 CLKBUF_X1 hold82 (.A(_173_),
    .Z(net82));
 CLKBUF_X1 hold83 (.A(net146),
    .Z(net83));
 CLKBUF_X1 hold84 (.A(_192_),
    .Z(net84));
 CLKBUF_X1 hold85 (.A(net100),
    .Z(net85));
 CLKBUF_X1 hold86 (.A(net97),
    .Z(net86));
 CLKBUF_X1 hold87 (.A(net108),
    .Z(net87));
 CLKBUF_X1 hold88 (.A(net111),
    .Z(net88));
 CLKBUF_X1 hold89 (.A(net117),
    .Z(net89));
 CLKBUF_X1 hold90 (.A(net128),
    .Z(net90));
 CLKBUF_X1 hold91 (.A(net123),
    .Z(net91));
 CLKBUF_X1 hold92 (.A(net120),
    .Z(net92));
 CLKBUF_X1 hold93 (.A(net133),
    .Z(net93));
 CLKBUF_X1 hold94 (.A(net135),
    .Z(net94));
 CLKBUF_X1 hold95 (.A(net142),
    .Z(net95));
 CLKBUF_X1 hold96 (.A(net130),
    .Z(net96));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_2_0_0_clk));
 CLKBUF_X3 clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_2_1_0_clk));
 CLKBUF_X3 clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .Z(clknet_2_2_0_clk));
 CLKBUF_X3 clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .Z(clknet_2_3_0_clk));
 CLKBUF_X3 clkbuf_3_0_0_clk (.A(clknet_2_0_0_clk),
    .Z(clknet_3_0_0_clk));
 CLKBUF_X3 clkbuf_3_1_0_clk (.A(clknet_2_0_0_clk),
    .Z(clknet_3_1_0_clk));
 CLKBUF_X3 clkbuf_3_2_0_clk (.A(clknet_2_1_0_clk),
    .Z(clknet_3_2_0_clk));
 CLKBUF_X3 clkbuf_3_3_0_clk (.A(clknet_2_1_0_clk),
    .Z(clknet_3_3_0_clk));
 CLKBUF_X3 clkbuf_3_4_0_clk (.A(clknet_2_2_0_clk),
    .Z(clknet_3_4_0_clk));
 CLKBUF_X3 clkbuf_3_5_0_clk (.A(clknet_2_2_0_clk),
    .Z(clknet_3_5_0_clk));
 CLKBUF_X3 clkbuf_3_6_0_clk (.A(clknet_2_3_0_clk),
    .Z(clknet_3_6_0_clk));
 CLKBUF_X3 clkbuf_3_7_0_clk (.A(clknet_2_3_0_clk),
    .Z(clknet_3_7_0_clk));
 INV_X2 clkload0 (.A(clknet_3_0_0_clk));
 INV_X2 clkload1 (.A(clknet_3_2_0_clk));
 INV_X1 clkload2 (.A(clknet_3_4_0_clk));
 INV_X2 clkload3 (.A(clknet_3_6_0_clk));
 CLKBUF_X1 hold1 (.A(_399_),
    .Z(net97));
 CLKBUF_X1 hold2 (.A(net86),
    .Z(net98));
 CLKBUF_X1 hold3 (.A(_117_),
    .Z(net99));
 CLKBUF_X1 hold4 (.A(_400_),
    .Z(net100));
 CLKBUF_X1 hold5 (.A(net85),
    .Z(net101));
 CLKBUF_X1 hold6 (.A(_118_),
    .Z(net102));
 CLKBUF_X1 hold7 (.A(_402_),
    .Z(net103));
 CLKBUF_X1 hold8 (.A(_278_),
    .Z(net104));
 CLKBUF_X1 hold9 (.A(_403_),
    .Z(net105));
 CLKBUF_X1 hold10 (.A(_280_),
    .Z(net106));
 CLKBUF_X1 hold11 (.A(net152),
    .Z(net107));
 CLKBUF_X1 hold12 (.A(_406_),
    .Z(net108));
 CLKBUF_X1 hold13 (.A(net87),
    .Z(net109));
 CLKBUF_X1 hold14 (.A(_172_),
    .Z(net110));
 CLKBUF_X1 hold15 (.A(_405_),
    .Z(net111));
 CLKBUF_X1 hold16 (.A(net88),
    .Z(net112));
 CLKBUF_X1 hold17 (.A(_171_),
    .Z(net113));
 CLKBUF_X1 hold18 (.A(curr_state[0]),
    .Z(net114));
 CLKBUF_X1 hold19 (.A(_251_),
    .Z(net115));
 CLKBUF_X1 hold20 (.A(_194_),
    .Z(net116));
 CLKBUF_X1 hold21 (.A(_404_),
    .Z(net117));
 CLKBUF_X1 hold22 (.A(net89),
    .Z(net118));
 CLKBUF_X1 hold23 (.A(_170_),
    .Z(net119));
 CLKBUF_X1 hold24 (.A(_401_),
    .Z(net120));
 CLKBUF_X1 hold25 (.A(net92),
    .Z(net121));
 CLKBUF_X1 hold26 (.A(net153),
    .Z(net122));
 CLKBUF_X1 hold27 (.A(addr_ptr[1]),
    .Z(net123));
 CLKBUF_X1 hold28 (.A(net91),
    .Z(net124));
 CLKBUF_X1 hold29 (.A(data_in_reg[1]),
    .Z(net125));
 CLKBUF_X1 hold30 (.A(data_in_reg[15]),
    .Z(net126));
 CLKBUF_X1 hold31 (.A(data_in_reg[14]),
    .Z(net127));
 CLKBUF_X1 hold32 (.A(addr_ptr[4]),
    .Z(net128));
 CLKBUF_X1 hold33 (.A(net90),
    .Z(net129));
 CLKBUF_X1 hold34 (.A(_408_),
    .Z(net130));
 CLKBUF_X1 hold35 (.A(net96),
    .Z(net131));
 CLKBUF_X1 hold36 (.A(_174_),
    .Z(net132));
 CLKBUF_X1 hold37 (.A(addr_ptr[2]),
    .Z(net133));
 CLKBUF_X1 hold38 (.A(net93),
    .Z(net134));
 CLKBUF_X1 hold39 (.A(addr_ptr[3]),
    .Z(net135));
 CLKBUF_X1 hold40 (.A(net94),
    .Z(net136));
 CLKBUF_X1 hold41 (.A(data_in_reg[12]),
    .Z(net137));
 CLKBUF_X1 hold42 (.A(data_in_reg[13]),
    .Z(net138));
 CLKBUF_X1 hold43 (.A(data_in_reg[11]),
    .Z(net139));
 CLKBUF_X1 hold44 (.A(data_in_reg[6]),
    .Z(net140));
 CLKBUF_X1 hold45 (.A(data_in_reg[7]),
    .Z(net141));
 CLKBUF_X1 hold46 (.A(addr_ptr[0]),
    .Z(net142));
 CLKBUF_X1 hold47 (.A(_407_),
    .Z(net143));
 CLKBUF_X1 hold48 (.A(data_in_reg[2]),
    .Z(net144));
 CLKBUF_X1 hold49 (.A(data_in_reg[3]),
    .Z(net145));
 CLKBUF_X1 hold50 (.A(_331_),
    .Z(net146));
 CLKBUF_X1 hold51 (.A(data_in_reg[4]),
    .Z(net147));
 CLKBUF_X1 hold52 (.A(data_in_reg[0]),
    .Z(net148));
 CLKBUF_X1 hold53 (.A(data_in_reg[8]),
    .Z(net149));
 CLKBUF_X1 hold54 (.A(data_in_reg[9]),
    .Z(net150));
 CLKBUF_X1 hold55 (.A(curr_state[2]),
    .Z(net151));
 CLKBUF_X1 hold56 (.A(data_in_reg[5]),
    .Z(net152));
 CLKBUF_X1 hold57 (.A(data_in_reg[10]),
    .Z(net153));
 FILLCELL_X4 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_8 ();
 FILLCELL_X16 FILLER_0_40 ();
 FILLCELL_X32 FILLER_0_59 ();
 FILLCELL_X32 FILLER_0_91 ();
 FILLCELL_X8 FILLER_0_123 ();
 FILLCELL_X2 FILLER_0_131 ();
 FILLCELL_X32 FILLER_0_136 ();
 FILLCELL_X32 FILLER_0_168 ();
 FILLCELL_X8 FILLER_0_200 ();
 FILLCELL_X4 FILLER_0_208 ();
 FILLCELL_X2 FILLER_0_212 ();
 FILLCELL_X1 FILLER_0_214 ();
 FILLCELL_X32 FILLER_0_218 ();
 FILLCELL_X32 FILLER_0_250 ();
 FILLCELL_X8 FILLER_0_282 ();
 FILLCELL_X2 FILLER_0_290 ();
 FILLCELL_X32 FILLER_0_295 ();
 FILLCELL_X32 FILLER_0_327 ();
 FILLCELL_X8 FILLER_0_359 ();
 FILLCELL_X4 FILLER_0_367 ();
 FILLCELL_X2 FILLER_0_371 ();
 FILLCELL_X1 FILLER_0_373 ();
 FILLCELL_X32 FILLER_0_377 ();
 FILLCELL_X32 FILLER_0_409 ();
 FILLCELL_X8 FILLER_0_441 ();
 FILLCELL_X2 FILLER_0_449 ();
 FILLCELL_X32 FILLER_0_454 ();
 FILLCELL_X32 FILLER_0_486 ();
 FILLCELL_X8 FILLER_0_518 ();
 FILLCELL_X2 FILLER_0_526 ();
 FILLCELL_X32 FILLER_0_531 ();
 FILLCELL_X32 FILLER_0_563 ();
 FILLCELL_X8 FILLER_0_595 ();
 FILLCELL_X4 FILLER_0_603 ();
 FILLCELL_X2 FILLER_0_607 ();
 FILLCELL_X1 FILLER_0_609 ();
 FILLCELL_X16 FILLER_0_613 ();
 FILLCELL_X2 FILLER_0_629 ();
 FILLCELL_X32 FILLER_0_632 ();
 FILLCELL_X16 FILLER_0_664 ();
 FILLCELL_X4 FILLER_0_680 ();
 FILLCELL_X2 FILLER_0_684 ();
 FILLCELL_X1 FILLER_0_686 ();
 FILLCELL_X32 FILLER_0_692 ();
 FILLCELL_X16 FILLER_0_724 ();
 FILLCELL_X2 FILLER_0_740 ();
 FILLCELL_X1 FILLER_0_742 ();
 FILLCELL_X16 FILLER_0_746 ();
 FILLCELL_X4 FILLER_0_762 ();
 FILLCELL_X2 FILLER_0_766 ();
 FILLCELL_X1 FILLER_0_768 ();
 FILLCELL_X8 FILLER_0_772 ();
 FILLCELL_X4 FILLER_0_780 ();
 FILLCELL_X2 FILLER_0_784 ();
 FILLCELL_X1 FILLER_0_786 ();
 FILLCELL_X4 FILLER_0_791 ();
 FILLCELL_X1 FILLER_0_795 ();
 FILLCELL_X4 FILLER_0_802 ();
 FILLCELL_X4 FILLER_0_809 ();
 FILLCELL_X2 FILLER_0_813 ();
 FILLCELL_X8 FILLER_0_817 ();
 FILLCELL_X4 FILLER_0_825 ();
 FILLCELL_X4 FILLER_0_833 ();
 FILLCELL_X4 FILLER_0_841 ();
 FILLCELL_X4 FILLER_0_848 ();
 FILLCELL_X4 FILLER_0_855 ();
 FILLCELL_X32 FILLER_0_862 ();
 FILLCELL_X8 FILLER_0_894 ();
 FILLCELL_X8 FILLER_0_912 ();
 FILLCELL_X4 FILLER_0_923 ();
 FILLCELL_X4 FILLER_0_931 ();
 FILLCELL_X2 FILLER_0_935 ();
 FILLCELL_X1 FILLER_0_937 ();
 FILLCELL_X4 FILLER_0_944 ();
 FILLCELL_X4 FILLER_0_954 ();
 FILLCELL_X4 FILLER_0_961 ();
 FILLCELL_X4 FILLER_0_967 ();
 FILLCELL_X1 FILLER_0_971 ();
 FILLCELL_X16 FILLER_0_975 ();
 FILLCELL_X4 FILLER_0_991 ();
 FILLCELL_X1 FILLER_0_995 ();
 FILLCELL_X4 FILLER_0_1000 ();
 FILLCELL_X1 FILLER_0_1004 ();
 FILLCELL_X16 FILLER_0_1008 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X32 FILLER_1_257 ();
 FILLCELL_X32 FILLER_1_289 ();
 FILLCELL_X32 FILLER_1_321 ();
 FILLCELL_X32 FILLER_1_353 ();
 FILLCELL_X32 FILLER_1_385 ();
 FILLCELL_X32 FILLER_1_417 ();
 FILLCELL_X32 FILLER_1_449 ();
 FILLCELL_X32 FILLER_1_481 ();
 FILLCELL_X32 FILLER_1_513 ();
 FILLCELL_X32 FILLER_1_545 ();
 FILLCELL_X32 FILLER_1_577 ();
 FILLCELL_X32 FILLER_1_609 ();
 FILLCELL_X32 FILLER_1_641 ();
 FILLCELL_X16 FILLER_1_673 ();
 FILLCELL_X2 FILLER_1_689 ();
 FILLCELL_X4 FILLER_1_693 ();
 FILLCELL_X4 FILLER_1_707 ();
 FILLCELL_X8 FILLER_1_714 ();
 FILLCELL_X4 FILLER_1_722 ();
 FILLCELL_X4 FILLER_1_735 ();
 FILLCELL_X4 FILLER_1_742 ();
 FILLCELL_X4 FILLER_1_755 ();
 FILLCELL_X4 FILLER_1_761 ();
 FILLCELL_X2 FILLER_1_765 ();
 FILLCELL_X1 FILLER_1_767 ();
 FILLCELL_X4 FILLER_1_771 ();
 FILLCELL_X8 FILLER_1_794 ();
 FILLCELL_X1 FILLER_1_802 ();
 FILLCELL_X8 FILLER_1_813 ();
 FILLCELL_X8 FILLER_1_827 ();
 FILLCELL_X4 FILLER_1_845 ();
 FILLCELL_X2 FILLER_1_849 ();
 FILLCELL_X1 FILLER_1_851 ();
 FILLCELL_X4 FILLER_1_856 ();
 FILLCELL_X4 FILLER_1_879 ();
 FILLCELL_X4 FILLER_1_902 ();
 FILLCELL_X1 FILLER_1_906 ();
 FILLCELL_X8 FILLER_1_909 ();
 FILLCELL_X8 FILLER_1_936 ();
 FILLCELL_X4 FILLER_1_951 ();
 FILLCELL_X4 FILLER_1_965 ();
 FILLCELL_X1 FILLER_1_969 ();
 FILLCELL_X8 FILLER_1_980 ();
 FILLCELL_X2 FILLER_1_988 ();
 FILLCELL_X4 FILLER_1_994 ();
 FILLCELL_X1 FILLER_1_998 ();
 FILLCELL_X4 FILLER_1_1018 ();
 FILLCELL_X2 FILLER_1_1022 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X32 FILLER_2_289 ();
 FILLCELL_X32 FILLER_2_321 ();
 FILLCELL_X32 FILLER_2_353 ();
 FILLCELL_X32 FILLER_2_385 ();
 FILLCELL_X32 FILLER_2_417 ();
 FILLCELL_X32 FILLER_2_449 ();
 FILLCELL_X32 FILLER_2_481 ();
 FILLCELL_X32 FILLER_2_513 ();
 FILLCELL_X32 FILLER_2_545 ();
 FILLCELL_X32 FILLER_2_577 ();
 FILLCELL_X16 FILLER_2_609 ();
 FILLCELL_X4 FILLER_2_625 ();
 FILLCELL_X2 FILLER_2_629 ();
 FILLCELL_X16 FILLER_2_632 ();
 FILLCELL_X8 FILLER_2_648 ();
 FILLCELL_X4 FILLER_2_666 ();
 FILLCELL_X16 FILLER_2_673 ();
 FILLCELL_X2 FILLER_2_689 ();
 FILLCELL_X1 FILLER_2_691 ();
 FILLCELL_X4 FILLER_2_695 ();
 FILLCELL_X4 FILLER_2_709 ();
 FILLCELL_X4 FILLER_2_720 ();
 FILLCELL_X8 FILLER_2_727 ();
 FILLCELL_X4 FILLER_2_735 ();
 FILLCELL_X1 FILLER_2_739 ();
 FILLCELL_X4 FILLER_2_743 ();
 FILLCELL_X4 FILLER_2_757 ();
 FILLCELL_X1 FILLER_2_761 ();
 FILLCELL_X4 FILLER_2_772 ();
 FILLCELL_X4 FILLER_2_782 ();
 FILLCELL_X4 FILLER_2_788 ();
 FILLCELL_X4 FILLER_2_798 ();
 FILLCELL_X4 FILLER_2_809 ();
 FILLCELL_X1 FILLER_2_813 ();
 FILLCELL_X8 FILLER_2_820 ();
 FILLCELL_X1 FILLER_2_828 ();
 FILLCELL_X4 FILLER_2_836 ();
 FILLCELL_X2 FILLER_2_840 ();
 FILLCELL_X4 FILLER_2_851 ();
 FILLCELL_X1 FILLER_2_855 ();
 FILLCELL_X4 FILLER_2_875 ();
 FILLCELL_X4 FILLER_2_883 ();
 FILLCELL_X8 FILLER_2_889 ();
 FILLCELL_X4 FILLER_2_897 ();
 FILLCELL_X2 FILLER_2_901 ();
 FILLCELL_X8 FILLER_2_906 ();
 FILLCELL_X2 FILLER_2_914 ();
 FILLCELL_X1 FILLER_2_916 ();
 FILLCELL_X4 FILLER_2_924 ();
 FILLCELL_X1 FILLER_2_928 ();
 FILLCELL_X4 FILLER_2_938 ();
 FILLCELL_X4 FILLER_2_945 ();
 FILLCELL_X16 FILLER_2_952 ();
 FILLCELL_X2 FILLER_2_968 ();
 FILLCELL_X1 FILLER_2_970 ();
 FILLCELL_X8 FILLER_2_975 ();
 FILLCELL_X2 FILLER_2_983 ();
 FILLCELL_X1 FILLER_2_985 ();
 FILLCELL_X4 FILLER_2_992 ();
 FILLCELL_X4 FILLER_2_1002 ();
 FILLCELL_X4 FILLER_2_1010 ();
 FILLCELL_X2 FILLER_2_1014 ();
 FILLCELL_X1 FILLER_2_1016 ();
 FILLCELL_X4 FILLER_2_1020 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X32 FILLER_3_289 ();
 FILLCELL_X32 FILLER_3_321 ();
 FILLCELL_X32 FILLER_3_353 ();
 FILLCELL_X32 FILLER_3_385 ();
 FILLCELL_X32 FILLER_3_417 ();
 FILLCELL_X32 FILLER_3_449 ();
 FILLCELL_X32 FILLER_3_481 ();
 FILLCELL_X32 FILLER_3_513 ();
 FILLCELL_X32 FILLER_3_545 ();
 FILLCELL_X32 FILLER_3_577 ();
 FILLCELL_X32 FILLER_3_609 ();
 FILLCELL_X2 FILLER_3_641 ();
 FILLCELL_X4 FILLER_3_646 ();
 FILLCELL_X4 FILLER_3_660 ();
 FILLCELL_X1 FILLER_3_664 ();
 FILLCELL_X4 FILLER_3_674 ();
 FILLCELL_X4 FILLER_3_681 ();
 FILLCELL_X4 FILLER_3_688 ();
 FILLCELL_X8 FILLER_3_695 ();
 FILLCELL_X1 FILLER_3_703 ();
 FILLCELL_X4 FILLER_3_713 ();
 FILLCELL_X4 FILLER_3_727 ();
 FILLCELL_X8 FILLER_3_738 ();
 FILLCELL_X1 FILLER_3_746 ();
 FILLCELL_X4 FILLER_3_750 ();
 FILLCELL_X4 FILLER_3_757 ();
 FILLCELL_X2 FILLER_3_761 ();
 FILLCELL_X1 FILLER_3_763 ();
 FILLCELL_X4 FILLER_3_771 ();
 FILLCELL_X4 FILLER_3_777 ();
 FILLCELL_X2 FILLER_3_781 ();
 FILLCELL_X4 FILLER_3_787 ();
 FILLCELL_X4 FILLER_3_797 ();
 FILLCELL_X4 FILLER_3_808 ();
 FILLCELL_X4 FILLER_3_822 ();
 FILLCELL_X4 FILLER_3_830 ();
 FILLCELL_X8 FILLER_3_837 ();
 FILLCELL_X4 FILLER_3_845 ();
 FILLCELL_X4 FILLER_3_853 ();
 FILLCELL_X16 FILLER_3_860 ();
 FILLCELL_X1 FILLER_3_876 ();
 FILLCELL_X4 FILLER_3_887 ();
 FILLCELL_X4 FILLER_3_898 ();
 FILLCELL_X4 FILLER_3_911 ();
 FILLCELL_X2 FILLER_3_915 ();
 FILLCELL_X4 FILLER_3_927 ();
 FILLCELL_X1 FILLER_3_931 ();
 FILLCELL_X8 FILLER_3_935 ();
 FILLCELL_X4 FILLER_3_953 ();
 FILLCELL_X2 FILLER_3_957 ();
 FILLCELL_X8 FILLER_3_966 ();
 FILLCELL_X4 FILLER_3_974 ();
 FILLCELL_X4 FILLER_3_987 ();
 FILLCELL_X1 FILLER_3_991 ();
 FILLCELL_X16 FILLER_3_999 ();
 FILLCELL_X8 FILLER_3_1015 ();
 FILLCELL_X1 FILLER_3_1023 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X32 FILLER_4_289 ();
 FILLCELL_X32 FILLER_4_321 ();
 FILLCELL_X32 FILLER_4_353 ();
 FILLCELL_X32 FILLER_4_385 ();
 FILLCELL_X32 FILLER_4_417 ();
 FILLCELL_X32 FILLER_4_449 ();
 FILLCELL_X32 FILLER_4_481 ();
 FILLCELL_X32 FILLER_4_513 ();
 FILLCELL_X32 FILLER_4_545 ();
 FILLCELL_X32 FILLER_4_577 ();
 FILLCELL_X8 FILLER_4_609 ();
 FILLCELL_X8 FILLER_4_619 ();
 FILLCELL_X4 FILLER_4_627 ();
 FILLCELL_X8 FILLER_4_632 ();
 FILLCELL_X4 FILLER_4_640 ();
 FILLCELL_X1 FILLER_4_644 ();
 FILLCELL_X8 FILLER_4_648 ();
 FILLCELL_X2 FILLER_4_656 ();
 FILLCELL_X4 FILLER_4_665 ();
 FILLCELL_X4 FILLER_4_671 ();
 FILLCELL_X2 FILLER_4_675 ();
 FILLCELL_X8 FILLER_4_686 ();
 FILLCELL_X4 FILLER_4_703 ();
 FILLCELL_X4 FILLER_4_716 ();
 FILLCELL_X4 FILLER_4_723 ();
 FILLCELL_X4 FILLER_4_737 ();
 FILLCELL_X2 FILLER_4_741 ();
 FILLCELL_X8 FILLER_4_752 ();
 FILLCELL_X1 FILLER_4_760 ();
 FILLCELL_X4 FILLER_4_771 ();
 FILLCELL_X4 FILLER_4_785 ();
 FILLCELL_X2 FILLER_4_789 ();
 FILLCELL_X1 FILLER_4_791 ();
 FILLCELL_X4 FILLER_4_796 ();
 FILLCELL_X16 FILLER_4_803 ();
 FILLCELL_X1 FILLER_4_819 ();
 FILLCELL_X4 FILLER_4_827 ();
 FILLCELL_X8 FILLER_4_840 ();
 FILLCELL_X4 FILLER_4_848 ();
 FILLCELL_X2 FILLER_4_852 ();
 FILLCELL_X16 FILLER_4_864 ();
 FILLCELL_X8 FILLER_4_880 ();
 FILLCELL_X4 FILLER_4_888 ();
 FILLCELL_X1 FILLER_4_892 ();
 FILLCELL_X4 FILLER_4_903 ();
 FILLCELL_X8 FILLER_4_910 ();
 FILLCELL_X4 FILLER_4_918 ();
 FILLCELL_X16 FILLER_4_925 ();
 FILLCELL_X2 FILLER_4_941 ();
 FILLCELL_X1 FILLER_4_943 ();
 FILLCELL_X4 FILLER_4_946 ();
 FILLCELL_X4 FILLER_4_953 ();
 FILLCELL_X4 FILLER_4_967 ();
 FILLCELL_X1 FILLER_4_971 ();
 FILLCELL_X4 FILLER_4_981 ();
 FILLCELL_X2 FILLER_4_985 ();
 FILLCELL_X1 FILLER_4_987 ();
 FILLCELL_X32 FILLER_4_991 ();
 FILLCELL_X1 FILLER_4_1023 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X4 FILLER_5_161 ();
 FILLCELL_X2 FILLER_5_165 ();
 FILLCELL_X1 FILLER_5_167 ();
 FILLCELL_X32 FILLER_5_172 ();
 FILLCELL_X32 FILLER_5_204 ();
 FILLCELL_X32 FILLER_5_236 ();
 FILLCELL_X32 FILLER_5_268 ();
 FILLCELL_X32 FILLER_5_300 ();
 FILLCELL_X32 FILLER_5_332 ();
 FILLCELL_X32 FILLER_5_364 ();
 FILLCELL_X32 FILLER_5_396 ();
 FILLCELL_X32 FILLER_5_428 ();
 FILLCELL_X32 FILLER_5_460 ();
 FILLCELL_X32 FILLER_5_492 ();
 FILLCELL_X32 FILLER_5_524 ();
 FILLCELL_X32 FILLER_5_556 ();
 FILLCELL_X16 FILLER_5_588 ();
 FILLCELL_X2 FILLER_5_604 ();
 FILLCELL_X4 FILLER_5_613 ();
 FILLCELL_X8 FILLER_5_627 ();
 FILLCELL_X4 FILLER_5_635 ();
 FILLCELL_X2 FILLER_5_639 ();
 FILLCELL_X4 FILLER_5_650 ();
 FILLCELL_X2 FILLER_5_654 ();
 FILLCELL_X1 FILLER_5_656 ();
 FILLCELL_X4 FILLER_5_661 ();
 FILLCELL_X4 FILLER_5_668 ();
 FILLCELL_X2 FILLER_5_672 ();
 FILLCELL_X4 FILLER_5_681 ();
 FILLCELL_X8 FILLER_5_687 ();
 FILLCELL_X1 FILLER_5_695 ();
 FILLCELL_X4 FILLER_5_700 ();
 FILLCELL_X8 FILLER_5_708 ();
 FILLCELL_X4 FILLER_5_720 ();
 FILLCELL_X4 FILLER_5_726 ();
 FILLCELL_X2 FILLER_5_730 ();
 FILLCELL_X8 FILLER_5_735 ();
 FILLCELL_X2 FILLER_5_743 ();
 FILLCELL_X1 FILLER_5_745 ();
 FILLCELL_X8 FILLER_5_749 ();
 FILLCELL_X2 FILLER_5_757 ();
 FILLCELL_X4 FILLER_5_762 ();
 FILLCELL_X8 FILLER_5_769 ();
 FILLCELL_X2 FILLER_5_777 ();
 FILLCELL_X1 FILLER_5_779 ();
 FILLCELL_X4 FILLER_5_784 ();
 FILLCELL_X1 FILLER_5_788 ();
 FILLCELL_X16 FILLER_5_796 ();
 FILLCELL_X8 FILLER_5_812 ();
 FILLCELL_X4 FILLER_5_820 ();
 FILLCELL_X1 FILLER_5_824 ();
 FILLCELL_X4 FILLER_5_828 ();
 FILLCELL_X8 FILLER_5_842 ();
 FILLCELL_X4 FILLER_5_850 ();
 FILLCELL_X2 FILLER_5_854 ();
 FILLCELL_X1 FILLER_5_856 ();
 FILLCELL_X4 FILLER_5_860 ();
 FILLCELL_X2 FILLER_5_864 ();
 FILLCELL_X4 FILLER_5_868 ();
 FILLCELL_X4 FILLER_5_875 ();
 FILLCELL_X4 FILLER_5_886 ();
 FILLCELL_X2 FILLER_5_890 ();
 FILLCELL_X1 FILLER_5_892 ();
 FILLCELL_X8 FILLER_5_897 ();
 FILLCELL_X1 FILLER_5_905 ();
 FILLCELL_X4 FILLER_5_915 ();
 FILLCELL_X4 FILLER_5_922 ();
 FILLCELL_X4 FILLER_5_929 ();
 FILLCELL_X8 FILLER_5_936 ();
 FILLCELL_X4 FILLER_5_944 ();
 FILLCELL_X2 FILLER_5_948 ();
 FILLCELL_X4 FILLER_5_953 ();
 FILLCELL_X1 FILLER_5_957 ();
 FILLCELL_X4 FILLER_5_967 ();
 FILLCELL_X4 FILLER_5_975 ();
 FILLCELL_X4 FILLER_5_982 ();
 FILLCELL_X8 FILLER_5_989 ();
 FILLCELL_X4 FILLER_5_997 ();
 FILLCELL_X4 FILLER_5_1020 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X8 FILLER_6_97 ();
 FILLCELL_X2 FILLER_6_105 ();
 FILLCELL_X32 FILLER_6_126 ();
 FILLCELL_X32 FILLER_6_158 ();
 FILLCELL_X32 FILLER_6_190 ();
 FILLCELL_X32 FILLER_6_222 ();
 FILLCELL_X32 FILLER_6_254 ();
 FILLCELL_X32 FILLER_6_286 ();
 FILLCELL_X32 FILLER_6_318 ();
 FILLCELL_X32 FILLER_6_350 ();
 FILLCELL_X32 FILLER_6_382 ();
 FILLCELL_X16 FILLER_6_414 ();
 FILLCELL_X4 FILLER_6_430 ();
 FILLCELL_X32 FILLER_6_453 ();
 FILLCELL_X32 FILLER_6_485 ();
 FILLCELL_X32 FILLER_6_517 ();
 FILLCELL_X32 FILLER_6_549 ();
 FILLCELL_X4 FILLER_6_581 ();
 FILLCELL_X2 FILLER_6_585 ();
 FILLCELL_X8 FILLER_6_592 ();
 FILLCELL_X2 FILLER_6_600 ();
 FILLCELL_X4 FILLER_6_612 ();
 FILLCELL_X8 FILLER_6_619 ();
 FILLCELL_X4 FILLER_6_627 ();
 FILLCELL_X4 FILLER_6_632 ();
 FILLCELL_X4 FILLER_6_645 ();
 FILLCELL_X4 FILLER_6_653 ();
 FILLCELL_X1 FILLER_6_657 ();
 FILLCELL_X4 FILLER_6_662 ();
 FILLCELL_X4 FILLER_6_671 ();
 FILLCELL_X4 FILLER_6_692 ();
 FILLCELL_X4 FILLER_6_700 ();
 FILLCELL_X32 FILLER_6_707 ();
 FILLCELL_X1 FILLER_6_739 ();
 FILLCELL_X4 FILLER_6_749 ();
 FILLCELL_X1 FILLER_6_753 ();
 FILLCELL_X4 FILLER_6_763 ();
 FILLCELL_X8 FILLER_6_770 ();
 FILLCELL_X4 FILLER_6_778 ();
 FILLCELL_X2 FILLER_6_782 ();
 FILLCELL_X4 FILLER_6_786 ();
 FILLCELL_X4 FILLER_6_800 ();
 FILLCELL_X4 FILLER_6_807 ();
 FILLCELL_X1 FILLER_6_811 ();
 FILLCELL_X8 FILLER_6_815 ();
 FILLCELL_X4 FILLER_6_823 ();
 FILLCELL_X1 FILLER_6_827 ();
 FILLCELL_X4 FILLER_6_831 ();
 FILLCELL_X8 FILLER_6_839 ();
 FILLCELL_X2 FILLER_6_847 ();
 FILLCELL_X1 FILLER_6_849 ();
 FILLCELL_X4 FILLER_6_859 ();
 FILLCELL_X4 FILLER_6_867 ();
 FILLCELL_X4 FILLER_6_874 ();
 FILLCELL_X1 FILLER_6_878 ();
 FILLCELL_X4 FILLER_6_889 ();
 FILLCELL_X8 FILLER_6_896 ();
 FILLCELL_X4 FILLER_6_908 ();
 FILLCELL_X4 FILLER_6_921 ();
 FILLCELL_X4 FILLER_6_935 ();
 FILLCELL_X8 FILLER_6_946 ();
 FILLCELL_X1 FILLER_6_954 ();
 FILLCELL_X4 FILLER_6_964 ();
 FILLCELL_X4 FILLER_6_972 ();
 FILLCELL_X8 FILLER_6_979 ();
 FILLCELL_X4 FILLER_6_987 ();
 FILLCELL_X1 FILLER_6_991 ();
 FILLCELL_X8 FILLER_6_998 ();
 FILLCELL_X2 FILLER_6_1006 ();
 FILLCELL_X8 FILLER_6_1012 ();
 FILLCELL_X4 FILLER_6_1020 ();
 FILLCELL_X4 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_8 ();
 FILLCELL_X32 FILLER_7_40 ();
 FILLCELL_X32 FILLER_7_72 ();
 FILLCELL_X32 FILLER_7_104 ();
 FILLCELL_X32 FILLER_7_136 ();
 FILLCELL_X32 FILLER_7_168 ();
 FILLCELL_X32 FILLER_7_200 ();
 FILLCELL_X8 FILLER_7_232 ();
 FILLCELL_X2 FILLER_7_240 ();
 FILLCELL_X1 FILLER_7_242 ();
 FILLCELL_X32 FILLER_7_262 ();
 FILLCELL_X32 FILLER_7_294 ();
 FILLCELL_X32 FILLER_7_326 ();
 FILLCELL_X32 FILLER_7_358 ();
 FILLCELL_X16 FILLER_7_390 ();
 FILLCELL_X8 FILLER_7_406 ();
 FILLCELL_X1 FILLER_7_414 ();
 FILLCELL_X16 FILLER_7_434 ();
 FILLCELL_X8 FILLER_7_450 ();
 FILLCELL_X4 FILLER_7_458 ();
 FILLCELL_X2 FILLER_7_462 ();
 FILLCELL_X32 FILLER_7_483 ();
 FILLCELL_X32 FILLER_7_515 ();
 FILLCELL_X32 FILLER_7_547 ();
 FILLCELL_X4 FILLER_7_579 ();
 FILLCELL_X2 FILLER_7_583 ();
 FILLCELL_X1 FILLER_7_585 ();
 FILLCELL_X8 FILLER_7_595 ();
 FILLCELL_X4 FILLER_7_603 ();
 FILLCELL_X2 FILLER_7_607 ();
 FILLCELL_X4 FILLER_7_613 ();
 FILLCELL_X4 FILLER_7_636 ();
 FILLCELL_X4 FILLER_7_644 ();
 FILLCELL_X8 FILLER_7_651 ();
 FILLCELL_X8 FILLER_7_662 ();
 FILLCELL_X4 FILLER_7_670 ();
 FILLCELL_X1 FILLER_7_674 ();
 FILLCELL_X4 FILLER_7_680 ();
 FILLCELL_X8 FILLER_7_688 ();
 FILLCELL_X1 FILLER_7_696 ();
 FILLCELL_X4 FILLER_7_707 ();
 FILLCELL_X4 FILLER_7_718 ();
 FILLCELL_X2 FILLER_7_722 ();
 FILLCELL_X1 FILLER_7_724 ();
 FILLCELL_X4 FILLER_7_729 ();
 FILLCELL_X2 FILLER_7_733 ();
 FILLCELL_X4 FILLER_7_739 ();
 FILLCELL_X16 FILLER_7_746 ();
 FILLCELL_X4 FILLER_7_762 ();
 FILLCELL_X1 FILLER_7_766 ();
 FILLCELL_X8 FILLER_7_777 ();
 FILLCELL_X4 FILLER_7_789 ();
 FILLCELL_X4 FILLER_7_803 ();
 FILLCELL_X4 FILLER_7_816 ();
 FILLCELL_X4 FILLER_7_829 ();
 FILLCELL_X4 FILLER_7_836 ();
 FILLCELL_X4 FILLER_7_844 ();
 FILLCELL_X1 FILLER_7_848 ();
 FILLCELL_X4 FILLER_7_853 ();
 FILLCELL_X8 FILLER_7_866 ();
 FILLCELL_X4 FILLER_7_874 ();
 FILLCELL_X4 FILLER_7_882 ();
 FILLCELL_X8 FILLER_7_895 ();
 FILLCELL_X4 FILLER_7_903 ();
 FILLCELL_X4 FILLER_7_910 ();
 FILLCELL_X4 FILLER_7_918 ();
 FILLCELL_X8 FILLER_7_926 ();
 FILLCELL_X4 FILLER_7_944 ();
 FILLCELL_X2 FILLER_7_948 ();
 FILLCELL_X1 FILLER_7_950 ();
 FILLCELL_X4 FILLER_7_955 ();
 FILLCELL_X8 FILLER_7_963 ();
 FILLCELL_X2 FILLER_7_971 ();
 FILLCELL_X4 FILLER_7_977 ();
 FILLCELL_X4 FILLER_7_986 ();
 FILLCELL_X4 FILLER_7_992 ();
 FILLCELL_X2 FILLER_7_996 ();
 FILLCELL_X4 FILLER_7_1004 ();
 FILLCELL_X8 FILLER_7_1010 ();
 FILLCELL_X4 FILLER_7_1018 ();
 FILLCELL_X2 FILLER_7_1022 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X16 FILLER_8_225 ();
 FILLCELL_X32 FILLER_8_245 ();
 FILLCELL_X32 FILLER_8_277 ();
 FILLCELL_X32 FILLER_8_309 ();
 FILLCELL_X32 FILLER_8_341 ();
 FILLCELL_X8 FILLER_8_373 ();
 FILLCELL_X4 FILLER_8_400 ();
 FILLCELL_X4 FILLER_8_408 ();
 FILLCELL_X4 FILLER_8_431 ();
 FILLCELL_X8 FILLER_8_439 ();
 FILLCELL_X4 FILLER_8_447 ();
 FILLCELL_X4 FILLER_8_470 ();
 FILLCELL_X32 FILLER_8_493 ();
 FILLCELL_X16 FILLER_8_525 ();
 FILLCELL_X8 FILLER_8_541 ();
 FILLCELL_X2 FILLER_8_549 ();
 FILLCELL_X16 FILLER_8_555 ();
 FILLCELL_X8 FILLER_8_571 ();
 FILLCELL_X1 FILLER_8_579 ();
 FILLCELL_X4 FILLER_8_589 ();
 FILLCELL_X4 FILLER_8_596 ();
 FILLCELL_X1 FILLER_8_600 ();
 FILLCELL_X16 FILLER_8_605 ();
 FILLCELL_X2 FILLER_8_621 ();
 FILLCELL_X4 FILLER_8_626 ();
 FILLCELL_X1 FILLER_8_630 ();
 FILLCELL_X4 FILLER_8_632 ();
 FILLCELL_X1 FILLER_8_636 ();
 FILLCELL_X4 FILLER_8_641 ();
 FILLCELL_X4 FILLER_8_649 ();
 FILLCELL_X4 FILLER_8_656 ();
 FILLCELL_X8 FILLER_8_663 ();
 FILLCELL_X4 FILLER_8_675 ();
 FILLCELL_X1 FILLER_8_679 ();
 FILLCELL_X8 FILLER_8_683 ();
 FILLCELL_X4 FILLER_8_693 ();
 FILLCELL_X4 FILLER_8_700 ();
 FILLCELL_X4 FILLER_8_707 ();
 FILLCELL_X8 FILLER_8_713 ();
 FILLCELL_X2 FILLER_8_721 ();
 FILLCELL_X4 FILLER_8_726 ();
 FILLCELL_X4 FILLER_8_739 ();
 FILLCELL_X4 FILLER_8_752 ();
 FILLCELL_X2 FILLER_8_756 ();
 FILLCELL_X1 FILLER_8_758 ();
 FILLCELL_X8 FILLER_8_776 ();
 FILLCELL_X1 FILLER_8_784 ();
 FILLCELL_X4 FILLER_8_792 ();
 FILLCELL_X16 FILLER_8_798 ();
 FILLCELL_X2 FILLER_8_814 ();
 FILLCELL_X4 FILLER_8_819 ();
 FILLCELL_X1 FILLER_8_823 ();
 FILLCELL_X4 FILLER_8_827 ();
 FILLCELL_X4 FILLER_8_838 ();
 FILLCELL_X8 FILLER_8_848 ();
 FILLCELL_X2 FILLER_8_856 ();
 FILLCELL_X8 FILLER_8_862 ();
 FILLCELL_X4 FILLER_8_870 ();
 FILLCELL_X1 FILLER_8_874 ();
 FILLCELL_X8 FILLER_8_882 ();
 FILLCELL_X4 FILLER_8_890 ();
 FILLCELL_X1 FILLER_8_894 ();
 FILLCELL_X16 FILLER_8_898 ();
 FILLCELL_X8 FILLER_8_914 ();
 FILLCELL_X2 FILLER_8_922 ();
 FILLCELL_X1 FILLER_8_924 ();
 FILLCELL_X4 FILLER_8_928 ();
 FILLCELL_X4 FILLER_8_936 ();
 FILLCELL_X8 FILLER_8_942 ();
 FILLCELL_X4 FILLER_8_950 ();
 FILLCELL_X2 FILLER_8_954 ();
 FILLCELL_X4 FILLER_8_959 ();
 FILLCELL_X4 FILLER_8_967 ();
 FILLCELL_X4 FILLER_8_978 ();
 FILLCELL_X4 FILLER_8_999 ();
 FILLCELL_X2 FILLER_8_1003 ();
 FILLCELL_X1 FILLER_8_1005 ();
 FILLCELL_X8 FILLER_8_1010 ();
 FILLCELL_X4 FILLER_8_1018 ();
 FILLCELL_X2 FILLER_8_1022 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X32 FILLER_9_257 ();
 FILLCELL_X32 FILLER_9_289 ();
 FILLCELL_X32 FILLER_9_321 ();
 FILLCELL_X16 FILLER_9_353 ();
 FILLCELL_X8 FILLER_9_369 ();
 FILLCELL_X4 FILLER_9_377 ();
 FILLCELL_X8 FILLER_9_385 ();
 FILLCELL_X16 FILLER_9_412 ();
 FILLCELL_X8 FILLER_9_428 ();
 FILLCELL_X4 FILLER_9_440 ();
 FILLCELL_X4 FILLER_9_463 ();
 FILLCELL_X8 FILLER_9_471 ();
 FILLCELL_X4 FILLER_9_479 ();
 FILLCELL_X2 FILLER_9_483 ();
 FILLCELL_X32 FILLER_9_504 ();
 FILLCELL_X16 FILLER_9_536 ();
 FILLCELL_X4 FILLER_9_552 ();
 FILLCELL_X1 FILLER_9_556 ();
 FILLCELL_X16 FILLER_9_561 ();
 FILLCELL_X4 FILLER_9_577 ();
 FILLCELL_X2 FILLER_9_581 ();
 FILLCELL_X4 FILLER_9_587 ();
 FILLCELL_X8 FILLER_9_594 ();
 FILLCELL_X2 FILLER_9_602 ();
 FILLCELL_X1 FILLER_9_604 ();
 FILLCELL_X4 FILLER_9_608 ();
 FILLCELL_X4 FILLER_9_616 ();
 FILLCELL_X8 FILLER_9_623 ();
 FILLCELL_X1 FILLER_9_631 ();
 FILLCELL_X4 FILLER_9_636 ();
 FILLCELL_X4 FILLER_9_649 ();
 FILLCELL_X8 FILLER_9_662 ();
 FILLCELL_X4 FILLER_9_674 ();
 FILLCELL_X4 FILLER_9_688 ();
 FILLCELL_X8 FILLER_9_699 ();
 FILLCELL_X4 FILLER_9_717 ();
 FILLCELL_X4 FILLER_9_725 ();
 FILLCELL_X4 FILLER_9_732 ();
 FILLCELL_X8 FILLER_9_739 ();
 FILLCELL_X2 FILLER_9_747 ();
 FILLCELL_X1 FILLER_9_749 ();
 FILLCELL_X4 FILLER_9_754 ();
 FILLCELL_X4 FILLER_9_765 ();
 FILLCELL_X8 FILLER_9_774 ();
 FILLCELL_X1 FILLER_9_782 ();
 FILLCELL_X4 FILLER_9_793 ();
 FILLCELL_X8 FILLER_9_800 ();
 FILLCELL_X4 FILLER_9_808 ();
 FILLCELL_X4 FILLER_9_815 ();
 FILLCELL_X4 FILLER_9_826 ();
 FILLCELL_X8 FILLER_9_840 ();
 FILLCELL_X2 FILLER_9_848 ();
 FILLCELL_X1 FILLER_9_850 ();
 FILLCELL_X4 FILLER_9_861 ();
 FILLCELL_X2 FILLER_9_865 ();
 FILLCELL_X1 FILLER_9_867 ();
 FILLCELL_X4 FILLER_9_872 ();
 FILLCELL_X4 FILLER_9_886 ();
 FILLCELL_X8 FILLER_9_893 ();
 FILLCELL_X4 FILLER_9_910 ();
 FILLCELL_X16 FILLER_9_917 ();
 FILLCELL_X4 FILLER_9_933 ();
 FILLCELL_X1 FILLER_9_937 ();
 FILLCELL_X4 FILLER_9_947 ();
 FILLCELL_X8 FILLER_9_954 ();
 FILLCELL_X8 FILLER_9_965 ();
 FILLCELL_X4 FILLER_9_973 ();
 FILLCELL_X2 FILLER_9_977 ();
 FILLCELL_X8 FILLER_9_984 ();
 FILLCELL_X2 FILLER_9_992 ();
 FILLCELL_X8 FILLER_9_1000 ();
 FILLCELL_X8 FILLER_9_1014 ();
 FILLCELL_X2 FILLER_9_1022 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X32 FILLER_10_257 ();
 FILLCELL_X32 FILLER_10_289 ();
 FILLCELL_X32 FILLER_10_321 ();
 FILLCELL_X4 FILLER_10_353 ();
 FILLCELL_X8 FILLER_10_361 ();
 FILLCELL_X1 FILLER_10_369 ();
 FILLCELL_X8 FILLER_10_389 ();
 FILLCELL_X2 FILLER_10_397 ();
 FILLCELL_X1 FILLER_10_399 ();
 FILLCELL_X4 FILLER_10_404 ();
 FILLCELL_X16 FILLER_10_412 ();
 FILLCELL_X4 FILLER_10_428 ();
 FILLCELL_X1 FILLER_10_432 ();
 FILLCELL_X4 FILLER_10_452 ();
 FILLCELL_X4 FILLER_10_460 ();
 FILLCELL_X16 FILLER_10_468 ();
 FILLCELL_X4 FILLER_10_484 ();
 FILLCELL_X4 FILLER_10_507 ();
 FILLCELL_X16 FILLER_10_530 ();
 FILLCELL_X8 FILLER_10_546 ();
 FILLCELL_X2 FILLER_10_554 ();
 FILLCELL_X4 FILLER_10_575 ();
 FILLCELL_X4 FILLER_10_583 ();
 FILLCELL_X4 FILLER_10_591 ();
 FILLCELL_X4 FILLER_10_599 ();
 FILLCELL_X4 FILLER_10_612 ();
 FILLCELL_X4 FILLER_10_625 ();
 FILLCELL_X2 FILLER_10_629 ();
 FILLCELL_X4 FILLER_10_632 ();
 FILLCELL_X4 FILLER_10_640 ();
 FILLCELL_X2 FILLER_10_644 ();
 FILLCELL_X4 FILLER_10_650 ();
 FILLCELL_X16 FILLER_10_657 ();
 FILLCELL_X8 FILLER_10_673 ();
 FILLCELL_X4 FILLER_10_681 ();
 FILLCELL_X2 FILLER_10_685 ();
 FILLCELL_X1 FILLER_10_687 ();
 FILLCELL_X4 FILLER_10_698 ();
 FILLCELL_X8 FILLER_10_711 ();
 FILLCELL_X1 FILLER_10_719 ();
 FILLCELL_X4 FILLER_10_730 ();
 FILLCELL_X8 FILLER_10_741 ();
 FILLCELL_X1 FILLER_10_749 ();
 FILLCELL_X8 FILLER_10_754 ();
 FILLCELL_X4 FILLER_10_767 ();
 FILLCELL_X2 FILLER_10_771 ();
 FILLCELL_X4 FILLER_10_777 ();
 FILLCELL_X8 FILLER_10_785 ();
 FILLCELL_X2 FILLER_10_793 ();
 FILLCELL_X1 FILLER_10_795 ();
 FILLCELL_X4 FILLER_10_805 ();
 FILLCELL_X4 FILLER_10_813 ();
 FILLCELL_X8 FILLER_10_820 ();
 FILLCELL_X4 FILLER_10_834 ();
 FILLCELL_X16 FILLER_10_841 ();
 FILLCELL_X4 FILLER_10_859 ();
 FILLCELL_X4 FILLER_10_867 ();
 FILLCELL_X8 FILLER_10_874 ();
 FILLCELL_X1 FILLER_10_882 ();
 FILLCELL_X4 FILLER_10_886 ();
 FILLCELL_X4 FILLER_10_899 ();
 FILLCELL_X2 FILLER_10_903 ();
 FILLCELL_X1 FILLER_10_905 ();
 FILLCELL_X8 FILLER_10_909 ();
 FILLCELL_X4 FILLER_10_917 ();
 FILLCELL_X2 FILLER_10_921 ();
 FILLCELL_X1 FILLER_10_923 ();
 FILLCELL_X4 FILLER_10_929 ();
 FILLCELL_X1 FILLER_10_933 ();
 FILLCELL_X4 FILLER_10_938 ();
 FILLCELL_X4 FILLER_10_946 ();
 FILLCELL_X8 FILLER_10_953 ();
 FILLCELL_X8 FILLER_10_971 ();
 FILLCELL_X4 FILLER_10_979 ();
 FILLCELL_X1 FILLER_10_983 ();
 FILLCELL_X4 FILLER_10_988 ();
 FILLCELL_X4 FILLER_10_996 ();
 FILLCELL_X8 FILLER_10_1003 ();
 FILLCELL_X1 FILLER_10_1011 ();
 FILLCELL_X8 FILLER_10_1016 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_11_193 ();
 FILLCELL_X32 FILLER_11_225 ();
 FILLCELL_X32 FILLER_11_257 ();
 FILLCELL_X32 FILLER_11_289 ();
 FILLCELL_X8 FILLER_11_321 ();
 FILLCELL_X2 FILLER_11_329 ();
 FILLCELL_X1 FILLER_11_331 ();
 FILLCELL_X4 FILLER_11_337 ();
 FILLCELL_X8 FILLER_11_344 ();
 FILLCELL_X2 FILLER_11_352 ();
 FILLCELL_X4 FILLER_11_373 ();
 FILLCELL_X8 FILLER_11_381 ();
 FILLCELL_X1 FILLER_11_389 ();
 FILLCELL_X4 FILLER_11_394 ();
 FILLCELL_X4 FILLER_11_403 ();
 FILLCELL_X4 FILLER_11_426 ();
 FILLCELL_X16 FILLER_11_434 ();
 FILLCELL_X8 FILLER_11_450 ();
 FILLCELL_X2 FILLER_11_458 ();
 FILLCELL_X8 FILLER_11_465 ();
 FILLCELL_X4 FILLER_11_477 ();
 FILLCELL_X2 FILLER_11_481 ();
 FILLCELL_X4 FILLER_11_487 ();
 FILLCELL_X1 FILLER_11_491 ();
 FILLCELL_X4 FILLER_11_495 ();
 FILLCELL_X8 FILLER_11_503 ();
 FILLCELL_X4 FILLER_11_511 ();
 FILLCELL_X2 FILLER_11_515 ();
 FILLCELL_X1 FILLER_11_517 ();
 FILLCELL_X16 FILLER_11_521 ();
 FILLCELL_X8 FILLER_11_537 ();
 FILLCELL_X1 FILLER_11_545 ();
 FILLCELL_X32 FILLER_11_549 ();
 FILLCELL_X16 FILLER_11_581 ();
 FILLCELL_X4 FILLER_11_597 ();
 FILLCELL_X16 FILLER_11_605 ();
 FILLCELL_X2 FILLER_11_621 ();
 FILLCELL_X1 FILLER_11_623 ();
 FILLCELL_X4 FILLER_11_627 ();
 FILLCELL_X8 FILLER_11_632 ();
 FILLCELL_X1 FILLER_11_640 ();
 FILLCELL_X16 FILLER_11_660 ();
 FILLCELL_X8 FILLER_11_676 ();
 FILLCELL_X2 FILLER_11_684 ();
 FILLCELL_X8 FILLER_11_689 ();
 FILLCELL_X4 FILLER_11_700 ();
 FILLCELL_X4 FILLER_11_707 ();
 FILLCELL_X1 FILLER_11_711 ();
 FILLCELL_X4 FILLER_11_721 ();
 FILLCELL_X4 FILLER_11_735 ();
 FILLCELL_X2 FILLER_11_739 ();
 FILLCELL_X8 FILLER_11_743 ();
 FILLCELL_X4 FILLER_11_751 ();
 FILLCELL_X1 FILLER_11_755 ();
 FILLCELL_X8 FILLER_11_760 ();
 FILLCELL_X1 FILLER_11_768 ();
 FILLCELL_X16 FILLER_11_771 ();
 FILLCELL_X4 FILLER_11_787 ();
 FILLCELL_X2 FILLER_11_791 ();
 FILLCELL_X4 FILLER_11_797 ();
 FILLCELL_X4 FILLER_11_810 ();
 FILLCELL_X4 FILLER_11_818 ();
 FILLCELL_X8 FILLER_11_825 ();
 FILLCELL_X4 FILLER_11_833 ();
 FILLCELL_X4 FILLER_11_840 ();
 FILLCELL_X8 FILLER_11_846 ();
 FILLCELL_X1 FILLER_11_854 ();
 FILLCELL_X4 FILLER_11_860 ();
 FILLCELL_X4 FILLER_11_873 ();
 FILLCELL_X8 FILLER_11_880 ();
 FILLCELL_X4 FILLER_11_892 ();
 FILLCELL_X4 FILLER_11_905 ();
 FILLCELL_X1 FILLER_11_909 ();
 FILLCELL_X8 FILLER_11_912 ();
 FILLCELL_X4 FILLER_11_937 ();
 FILLCELL_X4 FILLER_11_950 ();
 FILLCELL_X2 FILLER_11_954 ();
 FILLCELL_X4 FILLER_11_960 ();
 FILLCELL_X2 FILLER_11_964 ();
 FILLCELL_X1 FILLER_11_966 ();
 FILLCELL_X8 FILLER_11_974 ();
 FILLCELL_X4 FILLER_11_991 ();
 FILLCELL_X4 FILLER_11_998 ();
 FILLCELL_X4 FILLER_11_1005 ();
 FILLCELL_X8 FILLER_11_1012 ();
 FILLCELL_X4 FILLER_11_1020 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X8 FILLER_12_161 ();
 FILLCELL_X8 FILLER_12_819 ();
 FILLCELL_X4 FILLER_12_827 ();
 FILLCELL_X2 FILLER_12_831 ();
 FILLCELL_X1 FILLER_12_833 ();
 FILLCELL_X4 FILLER_12_844 ();
 FILLCELL_X4 FILLER_12_851 ();
 FILLCELL_X4 FILLER_12_858 ();
 FILLCELL_X2 FILLER_12_862 ();
 FILLCELL_X8 FILLER_12_868 ();
 FILLCELL_X1 FILLER_12_876 ();
 FILLCELL_X8 FILLER_12_886 ();
 FILLCELL_X1 FILLER_12_894 ();
 FILLCELL_X4 FILLER_12_899 ();
 FILLCELL_X4 FILLER_12_907 ();
 FILLCELL_X1 FILLER_12_911 ();
 FILLCELL_X4 FILLER_12_916 ();
 FILLCELL_X4 FILLER_12_927 ();
 FILLCELL_X4 FILLER_12_936 ();
 FILLCELL_X4 FILLER_12_944 ();
 FILLCELL_X2 FILLER_12_948 ();
 FILLCELL_X1 FILLER_12_950 ();
 FILLCELL_X4 FILLER_12_955 ();
 FILLCELL_X1 FILLER_12_959 ();
 FILLCELL_X8 FILLER_12_970 ();
 FILLCELL_X2 FILLER_12_978 ();
 FILLCELL_X4 FILLER_12_983 ();
 FILLCELL_X16 FILLER_12_996 ();
 FILLCELL_X8 FILLER_12_1012 ();
 FILLCELL_X4 FILLER_12_1020 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X8 FILLER_13_161 ();
 FILLCELL_X4 FILLER_13_819 ();
 FILLCELL_X4 FILLER_13_826 ();
 FILLCELL_X4 FILLER_13_833 ();
 FILLCELL_X2 FILLER_13_837 ();
 FILLCELL_X1 FILLER_13_839 ();
 FILLCELL_X4 FILLER_13_844 ();
 FILLCELL_X4 FILLER_13_857 ();
 FILLCELL_X4 FILLER_13_865 ();
 FILLCELL_X2 FILLER_13_869 ();
 FILLCELL_X8 FILLER_13_875 ();
 FILLCELL_X4 FILLER_13_883 ();
 FILLCELL_X4 FILLER_13_890 ();
 FILLCELL_X16 FILLER_13_898 ();
 FILLCELL_X4 FILLER_13_914 ();
 FILLCELL_X2 FILLER_13_918 ();
 FILLCELL_X4 FILLER_13_924 ();
 FILLCELL_X8 FILLER_13_932 ();
 FILLCELL_X2 FILLER_13_940 ();
 FILLCELL_X4 FILLER_13_945 ();
 FILLCELL_X2 FILLER_13_949 ();
 FILLCELL_X4 FILLER_13_960 ();
 FILLCELL_X16 FILLER_13_966 ();
 FILLCELL_X4 FILLER_13_982 ();
 FILLCELL_X2 FILLER_13_986 ();
 FILLCELL_X4 FILLER_13_991 ();
 FILLCELL_X2 FILLER_13_995 ();
 FILLCELL_X1 FILLER_13_997 ();
 FILLCELL_X8 FILLER_13_1008 ();
 FILLCELL_X1 FILLER_13_1016 ();
 FILLCELL_X4 FILLER_13_1020 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X8 FILLER_14_161 ();
 FILLCELL_X4 FILLER_14_819 ();
 FILLCELL_X4 FILLER_14_833 ();
 FILLCELL_X4 FILLER_14_846 ();
 FILLCELL_X2 FILLER_14_850 ();
 FILLCELL_X1 FILLER_14_852 ();
 FILLCELL_X4 FILLER_14_862 ();
 FILLCELL_X2 FILLER_14_866 ();
 FILLCELL_X8 FILLER_14_871 ();
 FILLCELL_X4 FILLER_14_879 ();
 FILLCELL_X2 FILLER_14_883 ();
 FILLCELL_X4 FILLER_14_888 ();
 FILLCELL_X32 FILLER_14_902 ();
 FILLCELL_X4 FILLER_14_934 ();
 FILLCELL_X2 FILLER_14_938 ();
 FILLCELL_X4 FILLER_14_949 ();
 FILLCELL_X16 FILLER_14_956 ();
 FILLCELL_X8 FILLER_14_976 ();
 FILLCELL_X1 FILLER_14_984 ();
 FILLCELL_X4 FILLER_14_995 ();
 FILLCELL_X4 FILLER_14_1003 ();
 FILLCELL_X4 FILLER_14_1011 ();
 FILLCELL_X4 FILLER_14_1017 ();
 FILLCELL_X2 FILLER_14_1021 ();
 FILLCELL_X1 FILLER_14_1023 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X8 FILLER_15_161 ();
 FILLCELL_X8 FILLER_15_819 ();
 FILLCELL_X1 FILLER_15_827 ();
 FILLCELL_X4 FILLER_15_835 ();
 FILLCELL_X4 FILLER_15_842 ();
 FILLCELL_X4 FILLER_15_850 ();
 FILLCELL_X2 FILLER_15_854 ();
 FILLCELL_X4 FILLER_15_859 ();
 FILLCELL_X4 FILLER_15_867 ();
 FILLCELL_X2 FILLER_15_871 ();
 FILLCELL_X8 FILLER_15_877 ();
 FILLCELL_X4 FILLER_15_885 ();
 FILLCELL_X2 FILLER_15_889 ();
 FILLCELL_X4 FILLER_15_898 ();
 FILLCELL_X8 FILLER_15_904 ();
 FILLCELL_X4 FILLER_15_912 ();
 FILLCELL_X1 FILLER_15_916 ();
 FILLCELL_X4 FILLER_15_921 ();
 FILLCELL_X4 FILLER_15_928 ();
 FILLCELL_X4 FILLER_15_936 ();
 FILLCELL_X4 FILLER_15_944 ();
 FILLCELL_X4 FILLER_15_951 ();
 FILLCELL_X16 FILLER_15_958 ();
 FILLCELL_X1 FILLER_15_974 ();
 FILLCELL_X4 FILLER_15_978 ();
 FILLCELL_X8 FILLER_15_1001 ();
 FILLCELL_X8 FILLER_15_1013 ();
 FILLCELL_X2 FILLER_15_1021 ();
 FILLCELL_X1 FILLER_15_1023 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X8 FILLER_16_161 ();
 FILLCELL_X4 FILLER_16_819 ();
 FILLCELL_X1 FILLER_16_823 ();
 FILLCELL_X4 FILLER_16_833 ();
 FILLCELL_X4 FILLER_16_840 ();
 FILLCELL_X8 FILLER_16_847 ();
 FILLCELL_X2 FILLER_16_855 ();
 FILLCELL_X1 FILLER_16_857 ();
 FILLCELL_X4 FILLER_16_862 ();
 FILLCELL_X4 FILLER_16_875 ();
 FILLCELL_X4 FILLER_16_888 ();
 FILLCELL_X2 FILLER_16_892 ();
 FILLCELL_X1 FILLER_16_894 ();
 FILLCELL_X4 FILLER_16_905 ();
 FILLCELL_X4 FILLER_16_913 ();
 FILLCELL_X4 FILLER_16_926 ();
 FILLCELL_X16 FILLER_16_934 ();
 FILLCELL_X8 FILLER_16_950 ();
 FILLCELL_X8 FILLER_16_962 ();
 FILLCELL_X2 FILLER_16_970 ();
 FILLCELL_X4 FILLER_16_976 ();
 FILLCELL_X8 FILLER_16_984 ();
 FILLCELL_X1 FILLER_16_992 ();
 FILLCELL_X4 FILLER_16_999 ();
 FILLCELL_X4 FILLER_16_1020 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X8 FILLER_17_161 ();
 FILLCELL_X4 FILLER_17_819 ();
 FILLCELL_X2 FILLER_17_823 ();
 FILLCELL_X1 FILLER_17_825 ();
 FILLCELL_X4 FILLER_17_831 ();
 FILLCELL_X4 FILLER_17_845 ();
 FILLCELL_X8 FILLER_17_851 ();
 FILLCELL_X1 FILLER_17_859 ();
 FILLCELL_X4 FILLER_17_863 ();
 FILLCELL_X8 FILLER_17_870 ();
 FILLCELL_X1 FILLER_17_878 ();
 FILLCELL_X4 FILLER_17_882 ();
 FILLCELL_X2 FILLER_17_886 ();
 FILLCELL_X4 FILLER_17_891 ();
 FILLCELL_X4 FILLER_17_905 ();
 FILLCELL_X8 FILLER_17_912 ();
 FILLCELL_X1 FILLER_17_920 ();
 FILLCELL_X4 FILLER_17_925 ();
 FILLCELL_X8 FILLER_17_932 ();
 FILLCELL_X4 FILLER_17_940 ();
 FILLCELL_X2 FILLER_17_944 ();
 FILLCELL_X4 FILLER_17_950 ();
 FILLCELL_X4 FILLER_17_958 ();
 FILLCELL_X2 FILLER_17_962 ();
 FILLCELL_X4 FILLER_17_970 ();
 FILLCELL_X4 FILLER_17_979 ();
 FILLCELL_X4 FILLER_17_987 ();
 FILLCELL_X4 FILLER_17_995 ();
 FILLCELL_X2 FILLER_17_999 ();
 FILLCELL_X4 FILLER_17_1007 ();
 FILLCELL_X8 FILLER_17_1015 ();
 FILLCELL_X1 FILLER_17_1023 ();
 FILLCELL_X4 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_8 ();
 FILLCELL_X32 FILLER_18_40 ();
 FILLCELL_X32 FILLER_18_72 ();
 FILLCELL_X32 FILLER_18_104 ();
 FILLCELL_X32 FILLER_18_136 ();
 FILLCELL_X1 FILLER_18_168 ();
 FILLCELL_X4 FILLER_18_819 ();
 FILLCELL_X2 FILLER_18_823 ();
 FILLCELL_X1 FILLER_18_825 ();
 FILLCELL_X8 FILLER_18_828 ();
 FILLCELL_X1 FILLER_18_836 ();
 FILLCELL_X8 FILLER_18_844 ();
 FILLCELL_X4 FILLER_18_852 ();
 FILLCELL_X2 FILLER_18_856 ();
 FILLCELL_X4 FILLER_18_861 ();
 FILLCELL_X8 FILLER_18_868 ();
 FILLCELL_X2 FILLER_18_876 ();
 FILLCELL_X8 FILLER_18_887 ();
 FILLCELL_X4 FILLER_18_902 ();
 FILLCELL_X8 FILLER_18_908 ();
 FILLCELL_X2 FILLER_18_916 ();
 FILLCELL_X1 FILLER_18_918 ();
 FILLCELL_X8 FILLER_18_928 ();
 FILLCELL_X4 FILLER_18_936 ();
 FILLCELL_X4 FILLER_18_950 ();
 FILLCELL_X4 FILLER_18_960 ();
 FILLCELL_X2 FILLER_18_964 ();
 FILLCELL_X4 FILLER_18_968 ();
 FILLCELL_X8 FILLER_18_981 ();
 FILLCELL_X2 FILLER_18_989 ();
 FILLCELL_X4 FILLER_18_997 ();
 FILLCELL_X4 FILLER_18_1020 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X8 FILLER_19_161 ();
 FILLCELL_X4 FILLER_19_819 ();
 FILLCELL_X1 FILLER_19_823 ();
 FILLCELL_X8 FILLER_19_830 ();
 FILLCELL_X8 FILLER_19_840 ();
 FILLCELL_X2 FILLER_19_848 ();
 FILLCELL_X1 FILLER_19_850 ();
 FILLCELL_X4 FILLER_19_855 ();
 FILLCELL_X8 FILLER_19_869 ();
 FILLCELL_X1 FILLER_19_877 ();
 FILLCELL_X8 FILLER_19_881 ();
 FILLCELL_X4 FILLER_19_889 ();
 FILLCELL_X4 FILLER_19_903 ();
 FILLCELL_X16 FILLER_19_910 ();
 FILLCELL_X8 FILLER_19_926 ();
 FILLCELL_X2 FILLER_19_934 ();
 FILLCELL_X4 FILLER_19_939 ();
 FILLCELL_X8 FILLER_19_945 ();
 FILLCELL_X4 FILLER_19_957 ();
 FILLCELL_X4 FILLER_19_965 ();
 FILLCELL_X1 FILLER_19_969 ();
 FILLCELL_X8 FILLER_19_975 ();
 FILLCELL_X2 FILLER_19_983 ();
 FILLCELL_X8 FILLER_19_991 ();
 FILLCELL_X2 FILLER_19_999 ();
 FILLCELL_X8 FILLER_19_1005 ();
 FILLCELL_X2 FILLER_19_1013 ();
 FILLCELL_X4 FILLER_19_1019 ();
 FILLCELL_X1 FILLER_19_1023 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X8 FILLER_20_161 ();
 FILLCELL_X4 FILLER_20_819 ();
 FILLCELL_X4 FILLER_20_830 ();
 FILLCELL_X1 FILLER_20_834 ();
 FILLCELL_X4 FILLER_20_845 ();
 FILLCELL_X2 FILLER_20_849 ();
 FILLCELL_X1 FILLER_20_851 ();
 FILLCELL_X4 FILLER_20_854 ();
 FILLCELL_X4 FILLER_20_867 ();
 FILLCELL_X4 FILLER_20_878 ();
 FILLCELL_X2 FILLER_20_882 ();
 FILLCELL_X4 FILLER_20_893 ();
 FILLCELL_X4 FILLER_20_900 ();
 FILLCELL_X4 FILLER_20_907 ();
 FILLCELL_X8 FILLER_20_915 ();
 FILLCELL_X4 FILLER_20_923 ();
 FILLCELL_X4 FILLER_20_931 ();
 FILLCELL_X4 FILLER_20_945 ();
 FILLCELL_X8 FILLER_20_956 ();
 FILLCELL_X2 FILLER_20_964 ();
 FILLCELL_X1 FILLER_20_966 ();
 FILLCELL_X4 FILLER_20_970 ();
 FILLCELL_X2 FILLER_20_974 ();
 FILLCELL_X1 FILLER_20_976 ();
 FILLCELL_X4 FILLER_20_981 ();
 FILLCELL_X4 FILLER_20_988 ();
 FILLCELL_X16 FILLER_20_995 ();
 FILLCELL_X8 FILLER_20_1011 ();
 FILLCELL_X4 FILLER_20_1019 ();
 FILLCELL_X1 FILLER_20_1023 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X8 FILLER_21_161 ();
 FILLCELL_X4 FILLER_21_819 ();
 FILLCELL_X4 FILLER_21_833 ();
 FILLCELL_X4 FILLER_21_841 ();
 FILLCELL_X16 FILLER_21_849 ();
 FILLCELL_X1 FILLER_21_865 ();
 FILLCELL_X4 FILLER_21_876 ();
 FILLCELL_X8 FILLER_21_883 ();
 FILLCELL_X4 FILLER_21_891 ();
 FILLCELL_X1 FILLER_21_895 ();
 FILLCELL_X4 FILLER_21_899 ();
 FILLCELL_X4 FILLER_21_907 ();
 FILLCELL_X4 FILLER_21_920 ();
 FILLCELL_X32 FILLER_21_928 ();
 FILLCELL_X4 FILLER_21_960 ();
 FILLCELL_X2 FILLER_21_964 ();
 FILLCELL_X4 FILLER_21_970 ();
 FILLCELL_X2 FILLER_21_974 ();
 FILLCELL_X4 FILLER_21_980 ();
 FILLCELL_X4 FILLER_21_987 ();
 FILLCELL_X4 FILLER_21_998 ();
 FILLCELL_X16 FILLER_21_1004 ();
 FILLCELL_X4 FILLER_21_1020 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X8 FILLER_22_161 ();
 FILLCELL_X4 FILLER_22_819 ();
 FILLCELL_X4 FILLER_22_829 ();
 FILLCELL_X1 FILLER_22_833 ();
 FILLCELL_X4 FILLER_22_841 ();
 FILLCELL_X4 FILLER_22_855 ();
 FILLCELL_X4 FILLER_22_862 ();
 FILLCELL_X4 FILLER_22_868 ();
 FILLCELL_X1 FILLER_22_872 ();
 FILLCELL_X16 FILLER_22_882 ();
 FILLCELL_X4 FILLER_22_898 ();
 FILLCELL_X2 FILLER_22_902 ();
 FILLCELL_X1 FILLER_22_904 ();
 FILLCELL_X8 FILLER_22_914 ();
 FILLCELL_X8 FILLER_22_926 ();
 FILLCELL_X8 FILLER_22_943 ();
 FILLCELL_X2 FILLER_22_951 ();
 FILLCELL_X4 FILLER_22_956 ();
 FILLCELL_X8 FILLER_22_964 ();
 FILLCELL_X2 FILLER_22_972 ();
 FILLCELL_X4 FILLER_22_983 ();
 FILLCELL_X4 FILLER_22_997 ();
 FILLCELL_X4 FILLER_22_1011 ();
 FILLCELL_X2 FILLER_22_1015 ();
 FILLCELL_X4 FILLER_22_1020 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X8 FILLER_23_161 ();
 FILLCELL_X8 FILLER_23_819 ();
 FILLCELL_X2 FILLER_23_827 ();
 FILLCELL_X4 FILLER_23_833 ();
 FILLCELL_X4 FILLER_23_840 ();
 FILLCELL_X4 FILLER_23_847 ();
 FILLCELL_X8 FILLER_23_854 ();
 FILLCELL_X1 FILLER_23_862 ();
 FILLCELL_X4 FILLER_23_867 ();
 FILLCELL_X4 FILLER_23_875 ();
 FILLCELL_X4 FILLER_23_882 ();
 FILLCELL_X2 FILLER_23_886 ();
 FILLCELL_X8 FILLER_23_891 ();
 FILLCELL_X8 FILLER_23_903 ();
 FILLCELL_X4 FILLER_23_911 ();
 FILLCELL_X4 FILLER_23_918 ();
 FILLCELL_X4 FILLER_23_932 ();
 FILLCELL_X4 FILLER_23_940 ();
 FILLCELL_X8 FILLER_23_948 ();
 FILLCELL_X2 FILLER_23_956 ();
 FILLCELL_X4 FILLER_23_964 ();
 FILLCELL_X4 FILLER_23_977 ();
 FILLCELL_X4 FILLER_23_984 ();
 FILLCELL_X2 FILLER_23_988 ();
 FILLCELL_X4 FILLER_23_994 ();
 FILLCELL_X2 FILLER_23_998 ();
 FILLCELL_X4 FILLER_23_1019 ();
 FILLCELL_X1 FILLER_23_1023 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X8 FILLER_24_161 ();
 FILLCELL_X4 FILLER_24_819 ();
 FILLCELL_X4 FILLER_24_826 ();
 FILLCELL_X8 FILLER_24_833 ();
 FILLCELL_X8 FILLER_24_851 ();
 FILLCELL_X4 FILLER_24_863 ();
 FILLCELL_X8 FILLER_24_876 ();
 FILLCELL_X2 FILLER_24_884 ();
 FILLCELL_X1 FILLER_24_886 ();
 FILLCELL_X4 FILLER_24_894 ();
 FILLCELL_X1 FILLER_24_898 ();
 FILLCELL_X4 FILLER_24_909 ();
 FILLCELL_X4 FILLER_24_916 ();
 FILLCELL_X4 FILLER_24_922 ();
 FILLCELL_X4 FILLER_24_930 ();
 FILLCELL_X4 FILLER_24_943 ();
 FILLCELL_X8 FILLER_24_950 ();
 FILLCELL_X4 FILLER_24_964 ();
 FILLCELL_X4 FILLER_24_972 ();
 FILLCELL_X4 FILLER_24_979 ();
 FILLCELL_X4 FILLER_24_986 ();
 FILLCELL_X4 FILLER_24_993 ();
 FILLCELL_X16 FILLER_24_999 ();
 FILLCELL_X8 FILLER_24_1015 ();
 FILLCELL_X1 FILLER_24_1023 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X8 FILLER_25_161 ();
 FILLCELL_X4 FILLER_25_819 ();
 FILLCELL_X4 FILLER_25_827 ();
 FILLCELL_X4 FILLER_25_841 ();
 FILLCELL_X4 FILLER_25_854 ();
 FILLCELL_X4 FILLER_25_861 ();
 FILLCELL_X4 FILLER_25_868 ();
 FILLCELL_X1 FILLER_25_872 ();
 FILLCELL_X4 FILLER_25_882 ();
 FILLCELL_X2 FILLER_25_886 ();
 FILLCELL_X4 FILLER_25_890 ();
 FILLCELL_X2 FILLER_25_894 ();
 FILLCELL_X4 FILLER_25_905 ();
 FILLCELL_X4 FILLER_25_912 ();
 FILLCELL_X2 FILLER_25_916 ();
 FILLCELL_X4 FILLER_25_925 ();
 FILLCELL_X4 FILLER_25_931 ();
 FILLCELL_X4 FILLER_25_938 ();
 FILLCELL_X2 FILLER_25_942 ();
 FILLCELL_X1 FILLER_25_944 ();
 FILLCELL_X4 FILLER_25_948 ();
 FILLCELL_X4 FILLER_25_955 ();
 FILLCELL_X8 FILLER_25_968 ();
 FILLCELL_X2 FILLER_25_976 ();
 FILLCELL_X1 FILLER_25_978 ();
 FILLCELL_X4 FILLER_25_988 ();
 FILLCELL_X4 FILLER_25_994 ();
 FILLCELL_X16 FILLER_25_1000 ();
 FILLCELL_X8 FILLER_25_1016 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X8 FILLER_26_161 ();
 FILLCELL_X8 FILLER_26_819 ();
 FILLCELL_X4 FILLER_26_829 ();
 FILLCELL_X4 FILLER_26_836 ();
 FILLCELL_X8 FILLER_26_849 ();
 FILLCELL_X4 FILLER_26_857 ();
 FILLCELL_X4 FILLER_26_863 ();
 FILLCELL_X8 FILLER_26_870 ();
 FILLCELL_X1 FILLER_26_878 ();
 FILLCELL_X8 FILLER_26_882 ();
 FILLCELL_X1 FILLER_26_890 ();
 FILLCELL_X4 FILLER_26_894 ();
 FILLCELL_X8 FILLER_26_908 ();
 FILLCELL_X4 FILLER_26_916 ();
 FILLCELL_X2 FILLER_26_920 ();
 FILLCELL_X1 FILLER_26_922 ();
 FILLCELL_X4 FILLER_26_933 ();
 FILLCELL_X4 FILLER_26_939 ();
 FILLCELL_X16 FILLER_26_945 ();
 FILLCELL_X4 FILLER_26_961 ();
 FILLCELL_X2 FILLER_26_965 ();
 FILLCELL_X4 FILLER_26_972 ();
 FILLCELL_X4 FILLER_26_980 ();
 FILLCELL_X32 FILLER_26_987 ();
 FILLCELL_X4 FILLER_26_1019 ();
 FILLCELL_X1 FILLER_26_1023 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X8 FILLER_27_161 ();
 FILLCELL_X8 FILLER_27_819 ();
 FILLCELL_X4 FILLER_27_827 ();
 FILLCELL_X1 FILLER_27_831 ();
 FILLCELL_X8 FILLER_27_842 ();
 FILLCELL_X4 FILLER_27_850 ();
 FILLCELL_X4 FILLER_27_861 ();
 FILLCELL_X4 FILLER_27_875 ();
 FILLCELL_X4 FILLER_27_883 ();
 FILLCELL_X2 FILLER_27_887 ();
 FILLCELL_X8 FILLER_27_898 ();
 FILLCELL_X4 FILLER_27_906 ();
 FILLCELL_X4 FILLER_27_913 ();
 FILLCELL_X4 FILLER_27_922 ();
 FILLCELL_X4 FILLER_27_929 ();
 FILLCELL_X16 FILLER_27_938 ();
 FILLCELL_X4 FILLER_27_958 ();
 FILLCELL_X4 FILLER_27_967 ();
 FILLCELL_X4 FILLER_27_980 ();
 FILLCELL_X32 FILLER_27_986 ();
 FILLCELL_X4 FILLER_27_1018 ();
 FILLCELL_X2 FILLER_27_1022 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X4 FILLER_28_129 ();
 FILLCELL_X2 FILLER_28_133 ();
 FILLCELL_X1 FILLER_28_135 ();
 FILLCELL_X8 FILLER_28_155 ();
 FILLCELL_X4 FILLER_28_163 ();
 FILLCELL_X2 FILLER_28_167 ();
 FILLCELL_X8 FILLER_28_819 ();
 FILLCELL_X4 FILLER_28_830 ();
 FILLCELL_X16 FILLER_28_837 ();
 FILLCELL_X4 FILLER_28_853 ();
 FILLCELL_X2 FILLER_28_857 ();
 FILLCELL_X8 FILLER_28_869 ();
 FILLCELL_X16 FILLER_28_887 ();
 FILLCELL_X1 FILLER_28_903 ();
 FILLCELL_X4 FILLER_28_907 ();
 FILLCELL_X8 FILLER_28_920 ();
 FILLCELL_X4 FILLER_28_928 ();
 FILLCELL_X8 FILLER_28_949 ();
 FILLCELL_X1 FILLER_28_957 ();
 FILLCELL_X4 FILLER_28_962 ();
 FILLCELL_X4 FILLER_28_970 ();
 FILLCELL_X8 FILLER_28_978 ();
 FILLCELL_X1 FILLER_28_986 ();
 FILLCELL_X32 FILLER_28_991 ();
 FILLCELL_X1 FILLER_28_1023 ();
 FILLCELL_X4 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_8 ();
 FILLCELL_X32 FILLER_29_40 ();
 FILLCELL_X32 FILLER_29_72 ();
 FILLCELL_X32 FILLER_29_104 ();
 FILLCELL_X32 FILLER_29_136 ();
 FILLCELL_X1 FILLER_29_168 ();
 FILLCELL_X4 FILLER_29_819 ();
 FILLCELL_X4 FILLER_29_829 ();
 FILLCELL_X4 FILLER_29_840 ();
 FILLCELL_X1 FILLER_29_844 ();
 FILLCELL_X4 FILLER_29_849 ();
 FILLCELL_X4 FILLER_29_857 ();
 FILLCELL_X8 FILLER_29_864 ();
 FILLCELL_X1 FILLER_29_872 ();
 FILLCELL_X8 FILLER_29_880 ();
 FILLCELL_X1 FILLER_29_888 ();
 FILLCELL_X4 FILLER_29_892 ();
 FILLCELL_X4 FILLER_29_906 ();
 FILLCELL_X2 FILLER_29_910 ();
 FILLCELL_X1 FILLER_29_912 ();
 FILLCELL_X4 FILLER_29_922 ();
 FILLCELL_X1 FILLER_29_926 ();
 FILLCELL_X4 FILLER_29_931 ();
 FILLCELL_X4 FILLER_29_942 ();
 FILLCELL_X4 FILLER_29_951 ();
 FILLCELL_X2 FILLER_29_955 ();
 FILLCELL_X1 FILLER_29_957 ();
 FILLCELL_X4 FILLER_29_961 ();
 FILLCELL_X16 FILLER_29_967 ();
 FILLCELL_X1 FILLER_29_983 ();
 FILLCELL_X16 FILLER_29_1003 ();
 FILLCELL_X4 FILLER_29_1019 ();
 FILLCELL_X1 FILLER_29_1023 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X8 FILLER_30_161 ();
 FILLCELL_X4 FILLER_30_819 ();
 FILLCELL_X2 FILLER_30_823 ();
 FILLCELL_X16 FILLER_30_831 ();
 FILLCELL_X2 FILLER_30_847 ();
 FILLCELL_X4 FILLER_30_858 ();
 FILLCELL_X4 FILLER_30_865 ();
 FILLCELL_X4 FILLER_30_872 ();
 FILLCELL_X2 FILLER_30_876 ();
 FILLCELL_X8 FILLER_30_880 ();
 FILLCELL_X4 FILLER_30_888 ();
 FILLCELL_X4 FILLER_30_896 ();
 FILLCELL_X4 FILLER_30_907 ();
 FILLCELL_X16 FILLER_30_913 ();
 FILLCELL_X4 FILLER_30_929 ();
 FILLCELL_X1 FILLER_30_933 ();
 FILLCELL_X4 FILLER_30_938 ();
 FILLCELL_X4 FILLER_30_946 ();
 FILLCELL_X2 FILLER_30_950 ();
 FILLCELL_X8 FILLER_30_955 ();
 FILLCELL_X1 FILLER_30_963 ();
 FILLCELL_X4 FILLER_30_968 ();
 FILLCELL_X32 FILLER_30_975 ();
 FILLCELL_X16 FILLER_30_1007 ();
 FILLCELL_X1 FILLER_30_1023 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X8 FILLER_31_161 ();
 FILLCELL_X4 FILLER_31_819 ();
 FILLCELL_X16 FILLER_31_826 ();
 FILLCELL_X4 FILLER_31_842 ();
 FILLCELL_X1 FILLER_31_846 ();
 FILLCELL_X4 FILLER_31_851 ();
 FILLCELL_X4 FILLER_31_864 ();
 FILLCELL_X2 FILLER_31_868 ();
 FILLCELL_X4 FILLER_31_873 ();
 FILLCELL_X4 FILLER_31_887 ();
 FILLCELL_X8 FILLER_31_894 ();
 FILLCELL_X4 FILLER_31_905 ();
 FILLCELL_X8 FILLER_31_919 ();
 FILLCELL_X1 FILLER_31_927 ();
 FILLCELL_X8 FILLER_31_931 ();
 FILLCELL_X4 FILLER_31_939 ();
 FILLCELL_X1 FILLER_31_943 ();
 FILLCELL_X4 FILLER_31_947 ();
 FILLCELL_X1 FILLER_31_951 ();
 FILLCELL_X4 FILLER_31_956 ();
 FILLCELL_X4 FILLER_31_969 ();
 FILLCELL_X8 FILLER_31_977 ();
 FILLCELL_X1 FILLER_31_985 ();
 FILLCELL_X32 FILLER_31_990 ();
 FILLCELL_X2 FILLER_31_1022 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X8 FILLER_32_161 ();
 FILLCELL_X8 FILLER_32_819 ();
 FILLCELL_X1 FILLER_32_827 ();
 FILLCELL_X8 FILLER_32_832 ();
 FILLCELL_X1 FILLER_32_840 ();
 FILLCELL_X4 FILLER_32_848 ();
 FILLCELL_X8 FILLER_32_862 ();
 FILLCELL_X4 FILLER_32_870 ();
 FILLCELL_X4 FILLER_32_883 ();
 FILLCELL_X2 FILLER_32_887 ();
 FILLCELL_X4 FILLER_32_898 ();
 FILLCELL_X4 FILLER_32_905 ();
 FILLCELL_X1 FILLER_32_909 ();
 FILLCELL_X4 FILLER_32_920 ();
 FILLCELL_X2 FILLER_32_924 ();
 FILLCELL_X4 FILLER_32_930 ();
 FILLCELL_X4 FILLER_32_938 ();
 FILLCELL_X4 FILLER_32_946 ();
 FILLCELL_X2 FILLER_32_950 ();
 FILLCELL_X4 FILLER_32_961 ();
 FILLCELL_X8 FILLER_32_968 ();
 FILLCELL_X4 FILLER_32_976 ();
 FILLCELL_X2 FILLER_32_980 ();
 FILLCELL_X1 FILLER_32_982 ();
 FILLCELL_X16 FILLER_32_1002 ();
 FILLCELL_X4 FILLER_32_1018 ();
 FILLCELL_X2 FILLER_32_1022 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X8 FILLER_33_161 ();
 FILLCELL_X4 FILLER_33_819 ();
 FILLCELL_X4 FILLER_33_842 ();
 FILLCELL_X2 FILLER_33_846 ();
 FILLCELL_X4 FILLER_33_850 ();
 FILLCELL_X16 FILLER_33_857 ();
 FILLCELL_X8 FILLER_33_873 ();
 FILLCELL_X4 FILLER_33_884 ();
 FILLCELL_X8 FILLER_33_891 ();
 FILLCELL_X1 FILLER_33_899 ();
 FILLCELL_X4 FILLER_33_902 ();
 FILLCELL_X4 FILLER_33_913 ();
 FILLCELL_X4 FILLER_33_919 ();
 FILLCELL_X1 FILLER_33_923 ();
 FILLCELL_X4 FILLER_33_933 ();
 FILLCELL_X8 FILLER_33_946 ();
 FILLCELL_X1 FILLER_33_954 ();
 FILLCELL_X4 FILLER_33_958 ();
 FILLCELL_X4 FILLER_33_966 ();
 FILLCELL_X32 FILLER_33_973 ();
 FILLCELL_X16 FILLER_33_1005 ();
 FILLCELL_X2 FILLER_33_1021 ();
 FILLCELL_X1 FILLER_33_1023 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X8 FILLER_34_161 ();
 FILLCELL_X4 FILLER_34_819 ();
 FILLCELL_X1 FILLER_34_823 ();
 FILLCELL_X8 FILLER_34_843 ();
 FILLCELL_X1 FILLER_34_851 ();
 FILLCELL_X4 FILLER_34_856 ();
 FILLCELL_X4 FILLER_34_870 ();
 FILLCELL_X8 FILLER_34_877 ();
 FILLCELL_X1 FILLER_34_885 ();
 FILLCELL_X8 FILLER_34_895 ();
 FILLCELL_X2 FILLER_34_903 ();
 FILLCELL_X16 FILLER_34_915 ();
 FILLCELL_X4 FILLER_34_931 ();
 FILLCELL_X1 FILLER_34_935 ();
 FILLCELL_X16 FILLER_34_939 ();
 FILLCELL_X4 FILLER_34_959 ();
 FILLCELL_X4 FILLER_34_972 ();
 FILLCELL_X32 FILLER_34_980 ();
 FILLCELL_X4 FILLER_34_1012 ();
 FILLCELL_X1 FILLER_34_1016 ();
 FILLCELL_X4 FILLER_34_1020 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X8 FILLER_35_161 ();
 FILLCELL_X4 FILLER_35_819 ();
 FILLCELL_X2 FILLER_35_823 ();
 FILLCELL_X1 FILLER_35_825 ();
 FILLCELL_X8 FILLER_35_830 ();
 FILLCELL_X4 FILLER_35_838 ();
 FILLCELL_X2 FILLER_35_842 ();
 FILLCELL_X8 FILLER_35_850 ();
 FILLCELL_X4 FILLER_35_858 ();
 FILLCELL_X2 FILLER_35_862 ();
 FILLCELL_X1 FILLER_35_864 ();
 FILLCELL_X4 FILLER_35_872 ();
 FILLCELL_X4 FILLER_35_880 ();
 FILLCELL_X1 FILLER_35_884 ();
 FILLCELL_X4 FILLER_35_895 ();
 FILLCELL_X4 FILLER_35_902 ();
 FILLCELL_X2 FILLER_35_906 ();
 FILLCELL_X4 FILLER_35_911 ();
 FILLCELL_X4 FILLER_35_918 ();
 FILLCELL_X16 FILLER_35_925 ();
 FILLCELL_X2 FILLER_35_941 ();
 FILLCELL_X8 FILLER_35_946 ();
 FILLCELL_X1 FILLER_35_954 ();
 FILLCELL_X4 FILLER_35_958 ();
 FILLCELL_X1 FILLER_35_962 ();
 FILLCELL_X32 FILLER_35_972 ();
 FILLCELL_X16 FILLER_35_1004 ();
 FILLCELL_X4 FILLER_35_1020 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X8 FILLER_36_161 ();
 FILLCELL_X16 FILLER_36_819 ();
 FILLCELL_X8 FILLER_36_839 ();
 FILLCELL_X8 FILLER_36_850 ();
 FILLCELL_X4 FILLER_36_860 ();
 FILLCELL_X8 FILLER_36_874 ();
 FILLCELL_X1 FILLER_36_882 ();
 FILLCELL_X4 FILLER_36_890 ();
 FILLCELL_X8 FILLER_36_904 ();
 FILLCELL_X1 FILLER_36_912 ();
 FILLCELL_X4 FILLER_36_922 ();
 FILLCELL_X4 FILLER_36_929 ();
 FILLCELL_X4 FILLER_36_937 ();
 FILLCELL_X8 FILLER_36_951 ();
 FILLCELL_X1 FILLER_36_959 ();
 FILLCELL_X4 FILLER_36_970 ();
 FILLCELL_X4 FILLER_36_978 ();
 FILLCELL_X32 FILLER_36_986 ();
 FILLCELL_X4 FILLER_36_1018 ();
 FILLCELL_X2 FILLER_36_1022 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X8 FILLER_37_161 ();
 FILLCELL_X4 FILLER_37_819 ();
 FILLCELL_X1 FILLER_37_823 ();
 FILLCELL_X4 FILLER_37_828 ();
 FILLCELL_X4 FILLER_37_839 ();
 FILLCELL_X4 FILLER_37_847 ();
 FILLCELL_X1 FILLER_37_851 ();
 FILLCELL_X4 FILLER_37_856 ();
 FILLCELL_X4 FILLER_37_863 ();
 FILLCELL_X4 FILLER_37_870 ();
 FILLCELL_X8 FILLER_37_876 ();
 FILLCELL_X2 FILLER_37_884 ();
 FILLCELL_X4 FILLER_37_888 ();
 FILLCELL_X8 FILLER_37_894 ();
 FILLCELL_X4 FILLER_37_902 ();
 FILLCELL_X2 FILLER_37_906 ();
 FILLCELL_X4 FILLER_37_917 ();
 FILLCELL_X4 FILLER_37_931 ();
 FILLCELL_X2 FILLER_37_935 ();
 FILLCELL_X1 FILLER_37_937 ();
 FILLCELL_X8 FILLER_37_945 ();
 FILLCELL_X1 FILLER_37_953 ();
 FILLCELL_X4 FILLER_37_961 ();
 FILLCELL_X32 FILLER_37_967 ();
 FILLCELL_X16 FILLER_37_999 ();
 FILLCELL_X8 FILLER_37_1015 ();
 FILLCELL_X1 FILLER_37_1023 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X4 FILLER_38_165 ();
 FILLCELL_X8 FILLER_38_819 ();
 FILLCELL_X2 FILLER_38_827 ();
 FILLCELL_X4 FILLER_38_839 ();
 FILLCELL_X1 FILLER_38_843 ();
 FILLCELL_X4 FILLER_38_853 ();
 FILLCELL_X4 FILLER_38_866 ();
 FILLCELL_X2 FILLER_38_870 ();
 FILLCELL_X1 FILLER_38_872 ();
 FILLCELL_X8 FILLER_38_877 ();
 FILLCELL_X2 FILLER_38_885 ();
 FILLCELL_X8 FILLER_38_890 ();
 FILLCELL_X4 FILLER_38_907 ();
 FILLCELL_X1 FILLER_38_911 ();
 FILLCELL_X4 FILLER_38_919 ();
 FILLCELL_X4 FILLER_38_925 ();
 FILLCELL_X2 FILLER_38_929 ();
 FILLCELL_X1 FILLER_38_931 ();
 FILLCELL_X4 FILLER_38_935 ();
 FILLCELL_X4 FILLER_38_949 ();
 FILLCELL_X4 FILLER_38_955 ();
 FILLCELL_X2 FILLER_38_959 ();
 FILLCELL_X1 FILLER_38_961 ();
 FILLCELL_X4 FILLER_38_966 ();
 FILLCELL_X4 FILLER_38_979 ();
 FILLCELL_X32 FILLER_38_986 ();
 FILLCELL_X4 FILLER_38_1018 ();
 FILLCELL_X2 FILLER_38_1022 ();
 FILLCELL_X4 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_8 ();
 FILLCELL_X32 FILLER_39_40 ();
 FILLCELL_X32 FILLER_39_72 ();
 FILLCELL_X32 FILLER_39_104 ();
 FILLCELL_X8 FILLER_39_136 ();
 FILLCELL_X4 FILLER_39_144 ();
 FILLCELL_X4 FILLER_39_165 ();
 FILLCELL_X4 FILLER_39_819 ();
 FILLCELL_X4 FILLER_39_826 ();
 FILLCELL_X2 FILLER_39_830 ();
 FILLCELL_X4 FILLER_39_838 ();
 FILLCELL_X16 FILLER_39_846 ();
 FILLCELL_X2 FILLER_39_862 ();
 FILLCELL_X4 FILLER_39_867 ();
 FILLCELL_X4 FILLER_39_881 ();
 FILLCELL_X4 FILLER_39_895 ();
 FILLCELL_X2 FILLER_39_899 ();
 FILLCELL_X1 FILLER_39_901 ();
 FILLCELL_X4 FILLER_39_905 ();
 FILLCELL_X4 FILLER_39_919 ();
 FILLCELL_X4 FILLER_39_925 ();
 FILLCELL_X8 FILLER_39_938 ();
 FILLCELL_X4 FILLER_39_946 ();
 FILLCELL_X1 FILLER_39_950 ();
 FILLCELL_X4 FILLER_39_961 ();
 FILLCELL_X4 FILLER_39_968 ();
 FILLCELL_X32 FILLER_39_975 ();
 FILLCELL_X16 FILLER_39_1007 ();
 FILLCELL_X1 FILLER_39_1023 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X32 FILLER_40_97 ();
 FILLCELL_X32 FILLER_40_129 ();
 FILLCELL_X1 FILLER_40_161 ();
 FILLCELL_X4 FILLER_40_165 ();
 FILLCELL_X4 FILLER_40_819 ();
 FILLCELL_X8 FILLER_40_826 ();
 FILLCELL_X4 FILLER_40_834 ();
 FILLCELL_X2 FILLER_40_838 ();
 FILLCELL_X1 FILLER_40_840 ();
 FILLCELL_X8 FILLER_40_844 ();
 FILLCELL_X4 FILLER_40_852 ();
 FILLCELL_X2 FILLER_40_856 ();
 FILLCELL_X4 FILLER_40_861 ();
 FILLCELL_X4 FILLER_40_867 ();
 FILLCELL_X1 FILLER_40_871 ();
 FILLCELL_X4 FILLER_40_874 ();
 FILLCELL_X2 FILLER_40_878 ();
 FILLCELL_X1 FILLER_40_880 ();
 FILLCELL_X4 FILLER_40_888 ();
 FILLCELL_X8 FILLER_40_894 ();
 FILLCELL_X4 FILLER_40_902 ();
 FILLCELL_X4 FILLER_40_909 ();
 FILLCELL_X8 FILLER_40_916 ();
 FILLCELL_X1 FILLER_40_924 ();
 FILLCELL_X4 FILLER_40_928 ();
 FILLCELL_X16 FILLER_40_942 ();
 FILLCELL_X2 FILLER_40_958 ();
 FILLCELL_X4 FILLER_40_969 ();
 FILLCELL_X4 FILLER_40_977 ();
 FILLCELL_X4 FILLER_40_984 ();
 FILLCELL_X32 FILLER_40_991 ();
 FILLCELL_X1 FILLER_40_1023 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X32 FILLER_41_97 ();
 FILLCELL_X16 FILLER_41_129 ();
 FILLCELL_X8 FILLER_41_145 ();
 FILLCELL_X4 FILLER_41_153 ();
 FILLCELL_X2 FILLER_41_157 ();
 FILLCELL_X1 FILLER_41_159 ();
 FILLCELL_X4 FILLER_41_165 ();
 FILLCELL_X4 FILLER_41_819 ();
 FILLCELL_X4 FILLER_41_827 ();
 FILLCELL_X4 FILLER_41_835 ();
 FILLCELL_X4 FILLER_41_842 ();
 FILLCELL_X2 FILLER_41_846 ();
 FILLCELL_X1 FILLER_41_848 ();
 FILLCELL_X4 FILLER_41_856 ();
 FILLCELL_X4 FILLER_41_863 ();
 FILLCELL_X1 FILLER_41_867 ();
 FILLCELL_X8 FILLER_41_878 ();
 FILLCELL_X1 FILLER_41_886 ();
 FILLCELL_X4 FILLER_41_890 ();
 FILLCELL_X4 FILLER_41_897 ();
 FILLCELL_X2 FILLER_41_901 ();
 FILLCELL_X4 FILLER_41_906 ();
 FILLCELL_X4 FILLER_41_919 ();
 FILLCELL_X16 FILLER_41_930 ();
 FILLCELL_X1 FILLER_41_946 ();
 FILLCELL_X8 FILLER_41_951 ();
 FILLCELL_X2 FILLER_41_959 ();
 FILLCELL_X1 FILLER_41_961 ();
 FILLCELL_X4 FILLER_41_965 ();
 FILLCELL_X4 FILLER_41_973 ();
 FILLCELL_X4 FILLER_41_986 ();
 FILLCELL_X16 FILLER_41_994 ();
 FILLCELL_X8 FILLER_41_1010 ();
 FILLCELL_X4 FILLER_41_1018 ();
 FILLCELL_X2 FILLER_41_1022 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X32 FILLER_42_65 ();
 FILLCELL_X32 FILLER_42_97 ();
 FILLCELL_X16 FILLER_42_129 ();
 FILLCELL_X8 FILLER_42_145 ();
 FILLCELL_X2 FILLER_42_153 ();
 FILLCELL_X4 FILLER_42_158 ();
 FILLCELL_X4 FILLER_42_165 ();
 FILLCELL_X8 FILLER_42_819 ();
 FILLCELL_X1 FILLER_42_827 ();
 FILLCELL_X4 FILLER_42_837 ();
 FILLCELL_X4 FILLER_42_845 ();
 FILLCELL_X4 FILLER_42_852 ();
 FILLCELL_X2 FILLER_42_856 ();
 FILLCELL_X1 FILLER_42_858 ();
 FILLCELL_X16 FILLER_42_865 ();
 FILLCELL_X4 FILLER_42_891 ();
 FILLCELL_X4 FILLER_42_904 ();
 FILLCELL_X2 FILLER_42_908 ();
 FILLCELL_X1 FILLER_42_910 ();
 FILLCELL_X8 FILLER_42_921 ();
 FILLCELL_X4 FILLER_42_929 ();
 FILLCELL_X2 FILLER_42_933 ();
 FILLCELL_X1 FILLER_42_935 ();
 FILLCELL_X4 FILLER_42_940 ();
 FILLCELL_X2 FILLER_42_944 ();
 FILLCELL_X4 FILLER_42_956 ();
 FILLCELL_X8 FILLER_42_963 ();
 FILLCELL_X2 FILLER_42_971 ();
 FILLCELL_X4 FILLER_42_982 ();
 FILLCELL_X32 FILLER_42_990 ();
 FILLCELL_X2 FILLER_42_1022 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X32 FILLER_43_65 ();
 FILLCELL_X32 FILLER_43_97 ();
 FILLCELL_X32 FILLER_43_129 ();
 FILLCELL_X1 FILLER_43_161 ();
 FILLCELL_X4 FILLER_43_165 ();
 FILLCELL_X4 FILLER_43_819 ();
 FILLCELL_X4 FILLER_43_826 ();
 FILLCELL_X2 FILLER_43_830 ();
 FILLCELL_X1 FILLER_43_832 ();
 FILLCELL_X4 FILLER_43_842 ();
 FILLCELL_X2 FILLER_43_846 ();
 FILLCELL_X4 FILLER_43_851 ();
 FILLCELL_X4 FILLER_43_862 ();
 FILLCELL_X8 FILLER_43_872 ();
 FILLCELL_X4 FILLER_43_880 ();
 FILLCELL_X4 FILLER_43_893 ();
 FILLCELL_X2 FILLER_43_897 ();
 FILLCELL_X1 FILLER_43_899 ();
 FILLCELL_X8 FILLER_43_903 ();
 FILLCELL_X1 FILLER_43_911 ();
 FILLCELL_X4 FILLER_43_921 ();
 FILLCELL_X8 FILLER_43_928 ();
 FILLCELL_X1 FILLER_43_936 ();
 FILLCELL_X8 FILLER_43_944 ();
 FILLCELL_X4 FILLER_43_952 ();
 FILLCELL_X2 FILLER_43_956 ();
 FILLCELL_X1 FILLER_43_958 ();
 FILLCELL_X32 FILLER_43_963 ();
 FILLCELL_X16 FILLER_43_995 ();
 FILLCELL_X8 FILLER_43_1011 ();
 FILLCELL_X4 FILLER_43_1019 ();
 FILLCELL_X1 FILLER_43_1023 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X32 FILLER_44_33 ();
 FILLCELL_X32 FILLER_44_65 ();
 FILLCELL_X32 FILLER_44_97 ();
 FILLCELL_X32 FILLER_44_129 ();
 FILLCELL_X8 FILLER_44_161 ();
 FILLCELL_X4 FILLER_44_819 ();
 FILLCELL_X8 FILLER_44_826 ();
 FILLCELL_X2 FILLER_44_834 ();
 FILLCELL_X1 FILLER_44_836 ();
 FILLCELL_X4 FILLER_44_841 ();
 FILLCELL_X4 FILLER_44_855 ();
 FILLCELL_X16 FILLER_44_869 ();
 FILLCELL_X8 FILLER_44_885 ();
 FILLCELL_X4 FILLER_44_893 ();
 FILLCELL_X4 FILLER_44_900 ();
 FILLCELL_X4 FILLER_44_911 ();
 FILLCELL_X4 FILLER_44_925 ();
 FILLCELL_X4 FILLER_44_932 ();
 FILLCELL_X4 FILLER_44_946 ();
 FILLCELL_X4 FILLER_44_953 ();
 FILLCELL_X4 FILLER_44_959 ();
 FILLCELL_X4 FILLER_44_966 ();
 FILLCELL_X32 FILLER_44_989 ();
 FILLCELL_X2 FILLER_44_1021 ();
 FILLCELL_X1 FILLER_44_1023 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X32 FILLER_45_33 ();
 FILLCELL_X32 FILLER_45_65 ();
 FILLCELL_X32 FILLER_45_97 ();
 FILLCELL_X32 FILLER_45_129 ();
 FILLCELL_X8 FILLER_45_161 ();
 FILLCELL_X4 FILLER_45_819 ();
 FILLCELL_X16 FILLER_45_828 ();
 FILLCELL_X8 FILLER_45_844 ();
 FILLCELL_X2 FILLER_45_852 ();
 FILLCELL_X8 FILLER_45_856 ();
 FILLCELL_X2 FILLER_45_864 ();
 FILLCELL_X1 FILLER_45_866 ();
 FILLCELL_X4 FILLER_45_877 ();
 FILLCELL_X4 FILLER_45_884 ();
 FILLCELL_X4 FILLER_45_891 ();
 FILLCELL_X1 FILLER_45_895 ();
 FILLCELL_X4 FILLER_45_905 ();
 FILLCELL_X16 FILLER_45_911 ();
 FILLCELL_X4 FILLER_45_930 ();
 FILLCELL_X4 FILLER_45_943 ();
 FILLCELL_X4 FILLER_45_951 ();
 FILLCELL_X4 FILLER_45_962 ();
 FILLCELL_X4 FILLER_45_976 ();
 FILLCELL_X4 FILLER_45_984 ();
 FILLCELL_X16 FILLER_45_990 ();
 FILLCELL_X8 FILLER_45_1006 ();
 FILLCELL_X2 FILLER_45_1014 ();
 FILLCELL_X1 FILLER_45_1016 ();
 FILLCELL_X4 FILLER_45_1020 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X32 FILLER_46_33 ();
 FILLCELL_X32 FILLER_46_65 ();
 FILLCELL_X32 FILLER_46_97 ();
 FILLCELL_X32 FILLER_46_129 ();
 FILLCELL_X8 FILLER_46_161 ();
 FILLCELL_X8 FILLER_46_819 ();
 FILLCELL_X4 FILLER_46_827 ();
 FILLCELL_X2 FILLER_46_831 ();
 FILLCELL_X4 FILLER_46_837 ();
 FILLCELL_X4 FILLER_46_844 ();
 FILLCELL_X4 FILLER_46_851 ();
 FILLCELL_X4 FILLER_46_858 ();
 FILLCELL_X4 FILLER_46_869 ();
 FILLCELL_X2 FILLER_46_873 ();
 FILLCELL_X1 FILLER_46_875 ();
 FILLCELL_X8 FILLER_46_885 ();
 FILLCELL_X4 FILLER_46_903 ();
 FILLCELL_X16 FILLER_46_917 ();
 FILLCELL_X4 FILLER_46_937 ();
 FILLCELL_X16 FILLER_46_944 ();
 FILLCELL_X8 FILLER_46_960 ();
 FILLCELL_X8 FILLER_46_978 ();
 FILLCELL_X4 FILLER_46_986 ();
 FILLCELL_X4 FILLER_46_994 ();
 FILLCELL_X4 FILLER_46_1001 ();
 FILLCELL_X16 FILLER_46_1008 ();
 FILLCELL_X32 FILLER_47_1 ();
 FILLCELL_X32 FILLER_47_33 ();
 FILLCELL_X32 FILLER_47_65 ();
 FILLCELL_X32 FILLER_47_97 ();
 FILLCELL_X2 FILLER_47_129 ();
 FILLCELL_X32 FILLER_47_134 ();
 FILLCELL_X2 FILLER_47_166 ();
 FILLCELL_X1 FILLER_47_168 ();
 FILLCELL_X4 FILLER_47_819 ();
 FILLCELL_X4 FILLER_47_827 ();
 FILLCELL_X4 FILLER_47_840 ();
 FILLCELL_X8 FILLER_47_848 ();
 FILLCELL_X4 FILLER_47_856 ();
 FILLCELL_X4 FILLER_47_862 ();
 FILLCELL_X4 FILLER_47_869 ();
 FILLCELL_X4 FILLER_47_876 ();
 FILLCELL_X4 FILLER_47_889 ();
 FILLCELL_X4 FILLER_47_900 ();
 FILLCELL_X16 FILLER_47_907 ();
 FILLCELL_X4 FILLER_47_925 ();
 FILLCELL_X8 FILLER_47_938 ();
 FILLCELL_X4 FILLER_47_946 ();
 FILLCELL_X4 FILLER_47_954 ();
 FILLCELL_X16 FILLER_47_961 ();
 FILLCELL_X4 FILLER_47_980 ();
 FILLCELL_X4 FILLER_47_988 ();
 FILLCELL_X4 FILLER_47_1001 ();
 FILLCELL_X8 FILLER_47_1009 ();
 FILLCELL_X4 FILLER_47_1017 ();
 FILLCELL_X2 FILLER_47_1021 ();
 FILLCELL_X1 FILLER_47_1023 ();
 FILLCELL_X32 FILLER_48_1 ();
 FILLCELL_X32 FILLER_48_33 ();
 FILLCELL_X32 FILLER_48_65 ();
 FILLCELL_X16 FILLER_48_97 ();
 FILLCELL_X4 FILLER_48_113 ();
 FILLCELL_X1 FILLER_48_117 ();
 FILLCELL_X4 FILLER_48_135 ();
 FILLCELL_X4 FILLER_48_144 ();
 FILLCELL_X16 FILLER_48_151 ();
 FILLCELL_X2 FILLER_48_167 ();
 FILLCELL_X4 FILLER_48_819 ();
 FILLCELL_X4 FILLER_48_828 ();
 FILLCELL_X8 FILLER_48_841 ();
 FILLCELL_X4 FILLER_48_849 ();
 FILLCELL_X2 FILLER_48_853 ();
 FILLCELL_X8 FILLER_48_865 ();
 FILLCELL_X8 FILLER_48_875 ();
 FILLCELL_X1 FILLER_48_883 ();
 FILLCELL_X8 FILLER_48_887 ();
 FILLCELL_X8 FILLER_48_904 ();
 FILLCELL_X2 FILLER_48_912 ();
 FILLCELL_X4 FILLER_48_918 ();
 FILLCELL_X4 FILLER_48_932 ();
 FILLCELL_X4 FILLER_48_939 ();
 FILLCELL_X4 FILLER_48_946 ();
 FILLCELL_X8 FILLER_48_954 ();
 FILLCELL_X2 FILLER_48_962 ();
 FILLCELL_X4 FILLER_48_968 ();
 FILLCELL_X2 FILLER_48_972 ();
 FILLCELL_X4 FILLER_48_978 ();
 FILLCELL_X4 FILLER_48_985 ();
 FILLCELL_X16 FILLER_48_998 ();
 FILLCELL_X8 FILLER_48_1014 ();
 FILLCELL_X2 FILLER_48_1022 ();
 FILLCELL_X32 FILLER_49_1 ();
 FILLCELL_X32 FILLER_49_33 ();
 FILLCELL_X32 FILLER_49_65 ();
 FILLCELL_X8 FILLER_49_97 ();
 FILLCELL_X4 FILLER_49_105 ();
 FILLCELL_X2 FILLER_49_109 ();
 FILLCELL_X4 FILLER_49_114 ();
 FILLCELL_X4 FILLER_49_121 ();
 FILLCELL_X4 FILLER_49_129 ();
 FILLCELL_X4 FILLER_49_137 ();
 FILLCELL_X2 FILLER_49_141 ();
 FILLCELL_X1 FILLER_49_143 ();
 FILLCELL_X4 FILLER_49_147 ();
 FILLCELL_X8 FILLER_49_154 ();
 FILLCELL_X4 FILLER_49_162 ();
 FILLCELL_X2 FILLER_49_166 ();
 FILLCELL_X1 FILLER_49_168 ();
 FILLCELL_X8 FILLER_49_819 ();
 FILLCELL_X4 FILLER_49_827 ();
 FILLCELL_X4 FILLER_49_836 ();
 FILLCELL_X16 FILLER_49_843 ();
 FILLCELL_X1 FILLER_49_859 ();
 FILLCELL_X4 FILLER_49_863 ();
 FILLCELL_X2 FILLER_49_867 ();
 FILLCELL_X8 FILLER_49_879 ();
 FILLCELL_X4 FILLER_49_894 ();
 FILLCELL_X8 FILLER_49_908 ();
 FILLCELL_X1 FILLER_49_916 ();
 FILLCELL_X8 FILLER_49_924 ();
 FILLCELL_X4 FILLER_49_932 ();
 FILLCELL_X2 FILLER_49_936 ();
 FILLCELL_X1 FILLER_49_938 ();
 FILLCELL_X4 FILLER_49_942 ();
 FILLCELL_X1 FILLER_49_946 ();
 FILLCELL_X8 FILLER_49_956 ();
 FILLCELL_X4 FILLER_49_964 ();
 FILLCELL_X1 FILLER_49_968 ();
 FILLCELL_X8 FILLER_49_972 ();
 FILLCELL_X1 FILLER_49_980 ();
 FILLCELL_X8 FILLER_49_991 ();
 FILLCELL_X2 FILLER_49_999 ();
 FILLCELL_X4 FILLER_49_1020 ();
 FILLCELL_X4 FILLER_50_1 ();
 FILLCELL_X32 FILLER_50_9 ();
 FILLCELL_X32 FILLER_50_41 ();
 FILLCELL_X32 FILLER_50_73 ();
 FILLCELL_X8 FILLER_50_105 ();
 FILLCELL_X1 FILLER_50_113 ();
 FILLCELL_X4 FILLER_50_117 ();
 FILLCELL_X4 FILLER_50_140 ();
 FILLCELL_X2 FILLER_50_144 ();
 FILLCELL_X4 FILLER_50_150 ();
 FILLCELL_X4 FILLER_50_157 ();
 FILLCELL_X4 FILLER_50_163 ();
 FILLCELL_X2 FILLER_50_167 ();
 FILLCELL_X8 FILLER_50_819 ();
 FILLCELL_X4 FILLER_50_827 ();
 FILLCELL_X4 FILLER_50_835 ();
 FILLCELL_X4 FILLER_50_846 ();
 FILLCELL_X4 FILLER_50_854 ();
 FILLCELL_X4 FILLER_50_867 ();
 FILLCELL_X4 FILLER_50_874 ();
 FILLCELL_X8 FILLER_50_881 ();
 FILLCELL_X2 FILLER_50_889 ();
 FILLCELL_X1 FILLER_50_891 ();
 FILLCELL_X4 FILLER_50_895 ();
 FILLCELL_X8 FILLER_50_901 ();
 FILLCELL_X1 FILLER_50_909 ();
 FILLCELL_X4 FILLER_50_913 ();
 FILLCELL_X1 FILLER_50_917 ();
 FILLCELL_X4 FILLER_50_928 ();
 FILLCELL_X2 FILLER_50_932 ();
 FILLCELL_X4 FILLER_50_938 ();
 FILLCELL_X4 FILLER_50_951 ();
 FILLCELL_X2 FILLER_50_955 ();
 FILLCELL_X4 FILLER_50_961 ();
 FILLCELL_X4 FILLER_50_974 ();
 FILLCELL_X2 FILLER_50_978 ();
 FILLCELL_X4 FILLER_50_990 ();
 FILLCELL_X2 FILLER_50_994 ();
 FILLCELL_X1 FILLER_50_996 ();
 FILLCELL_X16 FILLER_50_1001 ();
 FILLCELL_X4 FILLER_50_1017 ();
 FILLCELL_X2 FILLER_50_1021 ();
 FILLCELL_X1 FILLER_50_1023 ();
 FILLCELL_X32 FILLER_51_1 ();
 FILLCELL_X32 FILLER_51_33 ();
 FILLCELL_X16 FILLER_51_65 ();
 FILLCELL_X4 FILLER_51_81 ();
 FILLCELL_X2 FILLER_51_85 ();
 FILLCELL_X4 FILLER_51_90 ();
 FILLCELL_X2 FILLER_51_94 ();
 FILLCELL_X4 FILLER_51_100 ();
 FILLCELL_X4 FILLER_51_108 ();
 FILLCELL_X1 FILLER_51_112 ();
 FILLCELL_X4 FILLER_51_117 ();
 FILLCELL_X8 FILLER_51_125 ();
 FILLCELL_X1 FILLER_51_133 ();
 FILLCELL_X4 FILLER_51_137 ();
 FILLCELL_X8 FILLER_51_160 ();
 FILLCELL_X1 FILLER_51_168 ();
 FILLCELL_X4 FILLER_51_819 ();
 FILLCELL_X2 FILLER_51_823 ();
 FILLCELL_X4 FILLER_51_829 ();
 FILLCELL_X4 FILLER_51_843 ();
 FILLCELL_X4 FILLER_51_856 ();
 FILLCELL_X4 FILLER_51_869 ();
 FILLCELL_X8 FILLER_51_882 ();
 FILLCELL_X4 FILLER_51_900 ();
 FILLCELL_X4 FILLER_51_908 ();
 FILLCELL_X8 FILLER_51_915 ();
 FILLCELL_X2 FILLER_51_923 ();
 FILLCELL_X1 FILLER_51_925 ();
 FILLCELL_X8 FILLER_51_928 ();
 FILLCELL_X4 FILLER_51_936 ();
 FILLCELL_X8 FILLER_51_944 ();
 FILLCELL_X4 FILLER_51_952 ();
 FILLCELL_X2 FILLER_51_956 ();
 FILLCELL_X4 FILLER_51_961 ();
 FILLCELL_X8 FILLER_51_968 ();
 FILLCELL_X2 FILLER_51_976 ();
 FILLCELL_X4 FILLER_51_985 ();
 FILLCELL_X2 FILLER_51_989 ();
 FILLCELL_X1 FILLER_51_991 ();
 FILLCELL_X16 FILLER_51_994 ();
 FILLCELL_X8 FILLER_51_1010 ();
 FILLCELL_X4 FILLER_51_1018 ();
 FILLCELL_X2 FILLER_51_1022 ();
 FILLCELL_X32 FILLER_52_1 ();
 FILLCELL_X32 FILLER_52_33 ();
 FILLCELL_X8 FILLER_52_65 ();
 FILLCELL_X4 FILLER_52_73 ();
 FILLCELL_X2 FILLER_52_77 ();
 FILLCELL_X1 FILLER_52_79 ();
 FILLCELL_X4 FILLER_52_97 ();
 FILLCELL_X2 FILLER_52_101 ();
 FILLCELL_X4 FILLER_52_120 ();
 FILLCELL_X4 FILLER_52_127 ();
 FILLCELL_X4 FILLER_52_134 ();
 FILLCELL_X8 FILLER_52_141 ();
 FILLCELL_X4 FILLER_52_152 ();
 FILLCELL_X4 FILLER_52_165 ();
 FILLCELL_X8 FILLER_52_819 ();
 FILLCELL_X4 FILLER_52_827 ();
 FILLCELL_X2 FILLER_52_831 ();
 FILLCELL_X4 FILLER_52_837 ();
 FILLCELL_X4 FILLER_52_851 ();
 FILLCELL_X8 FILLER_52_858 ();
 FILLCELL_X2 FILLER_52_866 ();
 FILLCELL_X1 FILLER_52_868 ();
 FILLCELL_X4 FILLER_52_872 ();
 FILLCELL_X8 FILLER_52_886 ();
 FILLCELL_X1 FILLER_52_894 ();
 FILLCELL_X4 FILLER_52_898 ();
 FILLCELL_X8 FILLER_52_905 ();
 FILLCELL_X2 FILLER_52_913 ();
 FILLCELL_X4 FILLER_52_924 ();
 FILLCELL_X1 FILLER_52_928 ();
 FILLCELL_X4 FILLER_52_936 ();
 FILLCELL_X4 FILLER_52_950 ();
 FILLCELL_X4 FILLER_52_957 ();
 FILLCELL_X2 FILLER_52_961 ();
 FILLCELL_X1 FILLER_52_963 ();
 FILLCELL_X4 FILLER_52_968 ();
 FILLCELL_X4 FILLER_52_981 ();
 FILLCELL_X2 FILLER_52_985 ();
 FILLCELL_X4 FILLER_52_990 ();
 FILLCELL_X4 FILLER_52_998 ();
 FILLCELL_X4 FILLER_52_1005 ();
 FILLCELL_X8 FILLER_52_1012 ();
 FILLCELL_X4 FILLER_52_1020 ();
 FILLCELL_X32 FILLER_53_1 ();
 FILLCELL_X16 FILLER_53_33 ();
 FILLCELL_X8 FILLER_53_49 ();
 FILLCELL_X4 FILLER_53_57 ();
 FILLCELL_X2 FILLER_53_61 ();
 FILLCELL_X1 FILLER_53_63 ();
 FILLCELL_X4 FILLER_53_67 ();
 FILLCELL_X4 FILLER_53_74 ();
 FILLCELL_X4 FILLER_53_81 ();
 FILLCELL_X4 FILLER_53_90 ();
 FILLCELL_X4 FILLER_53_99 ();
 FILLCELL_X4 FILLER_53_106 ();
 FILLCELL_X4 FILLER_53_114 ();
 FILLCELL_X1 FILLER_53_118 ();
 FILLCELL_X4 FILLER_53_125 ();
 FILLCELL_X4 FILLER_53_134 ();
 FILLCELL_X1 FILLER_53_138 ();
 FILLCELL_X4 FILLER_53_142 ();
 FILLCELL_X8 FILLER_53_151 ();
 FILLCELL_X1 FILLER_53_159 ();
 FILLCELL_X4 FILLER_53_165 ();
 FILLCELL_X16 FILLER_53_819 ();
 FILLCELL_X8 FILLER_53_835 ();
 FILLCELL_X1 FILLER_53_843 ();
 FILLCELL_X16 FILLER_53_846 ();
 FILLCELL_X4 FILLER_53_862 ();
 FILLCELL_X4 FILLER_53_869 ();
 FILLCELL_X2 FILLER_53_873 ();
 FILLCELL_X1 FILLER_53_875 ();
 FILLCELL_X4 FILLER_53_883 ();
 FILLCELL_X8 FILLER_53_890 ();
 FILLCELL_X2 FILLER_53_898 ();
 FILLCELL_X8 FILLER_53_910 ();
 FILLCELL_X4 FILLER_53_927 ();
 FILLCELL_X4 FILLER_53_934 ();
 FILLCELL_X1 FILLER_53_938 ();
 FILLCELL_X4 FILLER_53_949 ();
 FILLCELL_X4 FILLER_53_955 ();
 FILLCELL_X4 FILLER_53_961 ();
 FILLCELL_X4 FILLER_53_969 ();
 FILLCELL_X4 FILLER_53_976 ();
 FILLCELL_X2 FILLER_53_980 ();
 FILLCELL_X1 FILLER_53_982 ();
 FILLCELL_X4 FILLER_53_987 ();
 FILLCELL_X4 FILLER_53_1000 ();
 FILLCELL_X8 FILLER_53_1013 ();
 FILLCELL_X2 FILLER_53_1021 ();
 FILLCELL_X1 FILLER_53_1023 ();
 FILLCELL_X32 FILLER_54_1 ();
 FILLCELL_X32 FILLER_54_33 ();
 FILLCELL_X8 FILLER_54_65 ();
 FILLCELL_X1 FILLER_54_73 ();
 FILLCELL_X4 FILLER_54_93 ();
 FILLCELL_X4 FILLER_54_103 ();
 FILLCELL_X4 FILLER_54_112 ();
 FILLCELL_X8 FILLER_54_121 ();
 FILLCELL_X1 FILLER_54_129 ();
 FILLCELL_X4 FILLER_54_135 ();
 FILLCELL_X4 FILLER_54_144 ();
 FILLCELL_X4 FILLER_54_152 ();
 FILLCELL_X4 FILLER_54_158 ();
 FILLCELL_X4 FILLER_54_165 ();
 FILLCELL_X4 FILLER_54_819 ();
 FILLCELL_X1 FILLER_54_823 ();
 FILLCELL_X4 FILLER_54_827 ();
 FILLCELL_X4 FILLER_54_835 ();
 FILLCELL_X1 FILLER_54_839 ();
 FILLCELL_X4 FILLER_54_844 ();
 FILLCELL_X16 FILLER_54_851 ();
 FILLCELL_X2 FILLER_54_867 ();
 FILLCELL_X4 FILLER_54_878 ();
 FILLCELL_X4 FILLER_54_891 ();
 FILLCELL_X8 FILLER_54_902 ();
 FILLCELL_X4 FILLER_54_917 ();
 FILLCELL_X4 FILLER_54_924 ();
 FILLCELL_X4 FILLER_54_931 ();
 FILLCELL_X8 FILLER_54_938 ();
 FILLCELL_X4 FILLER_54_946 ();
 FILLCELL_X2 FILLER_54_950 ();
 FILLCELL_X1 FILLER_54_952 ();
 FILLCELL_X4 FILLER_54_960 ();
 FILLCELL_X8 FILLER_54_974 ();
 FILLCELL_X4 FILLER_54_982 ();
 FILLCELL_X2 FILLER_54_986 ();
 FILLCELL_X1 FILLER_54_988 ();
 FILLCELL_X4 FILLER_54_993 ();
 FILLCELL_X16 FILLER_54_1001 ();
 FILLCELL_X4 FILLER_54_1017 ();
 FILLCELL_X2 FILLER_54_1021 ();
 FILLCELL_X1 FILLER_54_1023 ();
 FILLCELL_X32 FILLER_55_1 ();
 FILLCELL_X32 FILLER_55_33 ();
 FILLCELL_X4 FILLER_55_65 ();
 FILLCELL_X2 FILLER_55_69 ();
 FILLCELL_X4 FILLER_55_74 ();
 FILLCELL_X4 FILLER_55_81 ();
 FILLCELL_X4 FILLER_55_88 ();
 FILLCELL_X4 FILLER_55_97 ();
 FILLCELL_X8 FILLER_55_108 ();
 FILLCELL_X2 FILLER_55_116 ();
 FILLCELL_X4 FILLER_55_120 ();
 FILLCELL_X4 FILLER_55_131 ();
 FILLCELL_X2 FILLER_55_135 ();
 FILLCELL_X4 FILLER_55_154 ();
 FILLCELL_X2 FILLER_55_158 ();
 FILLCELL_X4 FILLER_55_163 ();
 FILLCELL_X2 FILLER_55_167 ();
 FILLCELL_X4 FILLER_55_819 ();
 FILLCELL_X1 FILLER_55_823 ();
 FILLCELL_X4 FILLER_55_828 ();
 FILLCELL_X4 FILLER_55_841 ();
 FILLCELL_X4 FILLER_55_854 ();
 FILLCELL_X4 FILLER_55_861 ();
 FILLCELL_X8 FILLER_55_868 ();
 FILLCELL_X2 FILLER_55_876 ();
 FILLCELL_X1 FILLER_55_878 ();
 FILLCELL_X4 FILLER_55_881 ();
 FILLCELL_X4 FILLER_55_887 ();
 FILLCELL_X2 FILLER_55_891 ();
 FILLCELL_X1 FILLER_55_893 ();
 FILLCELL_X4 FILLER_55_898 ();
 FILLCELL_X8 FILLER_55_912 ();
 FILLCELL_X1 FILLER_55_920 ();
 FILLCELL_X4 FILLER_55_931 ();
 FILLCELL_X4 FILLER_55_944 ();
 FILLCELL_X2 FILLER_55_948 ();
 FILLCELL_X1 FILLER_55_950 ();
 FILLCELL_X16 FILLER_55_961 ();
 FILLCELL_X2 FILLER_55_977 ();
 FILLCELL_X32 FILLER_55_982 ();
 FILLCELL_X2 FILLER_55_1014 ();
 FILLCELL_X1 FILLER_55_1016 ();
 FILLCELL_X4 FILLER_55_1020 ();
 FILLCELL_X32 FILLER_56_1 ();
 FILLCELL_X32 FILLER_56_33 ();
 FILLCELL_X16 FILLER_56_65 ();
 FILLCELL_X4 FILLER_56_85 ();
 FILLCELL_X8 FILLER_56_94 ();
 FILLCELL_X2 FILLER_56_102 ();
 FILLCELL_X4 FILLER_56_110 ();
 FILLCELL_X4 FILLER_56_118 ();
 FILLCELL_X1 FILLER_56_122 ();
 FILLCELL_X4 FILLER_56_125 ();
 FILLCELL_X4 FILLER_56_132 ();
 FILLCELL_X4 FILLER_56_141 ();
 FILLCELL_X4 FILLER_56_150 ();
 FILLCELL_X1 FILLER_56_154 ();
 FILLCELL_X4 FILLER_56_158 ();
 FILLCELL_X4 FILLER_56_165 ();
 FILLCELL_X16 FILLER_56_819 ();
 FILLCELL_X8 FILLER_56_835 ();
 FILLCELL_X8 FILLER_56_847 ();
 FILLCELL_X4 FILLER_56_855 ();
 FILLCELL_X2 FILLER_56_859 ();
 FILLCELL_X1 FILLER_56_861 ();
 FILLCELL_X4 FILLER_56_872 ();
 FILLCELL_X8 FILLER_56_886 ();
 FILLCELL_X2 FILLER_56_894 ();
 FILLCELL_X1 FILLER_56_896 ();
 FILLCELL_X8 FILLER_56_899 ();
 FILLCELL_X4 FILLER_56_907 ();
 FILLCELL_X2 FILLER_56_911 ();
 FILLCELL_X4 FILLER_56_915 ();
 FILLCELL_X8 FILLER_56_922 ();
 FILLCELL_X4 FILLER_56_930 ();
 FILLCELL_X1 FILLER_56_934 ();
 FILLCELL_X4 FILLER_56_938 ();
 FILLCELL_X16 FILLER_56_945 ();
 FILLCELL_X4 FILLER_56_965 ();
 FILLCELL_X4 FILLER_56_972 ();
 FILLCELL_X4 FILLER_56_979 ();
 FILLCELL_X1 FILLER_56_983 ();
 FILLCELL_X4 FILLER_56_994 ();
 FILLCELL_X4 FILLER_56_1002 ();
 FILLCELL_X8 FILLER_56_1010 ();
 FILLCELL_X4 FILLER_56_1018 ();
 FILLCELL_X2 FILLER_56_1022 ();
 FILLCELL_X32 FILLER_57_1 ();
 FILLCELL_X32 FILLER_57_33 ();
 FILLCELL_X4 FILLER_57_65 ();
 FILLCELL_X1 FILLER_57_69 ();
 FILLCELL_X4 FILLER_57_73 ();
 FILLCELL_X4 FILLER_57_94 ();
 FILLCELL_X4 FILLER_57_104 ();
 FILLCELL_X2 FILLER_57_108 ();
 FILLCELL_X4 FILLER_57_114 ();
 FILLCELL_X4 FILLER_57_121 ();
 FILLCELL_X2 FILLER_57_125 ();
 FILLCELL_X4 FILLER_57_129 ();
 FILLCELL_X4 FILLER_57_136 ();
 FILLCELL_X4 FILLER_57_143 ();
 FILLCELL_X4 FILLER_57_153 ();
 FILLCELL_X2 FILLER_57_157 ();
 FILLCELL_X1 FILLER_57_159 ();
 FILLCELL_X4 FILLER_57_165 ();
 FILLCELL_X16 FILLER_57_819 ();
 FILLCELL_X2 FILLER_57_835 ();
 FILLCELL_X4 FILLER_57_841 ();
 FILLCELL_X8 FILLER_57_852 ();
 FILLCELL_X4 FILLER_57_864 ();
 FILLCELL_X16 FILLER_57_870 ();
 FILLCELL_X4 FILLER_57_889 ();
 FILLCELL_X4 FILLER_57_903 ();
 FILLCELL_X4 FILLER_57_911 ();
 FILLCELL_X2 FILLER_57_915 ();
 FILLCELL_X1 FILLER_57_917 ();
 FILLCELL_X8 FILLER_57_922 ();
 FILLCELL_X4 FILLER_57_939 ();
 FILLCELL_X1 FILLER_57_943 ();
 FILLCELL_X4 FILLER_57_947 ();
 FILLCELL_X4 FILLER_57_955 ();
 FILLCELL_X4 FILLER_57_968 ();
 FILLCELL_X4 FILLER_57_976 ();
 FILLCELL_X8 FILLER_57_987 ();
 FILLCELL_X1 FILLER_57_995 ();
 FILLCELL_X4 FILLER_57_1005 ();
 FILLCELL_X8 FILLER_57_1012 ();
 FILLCELL_X4 FILLER_57_1020 ();
 FILLCELL_X32 FILLER_58_1 ();
 FILLCELL_X32 FILLER_58_33 ();
 FILLCELL_X16 FILLER_58_65 ();
 FILLCELL_X1 FILLER_58_81 ();
 FILLCELL_X4 FILLER_58_85 ();
 FILLCELL_X4 FILLER_58_92 ();
 FILLCELL_X4 FILLER_58_101 ();
 FILLCELL_X4 FILLER_58_109 ();
 FILLCELL_X4 FILLER_58_116 ();
 FILLCELL_X2 FILLER_58_120 ();
 FILLCELL_X4 FILLER_58_125 ();
 FILLCELL_X4 FILLER_58_132 ();
 FILLCELL_X4 FILLER_58_139 ();
 FILLCELL_X8 FILLER_58_160 ();
 FILLCELL_X1 FILLER_58_168 ();
 FILLCELL_X16 FILLER_58_819 ();
 FILLCELL_X8 FILLER_58_841 ();
 FILLCELL_X2 FILLER_58_849 ();
 FILLCELL_X1 FILLER_58_851 ();
 FILLCELL_X4 FILLER_58_855 ();
 FILLCELL_X4 FILLER_58_869 ();
 FILLCELL_X2 FILLER_58_873 ();
 FILLCELL_X4 FILLER_58_878 ();
 FILLCELL_X1 FILLER_58_882 ();
 FILLCELL_X4 FILLER_58_886 ();
 FILLCELL_X2 FILLER_58_890 ();
 FILLCELL_X4 FILLER_58_895 ();
 FILLCELL_X8 FILLER_58_902 ();
 FILLCELL_X4 FILLER_58_910 ();
 FILLCELL_X1 FILLER_58_914 ();
 FILLCELL_X4 FILLER_58_924 ();
 FILLCELL_X2 FILLER_58_928 ();
 FILLCELL_X4 FILLER_58_939 ();
 FILLCELL_X8 FILLER_58_946 ();
 FILLCELL_X2 FILLER_58_954 ();
 FILLCELL_X1 FILLER_58_956 ();
 FILLCELL_X8 FILLER_58_966 ();
 FILLCELL_X4 FILLER_58_974 ();
 FILLCELL_X1 FILLER_58_978 ();
 FILLCELL_X4 FILLER_58_981 ();
 FILLCELL_X4 FILLER_58_988 ();
 FILLCELL_X4 FILLER_58_1001 ();
 FILLCELL_X16 FILLER_58_1008 ();
 FILLCELL_X32 FILLER_59_1 ();
 FILLCELL_X32 FILLER_59_33 ();
 FILLCELL_X16 FILLER_59_65 ();
 FILLCELL_X4 FILLER_59_81 ();
 FILLCELL_X1 FILLER_59_85 ();
 FILLCELL_X4 FILLER_59_105 ();
 FILLCELL_X4 FILLER_59_112 ();
 FILLCELL_X8 FILLER_59_119 ();
 FILLCELL_X8 FILLER_59_133 ();
 FILLCELL_X1 FILLER_59_141 ();
 FILLCELL_X4 FILLER_59_149 ();
 FILLCELL_X4 FILLER_59_158 ();
 FILLCELL_X4 FILLER_59_165 ();
 FILLCELL_X8 FILLER_59_819 ();
 FILLCELL_X2 FILLER_59_827 ();
 FILLCELL_X1 FILLER_59_829 ();
 FILLCELL_X8 FILLER_59_840 ();
 FILLCELL_X1 FILLER_59_848 ();
 FILLCELL_X4 FILLER_59_856 ();
 FILLCELL_X4 FILLER_59_866 ();
 FILLCELL_X2 FILLER_59_870 ();
 FILLCELL_X4 FILLER_59_882 ();
 FILLCELL_X4 FILLER_59_895 ();
 FILLCELL_X8 FILLER_59_909 ();
 FILLCELL_X2 FILLER_59_917 ();
 FILLCELL_X16 FILLER_59_922 ();
 FILLCELL_X4 FILLER_59_938 ();
 FILLCELL_X4 FILLER_59_949 ();
 FILLCELL_X4 FILLER_59_963 ();
 FILLCELL_X8 FILLER_59_970 ();
 FILLCELL_X1 FILLER_59_978 ();
 FILLCELL_X4 FILLER_59_989 ();
 FILLCELL_X4 FILLER_59_997 ();
 FILLCELL_X4 FILLER_59_1020 ();
 FILLCELL_X32 FILLER_60_1 ();
 FILLCELL_X32 FILLER_60_33 ();
 FILLCELL_X16 FILLER_60_65 ();
 FILLCELL_X8 FILLER_60_81 ();
 FILLCELL_X4 FILLER_60_89 ();
 FILLCELL_X2 FILLER_60_93 ();
 FILLCELL_X8 FILLER_60_98 ();
 FILLCELL_X8 FILLER_60_109 ();
 FILLCELL_X2 FILLER_60_117 ();
 FILLCELL_X4 FILLER_60_136 ();
 FILLCELL_X4 FILLER_60_145 ();
 FILLCELL_X2 FILLER_60_149 ();
 FILLCELL_X1 FILLER_60_151 ();
 FILLCELL_X4 FILLER_60_156 ();
 FILLCELL_X4 FILLER_60_164 ();
 FILLCELL_X1 FILLER_60_168 ();
 FILLCELL_X16 FILLER_60_819 ();
 FILLCELL_X8 FILLER_60_835 ();
 FILLCELL_X2 FILLER_60_843 ();
 FILLCELL_X1 FILLER_60_845 ();
 FILLCELL_X4 FILLER_60_852 ();
 FILLCELL_X8 FILLER_60_859 ();
 FILLCELL_X16 FILLER_60_874 ();
 FILLCELL_X1 FILLER_60_890 ();
 FILLCELL_X4 FILLER_60_900 ();
 FILLCELL_X4 FILLER_60_911 ();
 FILLCELL_X2 FILLER_60_915 ();
 FILLCELL_X4 FILLER_60_919 ();
 FILLCELL_X8 FILLER_60_926 ();
 FILLCELL_X4 FILLER_60_934 ();
 FILLCELL_X1 FILLER_60_938 ();
 FILLCELL_X4 FILLER_60_942 ();
 FILLCELL_X4 FILLER_60_949 ();
 FILLCELL_X1 FILLER_60_953 ();
 FILLCELL_X4 FILLER_60_958 ();
 FILLCELL_X16 FILLER_60_964 ();
 FILLCELL_X8 FILLER_60_980 ();
 FILLCELL_X4 FILLER_60_988 ();
 FILLCELL_X4 FILLER_60_996 ();
 FILLCELL_X16 FILLER_60_1004 ();
 FILLCELL_X4 FILLER_60_1020 ();
 FILLCELL_X4 FILLER_61_1 ();
 FILLCELL_X32 FILLER_61_9 ();
 FILLCELL_X32 FILLER_61_41 ();
 FILLCELL_X32 FILLER_61_73 ();
 FILLCELL_X8 FILLER_61_105 ();
 FILLCELL_X1 FILLER_61_113 ();
 FILLCELL_X4 FILLER_61_117 ();
 FILLCELL_X4 FILLER_61_125 ();
 FILLCELL_X4 FILLER_61_135 ();
 FILLCELL_X4 FILLER_61_141 ();
 FILLCELL_X8 FILLER_61_150 ();
 FILLCELL_X8 FILLER_61_161 ();
 FILLCELL_X16 FILLER_61_819 ();
 FILLCELL_X4 FILLER_61_835 ();
 FILLCELL_X1 FILLER_61_839 ();
 FILLCELL_X16 FILLER_61_844 ();
 FILLCELL_X8 FILLER_61_860 ();
 FILLCELL_X1 FILLER_61_868 ();
 FILLCELL_X4 FILLER_61_875 ();
 FILLCELL_X4 FILLER_61_881 ();
 FILLCELL_X1 FILLER_61_885 ();
 FILLCELL_X4 FILLER_61_892 ();
 FILLCELL_X1 FILLER_61_896 ();
 FILLCELL_X8 FILLER_61_899 ();
 FILLCELL_X2 FILLER_61_907 ();
 FILLCELL_X1 FILLER_61_909 ();
 FILLCELL_X4 FILLER_61_917 ();
 FILLCELL_X4 FILLER_61_931 ();
 FILLCELL_X8 FILLER_61_939 ();
 FILLCELL_X2 FILLER_61_947 ();
 FILLCELL_X4 FILLER_61_959 ();
 FILLCELL_X4 FILLER_61_966 ();
 FILLCELL_X1 FILLER_61_970 ();
 FILLCELL_X4 FILLER_61_975 ();
 FILLCELL_X8 FILLER_61_982 ();
 FILLCELL_X4 FILLER_61_990 ();
 FILLCELL_X2 FILLER_61_994 ();
 FILLCELL_X1 FILLER_61_996 ();
 FILLCELL_X16 FILLER_61_1000 ();
 FILLCELL_X8 FILLER_61_1016 ();
 FILLCELL_X32 FILLER_62_1 ();
 FILLCELL_X32 FILLER_62_33 ();
 FILLCELL_X32 FILLER_62_65 ();
 FILLCELL_X16 FILLER_62_97 ();
 FILLCELL_X1 FILLER_62_113 ();
 FILLCELL_X4 FILLER_62_117 ();
 FILLCELL_X8 FILLER_62_138 ();
 FILLCELL_X4 FILLER_62_152 ();
 FILLCELL_X8 FILLER_62_161 ();
 FILLCELL_X8 FILLER_62_819 ();
 FILLCELL_X4 FILLER_62_827 ();
 FILLCELL_X1 FILLER_62_831 ();
 FILLCELL_X8 FILLER_62_851 ();
 FILLCELL_X2 FILLER_62_859 ();
 FILLCELL_X4 FILLER_62_865 ();
 FILLCELL_X4 FILLER_62_876 ();
 FILLCELL_X8 FILLER_62_886 ();
 FILLCELL_X1 FILLER_62_894 ();
 FILLCELL_X8 FILLER_62_905 ();
 FILLCELL_X1 FILLER_62_913 ();
 FILLCELL_X4 FILLER_62_924 ();
 FILLCELL_X1 FILLER_62_928 ();
 FILLCELL_X4 FILLER_62_938 ();
 FILLCELL_X8 FILLER_62_951 ();
 FILLCELL_X1 FILLER_62_959 ();
 FILLCELL_X4 FILLER_62_964 ();
 FILLCELL_X4 FILLER_62_977 ();
 FILLCELL_X4 FILLER_62_985 ();
 FILLCELL_X2 FILLER_62_989 ();
 FILLCELL_X4 FILLER_62_995 ();
 FILLCELL_X4 FILLER_62_1008 ();
 FILLCELL_X8 FILLER_62_1015 ();
 FILLCELL_X1 FILLER_62_1023 ();
 FILLCELL_X32 FILLER_63_1 ();
 FILLCELL_X32 FILLER_63_33 ();
 FILLCELL_X32 FILLER_63_65 ();
 FILLCELL_X32 FILLER_63_97 ();
 FILLCELL_X1 FILLER_63_129 ();
 FILLCELL_X4 FILLER_63_135 ();
 FILLCELL_X2 FILLER_63_139 ();
 FILLCELL_X4 FILLER_63_158 ();
 FILLCELL_X4 FILLER_63_165 ();
 FILLCELL_X4 FILLER_63_819 ();
 FILLCELL_X2 FILLER_63_823 ();
 FILLCELL_X4 FILLER_63_844 ();
 FILLCELL_X16 FILLER_63_852 ();
 FILLCELL_X2 FILLER_63_868 ();
 FILLCELL_X1 FILLER_63_870 ();
 FILLCELL_X4 FILLER_63_875 ();
 FILLCELL_X2 FILLER_63_879 ();
 FILLCELL_X4 FILLER_63_884 ();
 FILLCELL_X2 FILLER_63_888 ();
 FILLCELL_X1 FILLER_63_890 ();
 FILLCELL_X16 FILLER_63_900 ();
 FILLCELL_X1 FILLER_63_916 ();
 FILLCELL_X4 FILLER_63_920 ();
 FILLCELL_X4 FILLER_63_928 ();
 FILLCELL_X4 FILLER_63_936 ();
 FILLCELL_X2 FILLER_63_940 ();
 FILLCELL_X1 FILLER_63_942 ();
 FILLCELL_X8 FILLER_63_952 ();
 FILLCELL_X4 FILLER_63_960 ();
 FILLCELL_X4 FILLER_63_973 ();
 FILLCELL_X8 FILLER_63_980 ();
 FILLCELL_X4 FILLER_63_988 ();
 FILLCELL_X4 FILLER_63_995 ();
 FILLCELL_X4 FILLER_63_1009 ();
 FILLCELL_X4 FILLER_63_1017 ();
 FILLCELL_X2 FILLER_63_1021 ();
 FILLCELL_X1 FILLER_63_1023 ();
 FILLCELL_X32 FILLER_64_1 ();
 FILLCELL_X32 FILLER_64_33 ();
 FILLCELL_X32 FILLER_64_65 ();
 FILLCELL_X32 FILLER_64_97 ();
 FILLCELL_X4 FILLER_64_129 ();
 FILLCELL_X1 FILLER_64_133 ();
 FILLCELL_X8 FILLER_64_137 ();
 FILLCELL_X4 FILLER_64_148 ();
 FILLCELL_X4 FILLER_64_155 ();
 FILLCELL_X2 FILLER_64_159 ();
 FILLCELL_X4 FILLER_64_164 ();
 FILLCELL_X1 FILLER_64_168 ();
 FILLCELL_X8 FILLER_64_819 ();
 FILLCELL_X4 FILLER_64_831 ();
 FILLCELL_X1 FILLER_64_835 ();
 FILLCELL_X4 FILLER_64_853 ();
 FILLCELL_X1 FILLER_64_857 ();
 FILLCELL_X16 FILLER_64_862 ();
 FILLCELL_X8 FILLER_64_878 ();
 FILLCELL_X4 FILLER_64_889 ();
 FILLCELL_X4 FILLER_64_896 ();
 FILLCELL_X4 FILLER_64_910 ();
 FILLCELL_X8 FILLER_64_917 ();
 FILLCELL_X4 FILLER_64_929 ();
 FILLCELL_X2 FILLER_64_933 ();
 FILLCELL_X1 FILLER_64_935 ();
 FILLCELL_X16 FILLER_64_939 ();
 FILLCELL_X2 FILLER_64_955 ();
 FILLCELL_X1 FILLER_64_957 ();
 FILLCELL_X4 FILLER_64_962 ();
 FILLCELL_X2 FILLER_64_966 ();
 FILLCELL_X8 FILLER_64_970 ();
 FILLCELL_X4 FILLER_64_978 ();
 FILLCELL_X2 FILLER_64_982 ();
 FILLCELL_X4 FILLER_64_986 ();
 FILLCELL_X4 FILLER_64_997 ();
 FILLCELL_X4 FILLER_64_1020 ();
 FILLCELL_X32 FILLER_65_1 ();
 FILLCELL_X32 FILLER_65_33 ();
 FILLCELL_X32 FILLER_65_65 ();
 FILLCELL_X32 FILLER_65_97 ();
 FILLCELL_X8 FILLER_65_129 ();
 FILLCELL_X2 FILLER_65_137 ();
 FILLCELL_X1 FILLER_65_139 ();
 FILLCELL_X8 FILLER_65_144 ();
 FILLCELL_X8 FILLER_65_156 ();
 FILLCELL_X4 FILLER_65_164 ();
 FILLCELL_X1 FILLER_65_168 ();
 FILLCELL_X16 FILLER_65_819 ();
 FILLCELL_X8 FILLER_65_835 ();
 FILLCELL_X4 FILLER_65_843 ();
 FILLCELL_X4 FILLER_65_851 ();
 FILLCELL_X4 FILLER_65_861 ();
 FILLCELL_X8 FILLER_65_869 ();
 FILLCELL_X1 FILLER_65_877 ();
 FILLCELL_X4 FILLER_65_882 ();
 FILLCELL_X2 FILLER_65_886 ();
 FILLCELL_X1 FILLER_65_888 ();
 FILLCELL_X4 FILLER_65_892 ();
 FILLCELL_X4 FILLER_65_900 ();
 FILLCELL_X2 FILLER_65_904 ();
 FILLCELL_X1 FILLER_65_906 ();
 FILLCELL_X4 FILLER_65_910 ();
 FILLCELL_X4 FILLER_65_923 ();
 FILLCELL_X4 FILLER_65_931 ();
 FILLCELL_X8 FILLER_65_937 ();
 FILLCELL_X4 FILLER_65_945 ();
 FILLCELL_X2 FILLER_65_949 ();
 FILLCELL_X4 FILLER_65_955 ();
 FILLCELL_X4 FILLER_65_969 ();
 FILLCELL_X4 FILLER_65_976 ();
 FILLCELL_X4 FILLER_65_983 ();
 FILLCELL_X4 FILLER_65_997 ();
 FILLCELL_X4 FILLER_65_1005 ();
 FILLCELL_X4 FILLER_65_1012 ();
 FILLCELL_X4 FILLER_65_1019 ();
 FILLCELL_X1 FILLER_65_1023 ();
 FILLCELL_X32 FILLER_66_1 ();
 FILLCELL_X32 FILLER_66_33 ();
 FILLCELL_X32 FILLER_66_65 ();
 FILLCELL_X32 FILLER_66_97 ();
 FILLCELL_X4 FILLER_66_129 ();
 FILLCELL_X8 FILLER_66_152 ();
 FILLCELL_X2 FILLER_66_160 ();
 FILLCELL_X4 FILLER_66_165 ();
 FILLCELL_X16 FILLER_66_819 ();
 FILLCELL_X8 FILLER_66_835 ();
 FILLCELL_X4 FILLER_66_847 ();
 FILLCELL_X4 FILLER_66_860 ();
 FILLCELL_X4 FILLER_66_870 ();
 FILLCELL_X8 FILLER_66_878 ();
 FILLCELL_X1 FILLER_66_886 ();
 FILLCELL_X4 FILLER_66_896 ();
 FILLCELL_X2 FILLER_66_900 ();
 FILLCELL_X4 FILLER_66_911 ();
 FILLCELL_X8 FILLER_66_919 ();
 FILLCELL_X2 FILLER_66_927 ();
 FILLCELL_X4 FILLER_66_936 ();
 FILLCELL_X4 FILLER_66_950 ();
 FILLCELL_X4 FILLER_66_957 ();
 FILLCELL_X1 FILLER_66_961 ();
 FILLCELL_X4 FILLER_66_972 ();
 FILLCELL_X4 FILLER_66_985 ();
 FILLCELL_X2 FILLER_66_989 ();
 FILLCELL_X1 FILLER_66_991 ();
 FILLCELL_X4 FILLER_66_996 ();
 FILLCELL_X4 FILLER_66_1009 ();
 FILLCELL_X4 FILLER_66_1017 ();
 FILLCELL_X2 FILLER_66_1021 ();
 FILLCELL_X1 FILLER_66_1023 ();
 FILLCELL_X32 FILLER_67_1 ();
 FILLCELL_X32 FILLER_67_33 ();
 FILLCELL_X32 FILLER_67_65 ();
 FILLCELL_X32 FILLER_67_97 ();
 FILLCELL_X8 FILLER_67_129 ();
 FILLCELL_X4 FILLER_67_137 ();
 FILLCELL_X1 FILLER_67_141 ();
 FILLCELL_X8 FILLER_67_161 ();
 FILLCELL_X16 FILLER_67_819 ();
 FILLCELL_X4 FILLER_67_835 ();
 FILLCELL_X4 FILLER_67_843 ();
 FILLCELL_X4 FILLER_67_853 ();
 FILLCELL_X2 FILLER_67_857 ();
 FILLCELL_X4 FILLER_67_866 ();
 FILLCELL_X1 FILLER_67_870 ();
 FILLCELL_X4 FILLER_67_878 ();
 FILLCELL_X4 FILLER_67_892 ();
 FILLCELL_X8 FILLER_67_899 ();
 FILLCELL_X1 FILLER_67_907 ();
 FILLCELL_X8 FILLER_67_911 ();
 FILLCELL_X1 FILLER_67_919 ();
 FILLCELL_X4 FILLER_67_939 ();
 FILLCELL_X4 FILLER_67_945 ();
 FILLCELL_X4 FILLER_67_951 ();
 FILLCELL_X2 FILLER_67_955 ();
 FILLCELL_X8 FILLER_67_960 ();
 FILLCELL_X1 FILLER_67_968 ();
 FILLCELL_X4 FILLER_67_972 ();
 FILLCELL_X8 FILLER_67_979 ();
 FILLCELL_X2 FILLER_67_987 ();
 FILLCELL_X4 FILLER_67_996 ();
 FILLCELL_X8 FILLER_67_1004 ();
 FILLCELL_X8 FILLER_67_1015 ();
 FILLCELL_X1 FILLER_67_1023 ();
 FILLCELL_X32 FILLER_68_1 ();
 FILLCELL_X32 FILLER_68_33 ();
 FILLCELL_X32 FILLER_68_65 ();
 FILLCELL_X32 FILLER_68_97 ();
 FILLCELL_X16 FILLER_68_129 ();
 FILLCELL_X4 FILLER_68_145 ();
 FILLCELL_X4 FILLER_68_152 ();
 FILLCELL_X8 FILLER_68_159 ();
 FILLCELL_X2 FILLER_68_167 ();
 FILLCELL_X8 FILLER_68_819 ();
 FILLCELL_X4 FILLER_68_837 ();
 FILLCELL_X2 FILLER_68_841 ();
 FILLCELL_X1 FILLER_68_843 ();
 FILLCELL_X4 FILLER_68_851 ();
 FILLCELL_X4 FILLER_68_861 ();
 FILLCELL_X2 FILLER_68_865 ();
 FILLCELL_X1 FILLER_68_867 ();
 FILLCELL_X16 FILLER_68_870 ();
 FILLCELL_X2 FILLER_68_886 ();
 FILLCELL_X1 FILLER_68_888 ();
 FILLCELL_X8 FILLER_68_891 ();
 FILLCELL_X4 FILLER_68_903 ();
 FILLCELL_X4 FILLER_68_909 ();
 FILLCELL_X16 FILLER_68_918 ();
 FILLCELL_X4 FILLER_68_934 ();
 FILLCELL_X16 FILLER_68_944 ();
 FILLCELL_X4 FILLER_68_960 ();
 FILLCELL_X1 FILLER_68_964 ();
 FILLCELL_X4 FILLER_68_974 ();
 FILLCELL_X4 FILLER_68_982 ();
 FILLCELL_X4 FILLER_68_989 ();
 FILLCELL_X4 FILLER_68_1003 ();
 FILLCELL_X1 FILLER_68_1007 ();
 FILLCELL_X4 FILLER_68_1017 ();
 FILLCELL_X2 FILLER_68_1021 ();
 FILLCELL_X1 FILLER_68_1023 ();
 FILLCELL_X32 FILLER_69_1 ();
 FILLCELL_X32 FILLER_69_33 ();
 FILLCELL_X32 FILLER_69_65 ();
 FILLCELL_X16 FILLER_69_97 ();
 FILLCELL_X8 FILLER_69_113 ();
 FILLCELL_X4 FILLER_69_121 ();
 FILLCELL_X1 FILLER_69_125 ();
 FILLCELL_X4 FILLER_69_130 ();
 FILLCELL_X8 FILLER_69_153 ();
 FILLCELL_X1 FILLER_69_161 ();
 FILLCELL_X4 FILLER_69_165 ();
 FILLCELL_X16 FILLER_69_819 ();
 FILLCELL_X2 FILLER_69_835 ();
 FILLCELL_X1 FILLER_69_837 ();
 FILLCELL_X4 FILLER_69_841 ();
 FILLCELL_X4 FILLER_69_849 ();
 FILLCELL_X8 FILLER_69_856 ();
 FILLCELL_X2 FILLER_69_864 ();
 FILLCELL_X16 FILLER_69_869 ();
 FILLCELL_X2 FILLER_69_885 ();
 FILLCELL_X4 FILLER_69_897 ();
 FILLCELL_X4 FILLER_69_904 ();
 FILLCELL_X4 FILLER_69_918 ();
 FILLCELL_X2 FILLER_69_922 ();
 FILLCELL_X16 FILLER_69_927 ();
 FILLCELL_X2 FILLER_69_943 ();
 FILLCELL_X1 FILLER_69_945 ();
 FILLCELL_X4 FILLER_69_949 ();
 FILLCELL_X4 FILLER_69_963 ();
 FILLCELL_X4 FILLER_69_971 ();
 FILLCELL_X8 FILLER_69_979 ();
 FILLCELL_X1 FILLER_69_987 ();
 FILLCELL_X4 FILLER_69_998 ();
 FILLCELL_X2 FILLER_69_1002 ();
 FILLCELL_X8 FILLER_69_1008 ();
 FILLCELL_X1 FILLER_69_1016 ();
 FILLCELL_X4 FILLER_69_1020 ();
 FILLCELL_X32 FILLER_70_1 ();
 FILLCELL_X32 FILLER_70_33 ();
 FILLCELL_X32 FILLER_70_65 ();
 FILLCELL_X32 FILLER_70_97 ();
 FILLCELL_X16 FILLER_70_129 ();
 FILLCELL_X1 FILLER_70_145 ();
 FILLCELL_X4 FILLER_70_165 ();
 FILLCELL_X8 FILLER_70_819 ();
 FILLCELL_X2 FILLER_70_827 ();
 FILLCELL_X1 FILLER_70_829 ();
 FILLCELL_X4 FILLER_70_836 ();
 FILLCELL_X2 FILLER_70_840 ();
 FILLCELL_X4 FILLER_70_861 ();
 FILLCELL_X4 FILLER_70_875 ();
 FILLCELL_X2 FILLER_70_879 ();
 FILLCELL_X4 FILLER_70_884 ();
 FILLCELL_X2 FILLER_70_888 ();
 FILLCELL_X1 FILLER_70_890 ();
 FILLCELL_X8 FILLER_70_894 ();
 FILLCELL_X1 FILLER_70_902 ();
 FILLCELL_X4 FILLER_70_906 ();
 FILLCELL_X2 FILLER_70_910 ();
 FILLCELL_X1 FILLER_70_912 ();
 FILLCELL_X4 FILLER_70_922 ();
 FILLCELL_X2 FILLER_70_926 ();
 FILLCELL_X1 FILLER_70_928 ();
 FILLCELL_X4 FILLER_70_935 ();
 FILLCELL_X2 FILLER_70_939 ();
 FILLCELL_X4 FILLER_70_944 ();
 FILLCELL_X4 FILLER_70_955 ();
 FILLCELL_X8 FILLER_70_961 ();
 FILLCELL_X4 FILLER_70_978 ();
 FILLCELL_X8 FILLER_70_985 ();
 FILLCELL_X4 FILLER_70_995 ();
 FILLCELL_X4 FILLER_70_1003 ();
 FILLCELL_X8 FILLER_70_1016 ();
 FILLCELL_X4 FILLER_71_1 ();
 FILLCELL_X32 FILLER_71_8 ();
 FILLCELL_X32 FILLER_71_40 ();
 FILLCELL_X32 FILLER_71_72 ();
 FILLCELL_X32 FILLER_71_104 ();
 FILLCELL_X16 FILLER_71_136 ();
 FILLCELL_X2 FILLER_71_152 ();
 FILLCELL_X4 FILLER_71_158 ();
 FILLCELL_X4 FILLER_71_165 ();
 FILLCELL_X8 FILLER_71_819 ();
 FILLCELL_X4 FILLER_71_827 ();
 FILLCELL_X2 FILLER_71_831 ();
 FILLCELL_X4 FILLER_71_840 ();
 FILLCELL_X4 FILLER_71_848 ();
 FILLCELL_X4 FILLER_71_856 ();
 FILLCELL_X8 FILLER_71_863 ();
 FILLCELL_X4 FILLER_71_875 ();
 FILLCELL_X1 FILLER_71_879 ();
 FILLCELL_X4 FILLER_71_889 ();
 FILLCELL_X2 FILLER_71_893 ();
 FILLCELL_X1 FILLER_71_895 ();
 FILLCELL_X4 FILLER_71_906 ();
 FILLCELL_X2 FILLER_71_910 ();
 FILLCELL_X1 FILLER_71_912 ();
 FILLCELL_X4 FILLER_71_922 ();
 FILLCELL_X2 FILLER_71_926 ();
 FILLCELL_X4 FILLER_71_935 ();
 FILLCELL_X4 FILLER_71_942 ();
 FILLCELL_X4 FILLER_71_950 ();
 FILLCELL_X4 FILLER_71_964 ();
 FILLCELL_X1 FILLER_71_968 ();
 FILLCELL_X4 FILLER_71_971 ();
 FILLCELL_X1 FILLER_71_975 ();
 FILLCELL_X8 FILLER_71_985 ();
 FILLCELL_X4 FILLER_71_993 ();
 FILLCELL_X1 FILLER_71_997 ();
 FILLCELL_X4 FILLER_71_1000 ();
 FILLCELL_X8 FILLER_71_1014 ();
 FILLCELL_X2 FILLER_71_1022 ();
 FILLCELL_X32 FILLER_72_1 ();
 FILLCELL_X32 FILLER_72_33 ();
 FILLCELL_X32 FILLER_72_65 ();
 FILLCELL_X32 FILLER_72_97 ();
 FILLCELL_X4 FILLER_72_129 ();
 FILLCELL_X2 FILLER_72_133 ();
 FILLCELL_X1 FILLER_72_135 ();
 FILLCELL_X4 FILLER_72_140 ();
 FILLCELL_X4 FILLER_72_163 ();
 FILLCELL_X2 FILLER_72_167 ();
 FILLCELL_X8 FILLER_72_819 ();
 FILLCELL_X2 FILLER_72_827 ();
 FILLCELL_X1 FILLER_72_829 ();
 FILLCELL_X4 FILLER_72_832 ();
 FILLCELL_X8 FILLER_72_840 ();
 FILLCELL_X4 FILLER_72_858 ();
 FILLCELL_X2 FILLER_72_862 ();
 FILLCELL_X4 FILLER_72_868 ();
 FILLCELL_X4 FILLER_72_881 ();
 FILLCELL_X8 FILLER_72_889 ();
 FILLCELL_X4 FILLER_72_897 ();
 FILLCELL_X2 FILLER_72_901 ();
 FILLCELL_X4 FILLER_72_910 ();
 FILLCELL_X4 FILLER_72_917 ();
 FILLCELL_X2 FILLER_72_921 ();
 FILLCELL_X4 FILLER_72_925 ();
 FILLCELL_X4 FILLER_72_935 ();
 FILLCELL_X4 FILLER_72_943 ();
 FILLCELL_X4 FILLER_72_966 ();
 FILLCELL_X1 FILLER_72_970 ();
 FILLCELL_X4 FILLER_72_974 ();
 FILLCELL_X4 FILLER_72_981 ();
 FILLCELL_X2 FILLER_72_985 ();
 FILLCELL_X4 FILLER_72_989 ();
 FILLCELL_X4 FILLER_72_997 ();
 FILLCELL_X4 FILLER_72_1011 ();
 FILLCELL_X4 FILLER_72_1018 ();
 FILLCELL_X2 FILLER_72_1022 ();
 FILLCELL_X32 FILLER_73_1 ();
 FILLCELL_X32 FILLER_73_33 ();
 FILLCELL_X32 FILLER_73_65 ();
 FILLCELL_X32 FILLER_73_97 ();
 FILLCELL_X16 FILLER_73_129 ();
 FILLCELL_X8 FILLER_73_145 ();
 FILLCELL_X4 FILLER_73_153 ();
 FILLCELL_X1 FILLER_73_157 ();
 FILLCELL_X8 FILLER_73_161 ();
 FILLCELL_X16 FILLER_73_819 ();
 FILLCELL_X8 FILLER_73_835 ();
 FILLCELL_X4 FILLER_73_843 ();
 FILLCELL_X1 FILLER_73_847 ();
 FILLCELL_X4 FILLER_73_852 ();
 FILLCELL_X2 FILLER_73_856 ();
 FILLCELL_X8 FILLER_73_860 ();
 FILLCELL_X4 FILLER_73_868 ();
 FILLCELL_X1 FILLER_73_872 ();
 FILLCELL_X4 FILLER_73_878 ();
 FILLCELL_X16 FILLER_73_885 ();
 FILLCELL_X1 FILLER_73_901 ();
 FILLCELL_X4 FILLER_73_904 ();
 FILLCELL_X16 FILLER_73_918 ();
 FILLCELL_X4 FILLER_73_934 ();
 FILLCELL_X32 FILLER_73_941 ();
 FILLCELL_X4 FILLER_73_973 ();
 FILLCELL_X8 FILLER_73_986 ();
 FILLCELL_X4 FILLER_73_994 ();
 FILLCELL_X2 FILLER_73_998 ();
 FILLCELL_X4 FILLER_73_1019 ();
 FILLCELL_X1 FILLER_73_1023 ();
 FILLCELL_X32 FILLER_74_1 ();
 FILLCELL_X32 FILLER_74_33 ();
 FILLCELL_X32 FILLER_74_65 ();
 FILLCELL_X32 FILLER_74_97 ();
 FILLCELL_X32 FILLER_74_129 ();
 FILLCELL_X8 FILLER_74_161 ();
 FILLCELL_X4 FILLER_74_819 ();
 FILLCELL_X1 FILLER_74_823 ();
 FILLCELL_X4 FILLER_74_827 ();
 FILLCELL_X4 FILLER_74_835 ();
 FILLCELL_X4 FILLER_74_848 ();
 FILLCELL_X4 FILLER_74_858 ();
 FILLCELL_X1 FILLER_74_862 ();
 FILLCELL_X16 FILLER_74_866 ();
 FILLCELL_X1 FILLER_74_882 ();
 FILLCELL_X4 FILLER_74_887 ();
 FILLCELL_X4 FILLER_74_895 ();
 FILLCELL_X4 FILLER_74_902 ();
 FILLCELL_X2 FILLER_74_906 ();
 FILLCELL_X4 FILLER_74_912 ();
 FILLCELL_X1 FILLER_74_916 ();
 FILLCELL_X4 FILLER_74_920 ();
 FILLCELL_X4 FILLER_74_930 ();
 FILLCELL_X4 FILLER_74_943 ();
 FILLCELL_X8 FILLER_74_953 ();
 FILLCELL_X4 FILLER_74_961 ();
 FILLCELL_X2 FILLER_74_965 ();
 FILLCELL_X1 FILLER_74_967 ();
 FILLCELL_X4 FILLER_74_972 ();
 FILLCELL_X4 FILLER_74_986 ();
 FILLCELL_X1 FILLER_74_990 ();
 FILLCELL_X4 FILLER_74_998 ();
 FILLCELL_X8 FILLER_74_1006 ();
 FILLCELL_X2 FILLER_74_1014 ();
 FILLCELL_X4 FILLER_74_1019 ();
 FILLCELL_X1 FILLER_74_1023 ();
 FILLCELL_X32 FILLER_75_1 ();
 FILLCELL_X32 FILLER_75_33 ();
 FILLCELL_X32 FILLER_75_65 ();
 FILLCELL_X32 FILLER_75_97 ();
 FILLCELL_X32 FILLER_75_129 ();
 FILLCELL_X1 FILLER_75_161 ();
 FILLCELL_X4 FILLER_75_165 ();
 FILLCELL_X8 FILLER_75_819 ();
 FILLCELL_X4 FILLER_75_827 ();
 FILLCELL_X2 FILLER_75_831 ();
 FILLCELL_X4 FILLER_75_837 ();
 FILLCELL_X4 FILLER_75_844 ();
 FILLCELL_X4 FILLER_75_855 ();
 FILLCELL_X4 FILLER_75_863 ();
 FILLCELL_X1 FILLER_75_867 ();
 FILLCELL_X8 FILLER_75_872 ();
 FILLCELL_X4 FILLER_75_880 ();
 FILLCELL_X2 FILLER_75_884 ();
 FILLCELL_X4 FILLER_75_895 ();
 FILLCELL_X4 FILLER_75_908 ();
 FILLCELL_X4 FILLER_75_915 ();
 FILLCELL_X8 FILLER_75_922 ();
 FILLCELL_X8 FILLER_75_939 ();
 FILLCELL_X1 FILLER_75_947 ();
 FILLCELL_X4 FILLER_75_951 ();
 FILLCELL_X4 FILLER_75_965 ();
 FILLCELL_X1 FILLER_75_969 ();
 FILLCELL_X4 FILLER_75_972 ();
 FILLCELL_X4 FILLER_75_983 ();
 FILLCELL_X1 FILLER_75_987 ();
 FILLCELL_X8 FILLER_75_991 ();
 FILLCELL_X1 FILLER_75_999 ();
 FILLCELL_X4 FILLER_75_1003 ();
 FILLCELL_X4 FILLER_75_1011 ();
 FILLCELL_X2 FILLER_75_1015 ();
 FILLCELL_X4 FILLER_75_1020 ();
 FILLCELL_X32 FILLER_76_1 ();
 FILLCELL_X32 FILLER_76_33 ();
 FILLCELL_X32 FILLER_76_65 ();
 FILLCELL_X32 FILLER_76_97 ();
 FILLCELL_X16 FILLER_76_129 ();
 FILLCELL_X8 FILLER_76_145 ();
 FILLCELL_X4 FILLER_76_153 ();
 FILLCELL_X2 FILLER_76_157 ();
 FILLCELL_X4 FILLER_76_162 ();
 FILLCELL_X2 FILLER_76_166 ();
 FILLCELL_X1 FILLER_76_168 ();
 FILLCELL_X8 FILLER_76_819 ();
 FILLCELL_X1 FILLER_76_827 ();
 FILLCELL_X4 FILLER_76_832 ();
 FILLCELL_X4 FILLER_76_845 ();
 FILLCELL_X4 FILLER_76_852 ();
 FILLCELL_X1 FILLER_76_856 ();
 FILLCELL_X4 FILLER_76_867 ();
 FILLCELL_X4 FILLER_76_880 ();
 FILLCELL_X4 FILLER_76_887 ();
 FILLCELL_X1 FILLER_76_891 ();
 FILLCELL_X4 FILLER_76_896 ();
 FILLCELL_X4 FILLER_76_903 ();
 FILLCELL_X1 FILLER_76_907 ();
 FILLCELL_X4 FILLER_76_918 ();
 FILLCELL_X4 FILLER_76_929 ();
 FILLCELL_X8 FILLER_76_936 ();
 FILLCELL_X1 FILLER_76_944 ();
 FILLCELL_X8 FILLER_76_949 ();
 FILLCELL_X2 FILLER_76_957 ();
 FILLCELL_X16 FILLER_76_963 ();
 FILLCELL_X2 FILLER_76_979 ();
 FILLCELL_X1 FILLER_76_981 ();
 FILLCELL_X8 FILLER_76_992 ();
 FILLCELL_X2 FILLER_76_1000 ();
 FILLCELL_X4 FILLER_76_1006 ();
 FILLCELL_X8 FILLER_76_1014 ();
 FILLCELL_X2 FILLER_76_1022 ();
 FILLCELL_X32 FILLER_77_1 ();
 FILLCELL_X32 FILLER_77_33 ();
 FILLCELL_X32 FILLER_77_65 ();
 FILLCELL_X32 FILLER_77_97 ();
 FILLCELL_X16 FILLER_77_129 ();
 FILLCELL_X4 FILLER_77_162 ();
 FILLCELL_X2 FILLER_77_166 ();
 FILLCELL_X1 FILLER_77_168 ();
 FILLCELL_X16 FILLER_77_819 ();
 FILLCELL_X8 FILLER_77_835 ();
 FILLCELL_X2 FILLER_77_843 ();
 FILLCELL_X1 FILLER_77_845 ();
 FILLCELL_X4 FILLER_77_849 ();
 FILLCELL_X8 FILLER_77_855 ();
 FILLCELL_X4 FILLER_77_863 ();
 FILLCELL_X2 FILLER_77_867 ();
 FILLCELL_X4 FILLER_77_873 ();
 FILLCELL_X16 FILLER_77_886 ();
 FILLCELL_X8 FILLER_77_902 ();
 FILLCELL_X2 FILLER_77_910 ();
 FILLCELL_X1 FILLER_77_912 ();
 FILLCELL_X4 FILLER_77_915 ();
 FILLCELL_X4 FILLER_77_929 ();
 FILLCELL_X2 FILLER_77_933 ();
 FILLCELL_X1 FILLER_77_935 ();
 FILLCELL_X4 FILLER_77_942 ();
 FILLCELL_X8 FILLER_77_953 ();
 FILLCELL_X2 FILLER_77_961 ();
 FILLCELL_X1 FILLER_77_963 ();
 FILLCELL_X4 FILLER_77_974 ();
 FILLCELL_X2 FILLER_77_978 ();
 FILLCELL_X4 FILLER_77_983 ();
 FILLCELL_X4 FILLER_77_993 ();
 FILLCELL_X8 FILLER_77_1001 ();
 FILLCELL_X4 FILLER_77_1018 ();
 FILLCELL_X2 FILLER_77_1022 ();
 FILLCELL_X32 FILLER_78_1 ();
 FILLCELL_X32 FILLER_78_33 ();
 FILLCELL_X32 FILLER_78_65 ();
 FILLCELL_X32 FILLER_78_97 ();
 FILLCELL_X16 FILLER_78_129 ();
 FILLCELL_X2 FILLER_78_145 ();
 FILLCELL_X1 FILLER_78_147 ();
 FILLCELL_X4 FILLER_78_151 ();
 FILLCELL_X8 FILLER_78_159 ();
 FILLCELL_X2 FILLER_78_167 ();
 FILLCELL_X16 FILLER_78_819 ();
 FILLCELL_X1 FILLER_78_835 ();
 FILLCELL_X4 FILLER_78_842 ();
 FILLCELL_X4 FILLER_78_852 ();
 FILLCELL_X4 FILLER_78_859 ();
 FILLCELL_X8 FILLER_78_865 ();
 FILLCELL_X2 FILLER_78_873 ();
 FILLCELL_X1 FILLER_78_875 ();
 FILLCELL_X4 FILLER_78_879 ();
 FILLCELL_X16 FILLER_78_886 ();
 FILLCELL_X4 FILLER_78_902 ();
 FILLCELL_X2 FILLER_78_906 ();
 FILLCELL_X4 FILLER_78_912 ();
 FILLCELL_X8 FILLER_78_919 ();
 FILLCELL_X2 FILLER_78_927 ();
 FILLCELL_X8 FILLER_78_933 ();
 FILLCELL_X1 FILLER_78_941 ();
 FILLCELL_X4 FILLER_78_952 ();
 FILLCELL_X4 FILLER_78_960 ();
 FILLCELL_X4 FILLER_78_966 ();
 FILLCELL_X4 FILLER_78_973 ();
 FILLCELL_X4 FILLER_78_984 ();
 FILLCELL_X8 FILLER_78_994 ();
 FILLCELL_X4 FILLER_78_1005 ();
 FILLCELL_X4 FILLER_78_1018 ();
 FILLCELL_X2 FILLER_78_1022 ();
 FILLCELL_X32 FILLER_79_1 ();
 FILLCELL_X32 FILLER_79_33 ();
 FILLCELL_X32 FILLER_79_65 ();
 FILLCELL_X32 FILLER_79_97 ();
 FILLCELL_X32 FILLER_79_129 ();
 FILLCELL_X4 FILLER_79_165 ();
 FILLCELL_X8 FILLER_79_819 ();
 FILLCELL_X1 FILLER_79_827 ();
 FILLCELL_X4 FILLER_79_832 ();
 FILLCELL_X4 FILLER_79_846 ();
 FILLCELL_X4 FILLER_79_857 ();
 FILLCELL_X1 FILLER_79_861 ();
 FILLCELL_X8 FILLER_79_872 ();
 FILLCELL_X4 FILLER_79_880 ();
 FILLCELL_X8 FILLER_79_893 ();
 FILLCELL_X1 FILLER_79_901 ();
 FILLCELL_X4 FILLER_79_906 ();
 FILLCELL_X2 FILLER_79_910 ();
 FILLCELL_X1 FILLER_79_912 ();
 FILLCELL_X4 FILLER_79_922 ();
 FILLCELL_X4 FILLER_79_929 ();
 FILLCELL_X4 FILLER_79_936 ();
 FILLCELL_X16 FILLER_79_943 ();
 FILLCELL_X4 FILLER_79_959 ();
 FILLCELL_X4 FILLER_79_966 ();
 FILLCELL_X1 FILLER_79_970 ();
 FILLCELL_X4 FILLER_79_980 ();
 FILLCELL_X4 FILLER_79_987 ();
 FILLCELL_X4 FILLER_79_994 ();
 FILLCELL_X2 FILLER_79_998 ();
 FILLCELL_X1 FILLER_79_1000 ();
 FILLCELL_X4 FILLER_79_1004 ();
 FILLCELL_X4 FILLER_79_1017 ();
 FILLCELL_X2 FILLER_79_1021 ();
 FILLCELL_X1 FILLER_79_1023 ();
 FILLCELL_X32 FILLER_80_1 ();
 FILLCELL_X32 FILLER_80_33 ();
 FILLCELL_X32 FILLER_80_65 ();
 FILLCELL_X32 FILLER_80_97 ();
 FILLCELL_X32 FILLER_80_129 ();
 FILLCELL_X1 FILLER_80_161 ();
 FILLCELL_X4 FILLER_80_165 ();
 FILLCELL_X4 FILLER_80_819 ();
 FILLCELL_X2 FILLER_80_823 ();
 FILLCELL_X16 FILLER_80_844 ();
 FILLCELL_X2 FILLER_80_860 ();
 FILLCELL_X1 FILLER_80_862 ();
 FILLCELL_X4 FILLER_80_866 ();
 FILLCELL_X4 FILLER_80_880 ();
 FILLCELL_X4 FILLER_80_888 ();
 FILLCELL_X4 FILLER_80_896 ();
 FILLCELL_X4 FILLER_80_904 ();
 FILLCELL_X4 FILLER_80_912 ();
 FILLCELL_X1 FILLER_80_916 ();
 FILLCELL_X4 FILLER_80_921 ();
 FILLCELL_X8 FILLER_80_934 ();
 FILLCELL_X2 FILLER_80_942 ();
 FILLCELL_X8 FILLER_80_954 ();
 FILLCELL_X1 FILLER_80_962 ();
 FILLCELL_X4 FILLER_80_966 ();
 FILLCELL_X4 FILLER_80_979 ();
 FILLCELL_X4 FILLER_80_993 ();
 FILLCELL_X4 FILLER_80_1001 ();
 FILLCELL_X2 FILLER_80_1005 ();
 FILLCELL_X1 FILLER_80_1007 ();
 FILLCELL_X4 FILLER_80_1018 ();
 FILLCELL_X2 FILLER_80_1022 ();
 FILLCELL_X32 FILLER_81_1 ();
 FILLCELL_X32 FILLER_81_33 ();
 FILLCELL_X32 FILLER_81_65 ();
 FILLCELL_X32 FILLER_81_97 ();
 FILLCELL_X16 FILLER_81_129 ();
 FILLCELL_X2 FILLER_81_145 ();
 FILLCELL_X1 FILLER_81_147 ();
 FILLCELL_X4 FILLER_81_165 ();
 FILLCELL_X16 FILLER_81_819 ();
 FILLCELL_X4 FILLER_81_835 ();
 FILLCELL_X2 FILLER_81_839 ();
 FILLCELL_X1 FILLER_81_841 ();
 FILLCELL_X16 FILLER_81_848 ();
 FILLCELL_X2 FILLER_81_864 ();
 FILLCELL_X1 FILLER_81_866 ();
 FILLCELL_X8 FILLER_81_871 ();
 FILLCELL_X4 FILLER_81_879 ();
 FILLCELL_X16 FILLER_81_887 ();
 FILLCELL_X1 FILLER_81_903 ();
 FILLCELL_X8 FILLER_81_908 ();
 FILLCELL_X16 FILLER_81_919 ();
 FILLCELL_X4 FILLER_81_939 ();
 FILLCELL_X4 FILLER_81_946 ();
 FILLCELL_X2 FILLER_81_950 ();
 FILLCELL_X1 FILLER_81_952 ();
 FILLCELL_X4 FILLER_81_955 ();
 FILLCELL_X16 FILLER_81_966 ();
 FILLCELL_X8 FILLER_81_989 ();
 FILLCELL_X1 FILLER_81_997 ();
 FILLCELL_X4 FILLER_81_1001 ();
 FILLCELL_X2 FILLER_81_1005 ();
 FILLCELL_X4 FILLER_81_1014 ();
 FILLCELL_X4 FILLER_81_1020 ();
 FILLCELL_X4 FILLER_82_1 ();
 FILLCELL_X32 FILLER_82_8 ();
 FILLCELL_X32 FILLER_82_40 ();
 FILLCELL_X32 FILLER_82_72 ();
 FILLCELL_X32 FILLER_82_104 ();
 FILLCELL_X16 FILLER_82_136 ();
 FILLCELL_X8 FILLER_82_152 ();
 FILLCELL_X2 FILLER_82_160 ();
 FILLCELL_X4 FILLER_82_165 ();
 FILLCELL_X16 FILLER_82_819 ();
 FILLCELL_X8 FILLER_82_835 ();
 FILLCELL_X4 FILLER_82_843 ();
 FILLCELL_X4 FILLER_82_854 ();
 FILLCELL_X8 FILLER_82_862 ();
 FILLCELL_X4 FILLER_82_879 ();
 FILLCELL_X16 FILLER_82_886 ();
 FILLCELL_X2 FILLER_82_902 ();
 FILLCELL_X1 FILLER_82_904 ();
 FILLCELL_X8 FILLER_82_914 ();
 FILLCELL_X2 FILLER_82_922 ();
 FILLCELL_X4 FILLER_82_928 ();
 FILLCELL_X4 FILLER_82_936 ();
 FILLCELL_X4 FILLER_82_949 ();
 FILLCELL_X4 FILLER_82_956 ();
 FILLCELL_X8 FILLER_82_970 ();
 FILLCELL_X4 FILLER_82_978 ();
 FILLCELL_X1 FILLER_82_982 ();
 FILLCELL_X4 FILLER_82_986 ();
 FILLCELL_X2 FILLER_82_990 ();
 FILLCELL_X1 FILLER_82_992 ();
 FILLCELL_X4 FILLER_82_997 ();
 FILLCELL_X4 FILLER_82_1005 ();
 FILLCELL_X4 FILLER_82_1018 ();
 FILLCELL_X2 FILLER_82_1022 ();
 FILLCELL_X32 FILLER_83_1 ();
 FILLCELL_X32 FILLER_83_33 ();
 FILLCELL_X32 FILLER_83_65 ();
 FILLCELL_X32 FILLER_83_97 ();
 FILLCELL_X32 FILLER_83_129 ();
 FILLCELL_X8 FILLER_83_161 ();
 FILLCELL_X16 FILLER_83_819 ();
 FILLCELL_X8 FILLER_83_835 ();
 FILLCELL_X4 FILLER_83_843 ();
 FILLCELL_X2 FILLER_83_847 ();
 FILLCELL_X8 FILLER_83_853 ();
 FILLCELL_X1 FILLER_83_861 ();
 FILLCELL_X4 FILLER_83_866 ();
 FILLCELL_X4 FILLER_83_879 ();
 FILLCELL_X4 FILLER_83_887 ();
 FILLCELL_X4 FILLER_83_894 ();
 FILLCELL_X8 FILLER_83_901 ();
 FILLCELL_X4 FILLER_83_913 ();
 FILLCELL_X4 FILLER_83_921 ();
 FILLCELL_X4 FILLER_83_928 ();
 FILLCELL_X2 FILLER_83_932 ();
 FILLCELL_X1 FILLER_83_934 ();
 FILLCELL_X4 FILLER_83_939 ();
 FILLCELL_X4 FILLER_83_952 ();
 FILLCELL_X16 FILLER_83_959 ();
 FILLCELL_X2 FILLER_83_975 ();
 FILLCELL_X1 FILLER_83_977 ();
 FILLCELL_X4 FILLER_83_981 ();
 FILLCELL_X4 FILLER_83_987 ();
 FILLCELL_X8 FILLER_83_997 ();
 FILLCELL_X8 FILLER_83_1015 ();
 FILLCELL_X1 FILLER_83_1023 ();
 FILLCELL_X32 FILLER_84_1 ();
 FILLCELL_X32 FILLER_84_33 ();
 FILLCELL_X32 FILLER_84_65 ();
 FILLCELL_X32 FILLER_84_97 ();
 FILLCELL_X32 FILLER_84_129 ();
 FILLCELL_X8 FILLER_84_161 ();
 FILLCELL_X8 FILLER_84_819 ();
 FILLCELL_X4 FILLER_84_827 ();
 FILLCELL_X2 FILLER_84_831 ();
 FILLCELL_X1 FILLER_84_833 ();
 FILLCELL_X4 FILLER_84_838 ();
 FILLCELL_X4 FILLER_84_845 ();
 FILLCELL_X4 FILLER_84_855 ();
 FILLCELL_X4 FILLER_84_863 ();
 FILLCELL_X4 FILLER_84_869 ();
 FILLCELL_X4 FILLER_84_877 ();
 FILLCELL_X4 FILLER_84_888 ();
 FILLCELL_X4 FILLER_84_896 ();
 FILLCELL_X2 FILLER_84_900 ();
 FILLCELL_X4 FILLER_84_906 ();
 FILLCELL_X4 FILLER_84_919 ();
 FILLCELL_X2 FILLER_84_923 ();
 FILLCELL_X4 FILLER_84_929 ();
 FILLCELL_X16 FILLER_84_936 ();
 FILLCELL_X8 FILLER_84_952 ();
 FILLCELL_X4 FILLER_84_960 ();
 FILLCELL_X4 FILLER_84_966 ();
 FILLCELL_X1 FILLER_84_970 ();
 FILLCELL_X4 FILLER_84_974 ();
 FILLCELL_X4 FILLER_84_987 ();
 FILLCELL_X1 FILLER_84_991 ();
 FILLCELL_X4 FILLER_84_995 ();
 FILLCELL_X8 FILLER_84_1008 ();
 FILLCELL_X1 FILLER_84_1016 ();
 FILLCELL_X4 FILLER_84_1020 ();
 FILLCELL_X32 FILLER_85_1 ();
 FILLCELL_X32 FILLER_85_33 ();
 FILLCELL_X32 FILLER_85_65 ();
 FILLCELL_X32 FILLER_85_97 ();
 FILLCELL_X32 FILLER_85_129 ();
 FILLCELL_X1 FILLER_85_161 ();
 FILLCELL_X4 FILLER_85_165 ();
 FILLCELL_X4 FILLER_85_819 ();
 FILLCELL_X2 FILLER_85_823 ();
 FILLCELL_X1 FILLER_85_825 ();
 FILLCELL_X4 FILLER_85_830 ();
 FILLCELL_X8 FILLER_85_838 ();
 FILLCELL_X1 FILLER_85_846 ();
 FILLCELL_X4 FILLER_85_857 ();
 FILLCELL_X8 FILLER_85_868 ();
 FILLCELL_X1 FILLER_85_876 ();
 FILLCELL_X4 FILLER_85_881 ();
 FILLCELL_X8 FILLER_85_891 ();
 FILLCELL_X1 FILLER_85_899 ();
 FILLCELL_X4 FILLER_85_904 ();
 FILLCELL_X2 FILLER_85_908 ();
 FILLCELL_X16 FILLER_85_912 ();
 FILLCELL_X2 FILLER_85_928 ();
 FILLCELL_X8 FILLER_85_934 ();
 FILLCELL_X2 FILLER_85_942 ();
 FILLCELL_X1 FILLER_85_944 ();
 FILLCELL_X4 FILLER_85_955 ();
 FILLCELL_X4 FILLER_85_962 ();
 FILLCELL_X4 FILLER_85_973 ();
 FILLCELL_X4 FILLER_85_987 ();
 FILLCELL_X4 FILLER_85_995 ();
 FILLCELL_X16 FILLER_85_1002 ();
 FILLCELL_X4 FILLER_85_1018 ();
 FILLCELL_X2 FILLER_85_1022 ();
 FILLCELL_X32 FILLER_86_1 ();
 FILLCELL_X32 FILLER_86_33 ();
 FILLCELL_X32 FILLER_86_65 ();
 FILLCELL_X32 FILLER_86_97 ();
 FILLCELL_X32 FILLER_86_129 ();
 FILLCELL_X8 FILLER_86_161 ();
 FILLCELL_X4 FILLER_86_819 ();
 FILLCELL_X2 FILLER_86_823 ();
 FILLCELL_X4 FILLER_86_834 ();
 FILLCELL_X4 FILLER_86_842 ();
 FILLCELL_X4 FILLER_86_850 ();
 FILLCELL_X4 FILLER_86_858 ();
 FILLCELL_X4 FILLER_86_865 ();
 FILLCELL_X4 FILLER_86_872 ();
 FILLCELL_X4 FILLER_86_878 ();
 FILLCELL_X4 FILLER_86_884 ();
 FILLCELL_X2 FILLER_86_888 ();
 FILLCELL_X4 FILLER_86_896 ();
 FILLCELL_X4 FILLER_86_904 ();
 FILLCELL_X4 FILLER_86_912 ();
 FILLCELL_X4 FILLER_86_918 ();
 FILLCELL_X4 FILLER_86_926 ();
 FILLCELL_X4 FILLER_86_939 ();
 FILLCELL_X4 FILLER_86_946 ();
 FILLCELL_X4 FILLER_86_957 ();
 FILLCELL_X4 FILLER_86_971 ();
 FILLCELL_X4 FILLER_86_984 ();
 FILLCELL_X4 FILLER_86_991 ();
 FILLCELL_X16 FILLER_86_1005 ();
 FILLCELL_X2 FILLER_86_1021 ();
 FILLCELL_X1 FILLER_86_1023 ();
 FILLCELL_X32 FILLER_87_1 ();
 FILLCELL_X32 FILLER_87_33 ();
 FILLCELL_X32 FILLER_87_65 ();
 FILLCELL_X32 FILLER_87_97 ();
 FILLCELL_X32 FILLER_87_129 ();
 FILLCELL_X8 FILLER_87_161 ();
 FILLCELL_X8 FILLER_87_819 ();
 FILLCELL_X2 FILLER_87_827 ();
 FILLCELL_X4 FILLER_87_838 ();
 FILLCELL_X4 FILLER_87_845 ();
 FILLCELL_X4 FILLER_87_852 ();
 FILLCELL_X1 FILLER_87_856 ();
 FILLCELL_X8 FILLER_87_861 ();
 FILLCELL_X1 FILLER_87_869 ();
 FILLCELL_X4 FILLER_87_872 ();
 FILLCELL_X4 FILLER_87_880 ();
 FILLCELL_X8 FILLER_87_886 ();
 FILLCELL_X2 FILLER_87_894 ();
 FILLCELL_X1 FILLER_87_896 ();
 FILLCELL_X16 FILLER_87_899 ();
 FILLCELL_X1 FILLER_87_915 ();
 FILLCELL_X4 FILLER_87_920 ();
 FILLCELL_X4 FILLER_87_933 ();
 FILLCELL_X4 FILLER_87_940 ();
 FILLCELL_X2 FILLER_87_944 ();
 FILLCELL_X4 FILLER_87_949 ();
 FILLCELL_X32 FILLER_87_955 ();
 FILLCELL_X2 FILLER_87_987 ();
 FILLCELL_X4 FILLER_87_993 ();
 FILLCELL_X4 FILLER_87_1001 ();
 FILLCELL_X8 FILLER_87_1009 ();
 FILLCELL_X4 FILLER_87_1020 ();
 FILLCELL_X32 FILLER_88_1 ();
 FILLCELL_X32 FILLER_88_33 ();
 FILLCELL_X32 FILLER_88_65 ();
 FILLCELL_X32 FILLER_88_97 ();
 FILLCELL_X32 FILLER_88_129 ();
 FILLCELL_X8 FILLER_88_161 ();
 FILLCELL_X4 FILLER_88_819 ();
 FILLCELL_X2 FILLER_88_823 ();
 FILLCELL_X1 FILLER_88_825 ();
 FILLCELL_X4 FILLER_88_829 ();
 FILLCELL_X2 FILLER_88_833 ();
 FILLCELL_X4 FILLER_88_838 ();
 FILLCELL_X2 FILLER_88_842 ();
 FILLCELL_X1 FILLER_88_844 ();
 FILLCELL_X8 FILLER_88_855 ();
 FILLCELL_X4 FILLER_88_873 ();
 FILLCELL_X2 FILLER_88_877 ();
 FILLCELL_X4 FILLER_88_888 ();
 FILLCELL_X4 FILLER_88_895 ();
 FILLCELL_X2 FILLER_88_899 ();
 FILLCELL_X4 FILLER_88_907 ();
 FILLCELL_X4 FILLER_88_921 ();
 FILLCELL_X4 FILLER_88_928 ();
 FILLCELL_X2 FILLER_88_932 ();
 FILLCELL_X1 FILLER_88_934 ();
 FILLCELL_X8 FILLER_88_938 ();
 FILLCELL_X32 FILLER_88_956 ();
 FILLCELL_X4 FILLER_88_988 ();
 FILLCELL_X1 FILLER_88_992 ();
 FILLCELL_X4 FILLER_88_1000 ();
 FILLCELL_X8 FILLER_88_1010 ();
 FILLCELL_X4 FILLER_88_1018 ();
 FILLCELL_X2 FILLER_88_1022 ();
 FILLCELL_X32 FILLER_89_1 ();
 FILLCELL_X32 FILLER_89_33 ();
 FILLCELL_X32 FILLER_89_65 ();
 FILLCELL_X32 FILLER_89_97 ();
 FILLCELL_X32 FILLER_89_129 ();
 FILLCELL_X8 FILLER_89_161 ();
 FILLCELL_X16 FILLER_89_819 ();
 FILLCELL_X2 FILLER_89_835 ();
 FILLCELL_X4 FILLER_89_841 ();
 FILLCELL_X4 FILLER_89_854 ();
 FILLCELL_X8 FILLER_89_865 ();
 FILLCELL_X1 FILLER_89_873 ();
 FILLCELL_X4 FILLER_89_883 ();
 FILLCELL_X4 FILLER_89_890 ();
 FILLCELL_X4 FILLER_89_897 ();
 FILLCELL_X2 FILLER_89_901 ();
 FILLCELL_X1 FILLER_89_903 ();
 FILLCELL_X4 FILLER_89_911 ();
 FILLCELL_X4 FILLER_89_925 ();
 FILLCELL_X8 FILLER_89_935 ();
 FILLCELL_X2 FILLER_89_943 ();
 FILLCELL_X4 FILLER_89_954 ();
 FILLCELL_X4 FILLER_89_962 ();
 FILLCELL_X4 FILLER_89_969 ();
 FILLCELL_X4 FILLER_89_975 ();
 FILLCELL_X4 FILLER_89_989 ();
 FILLCELL_X2 FILLER_89_993 ();
 FILLCELL_X16 FILLER_89_1001 ();
 FILLCELL_X4 FILLER_89_1017 ();
 FILLCELL_X2 FILLER_89_1021 ();
 FILLCELL_X1 FILLER_89_1023 ();
 FILLCELL_X32 FILLER_90_1 ();
 FILLCELL_X32 FILLER_90_33 ();
 FILLCELL_X32 FILLER_90_65 ();
 FILLCELL_X32 FILLER_90_97 ();
 FILLCELL_X32 FILLER_90_129 ();
 FILLCELL_X8 FILLER_90_161 ();
 FILLCELL_X8 FILLER_90_819 ();
 FILLCELL_X1 FILLER_90_827 ();
 FILLCELL_X4 FILLER_90_830 ();
 FILLCELL_X8 FILLER_90_843 ();
 FILLCELL_X4 FILLER_90_854 ();
 FILLCELL_X4 FILLER_90_868 ();
 FILLCELL_X4 FILLER_90_875 ();
 FILLCELL_X4 FILLER_90_881 ();
 FILLCELL_X4 FILLER_90_887 ();
 FILLCELL_X1 FILLER_90_891 ();
 FILLCELL_X4 FILLER_90_902 ();
 FILLCELL_X8 FILLER_90_908 ();
 FILLCELL_X2 FILLER_90_916 ();
 FILLCELL_X4 FILLER_90_925 ();
 FILLCELL_X2 FILLER_90_929 ();
 FILLCELL_X4 FILLER_90_940 ();
 FILLCELL_X1 FILLER_90_944 ();
 FILLCELL_X4 FILLER_90_955 ();
 FILLCELL_X4 FILLER_90_978 ();
 FILLCELL_X16 FILLER_90_985 ();
 FILLCELL_X2 FILLER_90_1001 ();
 FILLCELL_X16 FILLER_90_1007 ();
 FILLCELL_X1 FILLER_90_1023 ();
 FILLCELL_X32 FILLER_91_1 ();
 FILLCELL_X32 FILLER_91_33 ();
 FILLCELL_X32 FILLER_91_65 ();
 FILLCELL_X32 FILLER_91_97 ();
 FILLCELL_X32 FILLER_91_129 ();
 FILLCELL_X8 FILLER_91_161 ();
 FILLCELL_X16 FILLER_91_819 ();
 FILLCELL_X4 FILLER_91_835 ();
 FILLCELL_X4 FILLER_91_849 ();
 FILLCELL_X2 FILLER_91_853 ();
 FILLCELL_X1 FILLER_91_855 ();
 FILLCELL_X4 FILLER_91_863 ();
 FILLCELL_X4 FILLER_91_870 ();
 FILLCELL_X8 FILLER_91_876 ();
 FILLCELL_X2 FILLER_91_884 ();
 FILLCELL_X8 FILLER_91_889 ();
 FILLCELL_X4 FILLER_91_897 ();
 FILLCELL_X8 FILLER_91_911 ();
 FILLCELL_X8 FILLER_91_923 ();
 FILLCELL_X4 FILLER_91_931 ();
 FILLCELL_X4 FILLER_91_938 ();
 FILLCELL_X4 FILLER_91_945 ();
 FILLCELL_X4 FILLER_91_952 ();
 FILLCELL_X8 FILLER_91_963 ();
 FILLCELL_X1 FILLER_91_971 ();
 FILLCELL_X4 FILLER_91_978 ();
 FILLCELL_X4 FILLER_91_989 ();
 FILLCELL_X4 FILLER_91_996 ();
 FILLCELL_X1 FILLER_91_1000 ();
 FILLCELL_X4 FILLER_91_1020 ();
 FILLCELL_X32 FILLER_92_1 ();
 FILLCELL_X32 FILLER_92_33 ();
 FILLCELL_X32 FILLER_92_65 ();
 FILLCELL_X32 FILLER_92_97 ();
 FILLCELL_X32 FILLER_92_129 ();
 FILLCELL_X8 FILLER_92_161 ();
 FILLCELL_X16 FILLER_92_819 ();
 FILLCELL_X2 FILLER_92_835 ();
 FILLCELL_X4 FILLER_92_846 ();
 FILLCELL_X4 FILLER_92_853 ();
 FILLCELL_X8 FILLER_92_860 ();
 FILLCELL_X1 FILLER_92_868 ();
 FILLCELL_X4 FILLER_92_878 ();
 FILLCELL_X2 FILLER_92_882 ();
 FILLCELL_X1 FILLER_92_884 ();
 FILLCELL_X4 FILLER_92_894 ();
 FILLCELL_X8 FILLER_92_902 ();
 FILLCELL_X2 FILLER_92_910 ();
 FILLCELL_X1 FILLER_92_912 ();
 FILLCELL_X16 FILLER_92_915 ();
 FILLCELL_X8 FILLER_92_931 ();
 FILLCELL_X2 FILLER_92_939 ();
 FILLCELL_X1 FILLER_92_941 ();
 FILLCELL_X4 FILLER_92_944 ();
 FILLCELL_X4 FILLER_92_954 ();
 FILLCELL_X1 FILLER_92_958 ();
 FILLCELL_X4 FILLER_92_963 ();
 FILLCELL_X8 FILLER_92_971 ();
 FILLCELL_X2 FILLER_92_979 ();
 FILLCELL_X1 FILLER_92_981 ();
 FILLCELL_X8 FILLER_92_988 ();
 FILLCELL_X8 FILLER_92_1015 ();
 FILLCELL_X1 FILLER_92_1023 ();
 FILLCELL_X4 FILLER_93_1 ();
 FILLCELL_X32 FILLER_93_8 ();
 FILLCELL_X32 FILLER_93_40 ();
 FILLCELL_X32 FILLER_93_72 ();
 FILLCELL_X32 FILLER_93_104 ();
 FILLCELL_X32 FILLER_93_136 ();
 FILLCELL_X1 FILLER_93_168 ();
 FILLCELL_X16 FILLER_93_819 ();
 FILLCELL_X1 FILLER_93_835 ();
 FILLCELL_X16 FILLER_93_840 ();
 FILLCELL_X4 FILLER_93_856 ();
 FILLCELL_X2 FILLER_93_860 ();
 FILLCELL_X4 FILLER_93_869 ();
 FILLCELL_X1 FILLER_93_873 ();
 FILLCELL_X4 FILLER_93_876 ();
 FILLCELL_X4 FILLER_93_884 ();
 FILLCELL_X4 FILLER_93_898 ();
 FILLCELL_X8 FILLER_93_905 ();
 FILLCELL_X4 FILLER_93_913 ();
 FILLCELL_X1 FILLER_93_917 ();
 FILLCELL_X8 FILLER_93_935 ();
 FILLCELL_X4 FILLER_93_943 ();
 FILLCELL_X2 FILLER_93_947 ();
 FILLCELL_X8 FILLER_93_955 ();
 FILLCELL_X1 FILLER_93_963 ();
 FILLCELL_X4 FILLER_93_971 ();
 FILLCELL_X8 FILLER_93_979 ();
 FILLCELL_X2 FILLER_93_987 ();
 FILLCELL_X1 FILLER_93_989 ();
 FILLCELL_X4 FILLER_93_994 ();
 FILLCELL_X2 FILLER_93_998 ();
 FILLCELL_X1 FILLER_93_1000 ();
 FILLCELL_X4 FILLER_93_1018 ();
 FILLCELL_X2 FILLER_93_1022 ();
 FILLCELL_X32 FILLER_94_1 ();
 FILLCELL_X32 FILLER_94_33 ();
 FILLCELL_X32 FILLER_94_65 ();
 FILLCELL_X32 FILLER_94_97 ();
 FILLCELL_X32 FILLER_94_129 ();
 FILLCELL_X8 FILLER_94_161 ();
 FILLCELL_X4 FILLER_94_819 ();
 FILLCELL_X2 FILLER_94_823 ();
 FILLCELL_X1 FILLER_94_825 ();
 FILLCELL_X4 FILLER_94_843 ();
 FILLCELL_X1 FILLER_94_847 ();
 FILLCELL_X4 FILLER_94_854 ();
 FILLCELL_X4 FILLER_94_864 ();
 FILLCELL_X1 FILLER_94_868 ();
 FILLCELL_X4 FILLER_94_879 ();
 FILLCELL_X2 FILLER_94_883 ();
 FILLCELL_X8 FILLER_94_888 ();
 FILLCELL_X2 FILLER_94_896 ();
 FILLCELL_X1 FILLER_94_898 ();
 FILLCELL_X16 FILLER_94_916 ();
 FILLCELL_X8 FILLER_94_932 ();
 FILLCELL_X4 FILLER_94_940 ();
 FILLCELL_X1 FILLER_94_944 ();
 FILLCELL_X32 FILLER_94_964 ();
 FILLCELL_X16 FILLER_94_996 ();
 FILLCELL_X8 FILLER_94_1012 ();
 FILLCELL_X4 FILLER_94_1020 ();
 FILLCELL_X32 FILLER_95_1 ();
 FILLCELL_X32 FILLER_95_33 ();
 FILLCELL_X32 FILLER_95_65 ();
 FILLCELL_X32 FILLER_95_97 ();
 FILLCELL_X32 FILLER_95_129 ();
 FILLCELL_X8 FILLER_95_161 ();
 FILLCELL_X32 FILLER_95_819 ();
 FILLCELL_X4 FILLER_95_851 ();
 FILLCELL_X2 FILLER_95_855 ();
 FILLCELL_X4 FILLER_95_860 ();
 FILLCELL_X32 FILLER_95_867 ();
 FILLCELL_X32 FILLER_95_899 ();
 FILLCELL_X16 FILLER_95_931 ();
 FILLCELL_X4 FILLER_95_947 ();
 FILLCELL_X32 FILLER_95_957 ();
 FILLCELL_X32 FILLER_95_989 ();
 FILLCELL_X2 FILLER_95_1021 ();
 FILLCELL_X1 FILLER_95_1023 ();
 FILLCELL_X32 FILLER_96_1 ();
 FILLCELL_X32 FILLER_96_33 ();
 FILLCELL_X32 FILLER_96_65 ();
 FILLCELL_X32 FILLER_96_97 ();
 FILLCELL_X32 FILLER_96_129 ();
 FILLCELL_X8 FILLER_96_161 ();
 FILLCELL_X32 FILLER_96_819 ();
 FILLCELL_X32 FILLER_96_851 ();
 FILLCELL_X32 FILLER_96_883 ();
 FILLCELL_X32 FILLER_96_915 ();
 FILLCELL_X32 FILLER_96_947 ();
 FILLCELL_X32 FILLER_96_979 ();
 FILLCELL_X8 FILLER_96_1011 ();
 FILLCELL_X4 FILLER_96_1019 ();
 FILLCELL_X1 FILLER_96_1023 ();
 FILLCELL_X32 FILLER_97_1 ();
 FILLCELL_X32 FILLER_97_33 ();
 FILLCELL_X32 FILLER_97_65 ();
 FILLCELL_X32 FILLER_97_97 ();
 FILLCELL_X32 FILLER_97_129 ();
 FILLCELL_X8 FILLER_97_161 ();
 FILLCELL_X32 FILLER_97_819 ();
 FILLCELL_X32 FILLER_97_851 ();
 FILLCELL_X32 FILLER_97_883 ();
 FILLCELL_X32 FILLER_97_915 ();
 FILLCELL_X32 FILLER_97_947 ();
 FILLCELL_X32 FILLER_97_979 ();
 FILLCELL_X8 FILLER_97_1011 ();
 FILLCELL_X4 FILLER_97_1019 ();
 FILLCELL_X1 FILLER_97_1023 ();
 FILLCELL_X32 FILLER_98_1 ();
 FILLCELL_X32 FILLER_98_33 ();
 FILLCELL_X32 FILLER_98_65 ();
 FILLCELL_X32 FILLER_98_97 ();
 FILLCELL_X32 FILLER_98_129 ();
 FILLCELL_X8 FILLER_98_161 ();
 FILLCELL_X32 FILLER_98_819 ();
 FILLCELL_X32 FILLER_98_851 ();
 FILLCELL_X32 FILLER_98_883 ();
 FILLCELL_X32 FILLER_98_915 ();
 FILLCELL_X32 FILLER_98_947 ();
 FILLCELL_X32 FILLER_98_979 ();
 FILLCELL_X4 FILLER_98_1011 ();
 FILLCELL_X2 FILLER_98_1015 ();
 FILLCELL_X4 FILLER_98_1020 ();
 FILLCELL_X32 FILLER_99_1 ();
 FILLCELL_X32 FILLER_99_33 ();
 FILLCELL_X32 FILLER_99_65 ();
 FILLCELL_X32 FILLER_99_97 ();
 FILLCELL_X32 FILLER_99_129 ();
 FILLCELL_X8 FILLER_99_161 ();
 FILLCELL_X32 FILLER_99_819 ();
 FILLCELL_X32 FILLER_99_851 ();
 FILLCELL_X32 FILLER_99_883 ();
 FILLCELL_X32 FILLER_99_915 ();
 FILLCELL_X32 FILLER_99_947 ();
 FILLCELL_X32 FILLER_99_979 ();
 FILLCELL_X8 FILLER_99_1011 ();
 FILLCELL_X4 FILLER_99_1019 ();
 FILLCELL_X1 FILLER_99_1023 ();
 FILLCELL_X32 FILLER_100_1 ();
 FILLCELL_X32 FILLER_100_33 ();
 FILLCELL_X32 FILLER_100_65 ();
 FILLCELL_X32 FILLER_100_97 ();
 FILLCELL_X32 FILLER_100_129 ();
 FILLCELL_X8 FILLER_100_161 ();
 FILLCELL_X32 FILLER_100_819 ();
 FILLCELL_X32 FILLER_100_851 ();
 FILLCELL_X32 FILLER_100_883 ();
 FILLCELL_X32 FILLER_100_915 ();
 FILLCELL_X32 FILLER_100_947 ();
 FILLCELL_X32 FILLER_100_979 ();
 FILLCELL_X8 FILLER_100_1011 ();
 FILLCELL_X4 FILLER_100_1019 ();
 FILLCELL_X1 FILLER_100_1023 ();
 FILLCELL_X32 FILLER_101_1 ();
 FILLCELL_X32 FILLER_101_33 ();
 FILLCELL_X32 FILLER_101_65 ();
 FILLCELL_X32 FILLER_101_97 ();
 FILLCELL_X32 FILLER_101_129 ();
 FILLCELL_X8 FILLER_101_161 ();
 FILLCELL_X32 FILLER_101_819 ();
 FILLCELL_X32 FILLER_101_851 ();
 FILLCELL_X32 FILLER_101_883 ();
 FILLCELL_X32 FILLER_101_915 ();
 FILLCELL_X32 FILLER_101_947 ();
 FILLCELL_X32 FILLER_101_979 ();
 FILLCELL_X8 FILLER_101_1011 ();
 FILLCELL_X4 FILLER_101_1019 ();
 FILLCELL_X1 FILLER_101_1023 ();
 FILLCELL_X32 FILLER_102_1 ();
 FILLCELL_X32 FILLER_102_33 ();
 FILLCELL_X32 FILLER_102_65 ();
 FILLCELL_X32 FILLER_102_97 ();
 FILLCELL_X32 FILLER_102_129 ();
 FILLCELL_X8 FILLER_102_161 ();
 FILLCELL_X32 FILLER_102_819 ();
 FILLCELL_X32 FILLER_102_851 ();
 FILLCELL_X32 FILLER_102_883 ();
 FILLCELL_X32 FILLER_102_915 ();
 FILLCELL_X32 FILLER_102_947 ();
 FILLCELL_X32 FILLER_102_979 ();
 FILLCELL_X8 FILLER_102_1011 ();
 FILLCELL_X4 FILLER_102_1019 ();
 FILLCELL_X1 FILLER_102_1023 ();
 FILLCELL_X32 FILLER_103_1 ();
 FILLCELL_X32 FILLER_103_33 ();
 FILLCELL_X32 FILLER_103_65 ();
 FILLCELL_X32 FILLER_103_97 ();
 FILLCELL_X32 FILLER_103_129 ();
 FILLCELL_X8 FILLER_103_161 ();
 FILLCELL_X32 FILLER_103_819 ();
 FILLCELL_X32 FILLER_103_851 ();
 FILLCELL_X32 FILLER_103_883 ();
 FILLCELL_X32 FILLER_103_915 ();
 FILLCELL_X32 FILLER_103_947 ();
 FILLCELL_X32 FILLER_103_979 ();
 FILLCELL_X8 FILLER_103_1011 ();
 FILLCELL_X4 FILLER_103_1019 ();
 FILLCELL_X1 FILLER_103_1023 ();
 FILLCELL_X32 FILLER_104_1 ();
 FILLCELL_X32 FILLER_104_33 ();
 FILLCELL_X32 FILLER_104_65 ();
 FILLCELL_X32 FILLER_104_97 ();
 FILLCELL_X32 FILLER_104_129 ();
 FILLCELL_X8 FILLER_104_161 ();
 FILLCELL_X32 FILLER_104_819 ();
 FILLCELL_X32 FILLER_104_851 ();
 FILLCELL_X32 FILLER_104_883 ();
 FILLCELL_X32 FILLER_104_915 ();
 FILLCELL_X32 FILLER_104_947 ();
 FILLCELL_X32 FILLER_104_979 ();
 FILLCELL_X8 FILLER_104_1011 ();
 FILLCELL_X4 FILLER_104_1019 ();
 FILLCELL_X1 FILLER_104_1023 ();
 FILLCELL_X32 FILLER_105_1 ();
 FILLCELL_X32 FILLER_105_33 ();
 FILLCELL_X32 FILLER_105_65 ();
 FILLCELL_X32 FILLER_105_97 ();
 FILLCELL_X32 FILLER_105_129 ();
 FILLCELL_X8 FILLER_105_161 ();
 FILLCELL_X32 FILLER_105_819 ();
 FILLCELL_X32 FILLER_105_851 ();
 FILLCELL_X32 FILLER_105_883 ();
 FILLCELL_X32 FILLER_105_915 ();
 FILLCELL_X32 FILLER_105_947 ();
 FILLCELL_X32 FILLER_105_979 ();
 FILLCELL_X8 FILLER_105_1011 ();
 FILLCELL_X4 FILLER_105_1019 ();
 FILLCELL_X1 FILLER_105_1023 ();
 FILLCELL_X32 FILLER_106_1 ();
 FILLCELL_X32 FILLER_106_33 ();
 FILLCELL_X32 FILLER_106_65 ();
 FILLCELL_X32 FILLER_106_97 ();
 FILLCELL_X32 FILLER_106_129 ();
 FILLCELL_X8 FILLER_106_161 ();
 FILLCELL_X32 FILLER_106_819 ();
 FILLCELL_X32 FILLER_106_851 ();
 FILLCELL_X32 FILLER_106_883 ();
 FILLCELL_X32 FILLER_106_915 ();
 FILLCELL_X32 FILLER_106_947 ();
 FILLCELL_X32 FILLER_106_979 ();
 FILLCELL_X8 FILLER_106_1011 ();
 FILLCELL_X4 FILLER_106_1019 ();
 FILLCELL_X1 FILLER_106_1023 ();
 FILLCELL_X32 FILLER_107_1 ();
 FILLCELL_X32 FILLER_107_33 ();
 FILLCELL_X32 FILLER_107_65 ();
 FILLCELL_X32 FILLER_107_97 ();
 FILLCELL_X32 FILLER_107_129 ();
 FILLCELL_X8 FILLER_107_161 ();
 FILLCELL_X32 FILLER_107_819 ();
 FILLCELL_X32 FILLER_107_851 ();
 FILLCELL_X32 FILLER_107_883 ();
 FILLCELL_X32 FILLER_107_915 ();
 FILLCELL_X32 FILLER_107_947 ();
 FILLCELL_X32 FILLER_107_979 ();
 FILLCELL_X8 FILLER_107_1011 ();
 FILLCELL_X4 FILLER_107_1019 ();
 FILLCELL_X1 FILLER_107_1023 ();
 FILLCELL_X32 FILLER_108_1 ();
 FILLCELL_X32 FILLER_108_33 ();
 FILLCELL_X32 FILLER_108_65 ();
 FILLCELL_X32 FILLER_108_97 ();
 FILLCELL_X32 FILLER_108_129 ();
 FILLCELL_X8 FILLER_108_161 ();
 FILLCELL_X32 FILLER_108_819 ();
 FILLCELL_X32 FILLER_108_851 ();
 FILLCELL_X32 FILLER_108_883 ();
 FILLCELL_X32 FILLER_108_915 ();
 FILLCELL_X32 FILLER_108_947 ();
 FILLCELL_X32 FILLER_108_979 ();
 FILLCELL_X8 FILLER_108_1011 ();
 FILLCELL_X4 FILLER_108_1019 ();
 FILLCELL_X1 FILLER_108_1023 ();
 FILLCELL_X32 FILLER_109_1 ();
 FILLCELL_X32 FILLER_109_33 ();
 FILLCELL_X32 FILLER_109_65 ();
 FILLCELL_X32 FILLER_109_97 ();
 FILLCELL_X32 FILLER_109_129 ();
 FILLCELL_X8 FILLER_109_161 ();
 FILLCELL_X32 FILLER_109_819 ();
 FILLCELL_X32 FILLER_109_851 ();
 FILLCELL_X32 FILLER_109_883 ();
 FILLCELL_X32 FILLER_109_915 ();
 FILLCELL_X32 FILLER_109_947 ();
 FILLCELL_X32 FILLER_109_979 ();
 FILLCELL_X4 FILLER_109_1011 ();
 FILLCELL_X2 FILLER_109_1015 ();
 FILLCELL_X4 FILLER_109_1020 ();
 FILLCELL_X32 FILLER_110_1 ();
 FILLCELL_X32 FILLER_110_33 ();
 FILLCELL_X32 FILLER_110_65 ();
 FILLCELL_X32 FILLER_110_97 ();
 FILLCELL_X32 FILLER_110_129 ();
 FILLCELL_X8 FILLER_110_161 ();
 FILLCELL_X32 FILLER_110_819 ();
 FILLCELL_X32 FILLER_110_851 ();
 FILLCELL_X32 FILLER_110_883 ();
 FILLCELL_X32 FILLER_110_915 ();
 FILLCELL_X32 FILLER_110_947 ();
 FILLCELL_X32 FILLER_110_979 ();
 FILLCELL_X8 FILLER_110_1011 ();
 FILLCELL_X4 FILLER_110_1019 ();
 FILLCELL_X1 FILLER_110_1023 ();
 FILLCELL_X32 FILLER_111_1 ();
 FILLCELL_X32 FILLER_111_33 ();
 FILLCELL_X32 FILLER_111_65 ();
 FILLCELL_X32 FILLER_111_97 ();
 FILLCELL_X32 FILLER_111_129 ();
 FILLCELL_X8 FILLER_111_161 ();
 FILLCELL_X32 FILLER_111_819 ();
 FILLCELL_X32 FILLER_111_851 ();
 FILLCELL_X32 FILLER_111_883 ();
 FILLCELL_X32 FILLER_111_915 ();
 FILLCELL_X32 FILLER_111_947 ();
 FILLCELL_X32 FILLER_111_979 ();
 FILLCELL_X8 FILLER_111_1011 ();
 FILLCELL_X4 FILLER_111_1019 ();
 FILLCELL_X1 FILLER_111_1023 ();
 FILLCELL_X32 FILLER_112_1 ();
 FILLCELL_X32 FILLER_112_33 ();
 FILLCELL_X32 FILLER_112_65 ();
 FILLCELL_X32 FILLER_112_97 ();
 FILLCELL_X32 FILLER_112_129 ();
 FILLCELL_X8 FILLER_112_161 ();
 FILLCELL_X32 FILLER_112_819 ();
 FILLCELL_X32 FILLER_112_851 ();
 FILLCELL_X32 FILLER_112_883 ();
 FILLCELL_X32 FILLER_112_915 ();
 FILLCELL_X32 FILLER_112_947 ();
 FILLCELL_X32 FILLER_112_979 ();
 FILLCELL_X8 FILLER_112_1011 ();
 FILLCELL_X4 FILLER_112_1019 ();
 FILLCELL_X1 FILLER_112_1023 ();
 FILLCELL_X32 FILLER_113_1 ();
 FILLCELL_X32 FILLER_113_33 ();
 FILLCELL_X32 FILLER_113_65 ();
 FILLCELL_X32 FILLER_113_97 ();
 FILLCELL_X32 FILLER_113_129 ();
 FILLCELL_X8 FILLER_113_161 ();
 FILLCELL_X32 FILLER_113_819 ();
 FILLCELL_X32 FILLER_113_851 ();
 FILLCELL_X32 FILLER_113_883 ();
 FILLCELL_X32 FILLER_113_915 ();
 FILLCELL_X32 FILLER_113_947 ();
 FILLCELL_X32 FILLER_113_979 ();
 FILLCELL_X8 FILLER_113_1011 ();
 FILLCELL_X4 FILLER_113_1019 ();
 FILLCELL_X1 FILLER_113_1023 ();
 FILLCELL_X4 FILLER_114_1 ();
 FILLCELL_X32 FILLER_114_8 ();
 FILLCELL_X32 FILLER_114_40 ();
 FILLCELL_X32 FILLER_114_72 ();
 FILLCELL_X32 FILLER_114_104 ();
 FILLCELL_X32 FILLER_114_136 ();
 FILLCELL_X1 FILLER_114_168 ();
 FILLCELL_X32 FILLER_114_819 ();
 FILLCELL_X32 FILLER_114_851 ();
 FILLCELL_X32 FILLER_114_883 ();
 FILLCELL_X32 FILLER_114_915 ();
 FILLCELL_X32 FILLER_114_947 ();
 FILLCELL_X32 FILLER_114_979 ();
 FILLCELL_X8 FILLER_114_1011 ();
 FILLCELL_X4 FILLER_114_1019 ();
 FILLCELL_X1 FILLER_114_1023 ();
 FILLCELL_X32 FILLER_115_1 ();
 FILLCELL_X32 FILLER_115_33 ();
 FILLCELL_X32 FILLER_115_65 ();
 FILLCELL_X32 FILLER_115_97 ();
 FILLCELL_X32 FILLER_115_129 ();
 FILLCELL_X8 FILLER_115_161 ();
 FILLCELL_X32 FILLER_115_819 ();
 FILLCELL_X32 FILLER_115_851 ();
 FILLCELL_X32 FILLER_115_883 ();
 FILLCELL_X32 FILLER_115_915 ();
 FILLCELL_X32 FILLER_115_947 ();
 FILLCELL_X32 FILLER_115_979 ();
 FILLCELL_X8 FILLER_115_1011 ();
 FILLCELL_X4 FILLER_115_1019 ();
 FILLCELL_X1 FILLER_115_1023 ();
 FILLCELL_X32 FILLER_116_1 ();
 FILLCELL_X32 FILLER_116_33 ();
 FILLCELL_X32 FILLER_116_65 ();
 FILLCELL_X32 FILLER_116_97 ();
 FILLCELL_X32 FILLER_116_129 ();
 FILLCELL_X8 FILLER_116_161 ();
 FILLCELL_X32 FILLER_116_819 ();
 FILLCELL_X32 FILLER_116_851 ();
 FILLCELL_X32 FILLER_116_883 ();
 FILLCELL_X32 FILLER_116_915 ();
 FILLCELL_X32 FILLER_116_947 ();
 FILLCELL_X32 FILLER_116_979 ();
 FILLCELL_X8 FILLER_116_1011 ();
 FILLCELL_X4 FILLER_116_1019 ();
 FILLCELL_X1 FILLER_116_1023 ();
 FILLCELL_X32 FILLER_117_1 ();
 FILLCELL_X32 FILLER_117_33 ();
 FILLCELL_X32 FILLER_117_65 ();
 FILLCELL_X32 FILLER_117_97 ();
 FILLCELL_X32 FILLER_117_129 ();
 FILLCELL_X32 FILLER_117_161 ();
 FILLCELL_X32 FILLER_117_193 ();
 FILLCELL_X32 FILLER_117_225 ();
 FILLCELL_X32 FILLER_117_257 ();
 FILLCELL_X32 FILLER_117_289 ();
 FILLCELL_X32 FILLER_117_321 ();
 FILLCELL_X32 FILLER_117_353 ();
 FILLCELL_X32 FILLER_117_385 ();
 FILLCELL_X32 FILLER_117_417 ();
 FILLCELL_X32 FILLER_117_449 ();
 FILLCELL_X32 FILLER_117_481 ();
 FILLCELL_X32 FILLER_117_513 ();
 FILLCELL_X32 FILLER_117_545 ();
 FILLCELL_X32 FILLER_117_577 ();
 FILLCELL_X16 FILLER_117_609 ();
 FILLCELL_X4 FILLER_117_625 ();
 FILLCELL_X2 FILLER_117_629 ();
 FILLCELL_X32 FILLER_117_632 ();
 FILLCELL_X32 FILLER_117_664 ();
 FILLCELL_X32 FILLER_117_696 ();
 FILLCELL_X32 FILLER_117_728 ();
 FILLCELL_X32 FILLER_117_760 ();
 FILLCELL_X32 FILLER_117_792 ();
 FILLCELL_X32 FILLER_117_824 ();
 FILLCELL_X32 FILLER_117_856 ();
 FILLCELL_X32 FILLER_117_888 ();
 FILLCELL_X32 FILLER_117_920 ();
 FILLCELL_X32 FILLER_117_952 ();
 FILLCELL_X32 FILLER_117_984 ();
 FILLCELL_X8 FILLER_117_1016 ();
 FILLCELL_X32 FILLER_118_1 ();
 FILLCELL_X32 FILLER_118_33 ();
 FILLCELL_X32 FILLER_118_65 ();
 FILLCELL_X32 FILLER_118_97 ();
 FILLCELL_X32 FILLER_118_129 ();
 FILLCELL_X32 FILLER_118_161 ();
 FILLCELL_X32 FILLER_118_193 ();
 FILLCELL_X32 FILLER_118_225 ();
 FILLCELL_X32 FILLER_118_257 ();
 FILLCELL_X32 FILLER_118_289 ();
 FILLCELL_X32 FILLER_118_321 ();
 FILLCELL_X32 FILLER_118_353 ();
 FILLCELL_X32 FILLER_118_385 ();
 FILLCELL_X32 FILLER_118_417 ();
 FILLCELL_X32 FILLER_118_449 ();
 FILLCELL_X32 FILLER_118_481 ();
 FILLCELL_X32 FILLER_118_513 ();
 FILLCELL_X32 FILLER_118_545 ();
 FILLCELL_X32 FILLER_118_577 ();
 FILLCELL_X16 FILLER_118_609 ();
 FILLCELL_X4 FILLER_118_625 ();
 FILLCELL_X2 FILLER_118_629 ();
 FILLCELL_X32 FILLER_118_632 ();
 FILLCELL_X32 FILLER_118_664 ();
 FILLCELL_X32 FILLER_118_696 ();
 FILLCELL_X32 FILLER_118_728 ();
 FILLCELL_X32 FILLER_118_760 ();
 FILLCELL_X32 FILLER_118_792 ();
 FILLCELL_X32 FILLER_118_824 ();
 FILLCELL_X32 FILLER_118_856 ();
 FILLCELL_X32 FILLER_118_888 ();
 FILLCELL_X32 FILLER_118_920 ();
 FILLCELL_X32 FILLER_118_952 ();
 FILLCELL_X32 FILLER_118_984 ();
 FILLCELL_X8 FILLER_118_1016 ();
 FILLCELL_X32 FILLER_119_1 ();
 FILLCELL_X32 FILLER_119_33 ();
 FILLCELL_X32 FILLER_119_65 ();
 FILLCELL_X32 FILLER_119_97 ();
 FILLCELL_X32 FILLER_119_129 ();
 FILLCELL_X32 FILLER_119_161 ();
 FILLCELL_X32 FILLER_119_193 ();
 FILLCELL_X32 FILLER_119_225 ();
 FILLCELL_X32 FILLER_119_257 ();
 FILLCELL_X32 FILLER_119_289 ();
 FILLCELL_X32 FILLER_119_321 ();
 FILLCELL_X32 FILLER_119_353 ();
 FILLCELL_X32 FILLER_119_385 ();
 FILLCELL_X32 FILLER_119_417 ();
 FILLCELL_X32 FILLER_119_449 ();
 FILLCELL_X32 FILLER_119_481 ();
 FILLCELL_X32 FILLER_119_513 ();
 FILLCELL_X32 FILLER_119_545 ();
 FILLCELL_X32 FILLER_119_577 ();
 FILLCELL_X32 FILLER_119_609 ();
 FILLCELL_X32 FILLER_119_641 ();
 FILLCELL_X32 FILLER_119_673 ();
 FILLCELL_X32 FILLER_119_705 ();
 FILLCELL_X32 FILLER_119_737 ();
 FILLCELL_X32 FILLER_119_769 ();
 FILLCELL_X32 FILLER_119_801 ();
 FILLCELL_X32 FILLER_119_833 ();
 FILLCELL_X32 FILLER_119_865 ();
 FILLCELL_X32 FILLER_119_897 ();
 FILLCELL_X32 FILLER_119_929 ();
 FILLCELL_X32 FILLER_119_961 ();
 FILLCELL_X16 FILLER_119_993 ();
 FILLCELL_X8 FILLER_119_1009 ();
 FILLCELL_X4 FILLER_119_1017 ();
 FILLCELL_X2 FILLER_119_1021 ();
 FILLCELL_X1 FILLER_119_1023 ();
 FILLCELL_X32 FILLER_120_1 ();
 FILLCELL_X32 FILLER_120_33 ();
 FILLCELL_X32 FILLER_120_65 ();
 FILLCELL_X32 FILLER_120_97 ();
 FILLCELL_X32 FILLER_120_129 ();
 FILLCELL_X32 FILLER_120_161 ();
 FILLCELL_X32 FILLER_120_193 ();
 FILLCELL_X32 FILLER_120_225 ();
 FILLCELL_X32 FILLER_120_257 ();
 FILLCELL_X32 FILLER_120_289 ();
 FILLCELL_X32 FILLER_120_321 ();
 FILLCELL_X32 FILLER_120_353 ();
 FILLCELL_X32 FILLER_120_385 ();
 FILLCELL_X32 FILLER_120_417 ();
 FILLCELL_X32 FILLER_120_449 ();
 FILLCELL_X32 FILLER_120_481 ();
 FILLCELL_X32 FILLER_120_513 ();
 FILLCELL_X32 FILLER_120_545 ();
 FILLCELL_X32 FILLER_120_577 ();
 FILLCELL_X16 FILLER_120_609 ();
 FILLCELL_X4 FILLER_120_625 ();
 FILLCELL_X2 FILLER_120_629 ();
 FILLCELL_X32 FILLER_120_632 ();
 FILLCELL_X32 FILLER_120_664 ();
 FILLCELL_X32 FILLER_120_696 ();
 FILLCELL_X32 FILLER_120_728 ();
 FILLCELL_X32 FILLER_120_760 ();
 FILLCELL_X32 FILLER_120_792 ();
 FILLCELL_X32 FILLER_120_824 ();
 FILLCELL_X32 FILLER_120_856 ();
 FILLCELL_X32 FILLER_120_888 ();
 FILLCELL_X32 FILLER_120_920 ();
 FILLCELL_X32 FILLER_120_952 ();
 FILLCELL_X32 FILLER_120_984 ();
 FILLCELL_X1 FILLER_120_1016 ();
 FILLCELL_X4 FILLER_120_1020 ();
 FILLCELL_X32 FILLER_121_1 ();
 FILLCELL_X32 FILLER_121_33 ();
 FILLCELL_X32 FILLER_121_65 ();
 FILLCELL_X32 FILLER_121_97 ();
 FILLCELL_X32 FILLER_121_129 ();
 FILLCELL_X32 FILLER_121_161 ();
 FILLCELL_X32 FILLER_121_193 ();
 FILLCELL_X32 FILLER_121_225 ();
 FILLCELL_X32 FILLER_121_257 ();
 FILLCELL_X32 FILLER_121_289 ();
 FILLCELL_X32 FILLER_121_321 ();
 FILLCELL_X32 FILLER_121_353 ();
 FILLCELL_X32 FILLER_121_385 ();
 FILLCELL_X32 FILLER_121_417 ();
 FILLCELL_X32 FILLER_121_449 ();
 FILLCELL_X32 FILLER_121_481 ();
 FILLCELL_X32 FILLER_121_513 ();
 FILLCELL_X32 FILLER_121_545 ();
 FILLCELL_X32 FILLER_121_577 ();
 FILLCELL_X32 FILLER_121_609 ();
 FILLCELL_X32 FILLER_121_641 ();
 FILLCELL_X32 FILLER_121_673 ();
 FILLCELL_X32 FILLER_121_705 ();
 FILLCELL_X32 FILLER_121_737 ();
 FILLCELL_X32 FILLER_121_769 ();
 FILLCELL_X32 FILLER_121_801 ();
 FILLCELL_X32 FILLER_121_833 ();
 FILLCELL_X32 FILLER_121_865 ();
 FILLCELL_X32 FILLER_121_897 ();
 FILLCELL_X32 FILLER_121_929 ();
 FILLCELL_X32 FILLER_121_961 ();
 FILLCELL_X16 FILLER_121_993 ();
 FILLCELL_X8 FILLER_121_1009 ();
 FILLCELL_X4 FILLER_121_1017 ();
 FILLCELL_X2 FILLER_121_1021 ();
 FILLCELL_X1 FILLER_121_1023 ();
 FILLCELL_X32 FILLER_122_1 ();
 FILLCELL_X32 FILLER_122_33 ();
 FILLCELL_X32 FILLER_122_65 ();
 FILLCELL_X32 FILLER_122_97 ();
 FILLCELL_X32 FILLER_122_129 ();
 FILLCELL_X32 FILLER_122_161 ();
 FILLCELL_X32 FILLER_122_193 ();
 FILLCELL_X32 FILLER_122_225 ();
 FILLCELL_X32 FILLER_122_257 ();
 FILLCELL_X32 FILLER_122_289 ();
 FILLCELL_X32 FILLER_122_321 ();
 FILLCELL_X32 FILLER_122_353 ();
 FILLCELL_X32 FILLER_122_385 ();
 FILLCELL_X32 FILLER_122_417 ();
 FILLCELL_X32 FILLER_122_449 ();
 FILLCELL_X32 FILLER_122_481 ();
 FILLCELL_X32 FILLER_122_513 ();
 FILLCELL_X32 FILLER_122_545 ();
 FILLCELL_X32 FILLER_122_577 ();
 FILLCELL_X16 FILLER_122_609 ();
 FILLCELL_X4 FILLER_122_625 ();
 FILLCELL_X2 FILLER_122_629 ();
 FILLCELL_X32 FILLER_122_632 ();
 FILLCELL_X32 FILLER_122_664 ();
 FILLCELL_X32 FILLER_122_696 ();
 FILLCELL_X32 FILLER_122_728 ();
 FILLCELL_X32 FILLER_122_760 ();
 FILLCELL_X32 FILLER_122_792 ();
 FILLCELL_X32 FILLER_122_824 ();
 FILLCELL_X32 FILLER_122_856 ();
 FILLCELL_X32 FILLER_122_888 ();
 FILLCELL_X32 FILLER_122_920 ();
 FILLCELL_X32 FILLER_122_952 ();
 FILLCELL_X32 FILLER_122_984 ();
 FILLCELL_X8 FILLER_122_1016 ();
 FILLCELL_X32 FILLER_123_1 ();
 FILLCELL_X32 FILLER_123_33 ();
 FILLCELL_X32 FILLER_123_65 ();
 FILLCELL_X32 FILLER_123_97 ();
 FILLCELL_X32 FILLER_123_129 ();
 FILLCELL_X32 FILLER_123_161 ();
 FILLCELL_X32 FILLER_123_193 ();
 FILLCELL_X32 FILLER_123_225 ();
 FILLCELL_X32 FILLER_123_257 ();
 FILLCELL_X32 FILLER_123_289 ();
 FILLCELL_X32 FILLER_123_321 ();
 FILLCELL_X32 FILLER_123_353 ();
 FILLCELL_X32 FILLER_123_385 ();
 FILLCELL_X32 FILLER_123_417 ();
 FILLCELL_X32 FILLER_123_449 ();
 FILLCELL_X32 FILLER_123_481 ();
 FILLCELL_X32 FILLER_123_513 ();
 FILLCELL_X32 FILLER_123_545 ();
 FILLCELL_X32 FILLER_123_577 ();
 FILLCELL_X32 FILLER_123_609 ();
 FILLCELL_X32 FILLER_123_641 ();
 FILLCELL_X32 FILLER_123_673 ();
 FILLCELL_X32 FILLER_123_705 ();
 FILLCELL_X32 FILLER_123_737 ();
 FILLCELL_X32 FILLER_123_769 ();
 FILLCELL_X32 FILLER_123_801 ();
 FILLCELL_X32 FILLER_123_833 ();
 FILLCELL_X32 FILLER_123_865 ();
 FILLCELL_X32 FILLER_123_897 ();
 FILLCELL_X32 FILLER_123_929 ();
 FILLCELL_X32 FILLER_123_961 ();
 FILLCELL_X16 FILLER_123_993 ();
 FILLCELL_X8 FILLER_123_1009 ();
 FILLCELL_X4 FILLER_123_1017 ();
 FILLCELL_X2 FILLER_123_1021 ();
 FILLCELL_X1 FILLER_123_1023 ();
 FILLCELL_X32 FILLER_124_1 ();
 FILLCELL_X32 FILLER_124_33 ();
 FILLCELL_X32 FILLER_124_65 ();
 FILLCELL_X32 FILLER_124_97 ();
 FILLCELL_X32 FILLER_124_129 ();
 FILLCELL_X32 FILLER_124_161 ();
 FILLCELL_X32 FILLER_124_193 ();
 FILLCELL_X32 FILLER_124_225 ();
 FILLCELL_X32 FILLER_124_257 ();
 FILLCELL_X32 FILLER_124_289 ();
 FILLCELL_X32 FILLER_124_321 ();
 FILLCELL_X32 FILLER_124_353 ();
 FILLCELL_X32 FILLER_124_385 ();
 FILLCELL_X32 FILLER_124_417 ();
 FILLCELL_X32 FILLER_124_449 ();
 FILLCELL_X32 FILLER_124_481 ();
 FILLCELL_X32 FILLER_124_513 ();
 FILLCELL_X32 FILLER_124_545 ();
 FILLCELL_X32 FILLER_124_577 ();
 FILLCELL_X16 FILLER_124_609 ();
 FILLCELL_X4 FILLER_124_625 ();
 FILLCELL_X2 FILLER_124_629 ();
 FILLCELL_X32 FILLER_124_632 ();
 FILLCELL_X32 FILLER_124_664 ();
 FILLCELL_X32 FILLER_124_696 ();
 FILLCELL_X32 FILLER_124_728 ();
 FILLCELL_X32 FILLER_124_760 ();
 FILLCELL_X32 FILLER_124_792 ();
 FILLCELL_X32 FILLER_124_824 ();
 FILLCELL_X32 FILLER_124_856 ();
 FILLCELL_X32 FILLER_124_888 ();
 FILLCELL_X32 FILLER_124_920 ();
 FILLCELL_X32 FILLER_124_952 ();
 FILLCELL_X32 FILLER_124_984 ();
 FILLCELL_X8 FILLER_124_1016 ();
 FILLCELL_X4 FILLER_125_1 ();
 FILLCELL_X32 FILLER_125_18 ();
 FILLCELL_X32 FILLER_125_50 ();
 FILLCELL_X32 FILLER_125_82 ();
 FILLCELL_X32 FILLER_125_114 ();
 FILLCELL_X32 FILLER_125_146 ();
 FILLCELL_X32 FILLER_125_178 ();
 FILLCELL_X32 FILLER_125_210 ();
 FILLCELL_X32 FILLER_125_242 ();
 FILLCELL_X32 FILLER_125_274 ();
 FILLCELL_X32 FILLER_125_306 ();
 FILLCELL_X32 FILLER_125_338 ();
 FILLCELL_X32 FILLER_125_370 ();
 FILLCELL_X32 FILLER_125_402 ();
 FILLCELL_X32 FILLER_125_434 ();
 FILLCELL_X32 FILLER_125_466 ();
 FILLCELL_X32 FILLER_125_498 ();
 FILLCELL_X32 FILLER_125_530 ();
 FILLCELL_X32 FILLER_125_562 ();
 FILLCELL_X32 FILLER_125_594 ();
 FILLCELL_X32 FILLER_125_626 ();
 FILLCELL_X32 FILLER_125_658 ();
 FILLCELL_X32 FILLER_125_690 ();
 FILLCELL_X32 FILLER_125_722 ();
 FILLCELL_X32 FILLER_125_754 ();
 FILLCELL_X32 FILLER_125_786 ();
 FILLCELL_X32 FILLER_125_818 ();
 FILLCELL_X32 FILLER_125_850 ();
 FILLCELL_X32 FILLER_125_882 ();
 FILLCELL_X32 FILLER_125_914 ();
 FILLCELL_X32 FILLER_125_946 ();
 FILLCELL_X32 FILLER_125_978 ();
 FILLCELL_X8 FILLER_125_1010 ();
 FILLCELL_X4 FILLER_125_1018 ();
 FILLCELL_X2 FILLER_125_1022 ();
 FILLCELL_X32 FILLER_126_1 ();
 FILLCELL_X32 FILLER_126_33 ();
 FILLCELL_X32 FILLER_126_65 ();
 FILLCELL_X32 FILLER_126_97 ();
 FILLCELL_X32 FILLER_126_129 ();
 FILLCELL_X32 FILLER_126_161 ();
 FILLCELL_X32 FILLER_126_193 ();
 FILLCELL_X32 FILLER_126_225 ();
 FILLCELL_X32 FILLER_126_257 ();
 FILLCELL_X32 FILLER_126_289 ();
 FILLCELL_X32 FILLER_126_321 ();
 FILLCELL_X32 FILLER_126_353 ();
 FILLCELL_X32 FILLER_126_385 ();
 FILLCELL_X32 FILLER_126_417 ();
 FILLCELL_X32 FILLER_126_449 ();
 FILLCELL_X32 FILLER_126_481 ();
 FILLCELL_X32 FILLER_126_513 ();
 FILLCELL_X32 FILLER_126_545 ();
 FILLCELL_X32 FILLER_126_577 ();
 FILLCELL_X16 FILLER_126_609 ();
 FILLCELL_X4 FILLER_126_625 ();
 FILLCELL_X2 FILLER_126_629 ();
 FILLCELL_X32 FILLER_126_632 ();
 FILLCELL_X32 FILLER_126_664 ();
 FILLCELL_X32 FILLER_126_696 ();
 FILLCELL_X32 FILLER_126_728 ();
 FILLCELL_X32 FILLER_126_760 ();
 FILLCELL_X32 FILLER_126_792 ();
 FILLCELL_X32 FILLER_126_824 ();
 FILLCELL_X32 FILLER_126_856 ();
 FILLCELL_X32 FILLER_126_888 ();
 FILLCELL_X32 FILLER_126_920 ();
 FILLCELL_X32 FILLER_126_952 ();
 FILLCELL_X32 FILLER_126_984 ();
 FILLCELL_X8 FILLER_126_1016 ();
 FILLCELL_X32 FILLER_127_1 ();
 FILLCELL_X32 FILLER_127_33 ();
 FILLCELL_X32 FILLER_127_65 ();
 FILLCELL_X32 FILLER_127_97 ();
 FILLCELL_X32 FILLER_127_129 ();
 FILLCELL_X32 FILLER_127_161 ();
 FILLCELL_X32 FILLER_127_193 ();
 FILLCELL_X32 FILLER_127_225 ();
 FILLCELL_X32 FILLER_127_257 ();
 FILLCELL_X32 FILLER_127_289 ();
 FILLCELL_X32 FILLER_127_321 ();
 FILLCELL_X32 FILLER_127_353 ();
 FILLCELL_X32 FILLER_127_385 ();
 FILLCELL_X32 FILLER_127_417 ();
 FILLCELL_X32 FILLER_127_449 ();
 FILLCELL_X32 FILLER_127_481 ();
 FILLCELL_X32 FILLER_127_513 ();
 FILLCELL_X32 FILLER_127_545 ();
 FILLCELL_X32 FILLER_127_577 ();
 FILLCELL_X32 FILLER_127_609 ();
 FILLCELL_X32 FILLER_127_641 ();
 FILLCELL_X32 FILLER_127_673 ();
 FILLCELL_X32 FILLER_127_705 ();
 FILLCELL_X32 FILLER_127_737 ();
 FILLCELL_X32 FILLER_127_769 ();
 FILLCELL_X32 FILLER_127_801 ();
 FILLCELL_X32 FILLER_127_833 ();
 FILLCELL_X32 FILLER_127_865 ();
 FILLCELL_X32 FILLER_127_897 ();
 FILLCELL_X32 FILLER_127_929 ();
 FILLCELL_X32 FILLER_127_961 ();
 FILLCELL_X16 FILLER_127_993 ();
 FILLCELL_X8 FILLER_127_1009 ();
 FILLCELL_X4 FILLER_127_1017 ();
 FILLCELL_X2 FILLER_127_1021 ();
 FILLCELL_X1 FILLER_127_1023 ();
 FILLCELL_X32 FILLER_128_1 ();
 FILLCELL_X32 FILLER_128_33 ();
 FILLCELL_X32 FILLER_128_65 ();
 FILLCELL_X32 FILLER_128_97 ();
 FILLCELL_X32 FILLER_128_129 ();
 FILLCELL_X32 FILLER_128_161 ();
 FILLCELL_X32 FILLER_128_193 ();
 FILLCELL_X32 FILLER_128_225 ();
 FILLCELL_X32 FILLER_128_257 ();
 FILLCELL_X32 FILLER_128_289 ();
 FILLCELL_X32 FILLER_128_321 ();
 FILLCELL_X32 FILLER_128_353 ();
 FILLCELL_X32 FILLER_128_385 ();
 FILLCELL_X32 FILLER_128_417 ();
 FILLCELL_X32 FILLER_128_449 ();
 FILLCELL_X32 FILLER_128_481 ();
 FILLCELL_X32 FILLER_128_513 ();
 FILLCELL_X32 FILLER_128_545 ();
 FILLCELL_X32 FILLER_128_577 ();
 FILLCELL_X16 FILLER_128_609 ();
 FILLCELL_X4 FILLER_128_625 ();
 FILLCELL_X2 FILLER_128_629 ();
 FILLCELL_X32 FILLER_128_632 ();
 FILLCELL_X32 FILLER_128_664 ();
 FILLCELL_X32 FILLER_128_696 ();
 FILLCELL_X32 FILLER_128_728 ();
 FILLCELL_X32 FILLER_128_760 ();
 FILLCELL_X32 FILLER_128_792 ();
 FILLCELL_X32 FILLER_128_824 ();
 FILLCELL_X32 FILLER_128_856 ();
 FILLCELL_X32 FILLER_128_888 ();
 FILLCELL_X32 FILLER_128_920 ();
 FILLCELL_X32 FILLER_128_952 ();
 FILLCELL_X32 FILLER_128_984 ();
 FILLCELL_X8 FILLER_128_1016 ();
 FILLCELL_X32 FILLER_129_1 ();
 FILLCELL_X32 FILLER_129_33 ();
 FILLCELL_X32 FILLER_129_65 ();
 FILLCELL_X32 FILLER_129_97 ();
 FILLCELL_X32 FILLER_129_129 ();
 FILLCELL_X32 FILLER_129_161 ();
 FILLCELL_X32 FILLER_129_193 ();
 FILLCELL_X32 FILLER_129_225 ();
 FILLCELL_X32 FILLER_129_257 ();
 FILLCELL_X32 FILLER_129_289 ();
 FILLCELL_X32 FILLER_129_321 ();
 FILLCELL_X32 FILLER_129_353 ();
 FILLCELL_X32 FILLER_129_385 ();
 FILLCELL_X32 FILLER_129_417 ();
 FILLCELL_X32 FILLER_129_449 ();
 FILLCELL_X32 FILLER_129_481 ();
 FILLCELL_X32 FILLER_129_513 ();
 FILLCELL_X32 FILLER_129_545 ();
 FILLCELL_X32 FILLER_129_577 ();
 FILLCELL_X32 FILLER_129_609 ();
 FILLCELL_X32 FILLER_129_641 ();
 FILLCELL_X32 FILLER_129_673 ();
 FILLCELL_X32 FILLER_129_705 ();
 FILLCELL_X32 FILLER_129_737 ();
 FILLCELL_X32 FILLER_129_769 ();
 FILLCELL_X32 FILLER_129_801 ();
 FILLCELL_X32 FILLER_129_833 ();
 FILLCELL_X32 FILLER_129_865 ();
 FILLCELL_X32 FILLER_129_897 ();
 FILLCELL_X32 FILLER_129_929 ();
 FILLCELL_X32 FILLER_129_961 ();
 FILLCELL_X16 FILLER_129_993 ();
 FILLCELL_X8 FILLER_129_1009 ();
 FILLCELL_X4 FILLER_129_1017 ();
 FILLCELL_X2 FILLER_129_1021 ();
 FILLCELL_X1 FILLER_129_1023 ();
 FILLCELL_X32 FILLER_130_1 ();
 FILLCELL_X32 FILLER_130_33 ();
 FILLCELL_X32 FILLER_130_65 ();
 FILLCELL_X32 FILLER_130_97 ();
 FILLCELL_X32 FILLER_130_129 ();
 FILLCELL_X32 FILLER_130_161 ();
 FILLCELL_X32 FILLER_130_193 ();
 FILLCELL_X32 FILLER_130_225 ();
 FILLCELL_X32 FILLER_130_257 ();
 FILLCELL_X32 FILLER_130_289 ();
 FILLCELL_X32 FILLER_130_321 ();
 FILLCELL_X32 FILLER_130_353 ();
 FILLCELL_X32 FILLER_130_385 ();
 FILLCELL_X32 FILLER_130_417 ();
 FILLCELL_X32 FILLER_130_449 ();
 FILLCELL_X32 FILLER_130_481 ();
 FILLCELL_X32 FILLER_130_513 ();
 FILLCELL_X32 FILLER_130_545 ();
 FILLCELL_X32 FILLER_130_577 ();
 FILLCELL_X16 FILLER_130_609 ();
 FILLCELL_X4 FILLER_130_625 ();
 FILLCELL_X2 FILLER_130_629 ();
 FILLCELL_X32 FILLER_130_632 ();
 FILLCELL_X32 FILLER_130_664 ();
 FILLCELL_X32 FILLER_130_696 ();
 FILLCELL_X32 FILLER_130_728 ();
 FILLCELL_X32 FILLER_130_760 ();
 FILLCELL_X32 FILLER_130_792 ();
 FILLCELL_X32 FILLER_130_824 ();
 FILLCELL_X32 FILLER_130_856 ();
 FILLCELL_X32 FILLER_130_888 ();
 FILLCELL_X32 FILLER_130_920 ();
 FILLCELL_X32 FILLER_130_952 ();
 FILLCELL_X32 FILLER_130_984 ();
 FILLCELL_X1 FILLER_130_1016 ();
 FILLCELL_X4 FILLER_130_1020 ();
 FILLCELL_X32 FILLER_131_1 ();
 FILLCELL_X32 FILLER_131_33 ();
 FILLCELL_X32 FILLER_131_65 ();
 FILLCELL_X32 FILLER_131_97 ();
 FILLCELL_X32 FILLER_131_129 ();
 FILLCELL_X32 FILLER_131_161 ();
 FILLCELL_X32 FILLER_131_193 ();
 FILLCELL_X32 FILLER_131_225 ();
 FILLCELL_X32 FILLER_131_257 ();
 FILLCELL_X32 FILLER_131_289 ();
 FILLCELL_X32 FILLER_131_321 ();
 FILLCELL_X32 FILLER_131_353 ();
 FILLCELL_X32 FILLER_131_385 ();
 FILLCELL_X32 FILLER_131_417 ();
 FILLCELL_X32 FILLER_131_449 ();
 FILLCELL_X32 FILLER_131_481 ();
 FILLCELL_X32 FILLER_131_513 ();
 FILLCELL_X32 FILLER_131_545 ();
 FILLCELL_X32 FILLER_131_577 ();
 FILLCELL_X32 FILLER_131_609 ();
 FILLCELL_X32 FILLER_131_641 ();
 FILLCELL_X32 FILLER_131_673 ();
 FILLCELL_X32 FILLER_131_705 ();
 FILLCELL_X32 FILLER_131_737 ();
 FILLCELL_X32 FILLER_131_769 ();
 FILLCELL_X32 FILLER_131_801 ();
 FILLCELL_X32 FILLER_131_833 ();
 FILLCELL_X32 FILLER_131_865 ();
 FILLCELL_X32 FILLER_131_897 ();
 FILLCELL_X32 FILLER_131_929 ();
 FILLCELL_X32 FILLER_131_961 ();
 FILLCELL_X16 FILLER_131_993 ();
 FILLCELL_X8 FILLER_131_1009 ();
 FILLCELL_X4 FILLER_131_1017 ();
 FILLCELL_X2 FILLER_131_1021 ();
 FILLCELL_X1 FILLER_131_1023 ();
 FILLCELL_X32 FILLER_132_1 ();
 FILLCELL_X32 FILLER_132_33 ();
 FILLCELL_X32 FILLER_132_65 ();
 FILLCELL_X32 FILLER_132_97 ();
 FILLCELL_X32 FILLER_132_129 ();
 FILLCELL_X32 FILLER_132_161 ();
 FILLCELL_X32 FILLER_132_193 ();
 FILLCELL_X32 FILLER_132_225 ();
 FILLCELL_X32 FILLER_132_257 ();
 FILLCELL_X32 FILLER_132_289 ();
 FILLCELL_X32 FILLER_132_321 ();
 FILLCELL_X32 FILLER_132_353 ();
 FILLCELL_X32 FILLER_132_385 ();
 FILLCELL_X32 FILLER_132_417 ();
 FILLCELL_X32 FILLER_132_449 ();
 FILLCELL_X32 FILLER_132_481 ();
 FILLCELL_X32 FILLER_132_513 ();
 FILLCELL_X32 FILLER_132_545 ();
 FILLCELL_X32 FILLER_132_577 ();
 FILLCELL_X16 FILLER_132_609 ();
 FILLCELL_X4 FILLER_132_625 ();
 FILLCELL_X2 FILLER_132_629 ();
 FILLCELL_X32 FILLER_132_632 ();
 FILLCELL_X32 FILLER_132_664 ();
 FILLCELL_X32 FILLER_132_696 ();
 FILLCELL_X32 FILLER_132_728 ();
 FILLCELL_X32 FILLER_132_760 ();
 FILLCELL_X32 FILLER_132_792 ();
 FILLCELL_X32 FILLER_132_824 ();
 FILLCELL_X32 FILLER_132_856 ();
 FILLCELL_X32 FILLER_132_888 ();
 FILLCELL_X32 FILLER_132_920 ();
 FILLCELL_X32 FILLER_132_952 ();
 FILLCELL_X32 FILLER_132_984 ();
 FILLCELL_X8 FILLER_132_1016 ();
 FILLCELL_X32 FILLER_133_1 ();
 FILLCELL_X32 FILLER_133_33 ();
 FILLCELL_X32 FILLER_133_65 ();
 FILLCELL_X32 FILLER_133_97 ();
 FILLCELL_X32 FILLER_133_129 ();
 FILLCELL_X32 FILLER_133_161 ();
 FILLCELL_X32 FILLER_133_193 ();
 FILLCELL_X32 FILLER_133_225 ();
 FILLCELL_X32 FILLER_133_257 ();
 FILLCELL_X32 FILLER_133_289 ();
 FILLCELL_X32 FILLER_133_321 ();
 FILLCELL_X32 FILLER_133_353 ();
 FILLCELL_X32 FILLER_133_385 ();
 FILLCELL_X32 FILLER_133_417 ();
 FILLCELL_X32 FILLER_133_449 ();
 FILLCELL_X32 FILLER_133_481 ();
 FILLCELL_X32 FILLER_133_513 ();
 FILLCELL_X32 FILLER_133_545 ();
 FILLCELL_X32 FILLER_133_577 ();
 FILLCELL_X32 FILLER_133_609 ();
 FILLCELL_X32 FILLER_133_641 ();
 FILLCELL_X32 FILLER_133_673 ();
 FILLCELL_X32 FILLER_133_705 ();
 FILLCELL_X32 FILLER_133_737 ();
 FILLCELL_X32 FILLER_133_769 ();
 FILLCELL_X32 FILLER_133_801 ();
 FILLCELL_X32 FILLER_133_833 ();
 FILLCELL_X32 FILLER_133_865 ();
 FILLCELL_X32 FILLER_133_897 ();
 FILLCELL_X32 FILLER_133_929 ();
 FILLCELL_X32 FILLER_133_961 ();
 FILLCELL_X16 FILLER_133_993 ();
 FILLCELL_X8 FILLER_133_1009 ();
 FILLCELL_X4 FILLER_133_1017 ();
 FILLCELL_X2 FILLER_133_1021 ();
 FILLCELL_X1 FILLER_133_1023 ();
 FILLCELL_X32 FILLER_134_1 ();
 FILLCELL_X32 FILLER_134_33 ();
 FILLCELL_X32 FILLER_134_65 ();
 FILLCELL_X32 FILLER_134_97 ();
 FILLCELL_X32 FILLER_134_129 ();
 FILLCELL_X32 FILLER_134_161 ();
 FILLCELL_X32 FILLER_134_193 ();
 FILLCELL_X32 FILLER_134_225 ();
 FILLCELL_X32 FILLER_134_257 ();
 FILLCELL_X32 FILLER_134_289 ();
 FILLCELL_X32 FILLER_134_321 ();
 FILLCELL_X32 FILLER_134_353 ();
 FILLCELL_X32 FILLER_134_385 ();
 FILLCELL_X32 FILLER_134_417 ();
 FILLCELL_X32 FILLER_134_449 ();
 FILLCELL_X32 FILLER_134_481 ();
 FILLCELL_X32 FILLER_134_513 ();
 FILLCELL_X32 FILLER_134_545 ();
 FILLCELL_X32 FILLER_134_577 ();
 FILLCELL_X16 FILLER_134_609 ();
 FILLCELL_X4 FILLER_134_625 ();
 FILLCELL_X2 FILLER_134_629 ();
 FILLCELL_X32 FILLER_134_632 ();
 FILLCELL_X32 FILLER_134_664 ();
 FILLCELL_X32 FILLER_134_696 ();
 FILLCELL_X32 FILLER_134_728 ();
 FILLCELL_X32 FILLER_134_760 ();
 FILLCELL_X32 FILLER_134_792 ();
 FILLCELL_X32 FILLER_134_824 ();
 FILLCELL_X32 FILLER_134_856 ();
 FILLCELL_X32 FILLER_134_888 ();
 FILLCELL_X32 FILLER_134_920 ();
 FILLCELL_X32 FILLER_134_952 ();
 FILLCELL_X32 FILLER_134_984 ();
 FILLCELL_X8 FILLER_134_1016 ();
 FILLCELL_X32 FILLER_135_1 ();
 FILLCELL_X32 FILLER_135_33 ();
 FILLCELL_X32 FILLER_135_65 ();
 FILLCELL_X32 FILLER_135_97 ();
 FILLCELL_X32 FILLER_135_129 ();
 FILLCELL_X32 FILLER_135_161 ();
 FILLCELL_X32 FILLER_135_193 ();
 FILLCELL_X32 FILLER_135_225 ();
 FILLCELL_X32 FILLER_135_257 ();
 FILLCELL_X32 FILLER_135_289 ();
 FILLCELL_X32 FILLER_135_321 ();
 FILLCELL_X32 FILLER_135_353 ();
 FILLCELL_X32 FILLER_135_385 ();
 FILLCELL_X32 FILLER_135_417 ();
 FILLCELL_X32 FILLER_135_449 ();
 FILLCELL_X32 FILLER_135_481 ();
 FILLCELL_X32 FILLER_135_513 ();
 FILLCELL_X32 FILLER_135_545 ();
 FILLCELL_X32 FILLER_135_577 ();
 FILLCELL_X32 FILLER_135_609 ();
 FILLCELL_X32 FILLER_135_641 ();
 FILLCELL_X32 FILLER_135_673 ();
 FILLCELL_X32 FILLER_135_705 ();
 FILLCELL_X32 FILLER_135_737 ();
 FILLCELL_X32 FILLER_135_769 ();
 FILLCELL_X32 FILLER_135_801 ();
 FILLCELL_X32 FILLER_135_833 ();
 FILLCELL_X32 FILLER_135_865 ();
 FILLCELL_X32 FILLER_135_897 ();
 FILLCELL_X32 FILLER_135_929 ();
 FILLCELL_X32 FILLER_135_961 ();
 FILLCELL_X16 FILLER_135_993 ();
 FILLCELL_X8 FILLER_135_1009 ();
 FILLCELL_X4 FILLER_135_1017 ();
 FILLCELL_X2 FILLER_135_1021 ();
 FILLCELL_X1 FILLER_135_1023 ();
 FILLCELL_X4 FILLER_136_1 ();
 FILLCELL_X32 FILLER_136_9 ();
 FILLCELL_X32 FILLER_136_41 ();
 FILLCELL_X32 FILLER_136_73 ();
 FILLCELL_X32 FILLER_136_105 ();
 FILLCELL_X32 FILLER_136_137 ();
 FILLCELL_X32 FILLER_136_169 ();
 FILLCELL_X32 FILLER_136_201 ();
 FILLCELL_X32 FILLER_136_233 ();
 FILLCELL_X32 FILLER_136_265 ();
 FILLCELL_X32 FILLER_136_297 ();
 FILLCELL_X32 FILLER_136_329 ();
 FILLCELL_X32 FILLER_136_361 ();
 FILLCELL_X32 FILLER_136_393 ();
 FILLCELL_X32 FILLER_136_425 ();
 FILLCELL_X32 FILLER_136_457 ();
 FILLCELL_X32 FILLER_136_489 ();
 FILLCELL_X32 FILLER_136_521 ();
 FILLCELL_X32 FILLER_136_553 ();
 FILLCELL_X32 FILLER_136_585 ();
 FILLCELL_X8 FILLER_136_617 ();
 FILLCELL_X4 FILLER_136_625 ();
 FILLCELL_X2 FILLER_136_629 ();
 FILLCELL_X32 FILLER_136_632 ();
 FILLCELL_X32 FILLER_136_664 ();
 FILLCELL_X32 FILLER_136_696 ();
 FILLCELL_X32 FILLER_136_728 ();
 FILLCELL_X32 FILLER_136_760 ();
 FILLCELL_X32 FILLER_136_792 ();
 FILLCELL_X32 FILLER_136_824 ();
 FILLCELL_X32 FILLER_136_856 ();
 FILLCELL_X32 FILLER_136_888 ();
 FILLCELL_X32 FILLER_136_920 ();
 FILLCELL_X32 FILLER_136_952 ();
 FILLCELL_X32 FILLER_136_984 ();
 FILLCELL_X8 FILLER_136_1016 ();
 FILLCELL_X8 FILLER_137_1 ();
 FILLCELL_X4 FILLER_137_9 ();
 FILLCELL_X2 FILLER_137_13 ();
 FILLCELL_X32 FILLER_137_19 ();
 FILLCELL_X32 FILLER_137_51 ();
 FILLCELL_X8 FILLER_137_83 ();
 FILLCELL_X4 FILLER_137_91 ();
 FILLCELL_X2 FILLER_137_95 ();
 FILLCELL_X32 FILLER_137_100 ();
 FILLCELL_X32 FILLER_137_132 ();
 FILLCELL_X8 FILLER_137_164 ();
 FILLCELL_X2 FILLER_137_172 ();
 FILLCELL_X32 FILLER_137_177 ();
 FILLCELL_X32 FILLER_137_209 ();
 FILLCELL_X8 FILLER_137_241 ();
 FILLCELL_X2 FILLER_137_249 ();
 FILLCELL_X32 FILLER_137_254 ();
 FILLCELL_X32 FILLER_137_286 ();
 FILLCELL_X8 FILLER_137_318 ();
 FILLCELL_X4 FILLER_137_326 ();
 FILLCELL_X2 FILLER_137_330 ();
 FILLCELL_X1 FILLER_137_332 ();
 FILLCELL_X32 FILLER_137_336 ();
 FILLCELL_X32 FILLER_137_368 ();
 FILLCELL_X8 FILLER_137_400 ();
 FILLCELL_X2 FILLER_137_408 ();
 FILLCELL_X32 FILLER_137_413 ();
 FILLCELL_X32 FILLER_137_445 ();
 FILLCELL_X8 FILLER_137_477 ();
 FILLCELL_X4 FILLER_137_485 ();
 FILLCELL_X2 FILLER_137_489 ();
 FILLCELL_X1 FILLER_137_491 ();
 FILLCELL_X32 FILLER_137_495 ();
 FILLCELL_X32 FILLER_137_527 ();
 FILLCELL_X8 FILLER_137_559 ();
 FILLCELL_X2 FILLER_137_567 ();
 FILLCELL_X32 FILLER_137_572 ();
 FILLCELL_X16 FILLER_137_604 ();
 FILLCELL_X8 FILLER_137_620 ();
 FILLCELL_X2 FILLER_137_628 ();
 FILLCELL_X1 FILLER_137_630 ();
 FILLCELL_X8 FILLER_137_632 ();
 FILLCELL_X4 FILLER_137_640 ();
 FILLCELL_X2 FILLER_137_644 ();
 FILLCELL_X32 FILLER_137_650 ();
 FILLCELL_X32 FILLER_137_682 ();
 FILLCELL_X8 FILLER_137_714 ();
 FILLCELL_X4 FILLER_137_722 ();
 FILLCELL_X2 FILLER_137_726 ();
 FILLCELL_X32 FILLER_137_731 ();
 FILLCELL_X32 FILLER_137_763 ();
 FILLCELL_X8 FILLER_137_795 ();
 FILLCELL_X2 FILLER_137_803 ();
 FILLCELL_X32 FILLER_137_809 ();
 FILLCELL_X32 FILLER_137_841 ();
 FILLCELL_X8 FILLER_137_873 ();
 FILLCELL_X4 FILLER_137_881 ();
 FILLCELL_X2 FILLER_137_885 ();
 FILLCELL_X32 FILLER_137_890 ();
 FILLCELL_X32 FILLER_137_922 ();
 FILLCELL_X8 FILLER_137_954 ();
 FILLCELL_X2 FILLER_137_962 ();
 FILLCELL_X32 FILLER_137_967 ();
 FILLCELL_X16 FILLER_137_999 ();
 FILLCELL_X2 FILLER_137_1015 ();
 FILLCELL_X4 FILLER_137_1020 ();
 assign init_done = curr_state[1];
 assign valid_out = valid_reg_out;
endmodule
