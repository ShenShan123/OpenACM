VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO SRAM_6T_CORE_64x32_MC_TB 
   CLASS BLOCK ;
   SIZE 211.78 BY 229.68 ;
   SYMMETRY X Y R90 ;
   PIN wd_in[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  26.03 0.0 26.18 0.15 ;
      END
   END wd_in[0]
   PIN wd_in[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  31.76 0.0 31.91 0.15 ;
      END
   END wd_in[1]
   PIN wd_in[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  37.48 0.0 37.63 0.15 ;
      END
   END wd_in[2]
   PIN wd_in[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  43.19 0.0 43.34 0.15 ;
      END
   END wd_in[3]
   PIN wd_in[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  48.91 0.0 49.06 0.15 ;
      END
   END wd_in[4]
   PIN wd_in[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  54.64 0.0 54.79 0.15 ;
      END
   END wd_in[5]
   PIN wd_in[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  60.36 0.0 60.51 0.15 ;
      END
   END wd_in[6]
   PIN wd_in[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  66.08 0.0 66.23 0.15 ;
      END
   END wd_in[7]
   PIN wd_in[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  71.8 0.0 71.95 0.15 ;
      END
   END wd_in[8]
   PIN wd_in[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  77.51 0.0 77.66 0.15 ;
      END
   END wd_in[9]
   PIN wd_in[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  83.23 0.0 83.38 0.15 ;
      END
   END wd_in[10]
   PIN wd_in[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  88.95 0.0 89.1 0.15 ;
      END
   END wd_in[11]
   PIN wd_in[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  94.67 0.0 94.82 0.15 ;
      END
   END wd_in[12]
   PIN wd_in[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  100.4 0.0 100.55 0.15 ;
      END
   END wd_in[13]
   PIN wd_in[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  106.12 0.0 106.27 0.15 ;
      END
   END wd_in[14]
   PIN wd_in[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  111.84 0.0 111.99 0.15 ;
      END
   END wd_in[15]
   PIN wd_in[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  117.56 0.0 117.71 0.15 ;
      END
   END wd_in[16]
   PIN wd_in[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  123.28 0.0 123.43 0.15 ;
      END
   END wd_in[17]
   PIN wd_in[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  129.0 0.0 129.15 0.15 ;
      END
   END wd_in[18]
   PIN wd_in[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  134.72 0.0 134.87 0.15 ;
      END
   END wd_in[19]
   PIN wd_in[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  140.44 0.0 140.59 0.15 ;
      END
   END wd_in[20]
   PIN wd_in[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  146.15 0.0 146.3 0.15 ;
      END
   END wd_in[21]
   PIN wd_in[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  151.87 0.0 152.02 0.15 ;
      END
   END wd_in[22]
   PIN wd_in[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  157.59 0.0 157.74 0.15 ;
      END
   END wd_in[23]
   PIN wd_in[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  163.32 0.0 163.47 0.15 ;
      END
   END wd_in[24]
   PIN wd_in[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  169.03 0.0 169.18 0.15 ;
      END
   END wd_in[25]
   PIN wd_in[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  174.76 0.0 174.91 0.15 ;
      END
   END wd_in[26]
   PIN wd_in[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  180.47 0.0 180.62 0.15 ;
      END
   END wd_in[27]
   PIN wd_in[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  186.2 0.0 186.35 0.15 ;
      END
   END wd_in[28]
   PIN wd_in[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  191.91 0.0 192.06 0.15 ;
      END
   END wd_in[29]
   PIN wd_in[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  197.64 0.0 197.79 0.15 ;
      END
   END wd_in[30]
   PIN wd_in[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  203.35 0.0 203.5 0.15 ;
      END
   END wd_in[31]
   PIN addr_in[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 94.57 0.15 94.72 ;
      END
   END addr_in[0]
   PIN addr_in[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 100.03 0.15 100.18 ;
      END
   END addr_in[1]
   PIN addr_in[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 104.45 0.15 104.6 ;
      END
   END addr_in[2]
   PIN addr_in[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 109.91 0.15 110.06 ;
      END
   END addr_in[3]
   PIN addr_in[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 114.33 0.15 114.48 ;
      END
   END addr_in[4]
   PIN addr_in[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 119.79 0.15 119.94 ;
      END
   END addr_in[5]
   PIN ce_in
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 5.52 0.15 5.67 ;
      END
   END ce_in
   PIN we_in
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 10.98 0.15 11.13 ;
      END
   END we_in
   PIN clk
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  12.61 0.0 12.76 0.15 ;
      END
   END clk
   PIN rd_out[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  36.2 0.0 36.35 0.15 ;
      END
   END rd_out[0]
   PIN rd_out[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  37.79 0.0 37.94 0.15 ;
      END
   END rd_out[1]
   PIN rd_out[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  39.14 0.0 39.29 0.15 ;
      END
   END rd_out[2]
   PIN rd_out[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  40.55 0.0 40.7 0.15 ;
      END
   END rd_out[3]
   PIN rd_out[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  41.92 0.0 42.07 0.15 ;
      END
   END rd_out[4]
   PIN rd_out[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  43.5 0.0 43.65 0.15 ;
      END
   END rd_out[5]
   PIN rd_out[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  44.78 0.0 44.93 0.15 ;
      END
   END rd_out[6]
   PIN rd_out[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  46.19 0.0 46.34 0.15 ;
      END
   END rd_out[7]
   PIN rd_out[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  47.6 0.0 47.75 0.15 ;
      END
   END rd_out[8]
   PIN rd_out[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  49.22 0.0 49.37 0.15 ;
      END
   END rd_out[9]
   PIN rd_out[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  50.42 0.0 50.57 0.15 ;
      END
   END rd_out[10]
   PIN rd_out[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  51.83 0.0 51.98 0.15 ;
      END
   END rd_out[11]
   PIN rd_out[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  53.25 0.0 53.4 0.15 ;
      END
   END rd_out[12]
   PIN rd_out[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  54.32 0.0 54.47 0.15 ;
      END
   END rd_out[13]
   PIN rd_out[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  56.06 0.0 56.21 0.15 ;
      END
   END rd_out[14]
   PIN rd_out[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  57.47 0.0 57.62 0.15 ;
      END
   END rd_out[15]
   PIN rd_out[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  58.88 0.0 59.03 0.15 ;
      END
   END rd_out[16]
   PIN rd_out[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  60.02 0.0 60.17 0.15 ;
      END
   END rd_out[17]
   PIN rd_out[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  61.7 0.0 61.85 0.15 ;
      END
   END rd_out[18]
   PIN rd_out[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  63.11 0.0 63.26 0.15 ;
      END
   END rd_out[19]
   PIN rd_out[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  64.52 0.0 64.67 0.15 ;
      END
   END rd_out[20]
   PIN rd_out[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  65.66 0.0 65.81 0.15 ;
      END
   END rd_out[21]
   PIN rd_out[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  67.34 0.0 67.49 0.15 ;
      END
   END rd_out[22]
   PIN rd_out[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  68.75 0.0 68.9 0.15 ;
      END
   END rd_out[23]
   PIN rd_out[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  70.16 0.0 70.31 0.15 ;
      END
   END rd_out[24]
   PIN rd_out[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  71.48 0.0 71.63 0.15 ;
      END
   END rd_out[25]
   PIN rd_out[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  72.98 0.0 73.13 0.15 ;
      END
   END rd_out[26]
   PIN rd_out[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  74.39 0.0 74.54 0.15 ;
      END
   END rd_out[27]
   PIN rd_out[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  75.8 0.0 75.95 0.15 ;
      END
   END rd_out[28]
   PIN rd_out[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  77.19 0.0 77.34 0.15 ;
      END
   END rd_out[29]
   PIN rd_out[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  78.62 0.0 78.77 0.15 ;
      END
   END rd_out[30]
   PIN rd_out[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  80.03 0.0 80.18 0.15 ;
      END
   END rd_out[31]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  0.0 0.0 0.73 229.68 ;
         LAYER metal3 ;
         RECT  0.0 0.0 211.78 0.73 ;
         LAYER metal3 ;
         RECT  0.0 228.95 211.78 229.68 ;
         LAYER metal4 ;
         RECT  211.05 0.0 211.78 229.68 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  209.59 1.46 210.32 228.22 ;
         LAYER metal3 ;
         RECT  1.46 227.49 210.32 228.22 ;
         LAYER metal4 ;
         RECT  1.46 1.46 2.19 228.22 ;
         LAYER metal3 ;
         RECT  1.46 1.46 210.32 2.19 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 211.64 229.54 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 211.64 229.54 ;
   LAYER  metal3 ;
      RECT  0.29 94.43 211.64 94.86 ;
      RECT  0.14 94.86 0.29 99.89 ;
      RECT  0.14 100.32 0.29 104.31 ;
      RECT  0.14 104.74 0.29 109.77 ;
      RECT  0.14 110.2 0.29 114.19 ;
      RECT  0.14 114.62 0.29 119.65 ;
      RECT  0.14 5.81 0.29 10.84 ;
      RECT  0.14 11.27 0.29 94.43 ;
      RECT  0.14 0.87 0.29 5.38 ;
      RECT  0.14 120.08 0.29 228.81 ;
      RECT  0.29 94.86 1.32 227.35 ;
      RECT  0.29 227.35 1.32 228.36 ;
      RECT  0.29 228.36 1.32 228.81 ;
      RECT  1.32 94.86 210.46 227.35 ;
      RECT  1.32 228.36 210.46 228.81 ;
      RECT  210.46 94.86 211.64 227.35 ;
      RECT  210.46 227.35 211.64 228.36 ;
      RECT  210.46 228.36 211.64 228.81 ;
      RECT  0.29 0.87 1.32 1.32 ;
      RECT  0.29 1.32 1.32 2.33 ;
      RECT  0.29 2.33 1.32 94.43 ;
      RECT  1.32 0.87 210.46 1.32 ;
      RECT  1.32 2.33 210.46 94.43 ;
      RECT  210.46 0.87 211.64 1.32 ;
      RECT  210.46 1.32 211.64 2.33 ;
      RECT  210.46 2.33 211.64 94.43 ;
   LAYER  metal4 ;
      RECT  25.75 0.43 26.46 229.54 ;
      RECT  26.46 0.14 31.48 0.43 ;
      RECT  83.66 0.14 88.67 0.43 ;
      RECT  89.38 0.14 94.39 0.43 ;
      RECT  95.1 0.14 100.12 0.43 ;
      RECT  100.83 0.14 105.84 0.43 ;
      RECT  106.55 0.14 111.56 0.43 ;
      RECT  112.27 0.14 117.28 0.43 ;
      RECT  117.99 0.14 123.0 0.43 ;
      RECT  123.71 0.14 128.72 0.43 ;
      RECT  129.43 0.14 134.44 0.43 ;
      RECT  135.15 0.14 140.16 0.43 ;
      RECT  140.87 0.14 145.87 0.43 ;
      RECT  146.58 0.14 151.59 0.43 ;
      RECT  152.3 0.14 157.31 0.43 ;
      RECT  158.02 0.14 163.04 0.43 ;
      RECT  163.75 0.14 168.75 0.43 ;
      RECT  169.46 0.14 174.48 0.43 ;
      RECT  175.19 0.14 180.19 0.43 ;
      RECT  180.9 0.14 185.92 0.43 ;
      RECT  186.63 0.14 191.63 0.43 ;
      RECT  192.34 0.14 197.36 0.43 ;
      RECT  198.07 0.14 203.07 0.43 ;
      RECT  13.04 0.14 25.75 0.43 ;
      RECT  32.19 0.14 35.92 0.43 ;
      RECT  36.63 0.14 37.2 0.43 ;
      RECT  38.22 0.14 38.86 0.43 ;
      RECT  39.57 0.14 40.27 0.43 ;
      RECT  40.98 0.14 41.64 0.43 ;
      RECT  42.35 0.14 42.91 0.43 ;
      RECT  43.93 0.14 44.5 0.43 ;
      RECT  45.21 0.14 45.91 0.43 ;
      RECT  46.62 0.14 47.32 0.43 ;
      RECT  48.03 0.14 48.63 0.43 ;
      RECT  49.65 0.14 50.14 0.43 ;
      RECT  50.85 0.14 51.55 0.43 ;
      RECT  52.26 0.14 52.97 0.43 ;
      RECT  53.68 0.14 54.04 0.43 ;
      RECT  55.07 0.14 55.78 0.43 ;
      RECT  56.49 0.14 57.19 0.43 ;
      RECT  57.9 0.14 58.6 0.43 ;
      RECT  59.31 0.14 59.74 0.43 ;
      RECT  60.79 0.14 61.42 0.43 ;
      RECT  62.13 0.14 62.83 0.43 ;
      RECT  63.54 0.14 64.24 0.43 ;
      RECT  64.95 0.14 65.38 0.43 ;
      RECT  66.51 0.14 67.06 0.43 ;
      RECT  67.77 0.14 68.47 0.43 ;
      RECT  69.18 0.14 69.88 0.43 ;
      RECT  70.59 0.14 71.2 0.43 ;
      RECT  72.23 0.14 72.7 0.43 ;
      RECT  73.41 0.14 74.11 0.43 ;
      RECT  74.82 0.14 75.52 0.43 ;
      RECT  76.23 0.14 76.91 0.43 ;
      RECT  77.94 0.14 78.34 0.43 ;
      RECT  79.05 0.14 79.75 0.43 ;
      RECT  80.46 0.14 82.95 0.43 ;
      RECT  1.01 0.14 12.33 0.43 ;
      RECT  203.78 0.14 210.77 0.43 ;
      RECT  26.46 0.43 209.31 1.18 ;
      RECT  26.46 1.18 209.31 228.5 ;
      RECT  26.46 228.5 209.31 229.54 ;
      RECT  209.31 0.43 210.6 1.18 ;
      RECT  209.31 228.5 210.6 229.54 ;
      RECT  210.6 0.43 210.77 1.18 ;
      RECT  210.6 1.18 210.77 228.5 ;
      RECT  210.6 228.5 210.77 229.54 ;
      RECT  1.01 0.43 1.18 1.18 ;
      RECT  1.01 1.18 1.18 228.5 ;
      RECT  1.01 228.5 1.18 229.54 ;
      RECT  1.18 0.43 2.47 1.18 ;
      RECT  1.18 228.5 2.47 229.54 ;
      RECT  2.47 0.43 25.75 1.18 ;
      RECT  2.47 1.18 25.75 228.5 ;
      RECT  2.47 228.5 25.75 229.54 ;
   END
END    SRAM_6T_CORE_64x32_MC_TB 
END    LIBRARY
