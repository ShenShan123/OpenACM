module sram_multiplier_system (clk,
    init_done,
    init_enable,
    pe_ce,
    rst_n,
    valid_out,
    data_in,
    data_out);
 input clk;
 output init_done;
 input init_enable;
 input pe_ce;
 input rst_n;
 output valid_out;
 input [31:0] data_in;
 output [63:0] data_out;

 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net161;
 wire net163;
 wire u_multiplier_pp1_0 ;
 wire u_multiplier_pp1_62 ;
 wire net132;
 wire u_multiplier_pp2_0 ;
 wire u_multiplier_pp2_62 ;
 wire net140;
 wire u_multiplier_pp3_0 ;
 wire u_multiplier_pp3_62 ;
 wire net147;
 wire u_multiplier_Final_add_Cout ;
 wire u_multiplier_Final_add_c1 ;
 wire u_multiplier_Final_add_cla1_c1 ;
 wire u_multiplier_Final_add_cla1_cla1_c1 ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_c1 ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__25_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__26_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__27_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__28_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__29_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__30_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__31_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__32_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__33_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__34_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__35_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__36_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__37_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__38_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__39_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__25_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__26_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__27_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__28_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__29_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__30_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__31_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__32_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__33_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__34_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__35_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__36_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__37_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__38_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__39_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_c1 ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__25_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__26_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__27_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__28_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__29_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__30_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__31_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__32_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__33_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__34_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__35_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__36_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__37_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__38_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__39_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__25_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__26_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__27_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__28_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__29_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__30_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__31_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__32_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__33_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__34_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__35_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__36_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__37_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__38_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__39_ ;
 wire u_multiplier_Final_add_cla1_cla2_c1 ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_c1 ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__25_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__26_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__27_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__28_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__29_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__30_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__31_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__32_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__33_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__34_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__35_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__36_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__37_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__38_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__39_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__25_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__26_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__27_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__28_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__29_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__30_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__31_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__32_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__33_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__34_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__35_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__36_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__37_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__38_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__39_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_c1 ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__25_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__26_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__27_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__28_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__29_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__30_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__31_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__32_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__33_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__34_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__35_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__36_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__37_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__38_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__39_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__25_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__26_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__27_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__28_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__29_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__30_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__31_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__32_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__33_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__34_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__35_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__36_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__37_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__38_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__39_ ;
 wire u_multiplier_Final_add_cla2_c1 ;
 wire u_multiplier_Final_add_cla2_cla1_c1 ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_c1 ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__25_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__26_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__27_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__28_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__29_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__30_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__31_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__32_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__33_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__34_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__35_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__36_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__37_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__38_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__39_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__25_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__26_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__27_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__28_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__29_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__30_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__31_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__32_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__33_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__34_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__35_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__36_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__37_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__38_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__39_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_c1 ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__25_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__26_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__27_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__28_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__29_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__30_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__31_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__32_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__33_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__34_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__35_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__36_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__37_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__38_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__39_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__25_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__26_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__27_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__28_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__29_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__30_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__31_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__32_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__33_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__34_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__35_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__36_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__37_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__38_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__39_ ;
 wire u_multiplier_Final_add_cla2_cla2_c1 ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_c1 ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__25_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__26_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__27_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__28_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__29_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__30_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__31_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__32_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__33_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__34_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__35_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__36_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__37_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__38_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__39_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__25_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__26_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__27_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__28_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__29_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__30_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__31_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__32_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__33_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__34_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__35_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__36_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__37_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__38_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__39_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_c1 ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__25_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__26_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__27_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__28_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__29_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__30_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__31_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__32_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__33_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__34_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__35_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__36_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__37_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__38_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__39_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__25_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__26_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__27_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__28_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__29_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__30_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__31_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__32_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__33_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__34_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__35_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__36_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__37_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__38_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__39_ ;
 wire u_multiplier_STAGE1__0607_ ;
 wire u_multiplier_STAGE1__0608_ ;
 wire u_multiplier_STAGE1__0609_ ;
 wire u_multiplier_STAGE1__0610_ ;
 wire u_multiplier_STAGE1__0611_ ;
 wire u_multiplier_STAGE1__0612_ ;
 wire u_multiplier_STAGE1__0613_ ;
 wire u_multiplier_STAGE1__0614_ ;
 wire u_multiplier_STAGE1__0615_ ;
 wire u_multiplier_STAGE1__0616_ ;
 wire u_multiplier_STAGE1__0617_ ;
 wire u_multiplier_STAGE1__0618_ ;
 wire u_multiplier_STAGE1__0619_ ;
 wire u_multiplier_STAGE1__0620_ ;
 wire u_multiplier_STAGE1__0621_ ;
 wire u_multiplier_STAGE1__0622_ ;
 wire u_multiplier_STAGE1__0623_ ;
 wire u_multiplier_STAGE1__0624_ ;
 wire u_multiplier_STAGE1__0625_ ;
 wire u_multiplier_STAGE1__0626_ ;
 wire u_multiplier_STAGE1__0627_ ;
 wire u_multiplier_STAGE1__0628_ ;
 wire u_multiplier_STAGE1__0629_ ;
 wire u_multiplier_STAGE1__0630_ ;
 wire u_multiplier_STAGE1__0631_ ;
 wire u_multiplier_STAGE1__0632_ ;
 wire u_multiplier_STAGE1__0633_ ;
 wire u_multiplier_STAGE1__0634_ ;
 wire u_multiplier_STAGE1__0635_ ;
 wire u_multiplier_STAGE1__0636_ ;
 wire u_multiplier_STAGE1__0637_ ;
 wire u_multiplier_STAGE1__0638_ ;
 wire u_multiplier_STAGE1__0639_ ;
 wire u_multiplier_STAGE1__0640_ ;
 wire u_multiplier_STAGE1__0641_ ;
 wire u_multiplier_STAGE1__0642_ ;
 wire u_multiplier_STAGE1__0643_ ;
 wire u_multiplier_STAGE1__0644_ ;
 wire u_multiplier_STAGE1__0645_ ;
 wire u_multiplier_STAGE1__0646_ ;
 wire u_multiplier_STAGE1__0647_ ;
 wire u_multiplier_STAGE1__0648_ ;
 wire u_multiplier_STAGE1__0649_ ;
 wire u_multiplier_STAGE1__0650_ ;
 wire u_multiplier_STAGE1__0651_ ;
 wire u_multiplier_STAGE1__0652_ ;
 wire u_multiplier_STAGE1__0653_ ;
 wire u_multiplier_STAGE1__0654_ ;
 wire u_multiplier_STAGE1__0655_ ;
 wire u_multiplier_STAGE1__0656_ ;
 wire u_multiplier_STAGE1__0657_ ;
 wire u_multiplier_STAGE1__0658_ ;
 wire u_multiplier_STAGE1__0659_ ;
 wire u_multiplier_STAGE1__0660_ ;
 wire u_multiplier_STAGE1__0661_ ;
 wire u_multiplier_STAGE1__0662_ ;
 wire u_multiplier_STAGE1__0663_ ;
 wire u_multiplier_STAGE1__0664_ ;
 wire u_multiplier_STAGE1__0665_ ;
 wire u_multiplier_STAGE1__0666_ ;
 wire u_multiplier_STAGE1__0667_ ;
 wire u_multiplier_STAGE1__0668_ ;
 wire u_multiplier_STAGE1__0669_ ;
 wire u_multiplier_STAGE1__0670_ ;
 wire u_multiplier_STAGE1__0671_ ;
 wire u_multiplier_STAGE1__0672_ ;
 wire u_multiplier_STAGE1__0673_ ;
 wire u_multiplier_STAGE1__0674_ ;
 wire u_multiplier_STAGE1__0675_ ;
 wire u_multiplier_STAGE1__0676_ ;
 wire u_multiplier_STAGE1__0677_ ;
 wire u_multiplier_STAGE1__0678_ ;
 wire u_multiplier_STAGE1__0679_ ;
 wire u_multiplier_STAGE1__0680_ ;
 wire u_multiplier_STAGE1__0681_ ;
 wire u_multiplier_STAGE1__0682_ ;
 wire u_multiplier_STAGE1__0683_ ;
 wire u_multiplier_STAGE1__0684_ ;
 wire u_multiplier_STAGE1__0685_ ;
 wire u_multiplier_STAGE1__0686_ ;
 wire u_multiplier_STAGE1__0687_ ;
 wire u_multiplier_STAGE1__0688_ ;
 wire u_multiplier_STAGE1__0689_ ;
 wire u_multiplier_STAGE1__0690_ ;
 wire u_multiplier_STAGE1__0691_ ;
 wire u_multiplier_STAGE1__0692_ ;
 wire u_multiplier_STAGE1__0693_ ;
 wire u_multiplier_STAGE1__0694_ ;
 wire u_multiplier_STAGE1__0695_ ;
 wire u_multiplier_STAGE1__0696_ ;
 wire u_multiplier_STAGE1__0697_ ;
 wire u_multiplier_STAGE1__0698_ ;
 wire u_multiplier_STAGE1__0699_ ;
 wire u_multiplier_STAGE1__0700_ ;
 wire u_multiplier_STAGE1__0701_ ;
 wire u_multiplier_STAGE1__0702_ ;
 wire u_multiplier_STAGE1__0703_ ;
 wire u_multiplier_STAGE1__0704_ ;
 wire u_multiplier_STAGE1__0705_ ;
 wire u_multiplier_STAGE1__0706_ ;
 wire u_multiplier_STAGE1__0707_ ;
 wire u_multiplier_STAGE1__0708_ ;
 wire u_multiplier_STAGE1__0709_ ;
 wire u_multiplier_STAGE1__0710_ ;
 wire u_multiplier_STAGE1__0711_ ;
 wire u_multiplier_STAGE1__0712_ ;
 wire u_multiplier_STAGE1__0713_ ;
 wire u_multiplier_STAGE1__0714_ ;
 wire u_multiplier_STAGE1__0715_ ;
 wire u_multiplier_STAGE1__0716_ ;
 wire u_multiplier_STAGE1__0717_ ;
 wire u_multiplier_STAGE1__0718_ ;
 wire u_multiplier_STAGE1__0719_ ;
 wire u_multiplier_STAGE1__0720_ ;
 wire u_multiplier_STAGE1__0721_ ;
 wire u_multiplier_STAGE1__0722_ ;
 wire u_multiplier_STAGE1__0723_ ;
 wire u_multiplier_STAGE1__0724_ ;
 wire u_multiplier_STAGE1__0725_ ;
 wire u_multiplier_STAGE1__0726_ ;
 wire u_multiplier_STAGE1__0727_ ;
 wire u_multiplier_STAGE1__0728_ ;
 wire u_multiplier_STAGE1__0729_ ;
 wire u_multiplier_STAGE1__0730_ ;
 wire u_multiplier_STAGE1__0731_ ;
 wire u_multiplier_STAGE1__0732_ ;
 wire u_multiplier_STAGE1__0733_ ;
 wire u_multiplier_STAGE1__0734_ ;
 wire u_multiplier_STAGE1__0735_ ;
 wire u_multiplier_STAGE1__0736_ ;
 wire u_multiplier_STAGE1__0737_ ;
 wire u_multiplier_STAGE1__0738_ ;
 wire u_multiplier_STAGE1__0739_ ;
 wire u_multiplier_STAGE1__0740_ ;
 wire u_multiplier_STAGE1__0741_ ;
 wire u_multiplier_STAGE1__0742_ ;
 wire u_multiplier_STAGE1__0743_ ;
 wire u_multiplier_STAGE1__0744_ ;
 wire u_multiplier_STAGE1__0745_ ;
 wire u_multiplier_STAGE1__0746_ ;
 wire u_multiplier_STAGE1__0747_ ;
 wire u_multiplier_STAGE1__0748_ ;
 wire u_multiplier_STAGE1__0749_ ;
 wire u_multiplier_STAGE1__0750_ ;
 wire u_multiplier_STAGE1__0751_ ;
 wire u_multiplier_STAGE1__0752_ ;
 wire u_multiplier_STAGE1__0753_ ;
 wire u_multiplier_STAGE1__0754_ ;
 wire u_multiplier_STAGE1__0755_ ;
 wire u_multiplier_STAGE1__0756_ ;
 wire u_multiplier_STAGE1__0757_ ;
 wire u_multiplier_STAGE1__0758_ ;
 wire u_multiplier_STAGE1__0759_ ;
 wire u_multiplier_STAGE1__0760_ ;
 wire u_multiplier_STAGE1__0761_ ;
 wire u_multiplier_STAGE1__0762_ ;
 wire u_multiplier_STAGE1__0763_ ;
 wire u_multiplier_STAGE1__0764_ ;
 wire u_multiplier_STAGE1__0765_ ;
 wire u_multiplier_STAGE1__0766_ ;
 wire u_multiplier_STAGE1__0767_ ;
 wire u_multiplier_STAGE1__0768_ ;
 wire u_multiplier_STAGE1__0769_ ;
 wire u_multiplier_STAGE1__0770_ ;
 wire u_multiplier_STAGE1__0771_ ;
 wire u_multiplier_STAGE1__0772_ ;
 wire u_multiplier_STAGE1__0773_ ;
 wire u_multiplier_STAGE1__0774_ ;
 wire u_multiplier_STAGE1__0775_ ;
 wire u_multiplier_STAGE1__0776_ ;
 wire u_multiplier_STAGE1__0777_ ;
 wire u_multiplier_STAGE1__0778_ ;
 wire u_multiplier_STAGE1__0779_ ;
 wire u_multiplier_STAGE1__0780_ ;
 wire u_multiplier_STAGE1__0781_ ;
 wire u_multiplier_STAGE1__0782_ ;
 wire u_multiplier_STAGE1__0783_ ;
 wire u_multiplier_STAGE1__0784_ ;
 wire u_multiplier_STAGE1__0785_ ;
 wire u_multiplier_STAGE1__0786_ ;
 wire u_multiplier_STAGE1__0787_ ;
 wire u_multiplier_STAGE1__0788_ ;
 wire u_multiplier_STAGE1__0789_ ;
 wire u_multiplier_STAGE1__0790_ ;
 wire u_multiplier_STAGE1__0791_ ;
 wire u_multiplier_STAGE1__0792_ ;
 wire u_multiplier_STAGE1__0793_ ;
 wire u_multiplier_STAGE1__0794_ ;
 wire u_multiplier_STAGE1__0795_ ;
 wire u_multiplier_STAGE1__0796_ ;
 wire u_multiplier_STAGE1__0797_ ;
 wire u_multiplier_STAGE1__0798_ ;
 wire u_multiplier_STAGE1__0799_ ;
 wire u_multiplier_STAGE1__0800_ ;
 wire u_multiplier_STAGE1__0801_ ;
 wire u_multiplier_STAGE1__0802_ ;
 wire u_multiplier_STAGE1__0803_ ;
 wire u_multiplier_STAGE1__0804_ ;
 wire u_multiplier_STAGE1__0805_ ;
 wire u_multiplier_STAGE1__0806_ ;
 wire u_multiplier_STAGE1__0807_ ;
 wire u_multiplier_STAGE1__0808_ ;
 wire u_multiplier_STAGE1__0809_ ;
 wire u_multiplier_STAGE1__0810_ ;
 wire u_multiplier_STAGE1__0811_ ;
 wire u_multiplier_STAGE1__0812_ ;
 wire u_multiplier_STAGE1__0813_ ;
 wire u_multiplier_STAGE1__0814_ ;
 wire u_multiplier_STAGE1__0815_ ;
 wire u_multiplier_STAGE1__0816_ ;
 wire u_multiplier_STAGE1__0817_ ;
 wire u_multiplier_STAGE1__0818_ ;
 wire u_multiplier_STAGE1__0819_ ;
 wire u_multiplier_STAGE1__0820_ ;
 wire u_multiplier_STAGE1__0821_ ;
 wire u_multiplier_STAGE1__0822_ ;
 wire u_multiplier_STAGE1__0823_ ;
 wire u_multiplier_STAGE1__0824_ ;
 wire u_multiplier_STAGE1__0825_ ;
 wire u_multiplier_STAGE1__0826_ ;
 wire u_multiplier_STAGE1__0827_ ;
 wire u_multiplier_STAGE1__0828_ ;
 wire u_multiplier_STAGE1__0829_ ;
 wire u_multiplier_STAGE1__0830_ ;
 wire u_multiplier_STAGE1__0831_ ;
 wire u_multiplier_STAGE1__0832_ ;
 wire u_multiplier_STAGE1__0833_ ;
 wire u_multiplier_STAGE1__0834_ ;
 wire u_multiplier_STAGE1__0835_ ;
 wire u_multiplier_STAGE1__0836_ ;
 wire u_multiplier_STAGE1__0837_ ;
 wire u_multiplier_STAGE1__0838_ ;
 wire u_multiplier_STAGE1__0839_ ;
 wire u_multiplier_STAGE1__0840_ ;
 wire u_multiplier_STAGE1__0841_ ;
 wire u_multiplier_STAGE1__0842_ ;
 wire u_multiplier_STAGE1__0843_ ;
 wire u_multiplier_STAGE1__0844_ ;
 wire u_multiplier_STAGE1__0845_ ;
 wire u_multiplier_STAGE1__0846_ ;
 wire u_multiplier_STAGE1__0847_ ;
 wire u_multiplier_STAGE1__0848_ ;
 wire u_multiplier_STAGE1__0849_ ;
 wire u_multiplier_STAGE1__0850_ ;
 wire u_multiplier_STAGE1__0851_ ;
 wire u_multiplier_STAGE1__0852_ ;
 wire u_multiplier_STAGE1__0853_ ;
 wire u_multiplier_STAGE1__0854_ ;
 wire u_multiplier_STAGE1__0855_ ;
 wire u_multiplier_STAGE1__0856_ ;
 wire u_multiplier_STAGE1__0857_ ;
 wire u_multiplier_STAGE1__0858_ ;
 wire u_multiplier_STAGE1__0859_ ;
 wire u_multiplier_STAGE1__0860_ ;
 wire u_multiplier_STAGE1__0861_ ;
 wire u_multiplier_STAGE1__0862_ ;
 wire u_multiplier_STAGE1__0863_ ;
 wire u_multiplier_STAGE1__0864_ ;
 wire u_multiplier_STAGE1__0865_ ;
 wire u_multiplier_STAGE1__0866_ ;
 wire u_multiplier_STAGE1__0867_ ;
 wire u_multiplier_STAGE1__0868_ ;
 wire u_multiplier_STAGE1__0869_ ;
 wire u_multiplier_STAGE1__0870_ ;
 wire u_multiplier_STAGE1__0871_ ;
 wire u_multiplier_STAGE1__0872_ ;
 wire u_multiplier_STAGE1__0873_ ;
 wire u_multiplier_STAGE1__0874_ ;
 wire u_multiplier_STAGE1__0875_ ;
 wire u_multiplier_STAGE1__0876_ ;
 wire u_multiplier_STAGE1__0877_ ;
 wire u_multiplier_STAGE1__0878_ ;
 wire u_multiplier_STAGE1__0879_ ;
 wire u_multiplier_STAGE1__0880_ ;
 wire u_multiplier_STAGE1__0881_ ;
 wire u_multiplier_STAGE1__0882_ ;
 wire u_multiplier_STAGE1__0883_ ;
 wire u_multiplier_STAGE1__0884_ ;
 wire u_multiplier_STAGE1__0885_ ;
 wire u_multiplier_STAGE1__0886_ ;
 wire u_multiplier_STAGE1__0887_ ;
 wire u_multiplier_STAGE1__0888_ ;
 wire u_multiplier_STAGE1__0889_ ;
 wire u_multiplier_STAGE1__0890_ ;
 wire u_multiplier_STAGE1__0891_ ;
 wire u_multiplier_STAGE1__0892_ ;
 wire u_multiplier_STAGE1__0893_ ;
 wire u_multiplier_STAGE1__0894_ ;
 wire u_multiplier_STAGE1__0895_ ;
 wire u_multiplier_STAGE1__0896_ ;
 wire u_multiplier_STAGE1__0897_ ;
 wire u_multiplier_STAGE1__0898_ ;
 wire u_multiplier_STAGE1__0899_ ;
 wire u_multiplier_STAGE1__0900_ ;
 wire u_multiplier_STAGE1__0901_ ;
 wire u_multiplier_STAGE1__0902_ ;
 wire u_multiplier_STAGE1__0903_ ;
 wire u_multiplier_STAGE1__0904_ ;
 wire u_multiplier_STAGE1__0905_ ;
 wire u_multiplier_STAGE1__0906_ ;
 wire u_multiplier_STAGE1__0907_ ;
 wire u_multiplier_STAGE1__0908_ ;
 wire u_multiplier_STAGE1__0909_ ;
 wire u_multiplier_STAGE1__0910_ ;
 wire u_multiplier_STAGE1__0911_ ;
 wire u_multiplier_STAGE1__0912_ ;
 wire u_multiplier_STAGE1__0913_ ;
 wire u_multiplier_STAGE1__0914_ ;
 wire u_multiplier_STAGE1__0915_ ;
 wire u_multiplier_STAGE1__0916_ ;
 wire u_multiplier_STAGE1__0917_ ;
 wire u_multiplier_STAGE1__0918_ ;
 wire u_multiplier_STAGE1__0919_ ;
 wire u_multiplier_STAGE1__0920_ ;
 wire u_multiplier_STAGE1__0921_ ;
 wire u_multiplier_STAGE1__0922_ ;
 wire u_multiplier_STAGE1__0923_ ;
 wire u_multiplier_STAGE1__0924_ ;
 wire u_multiplier_STAGE1__0925_ ;
 wire u_multiplier_STAGE1__0926_ ;
 wire u_multiplier_STAGE1__0927_ ;
 wire u_multiplier_STAGE1__0928_ ;
 wire u_multiplier_STAGE1__0929_ ;
 wire u_multiplier_STAGE1__0930_ ;
 wire u_multiplier_STAGE1__0931_ ;
 wire u_multiplier_STAGE1__0932_ ;
 wire u_multiplier_STAGE1__0933_ ;
 wire u_multiplier_STAGE1__0934_ ;
 wire u_multiplier_STAGE1__0935_ ;
 wire u_multiplier_STAGE1__0936_ ;
 wire u_multiplier_STAGE1__0937_ ;
 wire u_multiplier_STAGE1__0938_ ;
 wire u_multiplier_STAGE1__0939_ ;
 wire u_multiplier_STAGE1__0940_ ;
 wire u_multiplier_STAGE1__0941_ ;
 wire u_multiplier_STAGE1__0942_ ;
 wire u_multiplier_STAGE1__0943_ ;
 wire u_multiplier_STAGE1__0944_ ;
 wire u_multiplier_STAGE1__0945_ ;
 wire u_multiplier_STAGE1__0946_ ;
 wire u_multiplier_STAGE1__0947_ ;
 wire u_multiplier_STAGE1__0948_ ;
 wire u_multiplier_STAGE1__0949_ ;
 wire u_multiplier_STAGE1__0950_ ;
 wire u_multiplier_STAGE1__0951_ ;
 wire u_multiplier_STAGE1__0952_ ;
 wire u_multiplier_STAGE1__0953_ ;
 wire u_multiplier_STAGE1__0954_ ;
 wire u_multiplier_STAGE1__0955_ ;
 wire u_multiplier_STAGE1__0956_ ;
 wire u_multiplier_STAGE1__0957_ ;
 wire u_multiplier_STAGE1__0958_ ;
 wire u_multiplier_STAGE1__0959_ ;
 wire u_multiplier_STAGE1__0960_ ;
 wire u_multiplier_STAGE1__0961_ ;
 wire u_multiplier_STAGE1__0962_ ;
 wire u_multiplier_STAGE1__0963_ ;
 wire u_multiplier_STAGE1__0964_ ;
 wire u_multiplier_STAGE1__0965_ ;
 wire u_multiplier_STAGE1__0966_ ;
 wire u_multiplier_STAGE1__0967_ ;
 wire u_multiplier_STAGE1__0968_ ;
 wire u_multiplier_STAGE1__0969_ ;
 wire u_multiplier_STAGE1__0970_ ;
 wire u_multiplier_STAGE1__0971_ ;
 wire u_multiplier_STAGE1__0972_ ;
 wire u_multiplier_STAGE1__0973_ ;
 wire u_multiplier_STAGE1__0974_ ;
 wire u_multiplier_STAGE1__0975_ ;
 wire u_multiplier_STAGE1__0976_ ;
 wire u_multiplier_STAGE1__0977_ ;
 wire u_multiplier_STAGE1__0978_ ;
 wire u_multiplier_STAGE1__0979_ ;
 wire u_multiplier_STAGE1__0980_ ;
 wire u_multiplier_STAGE1__0981_ ;
 wire u_multiplier_STAGE1__0982_ ;
 wire u_multiplier_STAGE1__0983_ ;
 wire u_multiplier_STAGE1__0984_ ;
 wire u_multiplier_STAGE1__0985_ ;
 wire u_multiplier_STAGE1__0986_ ;
 wire u_multiplier_STAGE1__0987_ ;
 wire u_multiplier_STAGE1__0988_ ;
 wire u_multiplier_STAGE1__0989_ ;
 wire u_multiplier_STAGE1__0990_ ;
 wire u_multiplier_STAGE1__0991_ ;
 wire u_multiplier_STAGE1__0992_ ;
 wire u_multiplier_STAGE1__0993_ ;
 wire u_multiplier_STAGE1__0994_ ;
 wire u_multiplier_STAGE1__0995_ ;
 wire u_multiplier_STAGE1__0996_ ;
 wire u_multiplier_STAGE1__0997_ ;
 wire u_multiplier_STAGE1__0998_ ;
 wire u_multiplier_STAGE1__0999_ ;
 wire u_multiplier_STAGE1__1000_ ;
 wire u_multiplier_STAGE1__1001_ ;
 wire u_multiplier_STAGE1__1002_ ;
 wire u_multiplier_STAGE1__1003_ ;
 wire u_multiplier_STAGE1__1004_ ;
 wire u_multiplier_STAGE1__1005_ ;
 wire u_multiplier_STAGE1__1006_ ;
 wire u_multiplier_STAGE1__1007_ ;
 wire u_multiplier_STAGE1__1008_ ;
 wire u_multiplier_STAGE1__1009_ ;
 wire u_multiplier_STAGE1__1010_ ;
 wire u_multiplier_STAGE1__1011_ ;
 wire u_multiplier_STAGE1__1012_ ;
 wire u_multiplier_STAGE1__1013_ ;
 wire u_multiplier_STAGE1__1014_ ;
 wire u_multiplier_STAGE1__1015_ ;
 wire u_multiplier_STAGE1__1016_ ;
 wire u_multiplier_STAGE1__1017_ ;
 wire u_multiplier_STAGE1__1018_ ;
 wire u_multiplier_STAGE1__1019_ ;
 wire u_multiplier_STAGE1__1020_ ;
 wire u_multiplier_STAGE1__1021_ ;
 wire u_multiplier_STAGE1__1022_ ;
 wire u_multiplier_STAGE1__1023_ ;
 wire u_multiplier_STAGE1__1024_ ;
 wire u_multiplier_STAGE1__1025_ ;
 wire u_multiplier_STAGE1__1026_ ;
 wire u_multiplier_STAGE1__1027_ ;
 wire u_multiplier_STAGE1__1028_ ;
 wire u_multiplier_STAGE1__1029_ ;
 wire u_multiplier_STAGE1__1030_ ;
 wire u_multiplier_STAGE1__1031_ ;
 wire u_multiplier_STAGE1__1032_ ;
 wire u_multiplier_STAGE1__1033_ ;
 wire u_multiplier_STAGE1__1034_ ;
 wire u_multiplier_STAGE1__1035_ ;
 wire u_multiplier_STAGE1__1036_ ;
 wire u_multiplier_STAGE1__1037_ ;
 wire u_multiplier_STAGE1__1038_ ;
 wire u_multiplier_STAGE1__1039_ ;
 wire u_multiplier_STAGE1__1040_ ;
 wire u_multiplier_STAGE1__1041_ ;
 wire u_multiplier_STAGE1__1042_ ;
 wire u_multiplier_STAGE1__1043_ ;
 wire u_multiplier_STAGE1__1044_ ;
 wire u_multiplier_STAGE1__1045_ ;
 wire u_multiplier_STAGE1__1046_ ;
 wire u_multiplier_STAGE1__1047_ ;
 wire u_multiplier_STAGE1__1048_ ;
 wire u_multiplier_STAGE1__1049_ ;
 wire u_multiplier_STAGE1__1050_ ;
 wire u_multiplier_STAGE1__1051_ ;
 wire u_multiplier_STAGE1__1052_ ;
 wire u_multiplier_STAGE1__1053_ ;
 wire u_multiplier_STAGE1__1054_ ;
 wire u_multiplier_STAGE1__1055_ ;
 wire u_multiplier_STAGE1__1056_ ;
 wire u_multiplier_STAGE1__1057_ ;
 wire u_multiplier_STAGE1__1058_ ;
 wire u_multiplier_STAGE1__1059_ ;
 wire u_multiplier_STAGE1__1060_ ;
 wire u_multiplier_STAGE1__1061_ ;
 wire u_multiplier_STAGE1__1062_ ;
 wire u_multiplier_STAGE1__1063_ ;
 wire u_multiplier_STAGE1__1064_ ;
 wire u_multiplier_STAGE1__1065_ ;
 wire u_multiplier_STAGE1__1066_ ;
 wire u_multiplier_STAGE1__1067_ ;
 wire u_multiplier_STAGE1__1068_ ;
 wire u_multiplier_STAGE1__1069_ ;
 wire u_multiplier_STAGE1__1070_ ;
 wire u_multiplier_STAGE1__1071_ ;
 wire u_multiplier_STAGE1__1072_ ;
 wire u_multiplier_STAGE1__1073_ ;
 wire u_multiplier_STAGE1__1074_ ;
 wire u_multiplier_STAGE1__1075_ ;
 wire u_multiplier_STAGE1__1076_ ;
 wire u_multiplier_STAGE1__1077_ ;
 wire u_multiplier_STAGE1__1078_ ;
 wire u_multiplier_STAGE1__1079_ ;
 wire u_multiplier_STAGE1__1080_ ;
 wire u_multiplier_STAGE1__1081_ ;
 wire u_multiplier_STAGE1__1082_ ;
 wire u_multiplier_STAGE1__1083_ ;
 wire u_multiplier_STAGE1__1084_ ;
 wire u_multiplier_STAGE1__1085_ ;
 wire u_multiplier_STAGE1__1086_ ;
 wire u_multiplier_STAGE1__1087_ ;
 wire u_multiplier_STAGE1__1088_ ;
 wire u_multiplier_STAGE1__1089_ ;
 wire u_multiplier_STAGE1__1090_ ;
 wire u_multiplier_STAGE1__1091_ ;
 wire u_multiplier_STAGE1__1092_ ;
 wire u_multiplier_STAGE1__1093_ ;
 wire u_multiplier_STAGE1__1094_ ;
 wire u_multiplier_STAGE1__1095_ ;
 wire u_multiplier_STAGE1__1096_ ;
 wire u_multiplier_STAGE1__1097_ ;
 wire u_multiplier_STAGE1__1098_ ;
 wire u_multiplier_STAGE1__1099_ ;
 wire u_multiplier_STAGE1__1100_ ;
 wire u_multiplier_STAGE1__1101_ ;
 wire u_multiplier_STAGE1__1102_ ;
 wire u_multiplier_STAGE1__1103_ ;
 wire u_multiplier_STAGE1__1104_ ;
 wire u_multiplier_STAGE1__1105_ ;
 wire u_multiplier_STAGE1__1106_ ;
 wire u_multiplier_STAGE1__1107_ ;
 wire u_multiplier_STAGE1__1108_ ;
 wire u_multiplier_STAGE1__1109_ ;
 wire u_multiplier_STAGE1__1110_ ;
 wire u_multiplier_STAGE1__1111_ ;
 wire u_multiplier_STAGE1__1112_ ;
 wire u_multiplier_STAGE1__1113_ ;
 wire u_multiplier_STAGE1__1114_ ;
 wire u_multiplier_STAGE1__1115_ ;
 wire u_multiplier_STAGE1__1116_ ;
 wire u_multiplier_STAGE1__1117_ ;
 wire u_multiplier_STAGE1__1118_ ;
 wire u_multiplier_STAGE1__1119_ ;
 wire u_multiplier_STAGE1__1120_ ;
 wire u_multiplier_STAGE1__1121_ ;
 wire u_multiplier_STAGE1__1122_ ;
 wire u_multiplier_STAGE1__1123_ ;
 wire u_multiplier_STAGE1__1124_ ;
 wire u_multiplier_STAGE1__1125_ ;
 wire u_multiplier_STAGE1__1126_ ;
 wire u_multiplier_STAGE1__1127_ ;
 wire u_multiplier_STAGE1__1128_ ;
 wire u_multiplier_STAGE1__1129_ ;
 wire u_multiplier_STAGE1__1130_ ;
 wire u_multiplier_STAGE1__1131_ ;
 wire u_multiplier_STAGE1__1132_ ;
 wire u_multiplier_STAGE1__1133_ ;
 wire u_multiplier_STAGE1__1134_ ;
 wire u_multiplier_STAGE1__1135_ ;
 wire u_multiplier_STAGE1__1136_ ;
 wire u_multiplier_STAGE1__1137_ ;
 wire u_multiplier_STAGE1__1138_ ;
 wire u_multiplier_STAGE1__1139_ ;
 wire u_multiplier_STAGE1__1140_ ;
 wire u_multiplier_STAGE1__1141_ ;
 wire u_multiplier_STAGE1__1142_ ;
 wire u_multiplier_STAGE1__1143_ ;
 wire u_multiplier_STAGE1__1144_ ;
 wire u_multiplier_STAGE1__1145_ ;
 wire u_multiplier_STAGE1__1146_ ;
 wire u_multiplier_STAGE1__1147_ ;
 wire u_multiplier_STAGE1__1148_ ;
 wire u_multiplier_STAGE1__1149_ ;
 wire net133;
 wire u_multiplier_STAGE1_pp1_17_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_18_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_19_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_19_e42_2_cout ;
 wire u_multiplier_STAGE1_pp1_20_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_20_e42_2_cout ;
 wire u_multiplier_STAGE1_pp1_21_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_21_e42_2_cout ;
 wire u_multiplier_STAGE1_pp1_21_e42_3_cout ;
 wire u_multiplier_STAGE1_pp1_22_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_22_e42_2_cout ;
 wire u_multiplier_STAGE1_pp1_22_e42_3_cout ;
 wire u_multiplier_STAGE1_pp1_23_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_23_e42_2_cout ;
 wire u_multiplier_STAGE1_pp1_23_e42_3_cout ;
 wire u_multiplier_STAGE1_pp1_23_e42_4_cout ;
 wire u_multiplier_STAGE1_pp1_24_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_24_e42_2_cout ;
 wire u_multiplier_STAGE1_pp1_24_e42_3_cout ;
 wire u_multiplier_STAGE1_pp1_24_e42_4_cout ;
 wire u_multiplier_STAGE1_pp1_25_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_25_e42_2_cout ;
 wire u_multiplier_STAGE1_pp1_25_e42_3_cout ;
 wire u_multiplier_STAGE1_pp1_25_e42_4_cout ;
 wire u_multiplier_STAGE1_pp1_25_e42_5_cout ;
 wire u_multiplier_STAGE1_pp1_26_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_26_e42_2_cout ;
 wire u_multiplier_STAGE1_pp1_26_e42_3_cout ;
 wire u_multiplier_STAGE1_pp1_26_e42_4_cout ;
 wire u_multiplier_STAGE1_pp1_26_e42_5_cout ;
 wire u_multiplier_STAGE1_pp1_27_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_27_e42_2_cout ;
 wire u_multiplier_STAGE1_pp1_27_e42_3_cout ;
 wire u_multiplier_STAGE1_pp1_27_e42_4_cout ;
 wire u_multiplier_STAGE1_pp1_27_e42_5_cout ;
 wire u_multiplier_STAGE1_pp1_27_e42_6_cout ;
 wire u_multiplier_STAGE1_pp1_28_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_28_e42_2_cout ;
 wire u_multiplier_STAGE1_pp1_28_e42_3_cout ;
 wire u_multiplier_STAGE1_pp1_28_e42_4_cout ;
 wire u_multiplier_STAGE1_pp1_28_e42_5_cout ;
 wire u_multiplier_STAGE1_pp1_28_e42_6_cout ;
 wire u_multiplier_STAGE1_pp1_29_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_29_e42_2_cout ;
 wire u_multiplier_STAGE1_pp1_29_e42_3_cout ;
 wire u_multiplier_STAGE1_pp1_29_e42_4_cout ;
 wire u_multiplier_STAGE1_pp1_29_e42_5_cout ;
 wire u_multiplier_STAGE1_pp1_29_e42_6_cout ;
 wire u_multiplier_STAGE1_pp1_29_e42_7_cout ;
 wire u_multiplier_STAGE1_pp1_30_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_30_e42_2_cout ;
 wire u_multiplier_STAGE1_pp1_30_e42_3_cout ;
 wire u_multiplier_STAGE1_pp1_30_e42_4_cout ;
 wire u_multiplier_STAGE1_pp1_30_e42_5_cout ;
 wire u_multiplier_STAGE1_pp1_30_e42_6_cout ;
 wire u_multiplier_STAGE1_pp1_30_e42_7_cout ;
 wire u_multiplier_STAGE1_pp1_31_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_31_e42_2_cout ;
 wire u_multiplier_STAGE1_pp1_31_e42_3_cout ;
 wire u_multiplier_STAGE1_pp1_31_e42_4_cout ;
 wire u_multiplier_STAGE1_pp1_31_e42_5_cout ;
 wire u_multiplier_STAGE1_pp1_31_e42_6_cout ;
 wire u_multiplier_STAGE1_pp1_31_e42_7_cout ;
 wire u_multiplier_STAGE1_pp1_31_e42_8_cout ;
 wire u_multiplier_STAGE1_pp1_32_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_32_e42_2_cout ;
 wire u_multiplier_STAGE1_pp1_32_e42_3_cout ;
 wire u_multiplier_STAGE1_pp1_32_e42_4_cout ;
 wire u_multiplier_STAGE1_pp1_32_e42_5_cout ;
 wire u_multiplier_STAGE1_pp1_32_e42_6_cout ;
 wire u_multiplier_STAGE1_pp1_32_e42_7_cout ;
 wire u_multiplier_STAGE1_pp1_32_e42_8_cout ;
 wire u_multiplier_STAGE1_pp1_33_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_33_e42_2_cout ;
 wire u_multiplier_STAGE1_pp1_33_e42_3_cout ;
 wire u_multiplier_STAGE1_pp1_33_e42_4_cout ;
 wire u_multiplier_STAGE1_pp1_33_e42_5_cout ;
 wire u_multiplier_STAGE1_pp1_33_e42_6_cout ;
 wire u_multiplier_STAGE1_pp1_33_e42_7_cout ;
 wire u_multiplier_STAGE1_pp1_34_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_34_e42_2_cout ;
 wire u_multiplier_STAGE1_pp1_34_e42_3_cout ;
 wire u_multiplier_STAGE1_pp1_34_e42_4_cout ;
 wire u_multiplier_STAGE1_pp1_34_e42_5_cout ;
 wire u_multiplier_STAGE1_pp1_34_e42_6_cout ;
 wire u_multiplier_STAGE1_pp1_34_e42_7_cout ;
 wire u_multiplier_STAGE1_pp1_35_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_35_e42_2_cout ;
 wire u_multiplier_STAGE1_pp1_35_e42_3_cout ;
 wire u_multiplier_STAGE1_pp1_35_e42_4_cout ;
 wire u_multiplier_STAGE1_pp1_35_e42_5_cout ;
 wire u_multiplier_STAGE1_pp1_35_e42_6_cout ;
 wire u_multiplier_STAGE1_pp1_36_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_36_e42_2_cout ;
 wire u_multiplier_STAGE1_pp1_36_e42_3_cout ;
 wire u_multiplier_STAGE1_pp1_36_e42_4_cout ;
 wire u_multiplier_STAGE1_pp1_36_e42_5_cout ;
 wire u_multiplier_STAGE1_pp1_36_e42_6_cout ;
 wire u_multiplier_STAGE1_pp1_37_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_37_e42_2_cout ;
 wire u_multiplier_STAGE1_pp1_37_e42_3_cout ;
 wire u_multiplier_STAGE1_pp1_37_e42_4_cout ;
 wire u_multiplier_STAGE1_pp1_37_e42_5_cout ;
 wire u_multiplier_STAGE1_pp1_38_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_38_e42_2_cout ;
 wire u_multiplier_STAGE1_pp1_38_e42_3_cout ;
 wire u_multiplier_STAGE1_pp1_38_e42_4_cout ;
 wire u_multiplier_STAGE1_pp1_38_e42_5_cout ;
 wire u_multiplier_STAGE1_pp1_39_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_39_e42_2_cout ;
 wire u_multiplier_STAGE1_pp1_39_e42_3_cout ;
 wire u_multiplier_STAGE1_pp1_39_e42_4_cout ;
 wire u_multiplier_STAGE1_pp1_40_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_40_e42_2_cout ;
 wire u_multiplier_STAGE1_pp1_40_e42_3_cout ;
 wire u_multiplier_STAGE1_pp1_40_e42_4_cout ;
 wire u_multiplier_STAGE1_pp1_41_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_41_e42_2_cout ;
 wire u_multiplier_STAGE1_pp1_41_e42_3_cout ;
 wire u_multiplier_STAGE1_pp1_42_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_42_e42_2_cout ;
 wire u_multiplier_STAGE1_pp1_42_e42_3_cout ;
 wire u_multiplier_STAGE1_pp1_43_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_43_e42_2_cout ;
 wire u_multiplier_STAGE1_pp1_44_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_44_e42_2_cout ;
 wire u_multiplier_STAGE1_pp1_45_e42_1_cout ;
 wire u_multiplier_STAGE1_pp1_46_e42_1_cout ;
 wire u_multiplier_STAGE1_E_4_2_pp_17_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_17_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_17_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_17_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_17_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_17_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_17_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_18_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_18_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_18_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_18_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_18_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_18_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_18_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_19_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_19_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_19_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_19_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_19_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_19_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_19_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_19_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_19_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_19_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_19_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_19_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_19_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_19_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_20_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_20_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_20_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_20_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_20_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_20_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_20_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_20_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_20_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_20_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_20_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_20_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_20_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_20_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_21_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_21_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_21_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_21_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_21_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_21_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_21_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_21_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_21_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_21_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_21_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_21_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_21_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_21_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_21_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_21_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_21_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_21_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_21_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_21_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_21_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_22_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_22_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_22_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_22_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_22_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_22_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_22_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_22_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_22_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_22_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_22_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_22_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_22_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_22_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_22_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_22_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_22_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_22_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_22_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_22_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_22_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_4__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_4__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_4__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_4__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_4__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_4__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_23_4__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_4__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_4__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_4__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_4__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_4__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_4__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_24_4__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_4__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_4__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_4__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_4__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_4__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_4__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_4__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_5__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_5__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_5__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_5__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_5__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_5__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_25_5__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_4__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_4__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_4__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_4__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_4__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_4__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_4__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_5__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_5__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_5__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_5__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_5__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_5__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_26_5__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_4__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_4__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_4__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_4__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_4__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_4__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_4__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_5__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_5__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_5__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_5__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_5__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_5__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_5__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_6__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_6__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_6__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_6__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_6__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_6__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_27_6__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_4__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_4__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_4__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_4__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_4__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_4__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_4__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_5__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_5__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_5__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_5__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_5__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_5__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_5__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_6__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_6__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_6__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_6__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_6__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_6__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_28_6__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_4__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_4__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_4__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_4__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_4__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_4__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_4__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_5__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_5__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_5__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_5__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_5__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_5__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_5__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_6__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_6__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_6__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_6__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_6__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_6__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_6__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_7__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_7__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_7__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_7__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_7__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_7__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_29_7__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_4__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_4__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_4__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_4__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_4__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_4__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_4__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_5__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_5__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_5__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_5__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_5__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_5__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_5__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_6__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_6__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_6__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_6__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_6__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_6__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_6__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_7__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_7__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_7__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_7__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_7__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_7__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_30_7__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_4__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_4__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_4__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_4__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_4__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_4__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_4__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_5__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_5__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_5__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_5__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_5__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_5__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_5__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_6__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_6__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_6__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_6__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_6__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_6__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_6__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_7__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_7__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_7__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_7__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_7__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_7__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_7__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_8__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_8__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_8__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_8__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_8__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_8__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_31_8__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_4__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_4__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_4__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_4__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_4__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_4__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_4__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_5__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_5__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_5__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_5__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_5__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_5__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_5__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_6__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_6__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_6__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_6__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_6__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_6__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_6__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_7__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_7__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_7__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_7__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_7__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_7__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_7__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_8__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_8__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_8__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_8__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_8__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_8__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_8__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_4__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_4__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_4__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_4__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_4__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_4__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_4__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_5__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_5__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_5__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_5__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_5__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_5__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_5__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_6__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_6__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_6__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_6__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_6__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_6__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_6__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_7__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_7__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_7__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_7__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_7__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_7__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_7__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_4__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_4__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_4__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_4__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_4__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_4__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_4__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_5__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_5__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_5__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_5__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_5__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_5__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_5__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_6__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_6__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_6__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_6__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_6__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_6__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_6__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_7__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_7__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_7__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_7__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_7__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_7__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_7__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_4__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_4__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_4__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_4__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_4__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_4__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_4__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_5__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_5__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_5__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_5__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_5__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_5__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_5__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_6__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_6__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_6__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_6__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_6__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_6__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_6__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_4__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_4__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_4__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_4__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_4__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_4__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_4__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_5__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_5__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_5__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_5__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_5__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_5__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_5__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_6__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_6__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_6__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_6__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_6__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_6__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_6__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_4__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_4__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_4__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_4__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_4__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_4__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_4__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_5__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_5__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_5__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_5__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_5__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_5__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_5__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_4__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_4__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_4__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_4__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_4__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_4__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_4__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_5__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_5__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_5__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_5__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_5__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_5__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_5__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_4__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_4__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_4__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_4__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_4__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_4__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_4__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_4__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_4__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_4__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_4__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_4__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_4__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_4__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_45_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_45_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_45_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_45_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_45_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_45_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_45_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_46_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_46_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_46_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_46_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_46_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_46_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_46_1__17_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_33_1__08_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_33_1__09_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_33_1__10_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_33_1__11_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_35_1__08_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_35_1__09_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_35_1__10_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_35_1__11_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_37_1__08_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_37_1__09_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_37_1__10_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_37_1__11_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_39_1__08_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_39_1__09_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_39_1__10_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_39_1__11_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_41_1__08_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_41_1__09_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_41_1__10_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_41_1__11_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_43_1__08_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_43_1__09_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_43_1__10_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_43_1__11_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_45_1__08_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_45_1__09_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_45_1__10_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_45_1__11_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_47_1__08_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_47_1__09_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_47_1__10_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_47_1__11_ ;
 wire u_multiplier_STAGE2_pp2_10_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_11_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_11_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_12_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_12_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_13_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_13_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_13_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_14_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_14_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_14_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_15_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_15_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_15_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_15_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_16_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_16_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_16_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_16_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_17_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_17_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_17_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_17_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_18_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_18_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_18_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_18_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_19_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_19_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_19_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_19_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_20_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_20_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_20_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_20_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_21_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_21_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_21_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_21_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_22_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_22_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_22_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_22_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_23_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_23_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_23_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_23_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_24_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_24_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_24_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_24_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_25_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_25_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_25_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_25_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_26_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_26_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_26_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_26_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_27_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_27_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_27_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_27_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_28_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_28_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_28_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_28_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_29_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_29_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_29_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_29_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_30_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_30_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_30_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_30_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_31_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_31_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_31_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_31_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_32_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_32_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_32_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_32_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_33_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_33_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_33_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_33_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_34_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_34_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_34_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_34_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_35_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_35_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_35_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_35_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_36_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_36_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_36_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_36_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_37_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_37_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_37_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_37_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_38_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_38_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_38_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_38_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_39_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_39_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_39_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_39_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_40_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_40_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_40_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_40_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_41_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_41_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_41_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_41_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_42_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_42_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_42_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_42_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_43_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_43_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_43_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_43_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_44_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_44_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_44_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_44_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_45_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_45_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_45_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_45_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_46_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_46_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_46_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_46_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_47_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_47_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_47_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_47_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_48_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_48_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_48_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_48_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_49_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_49_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_49_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_50_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_50_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_50_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_51_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_51_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_52_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_52_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_53_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_54_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_9_e42_1_cout ;
 wire u_multiplier_STAGE2_E_4_2_pp2_10_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_10_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_10_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_10_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_10_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_10_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_10_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_11_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_11_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_11_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_11_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_11_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_11_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_11_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_11_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_11_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_11_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_11_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_11_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_11_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_11_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_12_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_12_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_12_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_12_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_12_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_12_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_12_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_12_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_12_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_12_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_12_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_12_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_12_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_12_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_13_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_13_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_13_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_13_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_13_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_13_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_13_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_13_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_13_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_13_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_13_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_13_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_13_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_13_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_13_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_13_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_13_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_13_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_13_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_13_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_13_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_14_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_14_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_14_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_14_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_14_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_14_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_14_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_14_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_14_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_14_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_14_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_14_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_14_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_14_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_14_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_14_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_14_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_14_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_14_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_14_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_14_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_15_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_16_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_17_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_18_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_19_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_20_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_21_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_22_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_23_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_24_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_25_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_26_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_27_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_28_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_29_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_30_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_31_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_53_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_53_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_53_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_53_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_53_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_53_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_53_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_54_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_54_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_54_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_54_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_54_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_54_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_54_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_9_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_9_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_9_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_9_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_9_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_9_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_9_1__17_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_49_1__08_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_49_1__09_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_49_1__10_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_49_1__11_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_51_1__08_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_51_1__09_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_51_1__10_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_51_1__11_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_53_1__08_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_53_1__09_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_53_1__10_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_53_1__11_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_55_1__08_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_55_1__09_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_55_1__10_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_55_1__11_ ;
 wire u_multiplier_STAGE3_pp3_10_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_10_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_11_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_11_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_12_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_12_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_13_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_13_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_14_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_14_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_15_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_15_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_16_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_16_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_17_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_17_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_18_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_18_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_19_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_19_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_20_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_20_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_21_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_21_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_22_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_22_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_23_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_23_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_24_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_24_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_25_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_25_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_26_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_26_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_27_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_27_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_28_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_28_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_29_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_29_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_30_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_30_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_31_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_31_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_32_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_32_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_33_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_33_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_34_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_34_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_35_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_35_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_36_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_36_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_37_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_37_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_38_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_38_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_39_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_39_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_40_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_40_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_41_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_41_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_42_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_42_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_43_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_43_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_44_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_44_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_45_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_45_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_46_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_46_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_47_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_47_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_48_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_48_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_49_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_49_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_50_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_50_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_51_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_51_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_52_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_52_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_53_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_53_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_54_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_54_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_55_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_55_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_56_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_56_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_57_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_58_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_5_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_6_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_7_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_7_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_8_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_8_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_9_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_9_e42_2_cout ;
 wire u_multiplier_STAGE3_E_4_2_pp3_10_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_10_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_10_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_10_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_10_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_10_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_10_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_10_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_10_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_10_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_10_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_10_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_10_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_10_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_11_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_11_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_11_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_11_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_11_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_11_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_11_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_11_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_11_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_11_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_11_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_11_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_11_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_11_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_12_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_12_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_12_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_12_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_12_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_12_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_12_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_12_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_12_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_12_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_12_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_12_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_12_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_12_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_13_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_13_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_13_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_13_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_13_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_13_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_13_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_13_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_13_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_13_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_13_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_13_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_13_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_13_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_14_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_14_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_14_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_14_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_14_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_14_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_14_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_14_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_14_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_14_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_14_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_14_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_14_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_14_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_15_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_15_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_15_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_15_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_15_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_15_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_15_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_15_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_15_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_15_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_15_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_15_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_15_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_15_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_16_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_16_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_16_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_16_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_16_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_16_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_16_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_16_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_16_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_16_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_16_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_16_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_16_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_16_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_17_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_17_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_17_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_17_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_17_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_17_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_17_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_17_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_17_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_17_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_17_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_17_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_17_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_17_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_18_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_18_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_18_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_18_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_18_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_18_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_18_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_18_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_18_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_18_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_18_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_18_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_18_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_18_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_19_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_19_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_19_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_19_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_19_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_19_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_19_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_19_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_19_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_19_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_19_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_19_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_19_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_19_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_20_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_20_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_20_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_20_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_20_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_20_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_20_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_20_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_20_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_20_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_20_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_20_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_20_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_20_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_21_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_21_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_21_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_21_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_21_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_21_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_21_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_21_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_21_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_21_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_21_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_21_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_21_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_21_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_22_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_22_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_22_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_22_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_22_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_22_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_22_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_22_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_22_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_22_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_22_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_22_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_22_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_22_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_23_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_23_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_23_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_23_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_23_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_23_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_23_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_23_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_23_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_23_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_23_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_23_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_23_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_23_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_24_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_24_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_24_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_24_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_24_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_24_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_24_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_24_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_24_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_24_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_24_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_24_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_24_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_24_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_25_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_25_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_25_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_25_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_25_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_25_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_25_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_25_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_25_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_25_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_25_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_25_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_25_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_25_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_26_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_26_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_26_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_26_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_26_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_26_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_26_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_26_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_26_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_26_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_26_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_26_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_26_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_26_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_27_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_27_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_27_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_27_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_27_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_27_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_27_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_27_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_27_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_27_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_27_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_27_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_27_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_27_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_28_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_28_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_28_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_28_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_28_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_28_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_28_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_28_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_28_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_28_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_28_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_28_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_28_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_28_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_29_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_29_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_29_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_29_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_29_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_29_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_29_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_29_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_29_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_29_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_29_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_29_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_29_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_29_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_30_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_30_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_30_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_30_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_30_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_30_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_30_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_30_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_30_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_30_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_30_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_30_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_30_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_30_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_31_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_31_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_31_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_31_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_31_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_31_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_31_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_31_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_31_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_31_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_31_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_31_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_31_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_31_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_57_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_57_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_57_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_57_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_57_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_57_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_57_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_58_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_58_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_58_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_58_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_58_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_58_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_58_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_5_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_5_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_5_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_5_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_5_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_5_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_5_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_6_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_6_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_6_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_6_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_6_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_6_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_6_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_7_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_7_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_7_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_7_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_7_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_7_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_7_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_7_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_7_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_7_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_7_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_7_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_7_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_7_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_8_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_8_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_8_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_8_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_8_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_8_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_8_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_8_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_8_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_8_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_8_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_8_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_8_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_8_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_9_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_9_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_9_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_9_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_9_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_9_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_9_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_9_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_9_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_9_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_9_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_9_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_9_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_9_2__17_ ;
 wire u_multiplier_STAGE3_Full_adder_pp3_57_1__08_ ;
 wire u_multiplier_STAGE3_Full_adder_pp3_57_1__09_ ;
 wire u_multiplier_STAGE3_Full_adder_pp3_57_1__10_ ;
 wire u_multiplier_STAGE3_Full_adder_pp3_57_1__11_ ;
 wire u_multiplier_STAGE3_Full_adder_pp3_59_1__08_ ;
 wire u_multiplier_STAGE3_Full_adder_pp3_59_1__09_ ;
 wire u_multiplier_STAGE3_Full_adder_pp3_59_1__10_ ;
 wire u_multiplier_STAGE3_Full_adder_pp3_59_1__11_ ;
 wire u_multiplier_STAGE4_pp4_10_cout ;
 wire u_multiplier_STAGE4_pp4_11_cout ;
 wire u_multiplier_STAGE4_pp4_12_cout ;
 wire u_multiplier_STAGE4_pp4_13_cout ;
 wire u_multiplier_STAGE4_pp4_14_cout ;
 wire u_multiplier_STAGE4_pp4_15_cout ;
 wire u_multiplier_STAGE4_pp4_16_cout ;
 wire u_multiplier_STAGE4_pp4_17_cout ;
 wire u_multiplier_STAGE4_pp4_18_cout ;
 wire u_multiplier_STAGE4_pp4_19_cout ;
 wire u_multiplier_STAGE4_pp4_1_ha_c ;
 wire u_multiplier_STAGE4_pp4_20_cout ;
 wire u_multiplier_STAGE4_pp4_21_cout ;
 wire u_multiplier_STAGE4_pp4_22_cout ;
 wire u_multiplier_STAGE4_pp4_23_cout ;
 wire u_multiplier_STAGE4_pp4_24_cout ;
 wire u_multiplier_STAGE4_pp4_25_cout ;
 wire u_multiplier_STAGE4_pp4_26_cout ;
 wire u_multiplier_STAGE4_pp4_27_cout ;
 wire u_multiplier_STAGE4_pp4_28_cout ;
 wire u_multiplier_STAGE4_pp4_29_cout ;
 wire u_multiplier_STAGE4_pp4_2_cout ;
 wire u_multiplier_STAGE4_pp4_30_cout ;
 wire u_multiplier_STAGE4_pp4_31_cout ;
 wire u_multiplier_STAGE4_pp4_32_cout ;
 wire u_multiplier_STAGE4_pp4_33_cout ;
 wire u_multiplier_STAGE4_pp4_34_cout ;
 wire u_multiplier_STAGE4_pp4_35_cout ;
 wire u_multiplier_STAGE4_pp4_36_cout ;
 wire u_multiplier_STAGE4_pp4_37_cout ;
 wire u_multiplier_STAGE4_pp4_38_cout ;
 wire u_multiplier_STAGE4_pp4_39_cout ;
 wire u_multiplier_STAGE4_pp4_3_cout ;
 wire u_multiplier_STAGE4_pp4_40_cout ;
 wire u_multiplier_STAGE4_pp4_41_cout ;
 wire u_multiplier_STAGE4_pp4_42_cout ;
 wire u_multiplier_STAGE4_pp4_43_cout ;
 wire u_multiplier_STAGE4_pp4_44_cout ;
 wire u_multiplier_STAGE4_pp4_45_cout ;
 wire u_multiplier_STAGE4_pp4_46_cout ;
 wire u_multiplier_STAGE4_pp4_47_cout ;
 wire u_multiplier_STAGE4_pp4_48_cout ;
 wire u_multiplier_STAGE4_pp4_49_cout ;
 wire u_multiplier_STAGE4_pp4_4_cout ;
 wire u_multiplier_STAGE4_pp4_50_cout ;
 wire u_multiplier_STAGE4_pp4_51_cout ;
 wire u_multiplier_STAGE4_pp4_52_cout ;
 wire u_multiplier_STAGE4_pp4_53_cout ;
 wire u_multiplier_STAGE4_pp4_54_cout ;
 wire u_multiplier_STAGE4_pp4_55_cout ;
 wire u_multiplier_STAGE4_pp4_56_cout ;
 wire u_multiplier_STAGE4_pp4_57_cout ;
 wire u_multiplier_STAGE4_pp4_58_cout ;
 wire u_multiplier_STAGE4_pp4_59_cout ;
 wire u_multiplier_STAGE4_pp4_5_cout ;
 wire u_multiplier_STAGE4_pp4_60_cout ;
 wire u_multiplier_STAGE4_pp4_6_cout ;
 wire u_multiplier_STAGE4_pp4_7_cout ;
 wire u_multiplier_STAGE4_pp4_8_cout ;
 wire u_multiplier_STAGE4_pp4_9_cout ;
 wire u_multiplier_STAGE4_E_4_2_pp4_10__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_10__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_10__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_10__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_10__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_10__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_10__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_11__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_11__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_11__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_11__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_11__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_11__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_11__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_12__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_12__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_12__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_12__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_12__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_12__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_12__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_13__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_13__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_13__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_13__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_13__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_13__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_13__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_14__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_14__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_14__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_14__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_14__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_14__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_14__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_15__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_15__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_15__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_15__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_15__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_15__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_15__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_16__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_16__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_16__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_16__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_16__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_16__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_16__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_17__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_17__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_17__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_17__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_17__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_17__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_17__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_18__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_18__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_18__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_18__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_18__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_18__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_18__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_19__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_19__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_19__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_19__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_19__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_19__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_19__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_2__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_2__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_2__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_2__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_2__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_2__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_2__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_20__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_20__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_20__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_20__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_20__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_20__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_20__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_21__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_21__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_21__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_21__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_21__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_21__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_21__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_22__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_22__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_22__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_22__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_22__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_22__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_22__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_23__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_23__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_23__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_23__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_23__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_23__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_23__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_24__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_24__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_24__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_24__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_24__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_24__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_24__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_25__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_25__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_25__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_25__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_25__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_25__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_25__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_26__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_26__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_26__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_26__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_26__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_26__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_26__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_27__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_27__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_27__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_27__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_27__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_27__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_27__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_28__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_28__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_28__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_28__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_28__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_28__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_28__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_29__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_29__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_29__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_29__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_29__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_29__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_29__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_3__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_3__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_3__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_3__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_3__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_3__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_3__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_30__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_30__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_30__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_30__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_30__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_30__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_30__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_31__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_31__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_31__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_31__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_31__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_31__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_31__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_32__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_32__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_32__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_32__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_32__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_32__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_32__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_33__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_33__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_33__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_33__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_33__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_33__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_33__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_34__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_34__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_34__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_34__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_34__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_34__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_34__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_35__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_35__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_35__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_35__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_35__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_35__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_35__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_36__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_36__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_36__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_36__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_36__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_36__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_36__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_37__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_37__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_37__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_37__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_37__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_37__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_37__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_38__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_38__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_38__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_38__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_38__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_38__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_38__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_39__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_39__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_39__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_39__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_39__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_39__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_39__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_4__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_4__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_4__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_4__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_4__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_4__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_4__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_40__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_40__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_40__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_40__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_40__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_40__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_40__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_41__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_41__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_41__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_41__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_41__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_41__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_41__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_42__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_42__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_42__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_42__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_42__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_42__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_42__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_43__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_43__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_43__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_43__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_43__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_43__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_43__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_44__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_44__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_44__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_44__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_44__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_44__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_44__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_45__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_45__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_45__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_45__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_45__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_45__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_45__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_46__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_46__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_46__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_46__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_46__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_46__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_46__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_47__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_47__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_47__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_47__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_47__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_47__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_47__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_48__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_48__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_48__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_48__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_48__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_48__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_48__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_49__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_49__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_49__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_49__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_49__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_49__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_49__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_5__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_5__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_5__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_5__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_5__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_5__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_5__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_50__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_50__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_50__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_50__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_50__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_50__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_50__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_51__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_51__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_51__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_51__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_51__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_51__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_51__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_52__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_52__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_52__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_52__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_52__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_52__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_52__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_53__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_53__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_53__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_53__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_53__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_53__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_53__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_54__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_54__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_54__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_54__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_54__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_54__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_54__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_55__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_55__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_55__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_55__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_55__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_55__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_55__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_56__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_56__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_56__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_56__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_56__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_56__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_56__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_57__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_57__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_57__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_57__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_57__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_57__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_57__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_58__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_58__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_58__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_58__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_58__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_58__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_58__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_59__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_59__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_59__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_59__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_59__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_59__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_59__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_6__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_6__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_6__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_6__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_6__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_6__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_6__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_60__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_60__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_60__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_60__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_60__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_60__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_60__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_7__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_7__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_7__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_7__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_7__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_7__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_7__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_8__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_8__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_8__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_8__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_8__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_8__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_8__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_9__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_9__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_9__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_9__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_9__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_9__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_9__17_ ;
 wire u_multiplier_STAGE4_Full_adder_pp4_61__08_ ;
 wire u_multiplier_STAGE4_Full_adder_pp4_61__09_ ;
 wire u_multiplier_STAGE4_Full_adder_pp4_61__10_ ;
 wire u_multiplier_STAGE4_Full_adder_pp4_61__11_ ;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire valid_reg_out;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net162;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire clknet_0_clk;
 wire clknet_1_0_0_clk;
 wire clknet_1_1_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_4_0__leaf_clk;
 wire clknet_4_1__leaf_clk;
 wire clknet_4_2__leaf_clk;
 wire clknet_4_3__leaf_clk;
 wire clknet_4_4__leaf_clk;
 wire clknet_4_5__leaf_clk;
 wire clknet_4_6__leaf_clk;
 wire clknet_4_7__leaf_clk;
 wire clknet_4_8__leaf_clk;
 wire clknet_4_9__leaf_clk;
 wire clknet_4_10__leaf_clk;
 wire clknet_4_11__leaf_clk;
 wire clknet_4_12__leaf_clk;
 wire clknet_4_13__leaf_clk;
 wire clknet_4_14__leaf_clk;
 wire clknet_4_15__leaf_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire [5:0] addr_ptr;
 wire [2:0] curr_state;
 wire [31:0] data_in_reg;
 wire [5:0] init_count;
 wire [63:0] product;
 wire [31:0] sram_rdata;
 wire [31:0] sram_rdata_reg;
 wire [63:0] u_multiplier_A ;
 wire [62:0] u_multiplier_B ;
 wire [1:0] u_multiplier_pp1_1 ;
 wire [10:0] u_multiplier_pp1_10 ;
 wire [11:0] u_multiplier_pp1_11 ;
 wire [12:0] u_multiplier_pp1_12 ;
 wire [13:0] u_multiplier_pp1_13 ;
 wire [14:0] u_multiplier_pp1_14 ;
 wire [15:0] u_multiplier_pp1_15 ;
 wire [15:0] u_multiplier_pp1_16 ;
 wire [15:0] u_multiplier_pp1_17 ;
 wire [15:0] u_multiplier_pp1_18 ;
 wire [15:0] u_multiplier_pp1_19 ;
 wire [2:0] u_multiplier_pp1_2 ;
 wire [15:0] u_multiplier_pp1_20 ;
 wire [15:0] u_multiplier_pp1_21 ;
 wire [15:0] u_multiplier_pp1_22 ;
 wire [15:0] u_multiplier_pp1_23 ;
 wire [15:0] u_multiplier_pp1_24 ;
 wire [15:0] u_multiplier_pp1_25 ;
 wire [15:0] u_multiplier_pp1_26 ;
 wire [15:0] u_multiplier_pp1_27 ;
 wire [15:0] u_multiplier_pp1_28 ;
 wire [15:0] u_multiplier_pp1_29 ;
 wire [3:0] u_multiplier_pp1_3 ;
 wire [15:0] u_multiplier_pp1_30 ;
 wire [15:0] u_multiplier_pp1_31 ;
 wire [15:0] u_multiplier_pp1_32 ;
 wire [15:0] u_multiplier_pp1_33 ;
 wire [15:0] u_multiplier_pp1_34 ;
 wire [15:0] u_multiplier_pp1_35 ;
 wire [15:0] u_multiplier_pp1_36 ;
 wire [15:0] u_multiplier_pp1_37 ;
 wire [15:0] u_multiplier_pp1_38 ;
 wire [15:0] u_multiplier_pp1_39 ;
 wire [4:0] u_multiplier_pp1_4 ;
 wire [15:0] u_multiplier_pp1_40 ;
 wire [15:0] u_multiplier_pp1_41 ;
 wire [15:0] u_multiplier_pp1_42 ;
 wire [15:0] u_multiplier_pp1_43 ;
 wire [15:0] u_multiplier_pp1_44 ;
 wire [15:0] u_multiplier_pp1_45 ;
 wire [15:0] u_multiplier_pp1_46 ;
 wire [15:0] u_multiplier_pp1_47 ;
 wire [15:0] u_multiplier_pp1_48 ;
 wire [13:0] u_multiplier_pp1_49 ;
 wire [5:0] u_multiplier_pp1_5 ;
 wire [12:0] u_multiplier_pp1_50 ;
 wire [11:0] u_multiplier_pp1_51 ;
 wire [10:0] u_multiplier_pp1_52 ;
 wire [9:0] u_multiplier_pp1_53 ;
 wire [8:0] u_multiplier_pp1_54 ;
 wire [7:0] u_multiplier_pp1_55 ;
 wire [6:0] u_multiplier_pp1_56 ;
 wire [5:0] u_multiplier_pp1_57 ;
 wire [4:0] u_multiplier_pp1_58 ;
 wire [3:0] u_multiplier_pp1_59 ;
 wire [6:0] u_multiplier_pp1_6 ;
 wire [2:0] u_multiplier_pp1_60 ;
 wire [1:0] u_multiplier_pp1_61 ;
 wire [7:0] u_multiplier_pp1_7 ;
 wire [8:0] u_multiplier_pp1_8 ;
 wire [9:0] u_multiplier_pp1_9 ;
 wire [1:0] u_multiplier_pp2_1 ;
 wire [7:0] u_multiplier_pp2_10 ;
 wire [7:0] u_multiplier_pp2_11 ;
 wire [7:0] u_multiplier_pp2_12 ;
 wire [7:0] u_multiplier_pp2_13 ;
 wire [7:0] u_multiplier_pp2_14 ;
 wire [7:0] u_multiplier_pp2_15 ;
 wire [7:0] u_multiplier_pp2_16 ;
 wire [7:0] u_multiplier_pp2_17 ;
 wire [7:0] u_multiplier_pp2_18 ;
 wire [7:0] u_multiplier_pp2_19 ;
 wire [2:0] u_multiplier_pp2_2 ;
 wire [7:0] u_multiplier_pp2_20 ;
 wire [7:0] u_multiplier_pp2_21 ;
 wire [7:0] u_multiplier_pp2_22 ;
 wire [7:0] u_multiplier_pp2_23 ;
 wire [7:0] u_multiplier_pp2_24 ;
 wire [7:0] u_multiplier_pp2_25 ;
 wire [7:0] u_multiplier_pp2_26 ;
 wire [7:0] u_multiplier_pp2_27 ;
 wire [7:0] u_multiplier_pp2_28 ;
 wire [7:0] u_multiplier_pp2_29 ;
 wire [3:0] u_multiplier_pp2_3 ;
 wire [7:0] u_multiplier_pp2_30 ;
 wire [7:0] u_multiplier_pp2_31 ;
 wire [7:0] u_multiplier_pp2_32 ;
 wire [7:0] u_multiplier_pp2_33 ;
 wire [7:0] u_multiplier_pp2_34 ;
 wire [7:0] u_multiplier_pp2_35 ;
 wire [7:0] u_multiplier_pp2_36 ;
 wire [7:0] u_multiplier_pp2_37 ;
 wire [7:0] u_multiplier_pp2_38 ;
 wire [7:0] u_multiplier_pp2_39 ;
 wire [4:0] u_multiplier_pp2_4 ;
 wire [7:0] u_multiplier_pp2_40 ;
 wire [7:0] u_multiplier_pp2_41 ;
 wire [7:0] u_multiplier_pp2_42 ;
 wire [7:0] u_multiplier_pp2_43 ;
 wire [7:0] u_multiplier_pp2_44 ;
 wire [7:0] u_multiplier_pp2_45 ;
 wire [7:0] u_multiplier_pp2_46 ;
 wire [7:0] u_multiplier_pp2_47 ;
 wire [7:0] u_multiplier_pp2_48 ;
 wire [7:0] u_multiplier_pp2_49 ;
 wire [5:0] u_multiplier_pp2_5 ;
 wire [7:0] u_multiplier_pp2_50 ;
 wire [7:0] u_multiplier_pp2_51 ;
 wire [7:0] u_multiplier_pp2_52 ;
 wire [7:0] u_multiplier_pp2_53 ;
 wire [7:0] u_multiplier_pp2_54 ;
 wire [7:0] u_multiplier_pp2_55 ;
 wire [7:0] u_multiplier_pp2_56 ;
 wire [5:0] u_multiplier_pp2_57 ;
 wire [4:0] u_multiplier_pp2_58 ;
 wire [3:0] u_multiplier_pp2_59 ;
 wire [6:0] u_multiplier_pp2_6 ;
 wire [2:0] u_multiplier_pp2_60 ;
 wire [1:0] u_multiplier_pp2_61 ;
 wire [7:0] u_multiplier_pp2_7 ;
 wire [7:0] u_multiplier_pp2_8 ;
 wire [7:0] u_multiplier_pp2_9 ;
 wire [1:0] u_multiplier_pp3_1 ;
 wire [3:0] u_multiplier_pp3_10 ;
 wire [3:0] u_multiplier_pp3_11 ;
 wire [3:0] u_multiplier_pp3_12 ;
 wire [3:0] u_multiplier_pp3_13 ;
 wire [3:0] u_multiplier_pp3_14 ;
 wire [3:0] u_multiplier_pp3_15 ;
 wire [3:0] u_multiplier_pp3_16 ;
 wire [3:0] u_multiplier_pp3_17 ;
 wire [3:0] u_multiplier_pp3_18 ;
 wire [3:0] u_multiplier_pp3_19 ;
 wire [2:0] u_multiplier_pp3_2 ;
 wire [3:0] u_multiplier_pp3_20 ;
 wire [3:0] u_multiplier_pp3_21 ;
 wire [3:0] u_multiplier_pp3_22 ;
 wire [3:0] u_multiplier_pp3_23 ;
 wire [3:0] u_multiplier_pp3_24 ;
 wire [3:0] u_multiplier_pp3_25 ;
 wire [3:0] u_multiplier_pp3_26 ;
 wire [3:0] u_multiplier_pp3_27 ;
 wire [3:0] u_multiplier_pp3_28 ;
 wire [3:0] u_multiplier_pp3_29 ;
 wire [3:0] u_multiplier_pp3_3 ;
 wire [3:0] u_multiplier_pp3_30 ;
 wire [3:0] u_multiplier_pp3_31 ;
 wire [3:0] u_multiplier_pp3_32 ;
 wire [3:0] u_multiplier_pp3_33 ;
 wire [3:0] u_multiplier_pp3_34 ;
 wire [3:0] u_multiplier_pp3_35 ;
 wire [3:0] u_multiplier_pp3_36 ;
 wire [3:0] u_multiplier_pp3_37 ;
 wire [3:0] u_multiplier_pp3_38 ;
 wire [3:0] u_multiplier_pp3_39 ;
 wire [3:0] u_multiplier_pp3_4 ;
 wire [3:0] u_multiplier_pp3_40 ;
 wire [3:0] u_multiplier_pp3_41 ;
 wire [3:0] u_multiplier_pp3_42 ;
 wire [3:0] u_multiplier_pp3_43 ;
 wire [3:0] u_multiplier_pp3_44 ;
 wire [3:0] u_multiplier_pp3_45 ;
 wire [3:0] u_multiplier_pp3_46 ;
 wire [3:0] u_multiplier_pp3_47 ;
 wire [3:0] u_multiplier_pp3_48 ;
 wire [3:0] u_multiplier_pp3_49 ;
 wire [3:0] u_multiplier_pp3_5 ;
 wire [3:0] u_multiplier_pp3_50 ;
 wire [3:0] u_multiplier_pp3_51 ;
 wire [3:0] u_multiplier_pp3_52 ;
 wire [3:0] u_multiplier_pp3_53 ;
 wire [3:0] u_multiplier_pp3_54 ;
 wire [3:0] u_multiplier_pp3_55 ;
 wire [3:0] u_multiplier_pp3_56 ;
 wire [3:0] u_multiplier_pp3_57 ;
 wire [3:0] u_multiplier_pp3_58 ;
 wire [3:0] u_multiplier_pp3_59 ;
 wire [3:0] u_multiplier_pp3_6 ;
 wire [3:0] u_multiplier_pp3_60 ;
 wire [1:0] u_multiplier_pp3_61 ;
 wire [3:0] u_multiplier_pp3_7 ;
 wire [3:0] u_multiplier_pp3_8 ;
 wire [3:0] u_multiplier_pp3_9 ;

 INV_X2 _0675_ (.A(net12),
    .ZN(_0370_));
 INV_X2 _0676_ (.A(net46),
    .ZN(_0307_));
 INV_X1 _0677_ (.A(init_count[5]),
    .ZN(_0371_));
 INV_X1 _0678_ (.A(curr_state[2]),
    .ZN(_0372_));
 INV_X1 _0679_ (.A(net48),
    .ZN(_0373_));
 INV_X1 _0680_ (.A(net180),
    .ZN(_0374_));
 NOR2_X4 _0681_ (.A1(_0370_),
    .A2(_0373_),
    .ZN(_0303_));
 NAND2_X2 _0682_ (.A1(net12),
    .A2(net220),
    .ZN(_0308_));
 NAND2_X1 _0683_ (.A1(init_count[1]),
    .A2(init_count[0]),
    .ZN(_0375_));
 AND4_X2 _0684_ (.A1(init_count[1]),
    .A2(init_count[0]),
    .A3(init_count[3]),
    .A4(init_count[2]),
    .ZN(_0376_));
 INV_X1 _0685_ (.A(_0376_),
    .ZN(_0377_));
 AND2_X1 _0686_ (.A1(init_count[5]),
    .A2(init_count[4]),
    .ZN(_0378_));
 AND3_X1 _0687_ (.A1(net46),
    .A2(_0376_),
    .A3(_0378_),
    .ZN(_0379_));
 NOR2_X2 _0688_ (.A1(_0370_),
    .A2(_0307_),
    .ZN(_0380_));
 NAND2_X2 _0689_ (.A1(net12),
    .A2(net46),
    .ZN(_0381_));
 AND3_X1 _0690_ (.A1(curr_state[2]),
    .A2(_0376_),
    .A3(_0378_),
    .ZN(_0382_));
 NAND2_X1 _0691_ (.A1(_0380_),
    .A2(_0382_),
    .ZN(_0383_));
 OAI21_X1 _0692_ (.A(_0383_),
    .B1(_0373_),
    .B2(_0370_),
    .ZN(_0305_));
 NAND3_X1 _0693_ (.A1(net45),
    .A2(net200),
    .A3(_0380_),
    .ZN(_0384_));
 OAI21_X1 _0694_ (.A(net201),
    .B1(_0379_),
    .B2(_0308_),
    .ZN(_0306_));
 AOI22_X1 _0695_ (.A1(net12),
    .A2(net163),
    .B1(_0380_),
    .B2(net45),
    .ZN(_0304_));
 AND2_X1 _0696_ (.A1(net11),
    .A2(sram_rdata[0]),
    .ZN(_0271_));
 AND2_X1 _0697_ (.A1(net11),
    .A2(sram_rdata[1]),
    .ZN(_0282_));
 AND2_X1 _0698_ (.A1(net11),
    .A2(sram_rdata[2]),
    .ZN(_0293_));
 AND2_X1 _0699_ (.A1(net11),
    .A2(sram_rdata[3]),
    .ZN(_0296_));
 AND2_X1 _0700_ (.A1(net11),
    .A2(sram_rdata[4]),
    .ZN(_0297_));
 AND2_X1 _0701_ (.A1(net11),
    .A2(sram_rdata[5]),
    .ZN(_0298_));
 AND2_X1 _0702_ (.A1(net11),
    .A2(sram_rdata[6]),
    .ZN(_0299_));
 AND2_X1 _0703_ (.A1(net11),
    .A2(sram_rdata[7]),
    .ZN(_0300_));
 AND2_X1 _0704_ (.A1(net11),
    .A2(sram_rdata[8]),
    .ZN(_0301_));
 AND2_X1 _0705_ (.A1(net11),
    .A2(sram_rdata[9]),
    .ZN(_0302_));
 AND2_X1 _0706_ (.A1(net11),
    .A2(sram_rdata[10]),
    .ZN(_0272_));
 AND2_X1 _0707_ (.A1(net11),
    .A2(sram_rdata[11]),
    .ZN(_0273_));
 AND2_X1 _0708_ (.A1(net11),
    .A2(sram_rdata[12]),
    .ZN(_0274_));
 AND2_X1 _0709_ (.A1(net11),
    .A2(sram_rdata[13]),
    .ZN(_0275_));
 AND2_X1 _0710_ (.A1(net11),
    .A2(sram_rdata[14]),
    .ZN(_0276_));
 AND2_X1 _0711_ (.A1(net11),
    .A2(sram_rdata[15]),
    .ZN(_0277_));
 AND2_X1 _0712_ (.A1(net11),
    .A2(sram_rdata[16]),
    .ZN(_0278_));
 AND2_X1 _0713_ (.A1(net11),
    .A2(sram_rdata[17]),
    .ZN(_0279_));
 AND2_X1 _0714_ (.A1(net11),
    .A2(sram_rdata[18]),
    .ZN(_0280_));
 AND2_X1 _0715_ (.A1(net11),
    .A2(sram_rdata[19]),
    .ZN(_0281_));
 AND2_X1 _0716_ (.A1(net11),
    .A2(sram_rdata[20]),
    .ZN(_0283_));
 AND2_X1 _0717_ (.A1(net11),
    .A2(sram_rdata[21]),
    .ZN(_0284_));
 AND2_X1 _0718_ (.A1(net11),
    .A2(sram_rdata[22]),
    .ZN(_0285_));
 AND2_X1 _0719_ (.A1(net11),
    .A2(sram_rdata[23]),
    .ZN(_0286_));
 AND2_X1 _0720_ (.A1(net11),
    .A2(sram_rdata[24]),
    .ZN(_0287_));
 AND2_X1 _0721_ (.A1(net11),
    .A2(sram_rdata[25]),
    .ZN(_0288_));
 AND2_X1 _0722_ (.A1(net11),
    .A2(sram_rdata[26]),
    .ZN(_0289_));
 AND2_X1 _0723_ (.A1(net11),
    .A2(sram_rdata[27]),
    .ZN(_0290_));
 AND2_X1 _0724_ (.A1(net11),
    .A2(sram_rdata[28]),
    .ZN(_0291_));
 AND2_X1 _0725_ (.A1(net11),
    .A2(sram_rdata[29]),
    .ZN(_0292_));
 AND2_X1 _0726_ (.A1(net11),
    .A2(sram_rdata[30]),
    .ZN(_0294_));
 AND2_X1 _0727_ (.A1(net11),
    .A2(sram_rdata[31]),
    .ZN(_0295_));
 AND2_X1 _0728_ (.A1(product[0]),
    .A2(net9),
    .ZN(_0201_));
 AND2_X1 _0729_ (.A1(product[1]),
    .A2(net9),
    .ZN(_0212_));
 AND2_X1 _0730_ (.A1(product[2]),
    .A2(net9),
    .ZN(_0223_));
 AND2_X1 _0731_ (.A1(product[3]),
    .A2(net9),
    .ZN(_0234_));
 AND2_X1 _0732_ (.A1(product[4]),
    .A2(_0303_),
    .ZN(_0245_));
 AND2_X1 _0733_ (.A1(product[5]),
    .A2(net9),
    .ZN(_0256_));
 AND2_X1 _0734_ (.A1(product[6]),
    .A2(net10),
    .ZN(_0261_));
 AND2_X1 _0735_ (.A1(product[7]),
    .A2(net10),
    .ZN(_0262_));
 AND2_X1 _0736_ (.A1(product[8]),
    .A2(_0303_),
    .ZN(_0263_));
 AND2_X1 _0737_ (.A1(product[9]),
    .A2(net10),
    .ZN(_0264_));
 AND2_X1 _0738_ (.A1(product[10]),
    .A2(net9),
    .ZN(_0202_));
 AND2_X1 _0739_ (.A1(product[11]),
    .A2(net10),
    .ZN(_0203_));
 AND2_X1 _0740_ (.A1(product[12]),
    .A2(net9),
    .ZN(_0204_));
 AND2_X1 _0741_ (.A1(product[13]),
    .A2(net9),
    .ZN(_0205_));
 AND2_X1 _0742_ (.A1(product[14]),
    .A2(net9),
    .ZN(_0206_));
 AND2_X1 _0743_ (.A1(product[15]),
    .A2(net9),
    .ZN(_0207_));
 AND2_X1 _0744_ (.A1(product[16]),
    .A2(net9),
    .ZN(_0208_));
 AND2_X1 _0745_ (.A1(product[17]),
    .A2(net9),
    .ZN(_0209_));
 AND2_X1 _0746_ (.A1(product[18]),
    .A2(net10),
    .ZN(_0210_));
 AND2_X1 _0747_ (.A1(product[19]),
    .A2(_0303_),
    .ZN(_0211_));
 AND2_X1 _0748_ (.A1(product[20]),
    .A2(net9),
    .ZN(_0213_));
 AND2_X1 _0749_ (.A1(product[21]),
    .A2(net9),
    .ZN(_0214_));
 AND2_X1 _0750_ (.A1(product[22]),
    .A2(_0303_),
    .ZN(_0215_));
 AND2_X1 _0751_ (.A1(product[23]),
    .A2(net10),
    .ZN(_0216_));
 AND2_X1 _0752_ (.A1(product[24]),
    .A2(net9),
    .ZN(_0217_));
 AND2_X1 _0753_ (.A1(product[25]),
    .A2(_0303_),
    .ZN(_0218_));
 AND2_X1 _0754_ (.A1(product[26]),
    .A2(_0303_),
    .ZN(_0219_));
 AND2_X1 _0755_ (.A1(product[27]),
    .A2(_0303_),
    .ZN(_0220_));
 AND2_X1 _0756_ (.A1(product[28]),
    .A2(_0303_),
    .ZN(_0221_));
 AND2_X1 _0757_ (.A1(product[29]),
    .A2(net9),
    .ZN(_0222_));
 AND2_X1 _0758_ (.A1(product[30]),
    .A2(_0303_),
    .ZN(_0224_));
 AND2_X1 _0759_ (.A1(product[31]),
    .A2(net10),
    .ZN(_0225_));
 AND2_X1 _0760_ (.A1(product[32]),
    .A2(net9),
    .ZN(_0226_));
 AND2_X1 _0761_ (.A1(product[33]),
    .A2(net9),
    .ZN(_0227_));
 AND2_X1 _0762_ (.A1(product[34]),
    .A2(net9),
    .ZN(_0228_));
 AND2_X1 _0763_ (.A1(product[35]),
    .A2(net9),
    .ZN(_0229_));
 AND2_X1 _0764_ (.A1(product[36]),
    .A2(_0303_),
    .ZN(_0230_));
 AND2_X1 _0765_ (.A1(product[37]),
    .A2(_0303_),
    .ZN(_0231_));
 AND2_X1 _0766_ (.A1(product[38]),
    .A2(net9),
    .ZN(_0232_));
 AND2_X1 _0767_ (.A1(product[39]),
    .A2(net10),
    .ZN(_0233_));
 AND2_X1 _0768_ (.A1(product[40]),
    .A2(net9),
    .ZN(_0235_));
 AND2_X1 _0769_ (.A1(product[41]),
    .A2(net9),
    .ZN(_0236_));
 AND2_X1 _0770_ (.A1(product[42]),
    .A2(net9),
    .ZN(_0237_));
 AND2_X1 _0771_ (.A1(product[43]),
    .A2(net10),
    .ZN(_0238_));
 AND2_X1 _0772_ (.A1(product[44]),
    .A2(_0303_),
    .ZN(_0239_));
 AND2_X1 _0773_ (.A1(product[45]),
    .A2(net9),
    .ZN(_0240_));
 AND2_X1 _0774_ (.A1(product[46]),
    .A2(_0303_),
    .ZN(_0241_));
 AND2_X1 _0775_ (.A1(product[47]),
    .A2(_0303_),
    .ZN(_0242_));
 AND2_X1 _0776_ (.A1(product[48]),
    .A2(_0303_),
    .ZN(_0243_));
 AND2_X1 _0777_ (.A1(product[49]),
    .A2(net10),
    .ZN(_0244_));
 AND2_X1 _0778_ (.A1(product[50]),
    .A2(_0303_),
    .ZN(_0246_));
 AND2_X1 _0779_ (.A1(product[51]),
    .A2(_0303_),
    .ZN(_0247_));
 AND2_X1 _0780_ (.A1(product[52]),
    .A2(_0303_),
    .ZN(_0248_));
 AND2_X1 _0781_ (.A1(product[53]),
    .A2(net9),
    .ZN(_0249_));
 AND2_X1 _0782_ (.A1(product[54]),
    .A2(net10),
    .ZN(_0250_));
 AND2_X1 _0783_ (.A1(product[55]),
    .A2(net9),
    .ZN(_0251_));
 AND2_X1 _0784_ (.A1(product[56]),
    .A2(net9),
    .ZN(_0252_));
 AND2_X1 _0785_ (.A1(product[57]),
    .A2(net9),
    .ZN(_0253_));
 AND2_X1 _0786_ (.A1(product[58]),
    .A2(net10),
    .ZN(_0254_));
 AND2_X1 _0787_ (.A1(product[59]),
    .A2(net9),
    .ZN(_0255_));
 AND2_X1 _0788_ (.A1(product[60]),
    .A2(net9),
    .ZN(_0257_));
 AND2_X1 _0789_ (.A1(product[61]),
    .A2(_0303_),
    .ZN(_0258_));
 AND2_X1 _0790_ (.A1(product[62]),
    .A2(net9),
    .ZN(_0259_));
 AND2_X1 _0791_ (.A1(product[63]),
    .A2(net9),
    .ZN(_0260_));
 AND2_X1 _0792_ (.A1(net11),
    .A2(net13),
    .ZN(_0169_));
 AND2_X1 _0793_ (.A1(net12),
    .A2(net24),
    .ZN(_0180_));
 AND2_X1 _0794_ (.A1(net12),
    .A2(net35),
    .ZN(_0191_));
 AND2_X1 _0795_ (.A1(net11),
    .A2(net38),
    .ZN(_0194_));
 AND2_X1 _0796_ (.A1(net11),
    .A2(net39),
    .ZN(_0195_));
 AND2_X1 _0797_ (.A1(net11),
    .A2(net40),
    .ZN(_0196_));
 AND2_X1 _0798_ (.A1(net12),
    .A2(net41),
    .ZN(_0197_));
 AND2_X1 _0799_ (.A1(net12),
    .A2(net42),
    .ZN(_0198_));
 AND2_X1 _0800_ (.A1(net11),
    .A2(net43),
    .ZN(_0199_));
 AND2_X1 _0801_ (.A1(net11),
    .A2(net44),
    .ZN(_0200_));
 AND2_X1 _0802_ (.A1(net11),
    .A2(net14),
    .ZN(_0170_));
 AND2_X1 _0803_ (.A1(net12),
    .A2(net15),
    .ZN(_0171_));
 AND2_X1 _0804_ (.A1(net12),
    .A2(net16),
    .ZN(_0172_));
 AND2_X1 _0805_ (.A1(net47),
    .A2(net17),
    .ZN(_0173_));
 AND2_X1 _0806_ (.A1(net11),
    .A2(net18),
    .ZN(_0174_));
 AND2_X1 _0807_ (.A1(net12),
    .A2(net19),
    .ZN(_0175_));
 AND2_X1 _0808_ (.A1(net12),
    .A2(net20),
    .ZN(_0176_));
 AND2_X1 _0809_ (.A1(net47),
    .A2(net21),
    .ZN(_0177_));
 AND2_X1 _0810_ (.A1(net12),
    .A2(net22),
    .ZN(_0178_));
 AND2_X1 _0811_ (.A1(net12),
    .A2(net23),
    .ZN(_0179_));
 AND2_X1 _0812_ (.A1(net12),
    .A2(net25),
    .ZN(_0181_));
 AND2_X1 _0813_ (.A1(net12),
    .A2(net26),
    .ZN(_0182_));
 AND2_X1 _0814_ (.A1(net11),
    .A2(net27),
    .ZN(_0183_));
 AND2_X1 _0815_ (.A1(net11),
    .A2(net28),
    .ZN(_0184_));
 AND2_X1 _0816_ (.A1(net12),
    .A2(net29),
    .ZN(_0185_));
 AND2_X1 _0817_ (.A1(net12),
    .A2(net30),
    .ZN(_0186_));
 AND2_X1 _0818_ (.A1(net47),
    .A2(net31),
    .ZN(_0187_));
 AND2_X1 _0819_ (.A1(net12),
    .A2(net32),
    .ZN(_0188_));
 AND2_X1 _0820_ (.A1(net12),
    .A2(net33),
    .ZN(_0189_));
 AND2_X1 _0821_ (.A1(net12),
    .A2(net34),
    .ZN(_0190_));
 AND2_X1 _0822_ (.A1(net12),
    .A2(net36),
    .ZN(_0192_));
 AND2_X1 _0823_ (.A1(net11),
    .A2(net37),
    .ZN(_0193_));
 NAND2_X2 _0824_ (.A1(net12),
    .A2(_0307_),
    .ZN(_0385_));
 OAI21_X1 _0825_ (.A(net12),
    .B1(_0307_),
    .B2(_0382_),
    .ZN(_0386_));
 AOI21_X4 _0826_ (.A(_0372_),
    .B1(_0376_),
    .B2(_0378_),
    .ZN(_0387_));
 AOI22_X1 _0827_ (.A1(init_count[0]),
    .A2(net48),
    .B1(net184),
    .B2(_0387_),
    .ZN(_0388_));
 OAI22_X1 _0828_ (.A1(net185),
    .A2(_0386_),
    .B1(_0388_),
    .B2(_0381_),
    .ZN(_0265_));
 AOI21_X1 _0829_ (.A(net48),
    .B1(_0375_),
    .B2(curr_state[2]),
    .ZN(_0389_));
 INV_X1 _0830_ (.A(_0389_),
    .ZN(_0390_));
 AOI21_X1 _0831_ (.A(init_count[1]),
    .B1(init_count[0]),
    .B2(curr_state[2]),
    .ZN(_0391_));
 OR3_X1 _0832_ (.A1(_0381_),
    .A2(_0389_),
    .A3(_0391_),
    .ZN(_0392_));
 OAI211_X1 _0833_ (.A(_0383_),
    .B(_0392_),
    .C1(_0385_),
    .C2(net199),
    .ZN(_0266_));
 NOR3_X1 _0834_ (.A1(init_count[2]),
    .A2(_0372_),
    .A3(_0375_),
    .ZN(_0393_));
 AOI211_X1 _0835_ (.A(_0382_),
    .B(_0393_),
    .C1(_0390_),
    .C2(init_count[2]),
    .ZN(_0394_));
 OAI22_X1 _0836_ (.A1(net193),
    .A2(_0385_),
    .B1(_0394_),
    .B2(_0381_),
    .ZN(_0267_));
 NOR2_X1 _0837_ (.A1(_0658_),
    .A2(_0375_),
    .ZN(_0395_));
 XOR2_X2 _0838_ (.A(init_count[3]),
    .B(_0395_),
    .Z(_0396_));
 AOI221_X2 _0839_ (.A(_0382_),
    .B1(_0396_),
    .B2(curr_state[2]),
    .C1(net48),
    .C2(init_count[3]),
    .ZN(_0397_));
 OAI22_X1 _0840_ (.A1(net204),
    .A2(_0385_),
    .B1(_0397_),
    .B2(_0381_),
    .ZN(_0268_));
 NAND3_X1 _0841_ (.A1(_0371_),
    .A2(init_count[4]),
    .A3(_0376_),
    .ZN(_0398_));
 OAI21_X1 _0842_ (.A(curr_state[2]),
    .B1(_0376_),
    .B2(init_count[4]),
    .ZN(_0399_));
 INV_X1 _0843_ (.A(_0399_),
    .ZN(_0400_));
 AOI22_X1 _0844_ (.A1(net234),
    .A2(net48),
    .B1(_0398_),
    .B2(_0400_),
    .ZN(_0401_));
 OAI22_X1 _0845_ (.A1(net196),
    .A2(_0385_),
    .B1(_0401_),
    .B2(_0381_),
    .ZN(_0269_));
 OAI21_X1 _0846_ (.A(net189),
    .B1(_0377_),
    .B2(_0660_),
    .ZN(_0402_));
 AOI22_X1 _0847_ (.A1(net233),
    .A2(net48),
    .B1(_0402_),
    .B2(curr_state[2]),
    .ZN(_0403_));
 OAI22_X1 _0848_ (.A1(net190),
    .A2(_0385_),
    .B1(_0403_),
    .B2(_0381_),
    .ZN(_0270_));
 NOR2_X1 _0849_ (.A1(_0373_),
    .A2(addr_ptr[0]),
    .ZN(_0404_));
 AOI21_X1 _0850_ (.A(_0404_),
    .B1(_0387_),
    .B2(net208),
    .ZN(_0405_));
 OAI22_X1 _0851_ (.A1(net176),
    .A2(_0385_),
    .B1(net209),
    .B2(_0381_),
    .ZN(_0163_));
 NAND2_X1 _0852_ (.A1(addr_ptr[0]),
    .A2(addr_ptr[1]),
    .ZN(_0406_));
 XOR2_X1 _0853_ (.A(addr_ptr[0]),
    .B(addr_ptr[1]),
    .Z(_0407_));
 OAI211_X1 _0854_ (.A(_0380_),
    .B(_0407_),
    .C1(_0387_),
    .C2(net48),
    .ZN(_0408_));
 OAI21_X1 _0855_ (.A(_0408_),
    .B1(_0385_),
    .B2(net2),
    .ZN(_0164_));
 AND4_X1 _0856_ (.A1(addr_ptr[0]),
    .A2(addr_ptr[1]),
    .A3(addr_ptr[3]),
    .A4(addr_ptr[2]),
    .ZN(_0409_));
 NAND3_X1 _0857_ (.A1(net187),
    .A2(net182),
    .A3(_0409_),
    .ZN(_0410_));
 AOI21_X2 _0858_ (.A(_0387_),
    .B1(_0410_),
    .B2(net48),
    .ZN(_0411_));
 AOI21_X1 _0859_ (.A(_0381_),
    .B1(_0406_),
    .B2(net213),
    .ZN(_0412_));
 OAI21_X1 _0860_ (.A(_0412_),
    .B1(_0406_),
    .B2(net213),
    .ZN(_0413_));
 OAI22_X1 _0861_ (.A1(net214),
    .A2(_0385_),
    .B1(_0411_),
    .B2(_0413_),
    .ZN(_0165_));
 NOR3_X1 _0862_ (.A1(_0307_),
    .A2(net213),
    .A3(_0406_),
    .ZN(_0414_));
 OAI21_X1 _0863_ (.A(net12),
    .B1(_0374_),
    .B2(_0414_),
    .ZN(_0415_));
 AOI221_X1 _0864_ (.A(_0415_),
    .B1(_0414_),
    .B2(_0374_),
    .C1(net46),
    .C2(_0411_),
    .ZN(_0166_));
 NAND2_X1 _0865_ (.A1(net46),
    .A2(_0409_),
    .ZN(_0416_));
 OR2_X1 _0866_ (.A1(_0654_),
    .A2(_0416_),
    .ZN(_0417_));
 XNOR2_X1 _0867_ (.A(net206),
    .B(_0416_),
    .ZN(_0418_));
 AOI211_X1 _0868_ (.A(_0370_),
    .B(net207),
    .C1(_0411_),
    .C2(net46),
    .ZN(_0167_));
 XNOR2_X1 _0869_ (.A(net7),
    .B(_0417_),
    .ZN(_0419_));
 AOI211_X1 _0870_ (.A(_0370_),
    .B(net8),
    .C1(_0411_),
    .C2(net46),
    .ZN(_0168_));
 DFF_X1 _0871_ (.D(net164),
    .CK(clknet_4_7__leaf_clk),
    .Q(curr_state[0]),
    .QN(_0518_));
 DFF_X2 _0872_ (.D(_0305_),
    .CK(clknet_4_7__leaf_clk),
    .Q(net48),
    .QN(_0519_));
 DFF_X2 _0873_ (.D(net202),
    .CK(clknet_4_6__leaf_clk),
    .Q(curr_state[2]),
    .QN(_0520_));
 DFF_X2 _0874_ (.D(_0201_),
    .CK(clknet_4_9__leaf_clk),
    .Q(net49),
    .QN(_0521_));
 DFF_X2 _0875_ (.D(_0212_),
    .CK(clknet_4_9__leaf_clk),
    .Q(net60),
    .QN(_0522_));
 DFF_X2 _0876_ (.D(_0223_),
    .CK(clknet_4_9__leaf_clk),
    .Q(net71),
    .QN(_0523_));
 DFF_X2 _0877_ (.D(_0234_),
    .CK(clknet_4_9__leaf_clk),
    .Q(net82),
    .QN(_0524_));
 DFF_X1 _0878_ (.D(_0245_),
    .CK(clknet_4_3__leaf_clk),
    .Q(net93),
    .QN(_0525_));
 DFF_X2 _0879_ (.D(_0256_),
    .CK(clknet_4_9__leaf_clk),
    .Q(net104),
    .QN(_0526_));
 DFF_X2 _0880_ (.D(_0261_),
    .CK(clknet_4_15__leaf_clk),
    .Q(net109),
    .QN(_0527_));
 DFF_X2 _0881_ (.D(_0262_),
    .CK(clknet_4_15__leaf_clk),
    .Q(net110),
    .QN(_0528_));
 DFF_X2 _0882_ (.D(_0263_),
    .CK(clknet_4_12__leaf_clk),
    .Q(net111),
    .QN(_0529_));
 DFF_X2 _0883_ (.D(_0264_),
    .CK(clknet_4_14__leaf_clk),
    .Q(net112),
    .QN(_0530_));
 DFF_X2 _0884_ (.D(_0202_),
    .CK(clknet_4_14__leaf_clk),
    .Q(net50),
    .QN(_0531_));
 DFF_X2 _0885_ (.D(_0203_),
    .CK(clknet_4_14__leaf_clk),
    .Q(net51),
    .QN(_0532_));
 DFF_X2 _0886_ (.D(_0204_),
    .CK(clknet_4_14__leaf_clk),
    .Q(net52),
    .QN(_0533_));
 DFF_X2 _0887_ (.D(_0205_),
    .CK(clknet_4_14__leaf_clk),
    .Q(net53),
    .QN(_0534_));
 DFF_X1 _0888_ (.D(_0206_),
    .CK(clknet_4_12__leaf_clk),
    .Q(net54),
    .QN(_0535_));
 DFF_X2 _0889_ (.D(_0207_),
    .CK(clknet_4_14__leaf_clk),
    .Q(net55),
    .QN(_0536_));
 DFF_X2 _0890_ (.D(_0208_),
    .CK(clknet_4_2__leaf_clk),
    .Q(net56),
    .QN(_0537_));
 DFF_X2 _0891_ (.D(_0209_),
    .CK(clknet_4_10__leaf_clk),
    .Q(net57),
    .QN(_0538_));
 DFF_X2 _0892_ (.D(_0210_),
    .CK(clknet_4_1__leaf_clk),
    .Q(net58),
    .QN(_0539_));
 DFF_X2 _0893_ (.D(_0211_),
    .CK(clknet_4_4__leaf_clk),
    .Q(net59),
    .QN(_0540_));
 DFF_X2 _0894_ (.D(_0213_),
    .CK(clknet_4_11__leaf_clk),
    .Q(net61),
    .QN(_0541_));
 DFF_X2 _0895_ (.D(_0214_),
    .CK(clknet_4_11__leaf_clk),
    .Q(net62),
    .QN(_0542_));
 DFF_X2 _0896_ (.D(_0215_),
    .CK(clknet_4_6__leaf_clk),
    .Q(net63),
    .QN(_0543_));
 DFF_X1 _0897_ (.D(_0216_),
    .CK(clknet_4_4__leaf_clk),
    .Q(net64),
    .QN(_0544_));
 DFF_X2 _0898_ (.D(_0217_),
    .CK(clknet_4_11__leaf_clk),
    .Q(net65),
    .QN(_0545_));
 DFF_X1 _0899_ (.D(_0218_),
    .CK(clknet_4_5__leaf_clk),
    .Q(net66),
    .QN(_0546_));
 DFF_X2 _0900_ (.D(_0219_),
    .CK(clknet_4_5__leaf_clk),
    .Q(net67),
    .QN(_0547_));
 DFF_X2 _0901_ (.D(_0220_),
    .CK(clknet_4_5__leaf_clk),
    .Q(net68),
    .QN(_0548_));
 DFF_X2 _0902_ (.D(_0221_),
    .CK(clknet_4_4__leaf_clk),
    .Q(net69),
    .QN(_0549_));
 DFF_X2 _0903_ (.D(_0222_),
    .CK(clknet_4_9__leaf_clk),
    .Q(net70),
    .QN(_0550_));
 DFF_X1 _0904_ (.D(_0224_),
    .CK(clknet_4_1__leaf_clk),
    .Q(net72),
    .QN(_0551_));
 DFF_X2 _0905_ (.D(_0225_),
    .CK(clknet_4_1__leaf_clk),
    .Q(net73),
    .QN(_0552_));
 DFF_X1 _0906_ (.D(_0226_),
    .CK(clknet_4_3__leaf_clk),
    .Q(net74),
    .QN(_0553_));
 DFF_X2 _0907_ (.D(_0227_),
    .CK(clknet_4_12__leaf_clk),
    .Q(net75),
    .QN(_0554_));
 DFF_X2 _0908_ (.D(_0228_),
    .CK(clknet_4_8__leaf_clk),
    .Q(net76),
    .QN(_0555_));
 DFF_X2 _0909_ (.D(_0229_),
    .CK(clknet_4_8__leaf_clk),
    .Q(net77),
    .QN(_0556_));
 DFF_X2 _0910_ (.D(_0230_),
    .CK(clknet_4_12__leaf_clk),
    .Q(net78),
    .QN(_0557_));
 DFF_X2 _0911_ (.D(_0231_),
    .CK(clknet_4_12__leaf_clk),
    .Q(net79),
    .QN(_0558_));
 DFF_X2 _0912_ (.D(_0232_),
    .CK(clknet_4_8__leaf_clk),
    .Q(net80),
    .QN(_0559_));
 DFF_X2 _0913_ (.D(_0233_),
    .CK(clknet_4_10__leaf_clk),
    .Q(net81),
    .QN(_0560_));
 DFF_X2 _0914_ (.D(_0235_),
    .CK(clknet_4_8__leaf_clk),
    .Q(net83),
    .QN(_0561_));
 DFF_X2 _0915_ (.D(_0236_),
    .CK(clknet_4_8__leaf_clk),
    .Q(net84),
    .QN(_0562_));
 DFF_X2 _0916_ (.D(_0237_),
    .CK(clknet_4_8__leaf_clk),
    .Q(net85),
    .QN(_0563_));
 DFF_X2 _0917_ (.D(_0238_),
    .CK(clknet_4_2__leaf_clk),
    .Q(net86),
    .QN(_0564_));
 DFF_X2 _0918_ (.D(_0239_),
    .CK(clknet_4_2__leaf_clk),
    .Q(net87),
    .QN(_0565_));
 DFF_X2 _0919_ (.D(_0240_),
    .CK(clknet_4_2__leaf_clk),
    .Q(net88),
    .QN(_0566_));
 DFF_X1 _0920_ (.D(_0241_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net89),
    .QN(_0567_));
 DFF_X2 _0921_ (.D(_0242_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net90),
    .QN(_0568_));
 DFF_X2 _0922_ (.D(_0243_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net91),
    .QN(_0569_));
 DFF_X2 _0923_ (.D(_0244_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net92),
    .QN(_0570_));
 DFF_X2 _0924_ (.D(_0246_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net94),
    .QN(_0571_));
 DFF_X1 _0925_ (.D(_0247_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net95),
    .QN(_0572_));
 DFF_X1 _0926_ (.D(_0248_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net96),
    .QN(_0573_));
 DFF_X2 _0927_ (.D(_0249_),
    .CK(clknet_4_2__leaf_clk),
    .Q(net97),
    .QN(_0574_));
 DFF_X2 _0928_ (.D(_0250_),
    .CK(clknet_4_12__leaf_clk),
    .Q(net98),
    .QN(_0575_));
 DFF_X1 _0929_ (.D(_0251_),
    .CK(clknet_4_14__leaf_clk),
    .Q(net99),
    .QN(_0576_));
 DFF_X2 _0930_ (.D(_0252_),
    .CK(clknet_4_10__leaf_clk),
    .Q(net100),
    .QN(_0577_));
 DFF_X1 _0931_ (.D(_0253_),
    .CK(clknet_4_10__leaf_clk),
    .Q(net101),
    .QN(_0578_));
 DFF_X2 _0932_ (.D(_0254_),
    .CK(clknet_4_10__leaf_clk),
    .Q(net102),
    .QN(_0579_));
 DFF_X2 _0933_ (.D(_0255_),
    .CK(clknet_4_11__leaf_clk),
    .Q(net103),
    .QN(_0580_));
 DFF_X2 _0934_ (.D(_0257_),
    .CK(clknet_4_11__leaf_clk),
    .Q(net105),
    .QN(_0581_));
 DFF_X2 _0935_ (.D(_0258_),
    .CK(clknet_4_15__leaf_clk),
    .Q(net106),
    .QN(_0582_));
 DFF_X2 _0936_ (.D(_0259_),
    .CK(clknet_4_11__leaf_clk),
    .Q(net107),
    .QN(_0583_));
 DFF_X1 _0937_ (.D(_0260_),
    .CK(clknet_4_9__leaf_clk),
    .Q(net108),
    .QN(_0584_));
 DFF_X2 _0938_ (.D(_0169_),
    .CK(clknet_4_14__leaf_clk),
    .Q(data_in_reg[0]),
    .QN(_0585_));
 DFF_X2 _0939_ (.D(_0180_),
    .CK(clknet_4_1__leaf_clk),
    .Q(data_in_reg[1]),
    .QN(_0586_));
 DFF_X2 _0940_ (.D(_0191_),
    .CK(clknet_4_9__leaf_clk),
    .Q(data_in_reg[2]),
    .QN(_0587_));
 DFF_X2 _0941_ (.D(_0194_),
    .CK(clknet_4_10__leaf_clk),
    .Q(data_in_reg[3]),
    .QN(_0588_));
 DFF_X2 _0942_ (.D(_0195_),
    .CK(clknet_4_0__leaf_clk),
    .Q(data_in_reg[4]),
    .QN(_0589_));
 DFF_X2 _0943_ (.D(_0196_),
    .CK(clknet_4_10__leaf_clk),
    .Q(data_in_reg[5]),
    .QN(_0590_));
 DFF_X2 _0944_ (.D(_0197_),
    .CK(clknet_4_12__leaf_clk),
    .Q(data_in_reg[6]),
    .QN(_0591_));
 DFF_X2 _0945_ (.D(_0198_),
    .CK(clknet_4_4__leaf_clk),
    .Q(data_in_reg[7]),
    .QN(_0592_));
 DFF_X2 _0946_ (.D(_0199_),
    .CK(clknet_4_10__leaf_clk),
    .Q(data_in_reg[8]),
    .QN(_0593_));
 DFF_X2 _0947_ (.D(_0200_),
    .CK(clknet_4_1__leaf_clk),
    .Q(data_in_reg[9]),
    .QN(_0594_));
 DFF_X2 _0948_ (.D(_0170_),
    .CK(clknet_4_10__leaf_clk),
    .Q(data_in_reg[10]),
    .QN(_0595_));
 DFF_X2 _0949_ (.D(_0171_),
    .CK(clknet_4_4__leaf_clk),
    .Q(data_in_reg[11]),
    .QN(_0596_));
 DFF_X2 _0950_ (.D(_0172_),
    .CK(clknet_4_14__leaf_clk),
    .Q(data_in_reg[12]),
    .QN(_0597_));
 DFF_X2 _0951_ (.D(_0173_),
    .CK(clknet_4_1__leaf_clk),
    .Q(data_in_reg[13]),
    .QN(_0598_));
 DFF_X2 _0952_ (.D(_0174_),
    .CK(clknet_4_10__leaf_clk),
    .Q(data_in_reg[14]),
    .QN(_0599_));
 DFF_X2 _0953_ (.D(_0175_),
    .CK(clknet_4_10__leaf_clk),
    .Q(data_in_reg[15]),
    .QN(_0600_));
 DFF_X2 _0954_ (.D(_0176_),
    .CK(clknet_4_1__leaf_clk),
    .Q(data_in_reg[16]),
    .QN(_0601_));
 DFF_X2 _0955_ (.D(_0177_),
    .CK(clknet_4_1__leaf_clk),
    .Q(data_in_reg[17]),
    .QN(_0602_));
 DFF_X2 _0956_ (.D(_0178_),
    .CK(clknet_4_2__leaf_clk),
    .Q(data_in_reg[18]),
    .QN(_0603_));
 DFF_X2 _0957_ (.D(_0179_),
    .CK(clknet_4_5__leaf_clk),
    .Q(data_in_reg[19]),
    .QN(_0604_));
 DFF_X2 _0958_ (.D(_0181_),
    .CK(clknet_4_5__leaf_clk),
    .Q(data_in_reg[20]),
    .QN(_0605_));
 DFF_X2 _0959_ (.D(_0182_),
    .CK(clknet_4_5__leaf_clk),
    .Q(data_in_reg[21]),
    .QN(_0606_));
 DFF_X2 _0960_ (.D(_0183_),
    .CK(clknet_4_10__leaf_clk),
    .Q(data_in_reg[22]),
    .QN(_0607_));
 DFF_X2 _0961_ (.D(_0184_),
    .CK(clknet_4_2__leaf_clk),
    .Q(data_in_reg[23]),
    .QN(_0608_));
 DFF_X2 _0962_ (.D(_0185_),
    .CK(clknet_4_10__leaf_clk),
    .Q(data_in_reg[24]),
    .QN(_0609_));
 DFF_X2 _0963_ (.D(_0186_),
    .CK(clknet_4_0__leaf_clk),
    .Q(data_in_reg[25]),
    .QN(_0610_));
 DFF_X2 _0964_ (.D(_0187_),
    .CK(clknet_4_3__leaf_clk),
    .Q(data_in_reg[26]),
    .QN(_0611_));
 DFF_X2 _0965_ (.D(_0188_),
    .CK(clknet_4_0__leaf_clk),
    .Q(data_in_reg[27]),
    .QN(_0612_));
 DFF_X2 _0966_ (.D(_0189_),
    .CK(clknet_4_14__leaf_clk),
    .Q(data_in_reg[28]),
    .QN(_0613_));
 DFF_X2 _0967_ (.D(_0190_),
    .CK(clknet_4_14__leaf_clk),
    .Q(data_in_reg[29]),
    .QN(_0614_));
 DFF_X2 _0968_ (.D(_0192_),
    .CK(clknet_4_0__leaf_clk),
    .Q(data_in_reg[30]),
    .QN(_0615_));
 DFF_X2 _0969_ (.D(_0193_),
    .CK(clknet_4_11__leaf_clk),
    .Q(data_in_reg[31]),
    .QN(_0616_));
 DFF_X2 _0970_ (.D(_0271_),
    .CK(clknet_4_3__leaf_clk),
    .Q(sram_rdata_reg[0]),
    .QN(_0617_));
 DFF_X2 _0971_ (.D(_0282_),
    .CK(clknet_4_12__leaf_clk),
    .Q(sram_rdata_reg[1]),
    .QN(_0618_));
 DFF_X2 _0972_ (.D(_0293_),
    .CK(clknet_4_12__leaf_clk),
    .Q(sram_rdata_reg[2]),
    .QN(_0619_));
 DFF_X2 _0973_ (.D(_0296_),
    .CK(clknet_4_12__leaf_clk),
    .Q(sram_rdata_reg[3]),
    .QN(_0620_));
 DFF_X2 _0974_ (.D(_0297_),
    .CK(clknet_4_12__leaf_clk),
    .Q(sram_rdata_reg[4]),
    .QN(_0621_));
 DFF_X2 _0975_ (.D(_0298_),
    .CK(clknet_4_12__leaf_clk),
    .Q(sram_rdata_reg[5]),
    .QN(_0622_));
 DFF_X2 _0976_ (.D(_0299_),
    .CK(clknet_4_12__leaf_clk),
    .Q(sram_rdata_reg[6]),
    .QN(_0623_));
 DFF_X2 _0977_ (.D(_0300_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[7]),
    .QN(_0624_));
 DFF_X2 _0978_ (.D(_0301_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[8]),
    .QN(_0625_));
 DFF_X2 _0979_ (.D(_0302_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[9]),
    .QN(_0626_));
 DFF_X2 _0980_ (.D(_0272_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[10]),
    .QN(_0627_));
 DFF_X2 _0981_ (.D(_0273_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[11]),
    .QN(_0628_));
 DFF_X2 _0982_ (.D(_0274_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[12]),
    .QN(_0629_));
 DFF_X2 _0983_ (.D(_0275_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[13]),
    .QN(_0630_));
 DFF_X2 _0984_ (.D(_0276_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[14]),
    .QN(_0631_));
 DFF_X2 _0985_ (.D(_0277_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[15]),
    .QN(_0632_));
 DFF_X2 _0986_ (.D(_0278_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[16]),
    .QN(_0633_));
 DFF_X2 _0987_ (.D(_0279_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[17]),
    .QN(_0634_));
 DFF_X2 _0988_ (.D(_0280_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[18]),
    .QN(_0635_));
 DFF_X2 _0989_ (.D(_0281_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[19]),
    .QN(_0636_));
 DFF_X2 _0990_ (.D(_0283_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[20]),
    .QN(_0637_));
 DFF_X2 _0991_ (.D(_0284_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[21]),
    .QN(_0638_));
 DFF_X2 _0992_ (.D(_0285_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[22]),
    .QN(_0639_));
 DFF_X2 _0993_ (.D(_0286_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[23]),
    .QN(_0640_));
 DFF_X2 _0994_ (.D(_0287_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[24]),
    .QN(_0641_));
 DFF_X2 _0995_ (.D(_0288_),
    .CK(clknet_4_15__leaf_clk),
    .Q(sram_rdata_reg[25]),
    .QN(_0642_));
 DFF_X2 _0996_ (.D(_0289_),
    .CK(clknet_4_15__leaf_clk),
    .Q(sram_rdata_reg[26]),
    .QN(_0643_));
 DFF_X2 _0997_ (.D(_0290_),
    .CK(clknet_4_15__leaf_clk),
    .Q(sram_rdata_reg[27]),
    .QN(_0644_));
 DFF_X2 _0998_ (.D(_0291_),
    .CK(clknet_4_15__leaf_clk),
    .Q(sram_rdata_reg[28]),
    .QN(_0645_));
 DFF_X2 _0999_ (.D(_0292_),
    .CK(clknet_4_15__leaf_clk),
    .Q(sram_rdata_reg[29]),
    .QN(_0646_));
 DFF_X2 _1000_ (.D(_0294_),
    .CK(clknet_4_15__leaf_clk),
    .Q(sram_rdata_reg[30]),
    .QN(_0647_));
 DFF_X2 _1001_ (.D(_0295_),
    .CK(clknet_4_15__leaf_clk),
    .Q(sram_rdata_reg[31]),
    .QN(_0648_));
 DFF_X2 _1002_ (.D(net9),
    .CK(clknet_4_11__leaf_clk),
    .Q(net113),
    .QN(_0649_));
 DFF_X2 _1003_ (.D(net210),
    .CK(clknet_4_7__leaf_clk),
    .Q(addr_ptr[0]),
    .QN(_0650_));
 DFF_X1 _1004_ (.D(_0164_),
    .CK(clknet_4_7__leaf_clk),
    .Q(addr_ptr[1]),
    .QN(_0651_));
 DFF_X1 _1005_ (.D(_0165_),
    .CK(clknet_4_7__leaf_clk),
    .Q(addr_ptr[2]),
    .QN(_0652_));
 DFF_X1 _1006_ (.D(_0166_),
    .CK(clknet_4_7__leaf_clk),
    .Q(addr_ptr[3]),
    .QN(_0653_));
 DFF_X1 _1007_ (.D(_0167_),
    .CK(clknet_4_7__leaf_clk),
    .Q(addr_ptr[4]),
    .QN(_0654_));
 DFF_X1 _1008_ (.D(net181),
    .CK(clknet_4_7__leaf_clk),
    .Q(addr_ptr[5]),
    .QN(_0655_));
 DFF_X1 _1009_ (.D(net186),
    .CK(clknet_4_6__leaf_clk),
    .Q(init_count[0]),
    .QN(_0656_));
 DFF_X1 _1010_ (.D(_0266_),
    .CK(clknet_4_6__leaf_clk),
    .Q(init_count[1]),
    .QN(_0657_));
 DFF_X1 _1011_ (.D(net194),
    .CK(clknet_4_6__leaf_clk),
    .Q(init_count[2]),
    .QN(_0658_));
 DFF_X2 _1012_ (.D(net205),
    .CK(clknet_4_6__leaf_clk),
    .Q(init_count[3]),
    .QN(_0659_));
 DFF_X1 _1013_ (.D(net197),
    .CK(clknet_4_6__leaf_clk),
    .Q(init_count[4]),
    .QN(_0660_));
 DFF_X1 _1014_ (.D(net191),
    .CK(clknet_4_6__leaf_clk),
    .Q(init_count[5]),
    .QN(_0661_));
 SRAM_6T_CORE_64x32_MC_TB sram_inst (.ce_in(_0307_),
    .we_in(_0308_),
    .clk(clknet_4_3__leaf_clk),
    .addr_in({net188,
    net183,
    net4,
    net6,
    net212,
    net179}),
    .rd_out({sram_rdata[31],
    sram_rdata[30],
    sram_rdata[29],
    sram_rdata[28],
    sram_rdata[27],
    sram_rdata[26],
    sram_rdata[25],
    sram_rdata[24],
    sram_rdata[23],
    sram_rdata[22],
    sram_rdata[21],
    sram_rdata[20],
    sram_rdata[19],
    sram_rdata[18],
    sram_rdata[17],
    sram_rdata[16],
    sram_rdata[15],
    sram_rdata[14],
    sram_rdata[13],
    sram_rdata[12],
    sram_rdata[11],
    sram_rdata[10],
    sram_rdata[9],
    sram_rdata[8],
    sram_rdata[7],
    sram_rdata[6],
    sram_rdata[5],
    sram_rdata[4],
    sram_rdata[3],
    sram_rdata[2],
    sram_rdata[1],
    sram_rdata[0]}),
    .wd_in({net224,
    data_in_reg[30],
    net231,
    net227,
    data_in_reg[27],
    data_in_reg[26],
    data_in_reg[25],
    net226,
    data_in_reg[23],
    net228,
    data_in_reg[21],
    data_in_reg[20],
    data_in_reg[19],
    net230,
    data_in_reg[17],
    data_in_reg[16],
    net218,
    net225,
    data_in_reg[13],
    net223,
    data_in_reg[11],
    net232,
    data_in_reg[9],
    data_in_reg[8],
    data_in_reg[7],
    net219,
    data_in_reg[5],
    data_in_reg[4],
    data_in_reg[3],
    net221,
    net229,
    net222}));
 AND2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__40_  (.A1(net147),
    .A2(u_multiplier_pp3_0 ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla1__25_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__41_  (.A1(net148),
    .A2(u_multiplier_pp3_0 ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla1__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__42_  (.A(net149),
    .B(u_multiplier_pp3_0 ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla1__27_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__43_  (.A(net161),
    .B(u_multiplier_Final_add_cla1_cla1_cla1_cla1__27_ ),
    .ZN(product[0]));
 AOI21_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__44_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla1__25_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla1_cla1__26_ ),
    .B2(net162),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla1__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__45_  (.A1(net150),
    .A2(u_multiplier_A [1]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla1__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__46_  (.A1(net151),
    .A2(u_multiplier_A [1]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla1__30_ ));
 XOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__47_  (.A(net152),
    .B(u_multiplier_A [1]),
    .Z(u_multiplier_Final_add_cla1_cla1_cla1_cla1__31_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__48_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla1__28_ ),
    .B(u_multiplier_Final_add_cla1_cla1_cla1_cla1__31_ ),
    .ZN(product[1]));
 OAI21_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__49_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla1__30_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla1_cla1__29_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla1_cla1__28_ ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla1__32_ ));
 AND2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__50_  (.A1(net153),
    .A2(u_multiplier_A [2]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla1__33_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__51_  (.A1(net154),
    .A2(u_multiplier_A [2]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla1__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__52_  (.A(net155),
    .B(u_multiplier_A [2]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla1__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__53_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla1__32_ ),
    .B(u_multiplier_Final_add_cla1_cla1_cla1_cla1__35_ ),
    .ZN(product[2]));
 AOI21_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__54_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla1__33_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla1_cla1__34_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla1_cla1__32_ ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla1__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__55_  (.A1(u_multiplier_B [3]),
    .A2(u_multiplier_A [3]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla1__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__56_  (.A1(u_multiplier_B [3]),
    .A2(u_multiplier_A [3]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla1__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__57_  (.A(u_multiplier_B [3]),
    .B(u_multiplier_A [3]),
    .Z(u_multiplier_Final_add_cla1_cla1_cla1_cla1__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__58_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla1__36_ ),
    .B(u_multiplier_Final_add_cla1_cla1_cla1_cla1__39_ ),
    .ZN(product[3]));
 OAI21_X2 u_multiplier_Final_add_cla1_cla1_cla1_cla1__59_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla1__38_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla1_cla1__37_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla1_cla1__36_ ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_c1 ));
 AND2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__40_  (.A1(u_multiplier_B [4]),
    .A2(u_multiplier_A [4]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla2__25_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__41_  (.A1(u_multiplier_B [4]),
    .A2(u_multiplier_A [4]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla2__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__42_  (.A(u_multiplier_B [4]),
    .B(u_multiplier_A [4]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla2__27_ ));
 XNOR2_X2 u_multiplier_Final_add_cla1_cla1_cla1_cla2__43_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_c1 ),
    .B(u_multiplier_Final_add_cla1_cla1_cla1_cla2__27_ ),
    .ZN(product[4]));
 AOI21_X2 u_multiplier_Final_add_cla1_cla1_cla1_cla2__44_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla2__25_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla1_cla2__26_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla1_c1 ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla2__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__45_  (.A1(u_multiplier_B [5]),
    .A2(u_multiplier_A [5]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla2__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__46_  (.A1(u_multiplier_B [5]),
    .A2(u_multiplier_A [5]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla2__30_ ));
 XOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__47_  (.A(u_multiplier_B [5]),
    .B(u_multiplier_A [5]),
    .Z(u_multiplier_Final_add_cla1_cla1_cla1_cla2__31_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__48_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla2__28_ ),
    .B(u_multiplier_Final_add_cla1_cla1_cla1_cla2__31_ ),
    .ZN(product[5]));
 OAI21_X2 u_multiplier_Final_add_cla1_cla1_cla1_cla2__49_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla2__30_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla1_cla2__29_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla1_cla2__28_ ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla2__32_ ));
 AND2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__50_  (.A1(u_multiplier_B [6]),
    .A2(u_multiplier_A [6]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla2__33_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__51_  (.A1(u_multiplier_B [6]),
    .A2(u_multiplier_A [6]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla2__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__52_  (.A(u_multiplier_B [6]),
    .B(u_multiplier_A [6]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla2__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__53_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla2__32_ ),
    .B(u_multiplier_Final_add_cla1_cla1_cla1_cla2__35_ ),
    .ZN(product[6]));
 AOI21_X2 u_multiplier_Final_add_cla1_cla1_cla1_cla2__54_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla2__33_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla1_cla2__34_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla1_cla2__32_ ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla2__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__55_  (.A1(u_multiplier_B [7]),
    .A2(u_multiplier_A [7]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla2__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__56_  (.A1(u_multiplier_B [7]),
    .A2(u_multiplier_A [7]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla2__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__57_  (.A(u_multiplier_B [7]),
    .B(u_multiplier_A [7]),
    .Z(u_multiplier_Final_add_cla1_cla1_cla1_cla2__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__58_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla2__36_ ),
    .B(u_multiplier_Final_add_cla1_cla1_cla1_cla2__39_ ),
    .ZN(product[7]));
 OAI21_X2 u_multiplier_Final_add_cla1_cla1_cla1_cla2__59_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla2__38_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla1_cla2__37_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla1_cla2__36_ ),
    .ZN(u_multiplier_Final_add_cla1_cla1_c1 ));
 AND2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__40_  (.A1(u_multiplier_B [8]),
    .A2(u_multiplier_A [8]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla1__25_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__41_  (.A1(u_multiplier_B [8]),
    .A2(u_multiplier_A [8]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla1__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__42_  (.A(u_multiplier_B [8]),
    .B(u_multiplier_A [8]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla1__27_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__43_  (.A(u_multiplier_Final_add_cla1_cla1_c1 ),
    .B(u_multiplier_Final_add_cla1_cla1_cla2_cla1__27_ ),
    .ZN(product[8]));
 AOI21_X2 u_multiplier_Final_add_cla1_cla1_cla2_cla1__44_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla1__25_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla2_cla1__26_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_c1 ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla1__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__45_  (.A1(u_multiplier_B [9]),
    .A2(u_multiplier_A [9]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla1__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__46_  (.A1(u_multiplier_B [9]),
    .A2(u_multiplier_A [9]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla1__30_ ));
 XOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__47_  (.A(u_multiplier_B [9]),
    .B(u_multiplier_A [9]),
    .Z(u_multiplier_Final_add_cla1_cla1_cla2_cla1__31_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__48_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla1__28_ ),
    .B(u_multiplier_Final_add_cla1_cla1_cla2_cla1__31_ ),
    .ZN(product[9]));
 OAI21_X2 u_multiplier_Final_add_cla1_cla1_cla2_cla1__49_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla1__30_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla2_cla1__29_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla2_cla1__28_ ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla1__32_ ));
 AND2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__50_  (.A1(u_multiplier_B [10]),
    .A2(u_multiplier_A [10]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla1__33_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__51_  (.A1(u_multiplier_B [10]),
    .A2(u_multiplier_A [10]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla1__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__52_  (.A(u_multiplier_B [10]),
    .B(u_multiplier_A [10]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla1__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__53_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla1__32_ ),
    .B(u_multiplier_Final_add_cla1_cla1_cla2_cla1__35_ ),
    .ZN(product[10]));
 AOI21_X2 u_multiplier_Final_add_cla1_cla1_cla2_cla1__54_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla1__33_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla2_cla1__34_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla2_cla1__32_ ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla1__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__55_  (.A1(u_multiplier_B [11]),
    .A2(u_multiplier_A [11]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla1__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__56_  (.A1(u_multiplier_B [11]),
    .A2(u_multiplier_A [11]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla1__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__57_  (.A(u_multiplier_B [11]),
    .B(u_multiplier_A [11]),
    .Z(u_multiplier_Final_add_cla1_cla1_cla2_cla1__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__58_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla1__36_ ),
    .B(u_multiplier_Final_add_cla1_cla1_cla2_cla1__39_ ),
    .ZN(product[11]));
 OAI21_X2 u_multiplier_Final_add_cla1_cla1_cla2_cla1__59_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla1__38_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla2_cla1__37_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla2_cla1__36_ ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_c1 ));
 AND2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__40_  (.A1(u_multiplier_B [12]),
    .A2(u_multiplier_A [12]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla2__25_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__41_  (.A1(u_multiplier_B [12]),
    .A2(u_multiplier_A [12]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla2__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__42_  (.A(u_multiplier_B [12]),
    .B(u_multiplier_A [12]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla2__27_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__43_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_c1 ),
    .B(u_multiplier_Final_add_cla1_cla1_cla2_cla2__27_ ),
    .ZN(product[12]));
 AOI21_X2 u_multiplier_Final_add_cla1_cla1_cla2_cla2__44_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla2__25_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla2_cla2__26_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla2_c1 ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla2__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__45_  (.A1(u_multiplier_B [13]),
    .A2(u_multiplier_A [13]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla2__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__46_  (.A1(u_multiplier_B [13]),
    .A2(u_multiplier_A [13]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla2__30_ ));
 XOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__47_  (.A(u_multiplier_B [13]),
    .B(u_multiplier_A [13]),
    .Z(u_multiplier_Final_add_cla1_cla1_cla2_cla2__31_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__48_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla2__28_ ),
    .B(u_multiplier_Final_add_cla1_cla1_cla2_cla2__31_ ),
    .ZN(product[13]));
 OAI21_X2 u_multiplier_Final_add_cla1_cla1_cla2_cla2__49_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla2__30_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla2_cla2__29_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla2_cla2__28_ ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla2__32_ ));
 AND2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__50_  (.A1(u_multiplier_B [14]),
    .A2(u_multiplier_A [14]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla2__33_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__51_  (.A1(u_multiplier_B [14]),
    .A2(u_multiplier_A [14]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla2__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__52_  (.A(u_multiplier_B [14]),
    .B(u_multiplier_A [14]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla2__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__53_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla2__32_ ),
    .B(u_multiplier_Final_add_cla1_cla1_cla2_cla2__35_ ),
    .ZN(product[14]));
 AOI21_X2 u_multiplier_Final_add_cla1_cla1_cla2_cla2__54_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla2__33_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla2_cla2__34_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla2_cla2__32_ ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla2__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__55_  (.A1(u_multiplier_B [15]),
    .A2(u_multiplier_A [15]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla2__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__56_  (.A1(u_multiplier_B [15]),
    .A2(u_multiplier_A [15]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla2__38_ ));
 XOR2_X2 u_multiplier_Final_add_cla1_cla1_cla2_cla2__57_  (.A(u_multiplier_B [15]),
    .B(u_multiplier_A [15]),
    .Z(u_multiplier_Final_add_cla1_cla1_cla2_cla2__39_ ));
 XNOR2_X2 u_multiplier_Final_add_cla1_cla1_cla2_cla2__58_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla2__36_ ),
    .B(u_multiplier_Final_add_cla1_cla1_cla2_cla2__39_ ),
    .ZN(product[15]));
 OAI21_X2 u_multiplier_Final_add_cla1_cla1_cla2_cla2__59_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla2__38_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla2_cla2__37_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla2_cla2__36_ ),
    .ZN(u_multiplier_Final_add_cla1_c1 ));
 AND2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__40_  (.A1(u_multiplier_B [16]),
    .A2(u_multiplier_A [16]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla1__25_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__41_  (.A1(u_multiplier_B [16]),
    .A2(u_multiplier_A [16]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla1__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__42_  (.A(u_multiplier_B [16]),
    .B(u_multiplier_A [16]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla1__27_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__43_  (.A(u_multiplier_Final_add_cla1_c1 ),
    .B(u_multiplier_Final_add_cla1_cla2_cla1_cla1__27_ ),
    .ZN(product[16]));
 AOI21_X2 u_multiplier_Final_add_cla1_cla2_cla1_cla1__44_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla1__25_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla1_cla1__26_ ),
    .B2(u_multiplier_Final_add_cla1_c1 ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla1__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__45_  (.A1(u_multiplier_B [17]),
    .A2(u_multiplier_A [17]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla1__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__46_  (.A1(u_multiplier_B [17]),
    .A2(u_multiplier_A [17]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla1__30_ ));
 XOR2_X2 u_multiplier_Final_add_cla1_cla2_cla1_cla1__47_  (.A(u_multiplier_B [17]),
    .B(u_multiplier_A [17]),
    .Z(u_multiplier_Final_add_cla1_cla2_cla1_cla1__31_ ));
 XNOR2_X2 u_multiplier_Final_add_cla1_cla2_cla1_cla1__48_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla1__28_ ),
    .B(u_multiplier_Final_add_cla1_cla2_cla1_cla1__31_ ),
    .ZN(product[17]));
 OAI21_X2 u_multiplier_Final_add_cla1_cla2_cla1_cla1__49_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla1__30_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla1_cla1__29_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla1_cla1__28_ ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla1__32_ ));
 AND2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__50_  (.A1(u_multiplier_B [18]),
    .A2(u_multiplier_A [18]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla1__33_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__51_  (.A1(u_multiplier_B [18]),
    .A2(u_multiplier_A [18]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla1__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__52_  (.A(u_multiplier_B [18]),
    .B(u_multiplier_A [18]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla1__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__53_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla1__32_ ),
    .B(u_multiplier_Final_add_cla1_cla2_cla1_cla1__35_ ),
    .ZN(product[18]));
 AOI21_X2 u_multiplier_Final_add_cla1_cla2_cla1_cla1__54_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla1__33_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla1_cla1__34_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla1_cla1__32_ ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla1__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__55_  (.A1(u_multiplier_B [19]),
    .A2(u_multiplier_A [19]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla1__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__56_  (.A1(u_multiplier_B [19]),
    .A2(u_multiplier_A [19]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla1__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__57_  (.A(u_multiplier_B [19]),
    .B(u_multiplier_A [19]),
    .Z(u_multiplier_Final_add_cla1_cla2_cla1_cla1__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__58_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla1__36_ ),
    .B(u_multiplier_Final_add_cla1_cla2_cla1_cla1__39_ ),
    .ZN(product[19]));
 OAI21_X2 u_multiplier_Final_add_cla1_cla2_cla1_cla1__59_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla1__38_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla1_cla1__37_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla1_cla1__36_ ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_c1 ));
 AND2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla2__40_  (.A1(u_multiplier_B [20]),
    .A2(u_multiplier_A [20]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla2__25_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla2__41_  (.A1(u_multiplier_B [20]),
    .A2(u_multiplier_A [20]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla2__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla2__42_  (.A(u_multiplier_B [20]),
    .B(u_multiplier_A [20]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla2__27_ ));
 XNOR2_X2 u_multiplier_Final_add_cla1_cla2_cla1_cla2__43_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_c1 ),
    .B(u_multiplier_Final_add_cla1_cla2_cla1_cla2__27_ ),
    .ZN(product[20]));
 AOI21_X2 u_multiplier_Final_add_cla1_cla2_cla1_cla2__44_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla2__25_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla1_cla2__26_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla1_c1 ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla2__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla2__45_  (.A1(u_multiplier_B [21]),
    .A2(u_multiplier_A [21]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla2__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla2__46_  (.A1(u_multiplier_B [21]),
    .A2(u_multiplier_A [21]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla2__30_ ));
 XOR2_X2 u_multiplier_Final_add_cla1_cla2_cla1_cla2__47_  (.A(u_multiplier_B [21]),
    .B(u_multiplier_A [21]),
    .Z(u_multiplier_Final_add_cla1_cla2_cla1_cla2__31_ ));
 XNOR2_X2 u_multiplier_Final_add_cla1_cla2_cla1_cla2__48_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla2__28_ ),
    .B(u_multiplier_Final_add_cla1_cla2_cla1_cla2__31_ ),
    .ZN(product[21]));
 OAI21_X2 u_multiplier_Final_add_cla1_cla2_cla1_cla2__49_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla2__30_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla1_cla2__29_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla1_cla2__28_ ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla2__32_ ));
 AND2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla2__50_  (.A1(u_multiplier_B [22]),
    .A2(u_multiplier_A [22]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla2__33_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla2__51_  (.A1(u_multiplier_B [22]),
    .A2(u_multiplier_A [22]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla2__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla2__52_  (.A(u_multiplier_B [22]),
    .B(u_multiplier_A [22]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla2__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla2__53_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla2__32_ ),
    .B(u_multiplier_Final_add_cla1_cla2_cla1_cla2__35_ ),
    .ZN(product[22]));
 AOI21_X2 u_multiplier_Final_add_cla1_cla2_cla1_cla2__54_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla2__33_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla1_cla2__34_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla1_cla2__32_ ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla2__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla2__55_  (.A1(u_multiplier_B [23]),
    .A2(u_multiplier_A [23]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla2__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla2__56_  (.A1(u_multiplier_B [23]),
    .A2(u_multiplier_A [23]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla2__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla2__57_  (.A(u_multiplier_B [23]),
    .B(u_multiplier_A [23]),
    .Z(u_multiplier_Final_add_cla1_cla2_cla1_cla2__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla2__58_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla2__36_ ),
    .B(u_multiplier_Final_add_cla1_cla2_cla1_cla2__39_ ),
    .ZN(product[23]));
 OAI21_X2 u_multiplier_Final_add_cla1_cla2_cla1_cla2__59_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla2__38_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla1_cla2__37_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla1_cla2__36_ ),
    .ZN(u_multiplier_Final_add_cla1_cla2_c1 ));
 AND2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__40_  (.A1(u_multiplier_B [24]),
    .A2(u_multiplier_A [24]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla1__25_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__41_  (.A1(u_multiplier_B [24]),
    .A2(u_multiplier_A [24]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla1__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__42_  (.A(u_multiplier_B [24]),
    .B(u_multiplier_A [24]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla1__27_ ));
 XNOR2_X2 u_multiplier_Final_add_cla1_cla2_cla2_cla1__43_  (.A(u_multiplier_Final_add_cla1_cla2_c1 ),
    .B(u_multiplier_Final_add_cla1_cla2_cla2_cla1__27_ ),
    .ZN(product[24]));
 AOI21_X2 u_multiplier_Final_add_cla1_cla2_cla2_cla1__44_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla1__25_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla2_cla1__26_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_c1 ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla1__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__45_  (.A1(u_multiplier_B [25]),
    .A2(u_multiplier_A [25]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla1__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__46_  (.A1(u_multiplier_B [25]),
    .A2(u_multiplier_A [25]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla1__30_ ));
 XOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__47_  (.A(u_multiplier_B [25]),
    .B(u_multiplier_A [25]),
    .Z(u_multiplier_Final_add_cla1_cla2_cla2_cla1__31_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__48_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla1__28_ ),
    .B(u_multiplier_Final_add_cla1_cla2_cla2_cla1__31_ ),
    .ZN(product[25]));
 OAI21_X2 u_multiplier_Final_add_cla1_cla2_cla2_cla1__49_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla1__30_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla2_cla1__29_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla2_cla1__28_ ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla1__32_ ));
 AND2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__50_  (.A1(u_multiplier_B [26]),
    .A2(u_multiplier_A [26]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla1__33_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__51_  (.A1(u_multiplier_B [26]),
    .A2(u_multiplier_A [26]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla1__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__52_  (.A(u_multiplier_B [26]),
    .B(u_multiplier_A [26]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla1__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__53_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla1__32_ ),
    .B(u_multiplier_Final_add_cla1_cla2_cla2_cla1__35_ ),
    .ZN(product[26]));
 AOI21_X2 u_multiplier_Final_add_cla1_cla2_cla2_cla1__54_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla1__33_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla2_cla1__34_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla2_cla1__32_ ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla1__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__55_  (.A1(u_multiplier_B [27]),
    .A2(u_multiplier_A [27]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla1__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__56_  (.A1(u_multiplier_B [27]),
    .A2(u_multiplier_A [27]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla1__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__57_  (.A(u_multiplier_B [27]),
    .B(u_multiplier_A [27]),
    .Z(u_multiplier_Final_add_cla1_cla2_cla2_cla1__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__58_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla1__36_ ),
    .B(u_multiplier_Final_add_cla1_cla2_cla2_cla1__39_ ),
    .ZN(product[27]));
 OAI21_X2 u_multiplier_Final_add_cla1_cla2_cla2_cla1__59_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla1__38_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla2_cla1__37_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla2_cla1__36_ ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_c1 ));
 AND2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__40_  (.A1(u_multiplier_B [28]),
    .A2(u_multiplier_A [28]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla2__25_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__41_  (.A1(u_multiplier_B [28]),
    .A2(u_multiplier_A [28]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla2__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__42_  (.A(u_multiplier_B [28]),
    .B(u_multiplier_A [28]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla2__27_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__43_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_c1 ),
    .B(u_multiplier_Final_add_cla1_cla2_cla2_cla2__27_ ),
    .ZN(product[28]));
 AOI21_X4 u_multiplier_Final_add_cla1_cla2_cla2_cla2__44_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla2__25_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla2_cla2__26_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla2_c1 ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla2__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__45_  (.A1(u_multiplier_B [29]),
    .A2(u_multiplier_A [29]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla2__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__46_  (.A1(u_multiplier_B [29]),
    .A2(u_multiplier_A [29]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla2__30_ ));
 XOR2_X2 u_multiplier_Final_add_cla1_cla2_cla2_cla2__47_  (.A(u_multiplier_B [29]),
    .B(u_multiplier_A [29]),
    .Z(u_multiplier_Final_add_cla1_cla2_cla2_cla2__31_ ));
 XNOR2_X2 u_multiplier_Final_add_cla1_cla2_cla2_cla2__48_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla2__28_ ),
    .B(u_multiplier_Final_add_cla1_cla2_cla2_cla2__31_ ),
    .ZN(product[29]));
 OAI21_X2 u_multiplier_Final_add_cla1_cla2_cla2_cla2__49_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla2__30_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla2_cla2__29_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla2_cla2__28_ ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla2__32_ ));
 AND2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__50_  (.A1(u_multiplier_B [30]),
    .A2(u_multiplier_A [30]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla2__33_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__51_  (.A1(u_multiplier_B [30]),
    .A2(u_multiplier_A [30]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla2__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__52_  (.A(u_multiplier_B [30]),
    .B(u_multiplier_A [30]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla2__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__53_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla2__32_ ),
    .B(u_multiplier_Final_add_cla1_cla2_cla2_cla2__35_ ),
    .ZN(product[30]));
 AOI21_X4 u_multiplier_Final_add_cla1_cla2_cla2_cla2__54_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla2__33_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla2_cla2__34_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla2_cla2__32_ ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla2__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__55_  (.A1(u_multiplier_B [31]),
    .A2(u_multiplier_A [31]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla2__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__56_  (.A1(u_multiplier_B [31]),
    .A2(u_multiplier_A [31]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla2__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__57_  (.A(u_multiplier_B [31]),
    .B(u_multiplier_A [31]),
    .Z(u_multiplier_Final_add_cla1_cla2_cla2_cla2__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__58_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla2__36_ ),
    .B(u_multiplier_Final_add_cla1_cla2_cla2_cla2__39_ ),
    .ZN(product[31]));
 OAI21_X4 u_multiplier_Final_add_cla1_cla2_cla2_cla2__59_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla2__38_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla2_cla2__37_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla2_cla2__36_ ),
    .ZN(u_multiplier_Final_add_c1 ));
 AND2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__40_  (.A1(u_multiplier_B [32]),
    .A2(u_multiplier_A [32]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla1__25_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__41_  (.A1(u_multiplier_B [32]),
    .A2(u_multiplier_A [32]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla1__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__42_  (.A(u_multiplier_B [32]),
    .B(u_multiplier_A [32]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla1__27_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__43_  (.A(u_multiplier_Final_add_c1 ),
    .B(u_multiplier_Final_add_cla2_cla1_cla1_cla1__27_ ),
    .ZN(product[32]));
 AOI21_X4 u_multiplier_Final_add_cla2_cla1_cla1_cla1__44_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla1__25_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla1_cla1__26_ ),
    .B2(u_multiplier_Final_add_c1 ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla1__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__45_  (.A1(u_multiplier_B [33]),
    .A2(u_multiplier_A [33]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla1__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__46_  (.A1(u_multiplier_B [33]),
    .A2(u_multiplier_A [33]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla1__30_ ));
 XOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__47_  (.A(u_multiplier_B [33]),
    .B(u_multiplier_A [33]),
    .Z(u_multiplier_Final_add_cla2_cla1_cla1_cla1__31_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__48_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla1__28_ ),
    .B(u_multiplier_Final_add_cla2_cla1_cla1_cla1__31_ ),
    .ZN(product[33]));
 OAI21_X4 u_multiplier_Final_add_cla2_cla1_cla1_cla1__49_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla1__30_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla1_cla1__29_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla1_cla1__28_ ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla1__32_ ));
 AND2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__50_  (.A1(u_multiplier_B [34]),
    .A2(u_multiplier_A [34]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla1__33_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__51_  (.A1(u_multiplier_B [34]),
    .A2(u_multiplier_A [34]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla1__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__52_  (.A(u_multiplier_B [34]),
    .B(u_multiplier_A [34]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla1__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__53_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla1__32_ ),
    .B(u_multiplier_Final_add_cla2_cla1_cla1_cla1__35_ ),
    .ZN(product[34]));
 AOI21_X2 u_multiplier_Final_add_cla2_cla1_cla1_cla1__54_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla1__33_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla1_cla1__34_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla1_cla1__32_ ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla1__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__55_  (.A1(u_multiplier_B [35]),
    .A2(u_multiplier_A [35]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla1__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__56_  (.A1(u_multiplier_B [35]),
    .A2(u_multiplier_A [35]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla1__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__57_  (.A(u_multiplier_B [35]),
    .B(u_multiplier_A [35]),
    .Z(u_multiplier_Final_add_cla2_cla1_cla1_cla1__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__58_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla1__36_ ),
    .B(u_multiplier_Final_add_cla2_cla1_cla1_cla1__39_ ),
    .ZN(product[35]));
 OAI21_X2 u_multiplier_Final_add_cla2_cla1_cla1_cla1__59_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla1__38_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla1_cla1__37_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla1_cla1__36_ ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_c1 ));
 AND2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla2__40_  (.A1(u_multiplier_B [36]),
    .A2(u_multiplier_A [36]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla2__25_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla2__41_  (.A1(u_multiplier_B [36]),
    .A2(u_multiplier_A [36]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla2__26_ ));
 XNOR2_X2 u_multiplier_Final_add_cla2_cla1_cla1_cla2__42_  (.A(u_multiplier_B [36]),
    .B(u_multiplier_A [36]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla2__27_ ));
 XNOR2_X2 u_multiplier_Final_add_cla2_cla1_cla1_cla2__43_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_c1 ),
    .B(u_multiplier_Final_add_cla2_cla1_cla1_cla2__27_ ),
    .ZN(product[36]));
 AOI21_X2 u_multiplier_Final_add_cla2_cla1_cla1_cla2__44_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla2__25_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla1_cla2__26_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla1_c1 ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla2__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla2__45_  (.A1(u_multiplier_B [37]),
    .A2(u_multiplier_A [37]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla2__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla2__46_  (.A1(u_multiplier_B [37]),
    .A2(u_multiplier_A [37]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla2__30_ ));
 XOR2_X2 u_multiplier_Final_add_cla2_cla1_cla1_cla2__47_  (.A(u_multiplier_B [37]),
    .B(u_multiplier_A [37]),
    .Z(u_multiplier_Final_add_cla2_cla1_cla1_cla2__31_ ));
 XNOR2_X2 u_multiplier_Final_add_cla2_cla1_cla1_cla2__48_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla2__28_ ),
    .B(u_multiplier_Final_add_cla2_cla1_cla1_cla2__31_ ),
    .ZN(product[37]));
 OAI21_X2 u_multiplier_Final_add_cla2_cla1_cla1_cla2__49_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla2__30_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla1_cla2__29_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla1_cla2__28_ ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla2__32_ ));
 AND2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla2__50_  (.A1(u_multiplier_B [38]),
    .A2(u_multiplier_A [38]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla2__33_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla2__51_  (.A1(u_multiplier_B [38]),
    .A2(u_multiplier_A [38]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla2__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla2__52_  (.A(u_multiplier_B [38]),
    .B(u_multiplier_A [38]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla2__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla2__53_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla2__32_ ),
    .B(u_multiplier_Final_add_cla2_cla1_cla1_cla2__35_ ),
    .ZN(product[38]));
 AOI21_X2 u_multiplier_Final_add_cla2_cla1_cla1_cla2__54_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla2__33_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla1_cla2__34_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla1_cla2__32_ ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla2__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla2__55_  (.A1(u_multiplier_B [39]),
    .A2(u_multiplier_A [39]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla2__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla2__56_  (.A1(u_multiplier_B [39]),
    .A2(u_multiplier_A [39]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla2__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla2__57_  (.A(u_multiplier_B [39]),
    .B(u_multiplier_A [39]),
    .Z(u_multiplier_Final_add_cla2_cla1_cla1_cla2__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla2__58_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla2__36_ ),
    .B(u_multiplier_Final_add_cla2_cla1_cla1_cla2__39_ ),
    .ZN(product[39]));
 OAI21_X2 u_multiplier_Final_add_cla2_cla1_cla1_cla2__59_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla2__38_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla1_cla2__37_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla1_cla2__36_ ),
    .ZN(u_multiplier_Final_add_cla2_cla1_c1 ));
 AND2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__40_  (.A1(u_multiplier_B [40]),
    .A2(u_multiplier_A [40]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla1__25_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__41_  (.A1(u_multiplier_B [40]),
    .A2(u_multiplier_A [40]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla1__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__42_  (.A(u_multiplier_B [40]),
    .B(u_multiplier_A [40]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla1__27_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__43_  (.A(u_multiplier_Final_add_cla2_cla1_c1 ),
    .B(u_multiplier_Final_add_cla2_cla1_cla2_cla1__27_ ),
    .ZN(product[40]));
 AOI21_X2 u_multiplier_Final_add_cla2_cla1_cla2_cla1__44_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla1__25_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla2_cla1__26_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_c1 ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla1__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__45_  (.A1(u_multiplier_B [41]),
    .A2(u_multiplier_A [41]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla1__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__46_  (.A1(u_multiplier_B [41]),
    .A2(u_multiplier_A [41]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla1__30_ ));
 XOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__47_  (.A(u_multiplier_B [41]),
    .B(u_multiplier_A [41]),
    .Z(u_multiplier_Final_add_cla2_cla1_cla2_cla1__31_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__48_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla1__28_ ),
    .B(u_multiplier_Final_add_cla2_cla1_cla2_cla1__31_ ),
    .ZN(product[41]));
 OAI21_X2 u_multiplier_Final_add_cla2_cla1_cla2_cla1__49_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla1__30_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla2_cla1__29_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla2_cla1__28_ ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla1__32_ ));
 AND2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__50_  (.A1(u_multiplier_B [42]),
    .A2(u_multiplier_A [42]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla1__33_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__51_  (.A1(u_multiplier_B [42]),
    .A2(u_multiplier_A [42]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla1__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__52_  (.A(u_multiplier_B [42]),
    .B(u_multiplier_A [42]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla1__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__53_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla1__32_ ),
    .B(u_multiplier_Final_add_cla2_cla1_cla2_cla1__35_ ),
    .ZN(product[42]));
 AOI21_X4 u_multiplier_Final_add_cla2_cla1_cla2_cla1__54_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla1__33_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla2_cla1__34_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla2_cla1__32_ ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla1__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__55_  (.A1(u_multiplier_B [43]),
    .A2(u_multiplier_A [43]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla1__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__56_  (.A1(u_multiplier_B [43]),
    .A2(u_multiplier_A [43]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla1__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__57_  (.A(u_multiplier_B [43]),
    .B(u_multiplier_A [43]),
    .Z(u_multiplier_Final_add_cla2_cla1_cla2_cla1__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__58_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla1__36_ ),
    .B(u_multiplier_Final_add_cla2_cla1_cla2_cla1__39_ ),
    .ZN(product[43]));
 OAI21_X2 u_multiplier_Final_add_cla2_cla1_cla2_cla1__59_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla1__38_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla2_cla1__37_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla2_cla1__36_ ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_c1 ));
 AND2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__40_  (.A1(u_multiplier_B [44]),
    .A2(u_multiplier_A [44]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla2__25_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__41_  (.A1(u_multiplier_B [44]),
    .A2(u_multiplier_A [44]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla2__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__42_  (.A(u_multiplier_B [44]),
    .B(u_multiplier_A [44]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla2__27_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__43_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_c1 ),
    .B(u_multiplier_Final_add_cla2_cla1_cla2_cla2__27_ ),
    .ZN(product[44]));
 AOI21_X2 u_multiplier_Final_add_cla2_cla1_cla2_cla2__44_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla2__25_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla2_cla2__26_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla2_c1 ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla2__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__45_  (.A1(u_multiplier_B [45]),
    .A2(u_multiplier_A [45]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla2__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__46_  (.A1(u_multiplier_B [45]),
    .A2(u_multiplier_A [45]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla2__30_ ));
 XOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__47_  (.A(u_multiplier_B [45]),
    .B(u_multiplier_A [45]),
    .Z(u_multiplier_Final_add_cla2_cla1_cla2_cla2__31_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__48_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla2__28_ ),
    .B(u_multiplier_Final_add_cla2_cla1_cla2_cla2__31_ ),
    .ZN(product[45]));
 OAI21_X2 u_multiplier_Final_add_cla2_cla1_cla2_cla2__49_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla2__30_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla2_cla2__29_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla2_cla2__28_ ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla2__32_ ));
 AND2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__50_  (.A1(u_multiplier_B [46]),
    .A2(u_multiplier_A [46]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla2__33_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__51_  (.A1(u_multiplier_B [46]),
    .A2(u_multiplier_A [46]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla2__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__52_  (.A(u_multiplier_B [46]),
    .B(u_multiplier_A [46]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla2__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__53_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla2__32_ ),
    .B(u_multiplier_Final_add_cla2_cla1_cla2_cla2__35_ ),
    .ZN(product[46]));
 AOI21_X2 u_multiplier_Final_add_cla2_cla1_cla2_cla2__54_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla2__33_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla2_cla2__34_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla2_cla2__32_ ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla2__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__55_  (.A1(u_multiplier_B [47]),
    .A2(u_multiplier_A [47]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla2__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__56_  (.A1(u_multiplier_B [47]),
    .A2(u_multiplier_A [47]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla2__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__57_  (.A(u_multiplier_B [47]),
    .B(u_multiplier_A [47]),
    .Z(u_multiplier_Final_add_cla2_cla1_cla2_cla2__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__58_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla2__36_ ),
    .B(u_multiplier_Final_add_cla2_cla1_cla2_cla2__39_ ),
    .ZN(product[47]));
 OAI21_X2 u_multiplier_Final_add_cla2_cla1_cla2_cla2__59_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla2__38_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla2_cla2__37_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla2_cla2__36_ ),
    .ZN(u_multiplier_Final_add_cla2_c1 ));
 AND2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__40_  (.A1(u_multiplier_B [48]),
    .A2(u_multiplier_A [48]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla1__25_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__41_  (.A1(u_multiplier_B [48]),
    .A2(u_multiplier_A [48]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla1__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__42_  (.A(u_multiplier_B [48]),
    .B(u_multiplier_A [48]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla1__27_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__43_  (.A(u_multiplier_Final_add_cla2_c1 ),
    .B(u_multiplier_Final_add_cla2_cla2_cla1_cla1__27_ ),
    .ZN(product[48]));
 AOI21_X2 u_multiplier_Final_add_cla2_cla2_cla1_cla1__44_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla1__25_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla1_cla1__26_ ),
    .B2(u_multiplier_Final_add_cla2_c1 ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla1__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__45_  (.A1(u_multiplier_B [49]),
    .A2(u_multiplier_A [49]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla1__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__46_  (.A1(u_multiplier_B [49]),
    .A2(u_multiplier_A [49]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla1__30_ ));
 XOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__47_  (.A(u_multiplier_B [49]),
    .B(u_multiplier_A [49]),
    .Z(u_multiplier_Final_add_cla2_cla2_cla1_cla1__31_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__48_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla1__28_ ),
    .B(u_multiplier_Final_add_cla2_cla2_cla1_cla1__31_ ),
    .ZN(product[49]));
 OAI21_X2 u_multiplier_Final_add_cla2_cla2_cla1_cla1__49_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla1__30_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla1_cla1__29_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla1_cla1__28_ ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla1__32_ ));
 AND2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__50_  (.A1(u_multiplier_B [50]),
    .A2(u_multiplier_A [50]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla1__33_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__51_  (.A1(u_multiplier_B [50]),
    .A2(u_multiplier_A [50]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla1__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__52_  (.A(u_multiplier_B [50]),
    .B(u_multiplier_A [50]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla1__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__53_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla1__32_ ),
    .B(u_multiplier_Final_add_cla2_cla2_cla1_cla1__35_ ),
    .ZN(product[50]));
 AOI21_X2 u_multiplier_Final_add_cla2_cla2_cla1_cla1__54_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla1__33_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla1_cla1__34_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla1_cla1__32_ ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla1__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__55_  (.A1(u_multiplier_B [51]),
    .A2(u_multiplier_A [51]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla1__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__56_  (.A1(u_multiplier_B [51]),
    .A2(u_multiplier_A [51]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla1__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__57_  (.A(u_multiplier_B [51]),
    .B(u_multiplier_A [51]),
    .Z(u_multiplier_Final_add_cla2_cla2_cla1_cla1__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__58_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla1__36_ ),
    .B(u_multiplier_Final_add_cla2_cla2_cla1_cla1__39_ ),
    .ZN(product[51]));
 OAI21_X2 u_multiplier_Final_add_cla2_cla2_cla1_cla1__59_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla1__38_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla1_cla1__37_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla1_cla1__36_ ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_c1 ));
 AND2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__40_  (.A1(u_multiplier_B [52]),
    .A2(u_multiplier_A [52]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla2__25_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__41_  (.A1(u_multiplier_B [52]),
    .A2(u_multiplier_A [52]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla2__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__42_  (.A(u_multiplier_B [52]),
    .B(u_multiplier_A [52]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla2__27_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__43_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_c1 ),
    .B(u_multiplier_Final_add_cla2_cla2_cla1_cla2__27_ ),
    .ZN(product[52]));
 AOI21_X4 u_multiplier_Final_add_cla2_cla2_cla1_cla2__44_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla2__25_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla1_cla2__26_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla1_c1 ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla2__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__45_  (.A1(u_multiplier_B [53]),
    .A2(u_multiplier_A [53]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla2__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__46_  (.A1(u_multiplier_B [53]),
    .A2(u_multiplier_A [53]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla2__30_ ));
 XOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__47_  (.A(u_multiplier_B [53]),
    .B(u_multiplier_A [53]),
    .Z(u_multiplier_Final_add_cla2_cla2_cla1_cla2__31_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__48_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla2__28_ ),
    .B(u_multiplier_Final_add_cla2_cla2_cla1_cla2__31_ ),
    .ZN(product[53]));
 OAI21_X4 u_multiplier_Final_add_cla2_cla2_cla1_cla2__49_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla2__30_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla1_cla2__29_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla1_cla2__28_ ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla2__32_ ));
 AND2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__50_  (.A1(u_multiplier_B [54]),
    .A2(u_multiplier_A [54]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla2__33_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__51_  (.A1(u_multiplier_B [54]),
    .A2(u_multiplier_A [54]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla2__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__52_  (.A(u_multiplier_B [54]),
    .B(u_multiplier_A [54]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla2__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__53_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla2__32_ ),
    .B(u_multiplier_Final_add_cla2_cla2_cla1_cla2__35_ ),
    .ZN(product[54]));
 AOI21_X4 u_multiplier_Final_add_cla2_cla2_cla1_cla2__54_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla2__33_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla1_cla2__34_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla1_cla2__32_ ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla2__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__55_  (.A1(u_multiplier_B [55]),
    .A2(u_multiplier_A [55]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla2__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__56_  (.A1(u_multiplier_B [55]),
    .A2(u_multiplier_A [55]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla2__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__57_  (.A(u_multiplier_B [55]),
    .B(u_multiplier_A [55]),
    .Z(u_multiplier_Final_add_cla2_cla2_cla1_cla2__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__58_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla2__36_ ),
    .B(u_multiplier_Final_add_cla2_cla2_cla1_cla2__39_ ),
    .ZN(product[55]));
 OAI21_X4 u_multiplier_Final_add_cla2_cla2_cla1_cla2__59_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla2__38_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla1_cla2__37_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla1_cla2__36_ ),
    .ZN(u_multiplier_Final_add_cla2_cla2_c1 ));
 AND2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__40_  (.A1(u_multiplier_B [56]),
    .A2(u_multiplier_A [56]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla1__25_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__41_  (.A1(u_multiplier_B [56]),
    .A2(u_multiplier_A [56]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla1__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__42_  (.A(u_multiplier_B [56]),
    .B(u_multiplier_A [56]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla1__27_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__43_  (.A(u_multiplier_Final_add_cla2_cla2_c1 ),
    .B(u_multiplier_Final_add_cla2_cla2_cla2_cla1__27_ ),
    .ZN(product[56]));
 AOI21_X2 u_multiplier_Final_add_cla2_cla2_cla2_cla1__44_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla1__25_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla2_cla1__26_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_c1 ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla1__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__45_  (.A1(u_multiplier_B [57]),
    .A2(u_multiplier_A [57]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla1__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__46_  (.A1(u_multiplier_B [57]),
    .A2(u_multiplier_A [57]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla1__30_ ));
 XOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__47_  (.A(u_multiplier_B [57]),
    .B(u_multiplier_A [57]),
    .Z(u_multiplier_Final_add_cla2_cla2_cla2_cla1__31_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__48_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla1__28_ ),
    .B(u_multiplier_Final_add_cla2_cla2_cla2_cla1__31_ ),
    .ZN(product[57]));
 OAI21_X2 u_multiplier_Final_add_cla2_cla2_cla2_cla1__49_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla1__30_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla2_cla1__29_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla2_cla1__28_ ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla1__32_ ));
 AND2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__50_  (.A1(u_multiplier_B [58]),
    .A2(u_multiplier_A [58]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla1__33_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__51_  (.A1(u_multiplier_B [58]),
    .A2(u_multiplier_A [58]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla1__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__52_  (.A(u_multiplier_B [58]),
    .B(u_multiplier_A [58]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla1__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__53_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla1__32_ ),
    .B(u_multiplier_Final_add_cla2_cla2_cla2_cla1__35_ ),
    .ZN(product[58]));
 AOI21_X2 u_multiplier_Final_add_cla2_cla2_cla2_cla1__54_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla1__33_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla2_cla1__34_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla2_cla1__32_ ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla1__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__55_  (.A1(u_multiplier_B [59]),
    .A2(u_multiplier_A [59]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla1__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__56_  (.A1(u_multiplier_B [59]),
    .A2(u_multiplier_A [59]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla1__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__57_  (.A(u_multiplier_B [59]),
    .B(u_multiplier_A [59]),
    .Z(u_multiplier_Final_add_cla2_cla2_cla2_cla1__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__58_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla1__36_ ),
    .B(u_multiplier_Final_add_cla2_cla2_cla2_cla1__39_ ),
    .ZN(product[59]));
 OAI21_X2 u_multiplier_Final_add_cla2_cla2_cla2_cla1__59_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla1__38_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla2_cla1__37_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla2_cla1__36_ ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_c1 ));
 AND2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__40_  (.A1(u_multiplier_B [60]),
    .A2(u_multiplier_A [60]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla2__25_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__41_  (.A1(u_multiplier_B [60]),
    .A2(u_multiplier_A [60]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla2__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__42_  (.A(u_multiplier_B [60]),
    .B(u_multiplier_A [60]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla2__27_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__43_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_c1 ),
    .B(u_multiplier_Final_add_cla2_cla2_cla2_cla2__27_ ),
    .ZN(product[60]));
 AOI21_X2 u_multiplier_Final_add_cla2_cla2_cla2_cla2__44_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla2__25_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla2_cla2__26_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla2_c1 ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla2__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__45_  (.A1(u_multiplier_B [61]),
    .A2(u_multiplier_A [61]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla2__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__46_  (.A1(u_multiplier_B [61]),
    .A2(u_multiplier_A [61]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla2__30_ ));
 XOR2_X2 u_multiplier_Final_add_cla2_cla2_cla2_cla2__47_  (.A(u_multiplier_B [61]),
    .B(u_multiplier_A [61]),
    .Z(u_multiplier_Final_add_cla2_cla2_cla2_cla2__31_ ));
 XNOR2_X2 u_multiplier_Final_add_cla2_cla2_cla2_cla2__48_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla2__28_ ),
    .B(u_multiplier_Final_add_cla2_cla2_cla2_cla2__31_ ),
    .ZN(product[61]));
 OAI21_X2 u_multiplier_Final_add_cla2_cla2_cla2_cla2__49_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla2__30_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla2_cla2__29_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla2_cla2__28_ ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla2__32_ ));
 AND2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__50_  (.A1(u_multiplier_B [62]),
    .A2(u_multiplier_pp3_62 ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla2__33_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__51_  (.A1(u_multiplier_B [62]),
    .A2(u_multiplier_pp3_62 ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla2__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__52_  (.A(u_multiplier_B [62]),
    .B(u_multiplier_pp3_62 ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla2__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__53_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla2__32_ ),
    .B(u_multiplier_Final_add_cla2_cla2_cla2_cla2__35_ ),
    .ZN(product[62]));
 AOI21_X4 u_multiplier_Final_add_cla2_cla2_cla2_cla2__54_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla2__33_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla2_cla2__34_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla2_cla2__32_ ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla2__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__55_  (.A1(net156),
    .A2(net140),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla2__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__56_  (.A1(net157),
    .A2(net141),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla2__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__57_  (.A(net158),
    .B(net142),
    .Z(u_multiplier_Final_add_cla2_cla2_cla2_cla2__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__58_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla2__36_ ),
    .B(u_multiplier_Final_add_cla2_cla2_cla2_cla2__39_ ),
    .ZN(product[63]));
 OAI21_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__59_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla2__38_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla2_cla2__37_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla2_cla2__36_ ),
    .ZN(u_multiplier_Final_add_Cout ));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_17_1__18_  (.A(net114),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_17_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_17_1__19_  (.A1(u_multiplier_STAGE1__0610_ ),
    .A2(u_multiplier_STAGE1__0609_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_17_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_17_1__20_  (.A(u_multiplier_STAGE1__0610_ ),
    .B(u_multiplier_STAGE1__0609_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_17_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_17_1__21_  (.A1(u_multiplier_STAGE1__0611_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_17_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_17_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_17_1__22_  (.A(u_multiplier_STAGE1__0611_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_17_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_17_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_17_1__23_  (.A1(u_multiplier_STAGE1__0612_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_17_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_17_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_17_1__24_  (.A(u_multiplier_STAGE1__0612_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_17_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_17_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_17_1__25_  (.A(net115),
    .B(u_multiplier_STAGE1_E_4_2_pp_17_1__16_ ),
    .ZN(u_multiplier_pp1_17 [0]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_17_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_17_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_17_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_17_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_17_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_17_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_17_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_17_1__17_ ),
    .ZN(u_multiplier_pp1_18 [2]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_18_1__18_  (.A(u_multiplier_STAGE1_pp1_17_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_18_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_18_1__19_  (.A1(u_multiplier_STAGE1__0614_ ),
    .A2(u_multiplier_STAGE1__0613_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_18_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_18_1__20_  (.A(u_multiplier_STAGE1__0614_ ),
    .B(u_multiplier_STAGE1__0613_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_18_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_18_1__21_  (.A1(u_multiplier_STAGE1__0615_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_18_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_18_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_18_1__22_  (.A(u_multiplier_STAGE1__0615_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_18_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_18_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_18_1__23_  (.A1(u_multiplier_STAGE1__0616_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_18_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_18_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_18_1__24_  (.A(u_multiplier_STAGE1__0616_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_18_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_18_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_18_1__25_  (.A(u_multiplier_STAGE1_pp1_17_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_18_1__16_ ),
    .ZN(u_multiplier_pp1_18 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_18_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_18_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_18_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_18_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_18_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_18_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_18_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_18_1__17_ ),
    .ZN(u_multiplier_pp1_19 [3]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_19_1__18_  (.A(u_multiplier_STAGE1_pp1_18_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_19_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_19_1__19_  (.A1(u_multiplier_STAGE1__0620_ ),
    .A2(u_multiplier_STAGE1__0619_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_19_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_19_1__20_  (.A(u_multiplier_STAGE1__0620_ ),
    .B(u_multiplier_STAGE1__0619_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_19_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_19_1__21_  (.A1(u_multiplier_STAGE1__0621_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_19_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_19_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_19_1__22_  (.A(u_multiplier_STAGE1__0621_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_19_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_19_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_19_1__23_  (.A1(u_multiplier_STAGE1__0622_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_19_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_19_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_19_1__24_  (.A(u_multiplier_STAGE1__0622_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_19_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_19_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_19_1__25_  (.A(u_multiplier_STAGE1_pp1_18_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_19_1__16_ ),
    .ZN(u_multiplier_pp1_19 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_19_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_19_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_19_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_19_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_19_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_19_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_19_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_19_1__17_ ),
    .ZN(u_multiplier_pp1_20 [4]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_19_2__18_  (.A(net116),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_19_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_19_2__19_  (.A1(u_multiplier_STAGE1__0624_ ),
    .A2(u_multiplier_STAGE1__0623_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_19_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_19_2__20_  (.A(u_multiplier_STAGE1__0624_ ),
    .B(u_multiplier_STAGE1__0623_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_19_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_19_2__21_  (.A1(u_multiplier_STAGE1__0625_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_19_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_19_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_19_2__22_  (.A(u_multiplier_STAGE1__0625_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_19_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_19_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_19_2__23_  (.A1(u_multiplier_STAGE1__0626_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_19_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_19_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_19_2__24_  (.A(u_multiplier_STAGE1__0626_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_19_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_19_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_19_2__25_  (.A(net117),
    .B(u_multiplier_STAGE1_E_4_2_pp_19_2__16_ ),
    .ZN(u_multiplier_pp1_19 [0]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_19_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_19_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_19_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_19_e42_2_cout ));
 OAI21_X1 u_multiplier_STAGE1_E_4_2_pp_19_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_19_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_19_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_19_2__17_ ),
    .ZN(u_multiplier_pp1_20 [3]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_20_1__18_  (.A(u_multiplier_STAGE1_pp1_19_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_20_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_20_1__19_  (.A1(u_multiplier_STAGE1__0628_ ),
    .A2(u_multiplier_STAGE1__0627_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_20_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_20_1__20_  (.A(u_multiplier_STAGE1__0628_ ),
    .B(u_multiplier_STAGE1__0627_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_20_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_20_1__21_  (.A1(u_multiplier_STAGE1__0629_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_20_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_20_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_20_1__22_  (.A(u_multiplier_STAGE1__0629_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_20_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_20_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_20_1__23_  (.A1(u_multiplier_STAGE1__0630_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_20_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_20_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_20_1__24_  (.A(u_multiplier_STAGE1__0630_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_20_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_20_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_20_1__25_  (.A(u_multiplier_STAGE1_pp1_19_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_20_1__16_ ),
    .ZN(u_multiplier_pp1_20 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_20_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_20_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_20_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_20_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_20_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_20_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_20_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_20_1__17_ ),
    .ZN(u_multiplier_pp1_21 [5]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_20_2__18_  (.A(u_multiplier_STAGE1_pp1_19_e42_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_20_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_20_2__19_  (.A1(u_multiplier_STAGE1__0632_ ),
    .A2(u_multiplier_STAGE1__0631_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_20_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_20_2__20_  (.A(u_multiplier_STAGE1__0632_ ),
    .B(u_multiplier_STAGE1__0631_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_20_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_20_2__21_  (.A1(u_multiplier_STAGE1__0633_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_20_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_20_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_20_2__22_  (.A(u_multiplier_STAGE1__0633_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_20_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_20_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_20_2__23_  (.A1(u_multiplier_STAGE1__0634_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_20_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_20_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_20_2__24_  (.A(u_multiplier_STAGE1__0634_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_20_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_20_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_20_2__25_  (.A(u_multiplier_STAGE1_pp1_19_e42_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_20_2__16_ ),
    .ZN(u_multiplier_pp1_20 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_20_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_20_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_20_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_20_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_20_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_20_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_20_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_20_2__17_ ),
    .ZN(u_multiplier_pp1_21 [4]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_21_1__18_  (.A(u_multiplier_STAGE1_pp1_20_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_21_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_21_1__19_  (.A1(u_multiplier_STAGE1__0638_ ),
    .A2(u_multiplier_STAGE1__0637_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_21_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_21_1__20_  (.A(u_multiplier_STAGE1__0638_ ),
    .B(u_multiplier_STAGE1__0637_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_21_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_21_1__21_  (.A1(u_multiplier_STAGE1__0639_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_21_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_21_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_21_1__22_  (.A(u_multiplier_STAGE1__0639_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_21_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_21_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_21_1__23_  (.A1(u_multiplier_STAGE1__0640_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_21_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_21_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_21_1__24_  (.A(u_multiplier_STAGE1__0640_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_21_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_21_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_21_1__25_  (.A(u_multiplier_STAGE1_pp1_20_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_21_1__16_ ),
    .ZN(u_multiplier_pp1_21 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_21_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_21_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_21_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_21_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_21_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_21_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_21_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_21_1__17_ ),
    .ZN(u_multiplier_pp1_22 [6]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_21_2__18_  (.A(u_multiplier_STAGE1_pp1_20_e42_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_21_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_21_2__19_  (.A1(u_multiplier_STAGE1__0642_ ),
    .A2(u_multiplier_STAGE1__0641_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_21_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_21_2__20_  (.A(u_multiplier_STAGE1__0642_ ),
    .B(u_multiplier_STAGE1__0641_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_21_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_21_2__21_  (.A1(u_multiplier_STAGE1__0643_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_21_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_21_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_21_2__22_  (.A(u_multiplier_STAGE1__0643_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_21_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_21_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_21_2__23_  (.A1(u_multiplier_STAGE1__0644_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_21_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_21_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_21_2__24_  (.A(u_multiplier_STAGE1__0644_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_21_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_21_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_21_2__25_  (.A(u_multiplier_STAGE1_pp1_20_e42_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_21_2__16_ ),
    .ZN(u_multiplier_pp1_21 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_21_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_21_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_21_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_21_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_21_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_21_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_21_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_21_2__17_ ),
    .ZN(u_multiplier_pp1_22 [5]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_21_3__18_  (.A(net118),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_21_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_21_3__19_  (.A1(u_multiplier_STAGE1__0646_ ),
    .A2(u_multiplier_STAGE1__0645_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_21_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_21_3__20_  (.A(u_multiplier_STAGE1__0646_ ),
    .B(u_multiplier_STAGE1__0645_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_21_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_21_3__21_  (.A1(u_multiplier_STAGE1__0647_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_21_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_21_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_21_3__22_  (.A(u_multiplier_STAGE1__0647_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_21_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_21_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_21_3__23_  (.A1(u_multiplier_STAGE1__0648_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_21_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_21_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_21_3__24_  (.A(u_multiplier_STAGE1__0648_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_21_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_21_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_21_3__25_  (.A(net119),
    .B(u_multiplier_STAGE1_E_4_2_pp_21_3__16_ ),
    .ZN(u_multiplier_pp1_21 [0]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_21_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_21_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_21_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_21_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_21_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_21_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_21_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_21_3__17_ ),
    .ZN(u_multiplier_pp1_22 [4]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_22_1__18_  (.A(u_multiplier_STAGE1_pp1_21_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_22_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_22_1__19_  (.A1(u_multiplier_STAGE1__0650_ ),
    .A2(u_multiplier_STAGE1__0649_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_22_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_22_1__20_  (.A(u_multiplier_STAGE1__0650_ ),
    .B(u_multiplier_STAGE1__0649_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_22_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_22_1__21_  (.A1(u_multiplier_STAGE1__0651_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_22_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_22_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_22_1__22_  (.A(u_multiplier_STAGE1__0651_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_22_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_22_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_22_1__23_  (.A1(u_multiplier_STAGE1__0652_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_22_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_22_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_22_1__24_  (.A(u_multiplier_STAGE1__0652_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_22_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_22_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_22_1__25_  (.A(u_multiplier_STAGE1_pp1_21_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_22_1__16_ ),
    .ZN(u_multiplier_pp1_22 [3]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_22_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_22_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_22_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_22_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_22_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_22_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_22_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_22_1__17_ ),
    .ZN(u_multiplier_pp1_23 [7]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_22_2__18_  (.A(u_multiplier_STAGE1_pp1_21_e42_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_22_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_22_2__19_  (.A1(u_multiplier_STAGE1__0654_ ),
    .A2(u_multiplier_STAGE1__0653_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_22_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_22_2__20_  (.A(u_multiplier_STAGE1__0654_ ),
    .B(u_multiplier_STAGE1__0653_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_22_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_22_2__21_  (.A1(u_multiplier_STAGE1__0655_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_22_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_22_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_22_2__22_  (.A(u_multiplier_STAGE1__0655_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_22_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_22_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_22_2__23_  (.A1(u_multiplier_STAGE1__0656_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_22_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_22_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_22_2__24_  (.A(u_multiplier_STAGE1__0656_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_22_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_22_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_22_2__25_  (.A(u_multiplier_STAGE1_pp1_21_e42_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_22_2__16_ ),
    .ZN(u_multiplier_pp1_22 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_22_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_22_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_22_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_22_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_22_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_22_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_22_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_22_2__17_ ),
    .ZN(u_multiplier_pp1_23 [6]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_22_3__18_  (.A(u_multiplier_STAGE1_pp1_21_e42_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_22_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_22_3__19_  (.A1(u_multiplier_STAGE1__0658_ ),
    .A2(u_multiplier_STAGE1__0657_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_22_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_22_3__20_  (.A(u_multiplier_STAGE1__0658_ ),
    .B(u_multiplier_STAGE1__0657_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_22_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_22_3__21_  (.A1(u_multiplier_STAGE1__0659_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_22_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_22_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_22_3__22_  (.A(u_multiplier_STAGE1__0659_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_22_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_22_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_22_3__23_  (.A1(u_multiplier_STAGE1__0660_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_22_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_22_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_22_3__24_  (.A(u_multiplier_STAGE1__0660_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_22_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_22_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_22_3__25_  (.A(u_multiplier_STAGE1_pp1_21_e42_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_22_3__16_ ),
    .ZN(u_multiplier_pp1_22 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_22_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_22_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_22_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_22_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_22_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_22_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_22_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_22_3__17_ ),
    .ZN(u_multiplier_pp1_23 [5]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_23_1__18_  (.A(u_multiplier_STAGE1_pp1_22_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_23_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_23_1__19_  (.A1(u_multiplier_STAGE1__0664_ ),
    .A2(u_multiplier_STAGE1__0663_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_23_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_23_1__20_  (.A(u_multiplier_STAGE1__0664_ ),
    .B(u_multiplier_STAGE1__0663_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_23_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_23_1__21_  (.A1(u_multiplier_STAGE1__0665_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_23_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_23_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_23_1__22_  (.A(u_multiplier_STAGE1__0665_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_23_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_23_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_23_1__23_  (.A1(u_multiplier_STAGE1__0666_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_23_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_23_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_23_1__24_  (.A(u_multiplier_STAGE1__0666_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_23_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_23_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_23_1__25_  (.A(u_multiplier_STAGE1_pp1_22_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_23_1__16_ ),
    .ZN(u_multiplier_pp1_23 [3]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_23_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_23_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_23_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_23_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_23_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_23_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_23_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_23_1__17_ ),
    .ZN(u_multiplier_pp1_24 [8]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_23_2__18_  (.A(u_multiplier_STAGE1_pp1_22_e42_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_23_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_23_2__19_  (.A1(u_multiplier_STAGE1__0668_ ),
    .A2(u_multiplier_STAGE1__0667_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_23_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_23_2__20_  (.A(u_multiplier_STAGE1__0668_ ),
    .B(u_multiplier_STAGE1__0667_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_23_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_23_2__21_  (.A1(u_multiplier_STAGE1__0669_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_23_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_23_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_23_2__22_  (.A(u_multiplier_STAGE1__0669_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_23_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_23_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_23_2__23_  (.A1(u_multiplier_STAGE1__0670_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_23_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_23_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_23_2__24_  (.A(u_multiplier_STAGE1__0670_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_23_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_23_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_23_2__25_  (.A(u_multiplier_STAGE1_pp1_22_e42_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_23_2__16_ ),
    .ZN(u_multiplier_pp1_23 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_23_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_23_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_23_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_23_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_23_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_23_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_23_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_23_2__17_ ),
    .ZN(u_multiplier_pp1_24 [7]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_23_3__18_  (.A(u_multiplier_STAGE1_pp1_22_e42_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_23_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_23_3__19_  (.A1(u_multiplier_STAGE1__0672_ ),
    .A2(u_multiplier_STAGE1__0671_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_23_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_23_3__20_  (.A(u_multiplier_STAGE1__0672_ ),
    .B(u_multiplier_STAGE1__0671_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_23_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_23_3__21_  (.A1(u_multiplier_STAGE1__0673_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_23_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_23_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_23_3__22_  (.A(u_multiplier_STAGE1__0673_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_23_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_23_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_23_3__23_  (.A1(u_multiplier_STAGE1__0674_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_23_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_23_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_23_3__24_  (.A(u_multiplier_STAGE1__0674_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_23_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_23_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_23_3__25_  (.A(u_multiplier_STAGE1_pp1_22_e42_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_23_3__16_ ),
    .ZN(u_multiplier_pp1_23 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_23_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_23_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_23_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_23_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_23_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_23_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_23_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_23_3__17_ ),
    .ZN(u_multiplier_pp1_24 [6]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_23_4__18_  (.A(net120),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_23_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_23_4__19_  (.A1(u_multiplier_STAGE1__0676_ ),
    .A2(u_multiplier_STAGE1__0675_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_23_4__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_23_4__20_  (.A(u_multiplier_STAGE1__0676_ ),
    .B(u_multiplier_STAGE1__0675_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_23_4__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_23_4__21_  (.A1(u_multiplier_STAGE1__0677_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_23_4__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_23_4__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_23_4__22_  (.A(u_multiplier_STAGE1__0677_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_23_4__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_23_4__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_23_4__23_  (.A1(u_multiplier_STAGE1__0678_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_23_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_23_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_23_4__24_  (.A(u_multiplier_STAGE1__0678_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_23_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_23_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_23_4__25_  (.A(net121),
    .B(u_multiplier_STAGE1_E_4_2_pp_23_4__16_ ),
    .ZN(u_multiplier_pp1_23 [0]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_23_4__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_23_4__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_23_4__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_23_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_23_4__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_23_4__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_23_4__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_23_4__17_ ),
    .ZN(u_multiplier_pp1_24 [5]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_24_1__18_  (.A(u_multiplier_STAGE1_pp1_23_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_24_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_24_1__19_  (.A1(u_multiplier_STAGE1__0680_ ),
    .A2(u_multiplier_STAGE1__0679_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_24_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_24_1__20_  (.A(u_multiplier_STAGE1__0680_ ),
    .B(u_multiplier_STAGE1__0679_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_24_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_24_1__21_  (.A1(u_multiplier_STAGE1__0681_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_24_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_24_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_24_1__22_  (.A(u_multiplier_STAGE1__0681_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_24_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_24_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_24_1__23_  (.A1(u_multiplier_STAGE1__0682_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_24_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_24_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_24_1__24_  (.A(u_multiplier_STAGE1__0682_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_24_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_24_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_24_1__25_  (.A(u_multiplier_STAGE1_pp1_23_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_24_1__16_ ),
    .ZN(u_multiplier_pp1_24 [4]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_24_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_24_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_24_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_24_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_24_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_24_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_24_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_24_1__17_ ),
    .ZN(u_multiplier_pp1_25 [9]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_24_2__18_  (.A(u_multiplier_STAGE1_pp1_23_e42_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_24_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_24_2__19_  (.A1(u_multiplier_STAGE1__0684_ ),
    .A2(u_multiplier_STAGE1__0683_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_24_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_24_2__20_  (.A(u_multiplier_STAGE1__0684_ ),
    .B(u_multiplier_STAGE1__0683_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_24_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_24_2__21_  (.A1(u_multiplier_STAGE1__0685_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_24_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_24_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_24_2__22_  (.A(u_multiplier_STAGE1__0685_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_24_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_24_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_24_2__23_  (.A1(u_multiplier_STAGE1__0686_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_24_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_24_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_24_2__24_  (.A(u_multiplier_STAGE1__0686_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_24_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_24_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_24_2__25_  (.A(u_multiplier_STAGE1_pp1_23_e42_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_24_2__16_ ),
    .ZN(u_multiplier_pp1_24 [3]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_24_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_24_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_24_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_24_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_24_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_24_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_24_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_24_2__17_ ),
    .ZN(u_multiplier_pp1_25 [8]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_24_3__18_  (.A(u_multiplier_STAGE1_pp1_23_e42_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_24_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_24_3__19_  (.A1(u_multiplier_STAGE1__0688_ ),
    .A2(u_multiplier_STAGE1__0687_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_24_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_24_3__20_  (.A(u_multiplier_STAGE1__0688_ ),
    .B(u_multiplier_STAGE1__0687_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_24_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_24_3__21_  (.A1(u_multiplier_STAGE1__0689_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_24_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_24_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_24_3__22_  (.A(u_multiplier_STAGE1__0689_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_24_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_24_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_24_3__23_  (.A1(u_multiplier_STAGE1__0690_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_24_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_24_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_24_3__24_  (.A(u_multiplier_STAGE1__0690_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_24_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_24_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_24_3__25_  (.A(u_multiplier_STAGE1_pp1_23_e42_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_24_3__16_ ),
    .ZN(u_multiplier_pp1_24 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_24_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_24_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_24_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_24_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_24_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_24_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_24_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_24_3__17_ ),
    .ZN(u_multiplier_pp1_25 [7]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_24_4__18_  (.A(u_multiplier_STAGE1_pp1_23_e42_4_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_24_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_24_4__19_  (.A1(u_multiplier_STAGE1__0692_ ),
    .A2(u_multiplier_STAGE1__0691_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_24_4__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_24_4__20_  (.A(u_multiplier_STAGE1__0692_ ),
    .B(u_multiplier_STAGE1__0691_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_24_4__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_24_4__21_  (.A1(u_multiplier_STAGE1__0693_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_24_4__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_24_4__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_24_4__22_  (.A(u_multiplier_STAGE1__0693_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_24_4__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_24_4__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_24_4__23_  (.A1(u_multiplier_STAGE1__0694_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_24_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_24_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_24_4__24_  (.A(u_multiplier_STAGE1__0694_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_24_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_24_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_24_4__25_  (.A(u_multiplier_STAGE1_pp1_23_e42_4_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_24_4__16_ ),
    .ZN(u_multiplier_pp1_24 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_24_4__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_24_4__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_24_4__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_24_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_24_4__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_24_4__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_24_4__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_24_4__17_ ),
    .ZN(u_multiplier_pp1_25 [6]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_25_1__18_  (.A(u_multiplier_STAGE1_pp1_24_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_25_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_25_1__19_  (.A1(u_multiplier_STAGE1__0698_ ),
    .A2(u_multiplier_STAGE1__0697_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_25_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_25_1__20_  (.A(u_multiplier_STAGE1__0698_ ),
    .B(u_multiplier_STAGE1__0697_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_25_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_25_1__21_  (.A1(u_multiplier_STAGE1__0699_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_25_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_25_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_25_1__22_  (.A(u_multiplier_STAGE1__0699_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_25_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_25_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_25_1__23_  (.A1(u_multiplier_STAGE1__0700_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_25_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_25_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_25_1__24_  (.A(u_multiplier_STAGE1__0700_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_25_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_25_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_25_1__25_  (.A(u_multiplier_STAGE1_pp1_24_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_25_1__16_ ),
    .ZN(u_multiplier_pp1_25 [4]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_25_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_25_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_25_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_25_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_25_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_25_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_25_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_25_1__17_ ),
    .ZN(u_multiplier_pp1_26 [10]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_25_2__18_  (.A(u_multiplier_STAGE1_pp1_24_e42_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_25_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_25_2__19_  (.A1(u_multiplier_STAGE1__0702_ ),
    .A2(u_multiplier_STAGE1__0701_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_25_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_25_2__20_  (.A(u_multiplier_STAGE1__0702_ ),
    .B(u_multiplier_STAGE1__0701_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_25_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_25_2__21_  (.A1(u_multiplier_STAGE1__0703_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_25_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_25_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_25_2__22_  (.A(u_multiplier_STAGE1__0703_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_25_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_25_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_25_2__23_  (.A1(u_multiplier_STAGE1__0704_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_25_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_25_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_25_2__24_  (.A(u_multiplier_STAGE1__0704_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_25_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_25_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_25_2__25_  (.A(u_multiplier_STAGE1_pp1_24_e42_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_25_2__16_ ),
    .ZN(u_multiplier_pp1_25 [3]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_25_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_25_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_25_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_25_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_25_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_25_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_25_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_25_2__17_ ),
    .ZN(u_multiplier_pp1_26 [9]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_25_3__18_  (.A(u_multiplier_STAGE1_pp1_24_e42_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_25_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_25_3__19_  (.A1(u_multiplier_STAGE1__0706_ ),
    .A2(u_multiplier_STAGE1__0705_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_25_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_25_3__20_  (.A(u_multiplier_STAGE1__0706_ ),
    .B(u_multiplier_STAGE1__0705_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_25_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_25_3__21_  (.A1(u_multiplier_STAGE1__0707_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_25_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_25_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_25_3__22_  (.A(u_multiplier_STAGE1__0707_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_25_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_25_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_25_3__23_  (.A1(u_multiplier_STAGE1__0708_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_25_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_25_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_25_3__24_  (.A(u_multiplier_STAGE1__0708_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_25_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_25_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_25_3__25_  (.A(u_multiplier_STAGE1_pp1_24_e42_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_25_3__16_ ),
    .ZN(u_multiplier_pp1_25 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_25_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_25_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_25_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_25_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_25_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_25_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_25_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_25_3__17_ ),
    .ZN(u_multiplier_pp1_26 [8]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_25_4__18_  (.A(u_multiplier_STAGE1_pp1_24_e42_4_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_25_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_25_4__19_  (.A1(u_multiplier_STAGE1__0710_ ),
    .A2(u_multiplier_STAGE1__0709_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_25_4__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_25_4__20_  (.A(u_multiplier_STAGE1__0710_ ),
    .B(u_multiplier_STAGE1__0709_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_25_4__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_25_4__21_  (.A1(u_multiplier_STAGE1__0711_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_25_4__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_25_4__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_25_4__22_  (.A(u_multiplier_STAGE1__0711_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_25_4__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_25_4__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_25_4__23_  (.A1(u_multiplier_STAGE1__0712_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_25_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_25_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_25_4__24_  (.A(u_multiplier_STAGE1__0712_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_25_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_25_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_25_4__25_  (.A(u_multiplier_STAGE1_pp1_24_e42_4_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_25_4__16_ ),
    .ZN(u_multiplier_pp1_25 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_25_4__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_25_4__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_25_4__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_25_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_25_4__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_25_4__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_25_4__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_25_4__17_ ),
    .ZN(u_multiplier_pp1_26 [7]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_25_5__18_  (.A(net122),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_25_5__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_25_5__19_  (.A1(u_multiplier_STAGE1__0714_ ),
    .A2(u_multiplier_STAGE1__0713_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_25_5__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_25_5__20_  (.A(u_multiplier_STAGE1__0714_ ),
    .B(u_multiplier_STAGE1__0713_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_25_5__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_25_5__21_  (.A1(u_multiplier_STAGE1__0715_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_25_5__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_25_5__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_25_5__22_  (.A(u_multiplier_STAGE1__0715_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_25_5__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_25_5__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_25_5__23_  (.A1(u_multiplier_STAGE1__0716_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_25_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_25_5__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_25_5__24_  (.A(u_multiplier_STAGE1__0716_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_25_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_25_5__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_25_5__25_  (.A(net123),
    .B(u_multiplier_STAGE1_E_4_2_pp_25_5__16_ ),
    .ZN(u_multiplier_pp1_25 [0]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_25_5__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_25_5__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_25_5__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_25_e42_5_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_25_5__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_25_5__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_25_5__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_25_5__17_ ),
    .ZN(u_multiplier_pp1_26 [6]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_26_1__18_  (.A(u_multiplier_STAGE1_pp1_25_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_26_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_26_1__19_  (.A1(u_multiplier_STAGE1__0718_ ),
    .A2(u_multiplier_STAGE1__0717_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_26_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_26_1__20_  (.A(u_multiplier_STAGE1__0718_ ),
    .B(u_multiplier_STAGE1__0717_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_26_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_26_1__21_  (.A1(u_multiplier_STAGE1__0719_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_26_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_26_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_26_1__22_  (.A(u_multiplier_STAGE1__0719_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_26_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_26_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_26_1__23_  (.A1(u_multiplier_STAGE1__0720_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_26_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_26_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_26_1__24_  (.A(u_multiplier_STAGE1__0720_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_26_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_26_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_26_1__25_  (.A(u_multiplier_STAGE1_pp1_25_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_26_1__16_ ),
    .ZN(u_multiplier_pp1_26 [5]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_26_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_26_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_26_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_26_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE1_E_4_2_pp_26_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_26_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_26_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_26_1__17_ ),
    .ZN(u_multiplier_pp1_27 [11]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_26_2__18_  (.A(u_multiplier_STAGE1_pp1_25_e42_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_26_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_26_2__19_  (.A1(u_multiplier_STAGE1__0722_ ),
    .A2(u_multiplier_STAGE1__0721_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_26_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_26_2__20_  (.A(u_multiplier_STAGE1__0722_ ),
    .B(u_multiplier_STAGE1__0721_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_26_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_26_2__21_  (.A1(u_multiplier_STAGE1__0723_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_26_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_26_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_26_2__22_  (.A(u_multiplier_STAGE1__0723_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_26_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_26_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_26_2__23_  (.A1(u_multiplier_STAGE1__0724_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_26_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_26_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_26_2__24_  (.A(u_multiplier_STAGE1__0724_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_26_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_26_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_26_2__25_  (.A(u_multiplier_STAGE1_pp1_25_e42_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_26_2__16_ ),
    .ZN(u_multiplier_pp1_26 [4]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_26_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_26_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_26_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_26_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_26_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_26_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_26_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_26_2__17_ ),
    .ZN(u_multiplier_pp1_27 [10]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_26_3__18_  (.A(u_multiplier_STAGE1_pp1_25_e42_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_26_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_26_3__19_  (.A1(u_multiplier_STAGE1__0726_ ),
    .A2(u_multiplier_STAGE1__0725_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_26_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_26_3__20_  (.A(u_multiplier_STAGE1__0726_ ),
    .B(u_multiplier_STAGE1__0725_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_26_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_26_3__21_  (.A1(u_multiplier_STAGE1__0727_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_26_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_26_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_26_3__22_  (.A(u_multiplier_STAGE1__0727_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_26_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_26_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_26_3__23_  (.A1(u_multiplier_STAGE1__0728_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_26_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_26_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_26_3__24_  (.A(u_multiplier_STAGE1__0728_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_26_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_26_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_26_3__25_  (.A(u_multiplier_STAGE1_pp1_25_e42_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_26_3__16_ ),
    .ZN(u_multiplier_pp1_26 [3]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_26_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_26_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_26_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_26_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_26_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_26_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_26_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_26_3__17_ ),
    .ZN(u_multiplier_pp1_27 [9]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_26_4__18_  (.A(u_multiplier_STAGE1_pp1_25_e42_4_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_26_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_26_4__19_  (.A1(u_multiplier_STAGE1__0730_ ),
    .A2(u_multiplier_STAGE1__0729_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_26_4__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_26_4__20_  (.A(u_multiplier_STAGE1__0730_ ),
    .B(u_multiplier_STAGE1__0729_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_26_4__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_26_4__21_  (.A1(u_multiplier_STAGE1__0731_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_26_4__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_26_4__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_26_4__22_  (.A(u_multiplier_STAGE1__0731_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_26_4__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_26_4__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_26_4__23_  (.A1(u_multiplier_STAGE1__0732_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_26_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_26_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_26_4__24_  (.A(u_multiplier_STAGE1__0732_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_26_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_26_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_26_4__25_  (.A(u_multiplier_STAGE1_pp1_25_e42_4_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_26_4__16_ ),
    .ZN(u_multiplier_pp1_26 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_26_4__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_26_4__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_26_4__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_26_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_26_4__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_26_4__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_26_4__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_26_4__17_ ),
    .ZN(u_multiplier_pp1_27 [8]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_26_5__18_  (.A(u_multiplier_STAGE1_pp1_25_e42_5_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_26_5__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_26_5__19_  (.A1(u_multiplier_STAGE1__0734_ ),
    .A2(u_multiplier_STAGE1__0733_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_26_5__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_26_5__20_  (.A(u_multiplier_STAGE1__0734_ ),
    .B(u_multiplier_STAGE1__0733_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_26_5__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_26_5__21_  (.A1(u_multiplier_STAGE1__0735_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_26_5__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_26_5__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_26_5__22_  (.A(u_multiplier_STAGE1__0735_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_26_5__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_26_5__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_26_5__23_  (.A1(u_multiplier_STAGE1__0736_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_26_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_26_5__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_26_5__24_  (.A(u_multiplier_STAGE1__0736_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_26_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_26_5__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_26_5__25_  (.A(u_multiplier_STAGE1_pp1_25_e42_5_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_26_5__16_ ),
    .ZN(u_multiplier_pp1_26 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_26_5__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_26_5__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_26_5__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_26_e42_5_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_26_5__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_26_5__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_26_5__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_26_5__17_ ),
    .ZN(u_multiplier_pp1_27 [7]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_27_1__18_  (.A(u_multiplier_STAGE1_pp1_26_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_27_1__19_  (.A1(u_multiplier_STAGE1__0740_ ),
    .A2(u_multiplier_STAGE1__0739_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_27_1__20_  (.A(u_multiplier_STAGE1__0740_ ),
    .B(u_multiplier_STAGE1__0739_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_27_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_27_1__21_  (.A1(u_multiplier_STAGE1__0741_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_27_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_27_1__22_  (.A(u_multiplier_STAGE1__0741_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_27_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_27_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_27_1__23_  (.A1(u_multiplier_STAGE1__0742_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_27_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_27_1__24_  (.A(u_multiplier_STAGE1__0742_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_27_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_27_1__25_  (.A(u_multiplier_STAGE1_pp1_26_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_27_1__16_ ),
    .ZN(u_multiplier_pp1_27 [5]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_27_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_27_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_27_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_27_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_27_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_27_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_27_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_27_1__17_ ),
    .ZN(u_multiplier_pp1_28 [12]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_27_2__18_  (.A(u_multiplier_STAGE1_pp1_26_e42_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_27_2__19_  (.A1(u_multiplier_STAGE1__0744_ ),
    .A2(u_multiplier_STAGE1__0743_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_27_2__20_  (.A(u_multiplier_STAGE1__0744_ ),
    .B(u_multiplier_STAGE1__0743_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_27_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_27_2__21_  (.A1(u_multiplier_STAGE1__0745_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_27_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_27_2__22_  (.A(u_multiplier_STAGE1__0745_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_27_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_27_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_27_2__23_  (.A1(u_multiplier_STAGE1__0746_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_27_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_27_2__24_  (.A(u_multiplier_STAGE1__0746_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_27_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_27_2__25_  (.A(u_multiplier_STAGE1_pp1_26_e42_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_27_2__16_ ),
    .ZN(u_multiplier_pp1_27 [4]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_27_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_27_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_27_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_27_e42_2_cout ));
 OAI21_X1 u_multiplier_STAGE1_E_4_2_pp_27_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_27_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_27_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_27_2__17_ ),
    .ZN(u_multiplier_pp1_28 [11]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_27_3__18_  (.A(u_multiplier_STAGE1_pp1_26_e42_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_27_3__19_  (.A1(u_multiplier_STAGE1__0748_ ),
    .A2(u_multiplier_STAGE1__0747_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_27_3__20_  (.A(u_multiplier_STAGE1__0748_ ),
    .B(u_multiplier_STAGE1__0747_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_27_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_27_3__21_  (.A1(u_multiplier_STAGE1__0749_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_27_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_27_3__22_  (.A(u_multiplier_STAGE1__0749_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_27_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_27_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_27_3__23_  (.A1(u_multiplier_STAGE1__0750_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_27_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_27_3__24_  (.A(u_multiplier_STAGE1__0750_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_27_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_27_3__25_  (.A(u_multiplier_STAGE1_pp1_26_e42_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_27_3__16_ ),
    .ZN(u_multiplier_pp1_27 [3]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_27_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_27_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_27_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_27_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_27_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_27_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_27_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_27_3__17_ ),
    .ZN(u_multiplier_pp1_28 [10]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_27_4__18_  (.A(u_multiplier_STAGE1_pp1_26_e42_4_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_27_4__19_  (.A1(u_multiplier_STAGE1__0752_ ),
    .A2(u_multiplier_STAGE1__0751_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_4__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_27_4__20_  (.A(u_multiplier_STAGE1__0752_ ),
    .B(u_multiplier_STAGE1__0751_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_27_4__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_27_4__21_  (.A1(u_multiplier_STAGE1__0753_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_27_4__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_4__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_27_4__22_  (.A(u_multiplier_STAGE1__0753_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_27_4__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_27_4__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_27_4__23_  (.A1(u_multiplier_STAGE1__0754_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_27_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_27_4__24_  (.A(u_multiplier_STAGE1__0754_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_27_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_27_4__25_  (.A(u_multiplier_STAGE1_pp1_26_e42_4_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_27_4__16_ ),
    .ZN(u_multiplier_pp1_27 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_27_4__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_27_4__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_27_4__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_27_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_27_4__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_27_4__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_27_4__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_27_4__17_ ),
    .ZN(u_multiplier_pp1_28 [9]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_27_5__18_  (.A(u_multiplier_STAGE1_pp1_26_e42_5_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_5__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_27_5__19_  (.A1(u_multiplier_STAGE1__0756_ ),
    .A2(u_multiplier_STAGE1__0755_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_5__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_27_5__20_  (.A(u_multiplier_STAGE1__0756_ ),
    .B(u_multiplier_STAGE1__0755_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_27_5__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_27_5__21_  (.A1(u_multiplier_STAGE1__0757_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_27_5__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_5__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_27_5__22_  (.A(u_multiplier_STAGE1__0757_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_27_5__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_27_5__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_27_5__23_  (.A1(u_multiplier_STAGE1__0758_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_27_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_5__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_27_5__24_  (.A(u_multiplier_STAGE1__0758_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_27_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_5__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_27_5__25_  (.A(u_multiplier_STAGE1_pp1_26_e42_5_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_27_5__16_ ),
    .ZN(u_multiplier_pp1_27 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_27_5__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_27_5__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_27_5__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_27_e42_5_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_27_5__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_27_5__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_27_5__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_27_5__17_ ),
    .ZN(u_multiplier_pp1_28 [8]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_27_6__18_  (.A(net124),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_6__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_27_6__19_  (.A1(u_multiplier_STAGE1__0760_ ),
    .A2(u_multiplier_STAGE1__0759_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_6__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_27_6__20_  (.A(u_multiplier_STAGE1__0760_ ),
    .B(u_multiplier_STAGE1__0759_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_27_6__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_27_6__21_  (.A1(u_multiplier_STAGE1__0761_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_27_6__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_6__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_27_6__22_  (.A(u_multiplier_STAGE1__0761_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_27_6__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_27_6__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_27_6__23_  (.A1(u_multiplier_STAGE1__0762_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_27_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_6__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_27_6__24_  (.A(u_multiplier_STAGE1__0762_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_27_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_27_6__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_27_6__25_  (.A(net125),
    .B(u_multiplier_STAGE1_E_4_2_pp_27_6__16_ ),
    .ZN(u_multiplier_pp1_27 [0]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_27_6__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_27_6__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_27_6__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_27_e42_6_cout ));
 OAI21_X1 u_multiplier_STAGE1_E_4_2_pp_27_6__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_27_6__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_27_6__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_27_6__17_ ),
    .ZN(u_multiplier_pp1_28 [7]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_28_1__18_  (.A(u_multiplier_STAGE1_pp1_27_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_28_1__19_  (.A1(u_multiplier_STAGE1__0764_ ),
    .A2(u_multiplier_STAGE1__0763_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_28_1__20_  (.A(u_multiplier_STAGE1__0764_ ),
    .B(u_multiplier_STAGE1__0763_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_28_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_28_1__21_  (.A1(u_multiplier_STAGE1__0765_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_28_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_28_1__22_  (.A(u_multiplier_STAGE1__0765_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_28_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_28_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_28_1__23_  (.A1(u_multiplier_STAGE1__0766_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_28_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_28_1__24_  (.A(u_multiplier_STAGE1__0766_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_28_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_28_1__25_  (.A(u_multiplier_STAGE1_pp1_27_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_28_1__16_ ),
    .ZN(u_multiplier_pp1_28 [6]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_28_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_28_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_28_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_28_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_28_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_28_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_28_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_28_1__17_ ),
    .ZN(u_multiplier_pp1_29 [13]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_28_2__18_  (.A(u_multiplier_STAGE1_pp1_27_e42_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_28_2__19_  (.A1(u_multiplier_STAGE1__0768_ ),
    .A2(u_multiplier_STAGE1__0767_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_28_2__20_  (.A(u_multiplier_STAGE1__0768_ ),
    .B(u_multiplier_STAGE1__0767_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_28_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_28_2__21_  (.A1(u_multiplier_STAGE1__0769_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_28_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_28_2__22_  (.A(u_multiplier_STAGE1__0769_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_28_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_28_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_28_2__23_  (.A1(u_multiplier_STAGE1__0770_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_28_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_28_2__24_  (.A(u_multiplier_STAGE1__0770_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_28_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_28_2__25_  (.A(u_multiplier_STAGE1_pp1_27_e42_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_28_2__16_ ),
    .ZN(u_multiplier_pp1_28 [5]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_28_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_28_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_28_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_28_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_28_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_28_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_28_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_28_2__17_ ),
    .ZN(u_multiplier_pp1_29 [12]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_28_3__18_  (.A(u_multiplier_STAGE1_pp1_27_e42_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_28_3__19_  (.A1(u_multiplier_STAGE1__0772_ ),
    .A2(u_multiplier_STAGE1__0771_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_28_3__20_  (.A(u_multiplier_STAGE1__0772_ ),
    .B(u_multiplier_STAGE1__0771_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_28_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_28_3__21_  (.A1(u_multiplier_STAGE1__0773_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_28_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_28_3__22_  (.A(u_multiplier_STAGE1__0773_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_28_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_28_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_28_3__23_  (.A1(u_multiplier_STAGE1__0774_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_28_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_28_3__24_  (.A(u_multiplier_STAGE1__0774_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_28_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_28_3__25_  (.A(u_multiplier_STAGE1_pp1_27_e42_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_28_3__16_ ),
    .ZN(u_multiplier_pp1_28 [4]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_28_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_28_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_28_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_28_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_28_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_28_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_28_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_28_3__17_ ),
    .ZN(u_multiplier_pp1_29 [11]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_28_4__18_  (.A(u_multiplier_STAGE1_pp1_27_e42_4_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_28_4__19_  (.A1(u_multiplier_STAGE1__0776_ ),
    .A2(u_multiplier_STAGE1__0775_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_4__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_28_4__20_  (.A(u_multiplier_STAGE1__0776_ ),
    .B(u_multiplier_STAGE1__0775_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_28_4__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_28_4__21_  (.A1(u_multiplier_STAGE1__0777_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_28_4__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_4__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_28_4__22_  (.A(u_multiplier_STAGE1__0777_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_28_4__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_28_4__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_28_4__23_  (.A1(u_multiplier_STAGE1__0778_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_28_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_28_4__24_  (.A(u_multiplier_STAGE1__0778_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_28_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_28_4__25_  (.A(u_multiplier_STAGE1_pp1_27_e42_4_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_28_4__16_ ),
    .ZN(u_multiplier_pp1_28 [3]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_28_4__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_28_4__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_28_4__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_28_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_28_4__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_28_4__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_28_4__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_28_4__17_ ),
    .ZN(u_multiplier_pp1_29 [10]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_28_5__18_  (.A(u_multiplier_STAGE1_pp1_27_e42_5_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_5__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_28_5__19_  (.A1(u_multiplier_STAGE1__0780_ ),
    .A2(u_multiplier_STAGE1__0779_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_5__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_28_5__20_  (.A(u_multiplier_STAGE1__0780_ ),
    .B(u_multiplier_STAGE1__0779_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_28_5__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_28_5__21_  (.A1(u_multiplier_STAGE1__0781_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_28_5__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_5__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_28_5__22_  (.A(u_multiplier_STAGE1__0781_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_28_5__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_28_5__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_28_5__23_  (.A1(u_multiplier_STAGE1__0782_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_28_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_5__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_28_5__24_  (.A(u_multiplier_STAGE1__0782_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_28_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_5__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_28_5__25_  (.A(u_multiplier_STAGE1_pp1_27_e42_5_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_28_5__16_ ),
    .ZN(u_multiplier_pp1_28 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_28_5__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_28_5__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_28_5__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_28_e42_5_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_28_5__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_28_5__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_28_5__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_28_5__17_ ),
    .ZN(u_multiplier_pp1_29 [9]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_28_6__18_  (.A(u_multiplier_STAGE1_pp1_27_e42_6_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_6__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_28_6__19_  (.A1(u_multiplier_STAGE1__0784_ ),
    .A2(u_multiplier_STAGE1__0783_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_6__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_28_6__20_  (.A(u_multiplier_STAGE1__0784_ ),
    .B(u_multiplier_STAGE1__0783_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_28_6__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_28_6__21_  (.A1(u_multiplier_STAGE1__0785_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_28_6__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_6__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_28_6__22_  (.A(u_multiplier_STAGE1__0785_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_28_6__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_28_6__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_28_6__23_  (.A1(u_multiplier_STAGE1__0786_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_28_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_6__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_28_6__24_  (.A(u_multiplier_STAGE1__0786_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_28_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_28_6__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_28_6__25_  (.A(u_multiplier_STAGE1_pp1_27_e42_6_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_28_6__16_ ),
    .ZN(u_multiplier_pp1_28 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_28_6__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_28_6__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_28_6__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_28_e42_6_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_28_6__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_28_6__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_28_6__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_28_6__17_ ),
    .ZN(u_multiplier_pp1_29 [8]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_29_1__18_  (.A(u_multiplier_STAGE1_pp1_28_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_29_1__19_  (.A1(u_multiplier_STAGE1__0790_ ),
    .A2(u_multiplier_STAGE1__0789_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_1__20_  (.A(u_multiplier_STAGE1__0790_ ),
    .B(u_multiplier_STAGE1__0789_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_29_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_29_1__21_  (.A1(u_multiplier_STAGE1__0791_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_29_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_1__22_  (.A(u_multiplier_STAGE1__0791_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_29_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_29_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_29_1__23_  (.A1(u_multiplier_STAGE1__0792_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_29_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_1__24_  (.A(u_multiplier_STAGE1__0792_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_29_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_1__25_  (.A(u_multiplier_STAGE1_pp1_28_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_29_1__16_ ),
    .ZN(u_multiplier_pp1_29 [6]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_29_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_29_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_29_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_29_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_29_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_29_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_29_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_29_1__17_ ),
    .ZN(u_multiplier_pp1_30 [14]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_29_2__18_  (.A(u_multiplier_STAGE1_pp1_28_e42_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_29_2__19_  (.A1(u_multiplier_STAGE1__0794_ ),
    .A2(u_multiplier_STAGE1__0793_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_2__20_  (.A(u_multiplier_STAGE1__0794_ ),
    .B(u_multiplier_STAGE1__0793_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_29_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_29_2__21_  (.A1(u_multiplier_STAGE1__0795_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_29_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_2__22_  (.A(u_multiplier_STAGE1__0795_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_29_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_29_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_29_2__23_  (.A1(u_multiplier_STAGE1__0796_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_29_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_2__24_  (.A(u_multiplier_STAGE1__0796_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_29_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_2__25_  (.A(u_multiplier_STAGE1_pp1_28_e42_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_29_2__16_ ),
    .ZN(u_multiplier_pp1_29 [5]));
 NAND2_X2 u_multiplier_STAGE1_E_4_2_pp_29_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_29_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_29_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_29_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_29_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_29_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_29_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_29_2__17_ ),
    .ZN(u_multiplier_pp1_30 [13]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_29_3__18_  (.A(u_multiplier_STAGE1_pp1_28_e42_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_29_3__19_  (.A1(u_multiplier_STAGE1__0798_ ),
    .A2(u_multiplier_STAGE1__0797_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_3__20_  (.A(u_multiplier_STAGE1__0798_ ),
    .B(u_multiplier_STAGE1__0797_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_29_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_29_3__21_  (.A1(u_multiplier_STAGE1__0799_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_29_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_3__22_  (.A(u_multiplier_STAGE1__0799_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_29_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_29_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_29_3__23_  (.A1(u_multiplier_STAGE1__0800_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_29_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_3__24_  (.A(u_multiplier_STAGE1__0800_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_29_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_3__25_  (.A(u_multiplier_STAGE1_pp1_28_e42_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_29_3__16_ ),
    .ZN(u_multiplier_pp1_29 [4]));
 NAND2_X2 u_multiplier_STAGE1_E_4_2_pp_29_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_29_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_29_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_29_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_29_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_29_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_29_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_29_3__17_ ),
    .ZN(u_multiplier_pp1_30 [12]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_29_4__18_  (.A(u_multiplier_STAGE1_pp1_28_e42_4_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_29_4__19_  (.A1(u_multiplier_STAGE1__0802_ ),
    .A2(u_multiplier_STAGE1__0801_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_4__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_4__20_  (.A(u_multiplier_STAGE1__0802_ ),
    .B(u_multiplier_STAGE1__0801_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_29_4__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_29_4__21_  (.A1(u_multiplier_STAGE1__0803_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_29_4__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_4__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_4__22_  (.A(u_multiplier_STAGE1__0803_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_29_4__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_29_4__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_29_4__23_  (.A1(u_multiplier_STAGE1__0804_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_29_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_4__24_  (.A(u_multiplier_STAGE1__0804_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_29_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_4__25_  (.A(u_multiplier_STAGE1_pp1_28_e42_4_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_29_4__16_ ),
    .ZN(u_multiplier_pp1_29 [3]));
 NAND2_X2 u_multiplier_STAGE1_E_4_2_pp_29_4__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_29_4__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_29_4__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_29_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_29_4__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_29_4__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_29_4__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_29_4__17_ ),
    .ZN(u_multiplier_pp1_30 [11]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_29_5__18_  (.A(u_multiplier_STAGE1_pp1_28_e42_5_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_5__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_29_5__19_  (.A1(u_multiplier_STAGE1__0806_ ),
    .A2(u_multiplier_STAGE1__0805_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_5__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_5__20_  (.A(u_multiplier_STAGE1__0806_ ),
    .B(u_multiplier_STAGE1__0805_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_29_5__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_29_5__21_  (.A1(u_multiplier_STAGE1__0807_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_29_5__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_5__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_5__22_  (.A(u_multiplier_STAGE1__0807_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_29_5__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_29_5__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_29_5__23_  (.A1(u_multiplier_STAGE1__0808_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_29_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_5__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_5__24_  (.A(u_multiplier_STAGE1__0808_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_29_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_5__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_5__25_  (.A(u_multiplier_STAGE1_pp1_28_e42_5_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_29_5__16_ ),
    .ZN(u_multiplier_pp1_29 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_29_5__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_29_5__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_29_5__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_29_e42_5_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_29_5__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_29_5__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_29_5__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_29_5__17_ ),
    .ZN(u_multiplier_pp1_30 [10]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_29_6__18_  (.A(u_multiplier_STAGE1_pp1_28_e42_6_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_6__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_29_6__19_  (.A1(u_multiplier_STAGE1__0810_ ),
    .A2(u_multiplier_STAGE1__0809_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_6__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_6__20_  (.A(u_multiplier_STAGE1__0810_ ),
    .B(u_multiplier_STAGE1__0809_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_29_6__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_29_6__21_  (.A1(u_multiplier_STAGE1__0811_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_29_6__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_6__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_6__22_  (.A(u_multiplier_STAGE1__0811_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_29_6__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_29_6__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_29_6__23_  (.A1(u_multiplier_STAGE1__0812_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_29_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_6__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_6__24_  (.A(u_multiplier_STAGE1__0812_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_29_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_6__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_6__25_  (.A(u_multiplier_STAGE1_pp1_28_e42_6_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_29_6__16_ ),
    .ZN(u_multiplier_pp1_29 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_29_6__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_29_6__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_29_6__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_29_e42_6_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_29_6__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_29_6__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_29_6__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_29_6__17_ ),
    .ZN(u_multiplier_pp1_30 [9]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_29_7__18_  (.A(net126),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_7__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_29_7__19_  (.A1(u_multiplier_STAGE1__0814_ ),
    .A2(u_multiplier_STAGE1__0813_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_7__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_7__20_  (.A(u_multiplier_STAGE1__0814_ ),
    .B(u_multiplier_STAGE1__0813_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_29_7__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_29_7__21_  (.A1(u_multiplier_STAGE1__0815_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_29_7__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_7__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_7__22_  (.A(u_multiplier_STAGE1__0815_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_29_7__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_29_7__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_29_7__23_  (.A1(u_multiplier_STAGE1__0816_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_29_7__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_7__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_7__24_  (.A(u_multiplier_STAGE1__0816_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_29_7__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_29_7__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_29_7__25_  (.A(net127),
    .B(u_multiplier_STAGE1_E_4_2_pp_29_7__16_ ),
    .ZN(u_multiplier_pp1_29 [0]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_29_7__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_29_7__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_29_7__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_29_e42_7_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_29_7__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_29_7__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_29_7__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_29_7__17_ ),
    .ZN(u_multiplier_pp1_30 [8]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_30_1__18_  (.A(u_multiplier_STAGE1_pp1_29_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_30_1__19_  (.A1(u_multiplier_STAGE1__0818_ ),
    .A2(u_multiplier_STAGE1__0817_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_1__20_  (.A(u_multiplier_STAGE1__0818_ ),
    .B(u_multiplier_STAGE1__0817_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_30_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_30_1__21_  (.A1(u_multiplier_STAGE1__0819_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_30_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_1__22_  (.A(u_multiplier_STAGE1__0819_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_30_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_30_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_30_1__23_  (.A1(u_multiplier_STAGE1__0820_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_30_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_1__24_  (.A(u_multiplier_STAGE1__0820_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_30_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_1__25_  (.A(u_multiplier_STAGE1_pp1_29_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_30_1__16_ ),
    .ZN(u_multiplier_pp1_30 [7]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_30_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_30_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_30_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_30_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_30_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_30_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_30_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_30_1__17_ ),
    .ZN(u_multiplier_pp1_31 [15]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_30_2__18_  (.A(u_multiplier_STAGE1_pp1_29_e42_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_30_2__19_  (.A1(u_multiplier_STAGE1__0822_ ),
    .A2(u_multiplier_STAGE1__0821_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_2__20_  (.A(u_multiplier_STAGE1__0822_ ),
    .B(u_multiplier_STAGE1__0821_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_30_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_30_2__21_  (.A1(u_multiplier_STAGE1__0823_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_30_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_2__22_  (.A(u_multiplier_STAGE1__0823_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_30_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_30_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_30_2__23_  (.A1(u_multiplier_STAGE1__0824_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_30_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_2__24_  (.A(u_multiplier_STAGE1__0824_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_30_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_2__25_  (.A(u_multiplier_STAGE1_pp1_29_e42_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_30_2__16_ ),
    .ZN(u_multiplier_pp1_30 [6]));
 NAND2_X2 u_multiplier_STAGE1_E_4_2_pp_30_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_30_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_30_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_30_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_30_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_30_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_30_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_30_2__17_ ),
    .ZN(u_multiplier_pp1_31 [14]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_30_3__18_  (.A(u_multiplier_STAGE1_pp1_29_e42_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_30_3__19_  (.A1(u_multiplier_STAGE1__0826_ ),
    .A2(u_multiplier_STAGE1__0825_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_3__20_  (.A(u_multiplier_STAGE1__0826_ ),
    .B(u_multiplier_STAGE1__0825_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_30_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_30_3__21_  (.A1(u_multiplier_STAGE1__0827_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_30_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_3__22_  (.A(u_multiplier_STAGE1__0827_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_30_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_30_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_30_3__23_  (.A1(u_multiplier_STAGE1__0828_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_30_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_3__24_  (.A(u_multiplier_STAGE1__0828_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_30_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_3__25_  (.A(u_multiplier_STAGE1_pp1_29_e42_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_30_3__16_ ),
    .ZN(u_multiplier_pp1_30 [5]));
 NAND2_X2 u_multiplier_STAGE1_E_4_2_pp_30_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_30_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_30_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_30_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_30_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_30_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_30_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_30_3__17_ ),
    .ZN(u_multiplier_pp1_31 [13]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_30_4__18_  (.A(u_multiplier_STAGE1_pp1_29_e42_4_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_30_4__19_  (.A1(u_multiplier_STAGE1__0830_ ),
    .A2(u_multiplier_STAGE1__0829_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_4__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_4__20_  (.A(u_multiplier_STAGE1__0830_ ),
    .B(u_multiplier_STAGE1__0829_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_30_4__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_30_4__21_  (.A1(u_multiplier_STAGE1__0831_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_30_4__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_4__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_4__22_  (.A(u_multiplier_STAGE1__0831_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_30_4__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_30_4__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_30_4__23_  (.A1(u_multiplier_STAGE1__0832_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_30_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_4__24_  (.A(u_multiplier_STAGE1__0832_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_30_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_4__25_  (.A(u_multiplier_STAGE1_pp1_29_e42_4_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_30_4__16_ ),
    .ZN(u_multiplier_pp1_30 [4]));
 NAND2_X2 u_multiplier_STAGE1_E_4_2_pp_30_4__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_30_4__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_30_4__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_30_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_30_4__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_30_4__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_30_4__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_30_4__17_ ),
    .ZN(u_multiplier_pp1_31 [12]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_30_5__18_  (.A(u_multiplier_STAGE1_pp1_29_e42_5_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_5__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_30_5__19_  (.A1(u_multiplier_STAGE1__0834_ ),
    .A2(u_multiplier_STAGE1__0833_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_5__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_5__20_  (.A(u_multiplier_STAGE1__0834_ ),
    .B(u_multiplier_STAGE1__0833_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_30_5__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_30_5__21_  (.A1(u_multiplier_STAGE1__0835_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_30_5__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_5__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_5__22_  (.A(u_multiplier_STAGE1__0835_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_30_5__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_30_5__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_30_5__23_  (.A1(u_multiplier_STAGE1__0836_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_30_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_5__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_5__24_  (.A(u_multiplier_STAGE1__0836_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_30_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_5__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_5__25_  (.A(u_multiplier_STAGE1_pp1_29_e42_5_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_30_5__16_ ),
    .ZN(u_multiplier_pp1_30 [3]));
 NAND2_X2 u_multiplier_STAGE1_E_4_2_pp_30_5__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_30_5__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_30_5__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_30_e42_5_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_30_5__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_30_5__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_30_5__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_30_5__17_ ),
    .ZN(u_multiplier_pp1_31 [11]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_30_6__18_  (.A(u_multiplier_STAGE1_pp1_29_e42_6_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_6__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_30_6__19_  (.A1(u_multiplier_STAGE1__0838_ ),
    .A2(u_multiplier_STAGE1__0837_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_6__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_6__20_  (.A(u_multiplier_STAGE1__0838_ ),
    .B(u_multiplier_STAGE1__0837_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_30_6__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_30_6__21_  (.A1(u_multiplier_STAGE1__0839_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_30_6__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_6__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_6__22_  (.A(u_multiplier_STAGE1__0839_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_30_6__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_30_6__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_30_6__23_  (.A1(u_multiplier_STAGE1__0840_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_30_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_6__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_6__24_  (.A(u_multiplier_STAGE1__0840_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_30_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_6__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_6__25_  (.A(u_multiplier_STAGE1_pp1_29_e42_6_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_30_6__16_ ),
    .ZN(u_multiplier_pp1_30 [2]));
 NAND2_X2 u_multiplier_STAGE1_E_4_2_pp_30_6__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_30_6__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_30_6__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_30_e42_6_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_30_6__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_30_6__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_30_6__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_30_6__17_ ),
    .ZN(u_multiplier_pp1_31 [10]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_30_7__18_  (.A(u_multiplier_STAGE1_pp1_29_e42_7_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_7__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_30_7__19_  (.A1(u_multiplier_STAGE1__0842_ ),
    .A2(u_multiplier_STAGE1__0841_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_7__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_7__20_  (.A(u_multiplier_STAGE1__0842_ ),
    .B(u_multiplier_STAGE1__0841_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_30_7__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_30_7__21_  (.A1(u_multiplier_STAGE1__0843_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_30_7__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_7__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_7__22_  (.A(u_multiplier_STAGE1__0843_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_30_7__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_30_7__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_30_7__23_  (.A1(u_multiplier_STAGE1__0844_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_30_7__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_7__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_7__24_  (.A(u_multiplier_STAGE1__0844_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_30_7__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_30_7__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_30_7__25_  (.A(u_multiplier_STAGE1_pp1_29_e42_7_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_30_7__16_ ),
    .ZN(u_multiplier_pp1_30 [1]));
 NAND2_X2 u_multiplier_STAGE1_E_4_2_pp_30_7__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_30_7__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_30_7__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_30_e42_7_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_30_7__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_30_7__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_30_7__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_30_7__17_ ),
    .ZN(u_multiplier_pp1_31 [9]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_31_1__18_  (.A(u_multiplier_STAGE1_pp1_30_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_1__19_  (.A1(u_multiplier_STAGE1__0848_ ),
    .A2(u_multiplier_STAGE1__0847_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_1__20_  (.A(u_multiplier_STAGE1__0848_ ),
    .B(u_multiplier_STAGE1__0847_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_31_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_1__21_  (.A1(u_multiplier_STAGE1__0849_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_31_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_1__22_  (.A(u_multiplier_STAGE1__0849_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_31_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_31_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_1__23_  (.A1(u_multiplier_STAGE1__0850_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_31_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_1__24_  (.A(u_multiplier_STAGE1__0850_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_31_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_1__25_  (.A(u_multiplier_STAGE1_pp1_30_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_31_1__16_ ),
    .ZN(u_multiplier_pp1_31 [7]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_31_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_31_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_31_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_31_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_31_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_31_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_31_1__17_ ),
    .ZN(u_multiplier_pp1_32 [15]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_31_2__18_  (.A(u_multiplier_STAGE1_pp1_30_e42_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_2__19_  (.A1(u_multiplier_STAGE1__0852_ ),
    .A2(u_multiplier_STAGE1__0851_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_2__20_  (.A(u_multiplier_STAGE1__0852_ ),
    .B(u_multiplier_STAGE1__0851_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_31_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_2__21_  (.A1(u_multiplier_STAGE1__0853_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_31_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_2__22_  (.A(u_multiplier_STAGE1__0853_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_31_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_31_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_2__23_  (.A1(u_multiplier_STAGE1__0854_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_31_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_2__24_  (.A(u_multiplier_STAGE1__0854_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_31_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_2__25_  (.A(u_multiplier_STAGE1_pp1_30_e42_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_31_2__16_ ),
    .ZN(u_multiplier_pp1_31 [6]));
 NAND2_X2 u_multiplier_STAGE1_E_4_2_pp_31_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_31_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_31_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_31_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_31_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_31_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_31_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_31_2__17_ ),
    .ZN(u_multiplier_pp1_32 [14]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_31_3__18_  (.A(u_multiplier_STAGE1_pp1_30_e42_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_3__19_  (.A1(u_multiplier_STAGE1__0856_ ),
    .A2(u_multiplier_STAGE1__0855_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_3__20_  (.A(u_multiplier_STAGE1__0856_ ),
    .B(u_multiplier_STAGE1__0855_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_31_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_3__21_  (.A1(u_multiplier_STAGE1__0857_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_31_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_3__22_  (.A(u_multiplier_STAGE1__0857_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_31_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_31_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_3__23_  (.A1(u_multiplier_STAGE1__0858_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_31_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_3__24_  (.A(u_multiplier_STAGE1__0858_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_31_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_3__25_  (.A(u_multiplier_STAGE1_pp1_30_e42_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_31_3__16_ ),
    .ZN(u_multiplier_pp1_31 [5]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_31_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_31_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_31_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_31_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_31_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_31_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_31_3__17_ ),
    .ZN(u_multiplier_pp1_32 [13]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_31_4__18_  (.A(u_multiplier_STAGE1_pp1_30_e42_4_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_4__19_  (.A1(u_multiplier_STAGE1__0860_ ),
    .A2(u_multiplier_STAGE1__0859_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_4__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_4__20_  (.A(u_multiplier_STAGE1__0860_ ),
    .B(u_multiplier_STAGE1__0859_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_31_4__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_4__21_  (.A1(u_multiplier_STAGE1__0861_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_31_4__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_4__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_4__22_  (.A(u_multiplier_STAGE1__0861_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_31_4__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_31_4__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_4__23_  (.A1(u_multiplier_STAGE1__0862_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_31_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_4__24_  (.A(u_multiplier_STAGE1__0862_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_31_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_4__25_  (.A(u_multiplier_STAGE1_pp1_30_e42_4_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_31_4__16_ ),
    .ZN(u_multiplier_pp1_31 [4]));
 NAND2_X2 u_multiplier_STAGE1_E_4_2_pp_31_4__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_31_4__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_31_4__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_31_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_31_4__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_31_4__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_31_4__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_31_4__17_ ),
    .ZN(u_multiplier_pp1_32 [12]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_31_5__18_  (.A(u_multiplier_STAGE1_pp1_30_e42_5_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_5__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_5__19_  (.A1(u_multiplier_STAGE1__0864_ ),
    .A2(u_multiplier_STAGE1__0863_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_5__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_5__20_  (.A(u_multiplier_STAGE1__0864_ ),
    .B(u_multiplier_STAGE1__0863_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_31_5__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_5__21_  (.A1(u_multiplier_STAGE1__0865_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_31_5__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_5__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_5__22_  (.A(u_multiplier_STAGE1__0865_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_31_5__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_31_5__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_5__23_  (.A1(u_multiplier_STAGE1__0866_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_31_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_5__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_5__24_  (.A(u_multiplier_STAGE1__0866_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_31_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_5__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_5__25_  (.A(u_multiplier_STAGE1_pp1_30_e42_5_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_31_5__16_ ),
    .ZN(u_multiplier_pp1_31 [3]));
 NAND2_X2 u_multiplier_STAGE1_E_4_2_pp_31_5__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_31_5__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_31_5__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_31_e42_5_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_31_5__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_31_5__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_31_5__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_31_5__17_ ),
    .ZN(u_multiplier_pp1_32 [11]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_31_6__18_  (.A(u_multiplier_STAGE1_pp1_30_e42_6_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_6__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_6__19_  (.A1(u_multiplier_STAGE1__0868_ ),
    .A2(u_multiplier_STAGE1__0867_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_6__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_6__20_  (.A(u_multiplier_STAGE1__0868_ ),
    .B(u_multiplier_STAGE1__0867_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_31_6__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_6__21_  (.A1(u_multiplier_STAGE1__0869_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_31_6__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_6__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_6__22_  (.A(u_multiplier_STAGE1__0869_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_31_6__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_31_6__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_6__23_  (.A1(u_multiplier_STAGE1__0870_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_31_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_6__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_6__24_  (.A(u_multiplier_STAGE1__0870_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_31_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_6__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_6__25_  (.A(u_multiplier_STAGE1_pp1_30_e42_6_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_31_6__16_ ),
    .ZN(u_multiplier_pp1_31 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_6__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_31_6__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_31_6__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_31_e42_6_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_31_6__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_31_6__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_31_6__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_31_6__17_ ),
    .ZN(u_multiplier_pp1_32 [10]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_31_7__18_  (.A(u_multiplier_STAGE1_pp1_30_e42_7_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_7__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_7__19_  (.A1(u_multiplier_STAGE1__0872_ ),
    .A2(u_multiplier_STAGE1__0871_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_7__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_7__20_  (.A(u_multiplier_STAGE1__0872_ ),
    .B(u_multiplier_STAGE1__0871_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_31_7__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_7__21_  (.A1(u_multiplier_STAGE1__0873_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_31_7__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_7__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_7__22_  (.A(u_multiplier_STAGE1__0873_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_31_7__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_31_7__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_7__23_  (.A1(u_multiplier_STAGE1__0874_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_31_7__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_7__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_7__24_  (.A(u_multiplier_STAGE1__0874_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_31_7__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_7__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_7__25_  (.A(u_multiplier_STAGE1_pp1_30_e42_7_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_31_7__16_ ),
    .ZN(u_multiplier_pp1_31 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_7__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_31_7__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_31_7__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_31_e42_7_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_31_7__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_31_7__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_31_7__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_31_7__17_ ),
    .ZN(u_multiplier_pp1_32 [9]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_31_8__18_  (.A(net128),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_8__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_8__19_  (.A1(u_multiplier_STAGE1__0876_ ),
    .A2(u_multiplier_STAGE1__0875_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_8__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_8__20_  (.A(u_multiplier_STAGE1__0876_ ),
    .B(u_multiplier_STAGE1__0875_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_31_8__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_8__21_  (.A1(u_multiplier_STAGE1__0877_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_31_8__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_8__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_8__22_  (.A(u_multiplier_STAGE1__0877_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_31_8__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_31_8__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_8__23_  (.A1(u_multiplier_STAGE1__0878_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_31_8__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_8__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_8__24_  (.A(u_multiplier_STAGE1__0878_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_31_8__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_31_8__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_31_8__25_  (.A(net129),
    .B(u_multiplier_STAGE1_E_4_2_pp_31_8__16_ ),
    .ZN(u_multiplier_pp1_31 [0]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_31_8__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_31_8__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_31_8__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_31_e42_8_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_31_8__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_31_8__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_31_8__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_31_8__17_ ),
    .ZN(u_multiplier_pp1_32 [8]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_32_1__18_  (.A(u_multiplier_STAGE1_pp1_31_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_1__19_  (.A1(u_multiplier_STAGE1__0880_ ),
    .A2(u_multiplier_STAGE1__0879_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_1__20_  (.A(u_multiplier_STAGE1__0880_ ),
    .B(u_multiplier_STAGE1__0879_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_1__21_  (.A1(u_multiplier_STAGE1__0881_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_1__22_  (.A(u_multiplier_STAGE1__0881_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_1__23_  (.A1(u_multiplier_STAGE1__0882_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_1__24_  (.A(u_multiplier_STAGE1__0882_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_1__25_  (.A(u_multiplier_STAGE1_pp1_31_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_1__16_ ),
    .ZN(u_multiplier_pp1_32 [7]));
 NAND2_X2 u_multiplier_STAGE1_E_4_2_pp_32_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_32_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_32_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_32_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_32_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_32_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_32_1__17_ ),
    .ZN(u_multiplier_pp1_33 [15]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_32_2__18_  (.A(u_multiplier_STAGE1_pp1_31_e42_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_2__19_  (.A1(u_multiplier_STAGE1__0884_ ),
    .A2(u_multiplier_STAGE1__0883_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_2__20_  (.A(u_multiplier_STAGE1__0884_ ),
    .B(u_multiplier_STAGE1__0883_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_2__21_  (.A1(u_multiplier_STAGE1__0885_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_2__22_  (.A(u_multiplier_STAGE1__0885_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_2__23_  (.A1(u_multiplier_STAGE1__0886_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_2__24_  (.A(u_multiplier_STAGE1__0886_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_2__25_  (.A(u_multiplier_STAGE1_pp1_31_e42_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_2__16_ ),
    .ZN(u_multiplier_pp1_32 [6]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_32_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_32_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_32_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_32_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_32_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_32_2__17_ ),
    .ZN(u_multiplier_pp1_33 [14]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_32_3__18_  (.A(u_multiplier_STAGE1_pp1_31_e42_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_3__19_  (.A1(u_multiplier_STAGE1__0888_ ),
    .A2(u_multiplier_STAGE1__0887_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_3__20_  (.A(u_multiplier_STAGE1__0888_ ),
    .B(u_multiplier_STAGE1__0887_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_3__21_  (.A1(u_multiplier_STAGE1__0889_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_3__22_  (.A(u_multiplier_STAGE1__0889_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_3__23_  (.A1(u_multiplier_STAGE1__0890_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_3__24_  (.A(u_multiplier_STAGE1__0890_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_3__25_  (.A(u_multiplier_STAGE1_pp1_31_e42_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_3__16_ ),
    .ZN(u_multiplier_pp1_32 [5]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_32_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_32_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_32_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_32_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_32_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_32_3__17_ ),
    .ZN(u_multiplier_pp1_33 [13]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_32_4__18_  (.A(u_multiplier_STAGE1_pp1_31_e42_4_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_4__19_  (.A1(u_multiplier_STAGE1__0892_ ),
    .A2(u_multiplier_STAGE1__0891_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_4__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_4__20_  (.A(u_multiplier_STAGE1__0892_ ),
    .B(u_multiplier_STAGE1__0891_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_4__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_4__21_  (.A1(u_multiplier_STAGE1__0893_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_4__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_4__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_4__22_  (.A(u_multiplier_STAGE1__0893_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_4__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_4__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_4__23_  (.A1(u_multiplier_STAGE1__0894_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_4__24_  (.A(u_multiplier_STAGE1__0894_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_4__25_  (.A(u_multiplier_STAGE1_pp1_31_e42_4_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_4__16_ ),
    .ZN(u_multiplier_pp1_32 [4]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_4__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_32_4__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_4__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_32_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_32_4__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_32_4__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_32_4__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_32_4__17_ ),
    .ZN(u_multiplier_pp1_33 [12]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_32_5__18_  (.A(u_multiplier_STAGE1_pp1_31_e42_5_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_5__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_5__19_  (.A1(u_multiplier_STAGE1__0896_ ),
    .A2(u_multiplier_STAGE1__0895_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_5__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_5__20_  (.A(u_multiplier_STAGE1__0896_ ),
    .B(u_multiplier_STAGE1__0895_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_5__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_5__21_  (.A1(u_multiplier_STAGE1__0897_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_5__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_5__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_5__22_  (.A(u_multiplier_STAGE1__0897_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_5__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_5__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_5__23_  (.A1(u_multiplier_STAGE1__0898_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_5__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_5__24_  (.A(u_multiplier_STAGE1__0898_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_5__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_5__25_  (.A(u_multiplier_STAGE1_pp1_31_e42_5_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_5__16_ ),
    .ZN(u_multiplier_pp1_32 [3]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_5__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_32_5__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_5__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_32_e42_5_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_32_5__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_32_5__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_32_5__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_32_5__17_ ),
    .ZN(u_multiplier_pp1_33 [11]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_32_6__18_  (.A(u_multiplier_STAGE1_pp1_31_e42_6_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_6__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_6__19_  (.A1(u_multiplier_STAGE1__0900_ ),
    .A2(u_multiplier_STAGE1__0899_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_6__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_6__20_  (.A(u_multiplier_STAGE1__0900_ ),
    .B(u_multiplier_STAGE1__0899_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_6__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_6__21_  (.A1(u_multiplier_STAGE1__0901_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_6__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_6__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_6__22_  (.A(u_multiplier_STAGE1__0901_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_6__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_6__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_6__23_  (.A1(u_multiplier_STAGE1__0902_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_6__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_6__24_  (.A(u_multiplier_STAGE1__0902_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_6__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_6__25_  (.A(u_multiplier_STAGE1_pp1_31_e42_6_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_6__16_ ),
    .ZN(u_multiplier_pp1_32 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_6__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_32_6__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_6__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_32_e42_6_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_32_6__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_32_6__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_32_6__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_32_6__17_ ),
    .ZN(u_multiplier_pp1_33 [10]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_32_7__18_  (.A(u_multiplier_STAGE1_pp1_31_e42_7_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_7__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_7__19_  (.A1(u_multiplier_STAGE1__0904_ ),
    .A2(u_multiplier_STAGE1__0903_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_7__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_7__20_  (.A(u_multiplier_STAGE1__0904_ ),
    .B(u_multiplier_STAGE1__0903_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_7__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_7__21_  (.A1(u_multiplier_STAGE1__0905_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_7__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_7__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_7__22_  (.A(u_multiplier_STAGE1__0905_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_7__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_7__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_7__23_  (.A1(u_multiplier_STAGE1__0906_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_7__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_7__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_7__24_  (.A(u_multiplier_STAGE1__0906_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_7__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_7__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_7__25_  (.A(u_multiplier_STAGE1_pp1_31_e42_7_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_7__16_ ),
    .ZN(u_multiplier_pp1_32 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_7__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_32_7__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_7__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_32_e42_7_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_32_7__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_32_7__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_32_7__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_32_7__17_ ),
    .ZN(u_multiplier_pp1_33 [9]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_32_8__18_  (.A(u_multiplier_STAGE1_pp1_31_e42_8_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_8__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_8__19_  (.A1(u_multiplier_STAGE1__0908_ ),
    .A2(u_multiplier_STAGE1__0907_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_8__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_8__20_  (.A(u_multiplier_STAGE1__0908_ ),
    .B(u_multiplier_STAGE1__0907_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_8__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_8__21_  (.A1(u_multiplier_STAGE1__0909_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_8__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_8__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_8__22_  (.A(u_multiplier_STAGE1__0909_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_8__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_8__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_8__23_  (.A1(net130),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_8__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_8__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_8__24_  (.A(net131),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_8__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_8__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_8__25_  (.A(u_multiplier_STAGE1_pp1_31_e42_8_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_8__16_ ),
    .ZN(u_multiplier_pp1_32 [0]));
 NAND2_X2 u_multiplier_STAGE1_E_4_2_pp_32_8__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_32_8__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_8__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_32_e42_8_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_32_8__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_32_8__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_32_8__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_32_8__17_ ),
    .ZN(u_multiplier_pp1_33 [8]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_33_1__18_  (.A(u_multiplier_STAGE1_pp1_32_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_1__19_  (.A1(u_multiplier_STAGE1__0911_ ),
    .A2(u_multiplier_STAGE1__0910_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_1__20_  (.A(u_multiplier_STAGE1__0911_ ),
    .B(u_multiplier_STAGE1__0910_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_1__21_  (.A1(u_multiplier_STAGE1__0912_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_1__22_  (.A(u_multiplier_STAGE1__0912_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_1__23_  (.A1(u_multiplier_STAGE1__0913_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_1__24_  (.A(u_multiplier_STAGE1__0913_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_1__25_  (.A(u_multiplier_STAGE1_pp1_32_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_1__16_ ),
    .ZN(u_multiplier_pp1_33 [7]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_33_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_33_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_33_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_33_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_33_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_33_1__17_ ),
    .ZN(u_multiplier_pp1_34 [14]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_33_2__18_  (.A(u_multiplier_STAGE1_pp1_32_e42_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_2__19_  (.A1(u_multiplier_STAGE1__0915_ ),
    .A2(u_multiplier_STAGE1__0914_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_2__20_  (.A(u_multiplier_STAGE1__0915_ ),
    .B(u_multiplier_STAGE1__0914_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_2__21_  (.A1(u_multiplier_STAGE1__0916_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_2__22_  (.A(u_multiplier_STAGE1__0916_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_2__23_  (.A1(u_multiplier_STAGE1__0917_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_2__24_  (.A(u_multiplier_STAGE1__0917_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_2__25_  (.A(u_multiplier_STAGE1_pp1_32_e42_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_2__16_ ),
    .ZN(u_multiplier_pp1_33 [6]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_33_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_33_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_33_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_33_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_33_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_33_2__17_ ),
    .ZN(u_multiplier_pp1_34 [13]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_33_3__18_  (.A(u_multiplier_STAGE1_pp1_32_e42_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_3__19_  (.A1(u_multiplier_STAGE1__0919_ ),
    .A2(u_multiplier_STAGE1__0918_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_3__20_  (.A(u_multiplier_STAGE1__0919_ ),
    .B(u_multiplier_STAGE1__0918_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_3__21_  (.A1(u_multiplier_STAGE1__0920_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_3__22_  (.A(u_multiplier_STAGE1__0920_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_3__23_  (.A1(u_multiplier_STAGE1__0921_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_3__24_  (.A(u_multiplier_STAGE1__0921_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_3__25_  (.A(u_multiplier_STAGE1_pp1_32_e42_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_3__16_ ),
    .ZN(u_multiplier_pp1_33 [5]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_33_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_33_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_33_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_33_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_33_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_33_3__17_ ),
    .ZN(u_multiplier_pp1_34 [12]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_33_4__18_  (.A(u_multiplier_STAGE1_pp1_32_e42_4_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_4__19_  (.A1(u_multiplier_STAGE1__0923_ ),
    .A2(u_multiplier_STAGE1__0922_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_4__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_4__20_  (.A(u_multiplier_STAGE1__0923_ ),
    .B(u_multiplier_STAGE1__0922_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_4__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_4__21_  (.A1(u_multiplier_STAGE1__0924_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_4__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_4__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_4__22_  (.A(u_multiplier_STAGE1__0924_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_4__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_4__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_4__23_  (.A1(u_multiplier_STAGE1__0925_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_4__24_  (.A(u_multiplier_STAGE1__0925_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_4__25_  (.A(u_multiplier_STAGE1_pp1_32_e42_4_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_4__16_ ),
    .ZN(u_multiplier_pp1_33 [4]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_4__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_33_4__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_4__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_33_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_33_4__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_33_4__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_33_4__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_33_4__17_ ),
    .ZN(u_multiplier_pp1_34 [11]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_33_5__18_  (.A(u_multiplier_STAGE1_pp1_32_e42_5_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_5__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_5__19_  (.A1(u_multiplier_STAGE1__0927_ ),
    .A2(u_multiplier_STAGE1__0926_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_5__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_5__20_  (.A(u_multiplier_STAGE1__0927_ ),
    .B(u_multiplier_STAGE1__0926_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_5__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_5__21_  (.A1(u_multiplier_STAGE1__0928_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_5__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_5__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_5__22_  (.A(u_multiplier_STAGE1__0928_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_5__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_5__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_5__23_  (.A1(u_multiplier_STAGE1__0929_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_5__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_5__24_  (.A(u_multiplier_STAGE1__0929_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_5__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_5__25_  (.A(u_multiplier_STAGE1_pp1_32_e42_5_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_5__16_ ),
    .ZN(u_multiplier_pp1_33 [3]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_5__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_33_5__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_5__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_33_e42_5_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_33_5__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_33_5__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_33_5__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_33_5__17_ ),
    .ZN(u_multiplier_pp1_34 [10]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_33_6__18_  (.A(u_multiplier_STAGE1_pp1_32_e42_6_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_6__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_6__19_  (.A1(u_multiplier_STAGE1__0931_ ),
    .A2(u_multiplier_STAGE1__0930_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_6__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_6__20_  (.A(u_multiplier_STAGE1__0931_ ),
    .B(u_multiplier_STAGE1__0930_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_6__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_6__21_  (.A1(u_multiplier_STAGE1__0932_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_6__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_6__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_6__22_  (.A(u_multiplier_STAGE1__0932_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_6__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_6__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_6__23_  (.A1(u_multiplier_STAGE1__0933_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_6__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_6__24_  (.A(u_multiplier_STAGE1__0933_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_6__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_6__25_  (.A(u_multiplier_STAGE1_pp1_32_e42_6_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_6__16_ ),
    .ZN(u_multiplier_pp1_33 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_6__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_33_6__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_6__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_33_e42_6_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_33_6__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_33_6__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_33_6__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_33_6__17_ ),
    .ZN(u_multiplier_pp1_34 [9]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_33_7__18_  (.A(u_multiplier_STAGE1_pp1_32_e42_7_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_7__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_7__19_  (.A1(u_multiplier_STAGE1__0935_ ),
    .A2(u_multiplier_STAGE1__0934_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_7__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_7__20_  (.A(u_multiplier_STAGE1__0935_ ),
    .B(u_multiplier_STAGE1__0934_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_7__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_7__21_  (.A1(u_multiplier_STAGE1__0936_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_7__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_7__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_7__22_  (.A(u_multiplier_STAGE1__0936_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_7__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_7__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_7__23_  (.A1(u_multiplier_STAGE1__0937_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_7__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_7__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_7__24_  (.A(u_multiplier_STAGE1__0937_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_7__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_7__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_7__25_  (.A(u_multiplier_STAGE1_pp1_32_e42_7_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_7__16_ ),
    .ZN(u_multiplier_pp1_33 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_7__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_33_7__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_7__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_33_e42_7_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_33_7__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_33_7__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_33_7__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_33_7__17_ ),
    .ZN(u_multiplier_pp1_34 [8]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_34_1__18_  (.A(u_multiplier_STAGE1_pp1_33_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_1__19_  (.A1(u_multiplier_STAGE1__0941_ ),
    .A2(u_multiplier_STAGE1__0940_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_1__20_  (.A(u_multiplier_STAGE1__0941_ ),
    .B(u_multiplier_STAGE1__0940_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_1__21_  (.A1(u_multiplier_STAGE1__0942_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_1__22_  (.A(u_multiplier_STAGE1__0942_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_1__23_  (.A1(u_multiplier_STAGE1__0943_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_1__24_  (.A(u_multiplier_STAGE1__0943_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_1__25_  (.A(u_multiplier_STAGE1_pp1_33_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_1__16_ ),
    .ZN(u_multiplier_pp1_34 [6]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_34_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_34_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_34_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_34_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_34_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_34_1__17_ ),
    .ZN(u_multiplier_pp1_35 [13]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_34_2__18_  (.A(u_multiplier_STAGE1_pp1_33_e42_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_2__19_  (.A1(u_multiplier_STAGE1__0945_ ),
    .A2(u_multiplier_STAGE1__0944_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_2__20_  (.A(u_multiplier_STAGE1__0945_ ),
    .B(u_multiplier_STAGE1__0944_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_2__21_  (.A1(u_multiplier_STAGE1__0946_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_2__22_  (.A(u_multiplier_STAGE1__0946_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_2__23_  (.A1(u_multiplier_STAGE1__0947_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_2__24_  (.A(u_multiplier_STAGE1__0947_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_2__25_  (.A(u_multiplier_STAGE1_pp1_33_e42_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_2__16_ ),
    .ZN(u_multiplier_pp1_34 [5]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_34_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_34_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_34_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_34_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_34_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_34_2__17_ ),
    .ZN(u_multiplier_pp1_35 [12]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_34_3__18_  (.A(u_multiplier_STAGE1_pp1_33_e42_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_3__19_  (.A1(u_multiplier_STAGE1__0949_ ),
    .A2(u_multiplier_STAGE1__0948_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_3__20_  (.A(u_multiplier_STAGE1__0949_ ),
    .B(u_multiplier_STAGE1__0948_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_3__21_  (.A1(u_multiplier_STAGE1__0950_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_3__22_  (.A(u_multiplier_STAGE1__0950_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_3__23_  (.A1(u_multiplier_STAGE1__0951_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_3__24_  (.A(u_multiplier_STAGE1__0951_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_3__25_  (.A(u_multiplier_STAGE1_pp1_33_e42_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_3__16_ ),
    .ZN(u_multiplier_pp1_34 [4]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_34_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_34_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_34_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_34_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_34_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_34_3__17_ ),
    .ZN(u_multiplier_pp1_35 [11]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_34_4__18_  (.A(u_multiplier_STAGE1_pp1_33_e42_4_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_4__19_  (.A1(u_multiplier_STAGE1__0953_ ),
    .A2(u_multiplier_STAGE1__0952_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_4__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_4__20_  (.A(u_multiplier_STAGE1__0953_ ),
    .B(u_multiplier_STAGE1__0952_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_4__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_4__21_  (.A1(u_multiplier_STAGE1__0954_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_4__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_4__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_4__22_  (.A(u_multiplier_STAGE1__0954_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_4__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_4__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_4__23_  (.A1(u_multiplier_STAGE1__0955_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_4__24_  (.A(u_multiplier_STAGE1__0955_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_4__25_  (.A(u_multiplier_STAGE1_pp1_33_e42_4_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_4__16_ ),
    .ZN(u_multiplier_pp1_34 [3]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_4__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_34_4__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_4__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_34_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_34_4__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_34_4__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_34_4__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_34_4__17_ ),
    .ZN(u_multiplier_pp1_35 [10]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_34_5__18_  (.A(u_multiplier_STAGE1_pp1_33_e42_5_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_5__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_5__19_  (.A1(u_multiplier_STAGE1__0957_ ),
    .A2(u_multiplier_STAGE1__0956_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_5__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_5__20_  (.A(u_multiplier_STAGE1__0957_ ),
    .B(u_multiplier_STAGE1__0956_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_5__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_5__21_  (.A1(u_multiplier_STAGE1__0958_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_5__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_5__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_5__22_  (.A(u_multiplier_STAGE1__0958_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_5__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_5__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_5__23_  (.A1(u_multiplier_STAGE1__0959_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_5__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_5__24_  (.A(u_multiplier_STAGE1__0959_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_5__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_5__25_  (.A(u_multiplier_STAGE1_pp1_33_e42_5_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_5__16_ ),
    .ZN(u_multiplier_pp1_34 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_5__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_34_5__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_5__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_34_e42_5_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_34_5__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_34_5__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_34_5__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_34_5__17_ ),
    .ZN(u_multiplier_pp1_35 [9]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_34_6__18_  (.A(u_multiplier_STAGE1_pp1_33_e42_6_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_6__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_6__19_  (.A1(u_multiplier_STAGE1__0961_ ),
    .A2(u_multiplier_STAGE1__0960_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_6__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_6__20_  (.A(u_multiplier_STAGE1__0961_ ),
    .B(u_multiplier_STAGE1__0960_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_6__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_6__21_  (.A1(u_multiplier_STAGE1__0962_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_6__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_6__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_6__22_  (.A(u_multiplier_STAGE1__0962_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_6__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_6__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_6__23_  (.A1(u_multiplier_STAGE1__0963_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_6__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_6__24_  (.A(u_multiplier_STAGE1__0963_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_6__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_6__25_  (.A(u_multiplier_STAGE1_pp1_33_e42_6_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_6__16_ ),
    .ZN(u_multiplier_pp1_34 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_6__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_34_6__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_6__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_34_e42_6_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_34_6__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_34_6__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_34_6__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_34_6__17_ ),
    .ZN(u_multiplier_pp1_35 [8]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_34_7__18_  (.A(u_multiplier_STAGE1_pp1_33_e42_7_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_7__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_7__19_  (.A1(u_multiplier_STAGE1__0965_ ),
    .A2(u_multiplier_STAGE1__0964_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_7__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_7__20_  (.A(u_multiplier_STAGE1__0965_ ),
    .B(u_multiplier_STAGE1__0964_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_7__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_7__21_  (.A1(u_multiplier_STAGE1__0966_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_7__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_7__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_7__22_  (.A(u_multiplier_STAGE1__0966_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_7__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_7__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_7__23_  (.A1(u_multiplier_STAGE1__0967_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_7__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_7__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_7__24_  (.A(u_multiplier_STAGE1__0967_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_7__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_7__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_7__25_  (.A(u_multiplier_STAGE1_pp1_33_e42_7_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_7__16_ ),
    .ZN(u_multiplier_pp1_34 [0]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_7__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_34_7__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_7__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_34_e42_7_cout ));
 OAI21_X1 u_multiplier_STAGE1_E_4_2_pp_34_7__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_34_7__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_34_7__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_34_7__17_ ),
    .ZN(u_multiplier_pp1_35 [7]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_35_1__18_  (.A(u_multiplier_STAGE1_pp1_34_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_1__19_  (.A1(u_multiplier_STAGE1__0969_ ),
    .A2(u_multiplier_STAGE1__0968_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_1__20_  (.A(u_multiplier_STAGE1__0969_ ),
    .B(u_multiplier_STAGE1__0968_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_35_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_1__21_  (.A1(u_multiplier_STAGE1__0970_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_1__22_  (.A(u_multiplier_STAGE1__0970_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_35_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_1__23_  (.A1(u_multiplier_STAGE1__0971_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_1__24_  (.A(u_multiplier_STAGE1__0971_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_1__25_  (.A(u_multiplier_STAGE1_pp1_34_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_1__16_ ),
    .ZN(u_multiplier_pp1_35 [6]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_35_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_35_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_35_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_35_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_35_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_35_1__17_ ),
    .ZN(u_multiplier_pp1_36 [12]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_35_2__18_  (.A(u_multiplier_STAGE1_pp1_34_e42_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_2__19_  (.A1(u_multiplier_STAGE1__0973_ ),
    .A2(u_multiplier_STAGE1__0972_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_2__20_  (.A(u_multiplier_STAGE1__0973_ ),
    .B(u_multiplier_STAGE1__0972_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_35_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_2__21_  (.A1(u_multiplier_STAGE1__0974_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_2__22_  (.A(u_multiplier_STAGE1__0974_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_35_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_2__23_  (.A1(u_multiplier_STAGE1__0975_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_2__24_  (.A(u_multiplier_STAGE1__0975_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_2__25_  (.A(u_multiplier_STAGE1_pp1_34_e42_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_2__16_ ),
    .ZN(u_multiplier_pp1_35 [5]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_35_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_35_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_35_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_35_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_35_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_35_2__17_ ),
    .ZN(u_multiplier_pp1_36 [11]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_35_3__18_  (.A(u_multiplier_STAGE1_pp1_34_e42_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_3__19_  (.A1(u_multiplier_STAGE1__0977_ ),
    .A2(u_multiplier_STAGE1__0976_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_3__20_  (.A(u_multiplier_STAGE1__0977_ ),
    .B(u_multiplier_STAGE1__0976_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_35_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_3__21_  (.A1(u_multiplier_STAGE1__0978_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_3__22_  (.A(u_multiplier_STAGE1__0978_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_35_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_3__23_  (.A1(u_multiplier_STAGE1__0979_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_3__24_  (.A(u_multiplier_STAGE1__0979_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_3__25_  (.A(u_multiplier_STAGE1_pp1_34_e42_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_3__16_ ),
    .ZN(u_multiplier_pp1_35 [4]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_35_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_35_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_35_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_35_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_35_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_35_3__17_ ),
    .ZN(u_multiplier_pp1_36 [10]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_35_4__18_  (.A(u_multiplier_STAGE1_pp1_34_e42_4_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_4__19_  (.A1(u_multiplier_STAGE1__0981_ ),
    .A2(u_multiplier_STAGE1__0980_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_4__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_4__20_  (.A(u_multiplier_STAGE1__0981_ ),
    .B(u_multiplier_STAGE1__0980_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_35_4__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_4__21_  (.A1(u_multiplier_STAGE1__0982_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_4__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_4__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_4__22_  (.A(u_multiplier_STAGE1__0982_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_4__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_35_4__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_4__23_  (.A1(u_multiplier_STAGE1__0983_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_4__24_  (.A(u_multiplier_STAGE1__0983_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_4__25_  (.A(u_multiplier_STAGE1_pp1_34_e42_4_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_4__16_ ),
    .ZN(u_multiplier_pp1_35 [3]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_4__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_35_4__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_4__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_35_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_35_4__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_35_4__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_35_4__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_35_4__17_ ),
    .ZN(u_multiplier_pp1_36 [9]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_35_5__18_  (.A(u_multiplier_STAGE1_pp1_34_e42_5_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_5__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_5__19_  (.A1(u_multiplier_STAGE1__0985_ ),
    .A2(u_multiplier_STAGE1__0984_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_5__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_5__20_  (.A(u_multiplier_STAGE1__0985_ ),
    .B(u_multiplier_STAGE1__0984_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_35_5__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_5__21_  (.A1(u_multiplier_STAGE1__0986_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_5__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_5__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_5__22_  (.A(u_multiplier_STAGE1__0986_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_5__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_35_5__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_5__23_  (.A1(u_multiplier_STAGE1__0987_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_5__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_5__24_  (.A(u_multiplier_STAGE1__0987_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_5__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_5__25_  (.A(u_multiplier_STAGE1_pp1_34_e42_5_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_5__16_ ),
    .ZN(u_multiplier_pp1_35 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_5__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_35_5__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_5__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_35_e42_5_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_35_5__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_35_5__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_35_5__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_35_5__17_ ),
    .ZN(u_multiplier_pp1_36 [8]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_35_6__18_  (.A(u_multiplier_STAGE1_pp1_34_e42_6_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_6__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_6__19_  (.A1(u_multiplier_STAGE1__0989_ ),
    .A2(u_multiplier_STAGE1__0988_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_6__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_6__20_  (.A(u_multiplier_STAGE1__0989_ ),
    .B(u_multiplier_STAGE1__0988_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_35_6__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_6__21_  (.A1(u_multiplier_STAGE1__0990_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_6__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_6__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_6__22_  (.A(u_multiplier_STAGE1__0990_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_6__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_35_6__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_6__23_  (.A1(u_multiplier_STAGE1__0991_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_6__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_6__24_  (.A(u_multiplier_STAGE1__0991_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_6__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_6__25_  (.A(u_multiplier_STAGE1_pp1_34_e42_6_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_6__16_ ),
    .ZN(u_multiplier_pp1_35 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_6__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_35_6__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_6__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_35_e42_6_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_35_6__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_35_6__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_35_6__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_35_6__17_ ),
    .ZN(u_multiplier_pp1_36 [7]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_36_1__18_  (.A(u_multiplier_STAGE1_pp1_35_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_1__19_  (.A1(u_multiplier_STAGE1__0995_ ),
    .A2(u_multiplier_STAGE1__0994_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_1__20_  (.A(u_multiplier_STAGE1__0995_ ),
    .B(u_multiplier_STAGE1__0994_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_36_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_1__21_  (.A1(u_multiplier_STAGE1__0996_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_1__22_  (.A(u_multiplier_STAGE1__0996_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_36_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_1__23_  (.A1(u_multiplier_STAGE1__0997_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_1__24_  (.A(u_multiplier_STAGE1__0997_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_1__25_  (.A(u_multiplier_STAGE1_pp1_35_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_1__16_ ),
    .ZN(u_multiplier_pp1_36 [5]));
 NAND2_X2 u_multiplier_STAGE1_E_4_2_pp_36_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_36_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_36_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_36_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_36_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_36_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_36_1__17_ ),
    .ZN(u_multiplier_pp1_37 [11]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_36_2__18_  (.A(u_multiplier_STAGE1_pp1_35_e42_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_2__19_  (.A1(u_multiplier_STAGE1__0999_ ),
    .A2(u_multiplier_STAGE1__0998_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_2__20_  (.A(u_multiplier_STAGE1__0999_ ),
    .B(u_multiplier_STAGE1__0998_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_36_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_2__21_  (.A1(u_multiplier_STAGE1__1000_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_2__22_  (.A(u_multiplier_STAGE1__1000_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_36_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_2__23_  (.A1(u_multiplier_STAGE1__1001_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_2__24_  (.A(u_multiplier_STAGE1__1001_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_2__25_  (.A(u_multiplier_STAGE1_pp1_35_e42_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_2__16_ ),
    .ZN(u_multiplier_pp1_36 [4]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_36_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_36_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_36_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_36_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_36_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_36_2__17_ ),
    .ZN(u_multiplier_pp1_37 [10]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_36_3__18_  (.A(u_multiplier_STAGE1_pp1_35_e42_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_3__19_  (.A1(u_multiplier_STAGE1__1003_ ),
    .A2(u_multiplier_STAGE1__1002_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_3__20_  (.A(u_multiplier_STAGE1__1003_ ),
    .B(u_multiplier_STAGE1__1002_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_36_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_3__21_  (.A1(u_multiplier_STAGE1__1004_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_3__22_  (.A(u_multiplier_STAGE1__1004_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_36_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_3__23_  (.A1(u_multiplier_STAGE1__1005_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_3__24_  (.A(u_multiplier_STAGE1__1005_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_3__25_  (.A(u_multiplier_STAGE1_pp1_35_e42_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_3__16_ ),
    .ZN(u_multiplier_pp1_36 [3]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_36_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_36_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_36_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_36_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_36_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_36_3__17_ ),
    .ZN(u_multiplier_pp1_37 [9]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_36_4__18_  (.A(u_multiplier_STAGE1_pp1_35_e42_4_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_4__19_  (.A1(u_multiplier_STAGE1__1007_ ),
    .A2(u_multiplier_STAGE1__1006_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_4__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_4__20_  (.A(u_multiplier_STAGE1__1007_ ),
    .B(u_multiplier_STAGE1__1006_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_36_4__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_4__21_  (.A1(u_multiplier_STAGE1__1008_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_4__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_4__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_4__22_  (.A(u_multiplier_STAGE1__1008_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_4__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_36_4__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_4__23_  (.A1(u_multiplier_STAGE1__1009_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_4__24_  (.A(u_multiplier_STAGE1__1009_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_4__25_  (.A(u_multiplier_STAGE1_pp1_35_e42_4_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_4__16_ ),
    .ZN(u_multiplier_pp1_36 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_4__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_36_4__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_4__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_36_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_36_4__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_36_4__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_36_4__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_36_4__17_ ),
    .ZN(u_multiplier_pp1_37 [8]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_36_5__18_  (.A(u_multiplier_STAGE1_pp1_35_e42_5_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_5__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_5__19_  (.A1(u_multiplier_STAGE1__1011_ ),
    .A2(u_multiplier_STAGE1__1010_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_5__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_5__20_  (.A(u_multiplier_STAGE1__1011_ ),
    .B(u_multiplier_STAGE1__1010_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_36_5__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_5__21_  (.A1(u_multiplier_STAGE1__1012_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_5__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_5__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_5__22_  (.A(u_multiplier_STAGE1__1012_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_5__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_36_5__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_5__23_  (.A1(u_multiplier_STAGE1__1013_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_5__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_5__24_  (.A(u_multiplier_STAGE1__1013_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_5__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_5__25_  (.A(u_multiplier_STAGE1_pp1_35_e42_5_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_5__16_ ),
    .ZN(u_multiplier_pp1_36 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_5__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_36_5__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_5__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_36_e42_5_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_36_5__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_36_5__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_36_5__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_36_5__17_ ),
    .ZN(u_multiplier_pp1_37 [7]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_36_6__18_  (.A(u_multiplier_STAGE1_pp1_35_e42_6_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_6__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_6__19_  (.A1(u_multiplier_STAGE1__1015_ ),
    .A2(u_multiplier_STAGE1__1014_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_6__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_6__20_  (.A(u_multiplier_STAGE1__1015_ ),
    .B(u_multiplier_STAGE1__1014_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_36_6__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_6__21_  (.A1(u_multiplier_STAGE1__1016_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_6__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_6__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_6__22_  (.A(u_multiplier_STAGE1__1016_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_6__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_36_6__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_6__23_  (.A1(u_multiplier_STAGE1__1017_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_6__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_6__24_  (.A(u_multiplier_STAGE1__1017_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_6__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_6__25_  (.A(u_multiplier_STAGE1_pp1_35_e42_6_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_6__16_ ),
    .ZN(u_multiplier_pp1_36 [0]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_6__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_36_6__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_6__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_36_e42_6_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_36_6__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_36_6__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_36_6__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_36_6__17_ ),
    .ZN(u_multiplier_pp1_37 [6]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_37_1__18_  (.A(u_multiplier_STAGE1_pp1_36_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_1__19_  (.A1(u_multiplier_STAGE1__1019_ ),
    .A2(u_multiplier_STAGE1__1018_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_1__20_  (.A(u_multiplier_STAGE1__1019_ ),
    .B(u_multiplier_STAGE1__1018_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_37_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_1__21_  (.A1(u_multiplier_STAGE1__1020_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_1__22_  (.A(u_multiplier_STAGE1__1020_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_37_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_1__23_  (.A1(u_multiplier_STAGE1__1021_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_1__24_  (.A(u_multiplier_STAGE1__1021_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_1__25_  (.A(u_multiplier_STAGE1_pp1_36_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_1__16_ ),
    .ZN(u_multiplier_pp1_37 [5]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_37_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_37_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_37_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_37_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_37_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_37_1__17_ ),
    .ZN(u_multiplier_pp1_38 [10]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_37_2__18_  (.A(u_multiplier_STAGE1_pp1_36_e42_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_2__19_  (.A1(u_multiplier_STAGE1__1023_ ),
    .A2(u_multiplier_STAGE1__1022_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_2__20_  (.A(u_multiplier_STAGE1__1023_ ),
    .B(u_multiplier_STAGE1__1022_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_37_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_2__21_  (.A1(u_multiplier_STAGE1__1024_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_2__22_  (.A(u_multiplier_STAGE1__1024_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_37_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_2__23_  (.A1(u_multiplier_STAGE1__1025_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_2__24_  (.A(u_multiplier_STAGE1__1025_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_2__25_  (.A(u_multiplier_STAGE1_pp1_36_e42_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_2__16_ ),
    .ZN(u_multiplier_pp1_37 [4]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_37_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_37_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_37_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_37_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_37_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_37_2__17_ ),
    .ZN(u_multiplier_pp1_38 [9]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_37_3__18_  (.A(u_multiplier_STAGE1_pp1_36_e42_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_3__19_  (.A1(u_multiplier_STAGE1__1027_ ),
    .A2(u_multiplier_STAGE1__1026_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_3__20_  (.A(u_multiplier_STAGE1__1027_ ),
    .B(u_multiplier_STAGE1__1026_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_37_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_3__21_  (.A1(u_multiplier_STAGE1__1028_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_3__22_  (.A(u_multiplier_STAGE1__1028_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_37_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_3__23_  (.A1(u_multiplier_STAGE1__1029_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_3__24_  (.A(u_multiplier_STAGE1__1029_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_3__25_  (.A(u_multiplier_STAGE1_pp1_36_e42_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_3__16_ ),
    .ZN(u_multiplier_pp1_37 [3]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_37_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_37_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_37_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_37_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_37_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_37_3__17_ ),
    .ZN(u_multiplier_pp1_38 [8]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_37_4__18_  (.A(u_multiplier_STAGE1_pp1_36_e42_4_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_4__19_  (.A1(u_multiplier_STAGE1__1031_ ),
    .A2(u_multiplier_STAGE1__1030_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_4__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_4__20_  (.A(u_multiplier_STAGE1__1031_ ),
    .B(u_multiplier_STAGE1__1030_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_37_4__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_4__21_  (.A1(u_multiplier_STAGE1__1032_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_4__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_4__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_4__22_  (.A(u_multiplier_STAGE1__1032_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_4__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_37_4__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_4__23_  (.A1(u_multiplier_STAGE1__1033_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_4__24_  (.A(u_multiplier_STAGE1__1033_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_4__25_  (.A(u_multiplier_STAGE1_pp1_36_e42_4_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_4__16_ ),
    .ZN(u_multiplier_pp1_37 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_4__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_37_4__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_4__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_37_e42_4_cout ));
 OAI21_X1 u_multiplier_STAGE1_E_4_2_pp_37_4__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_37_4__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_37_4__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_37_4__17_ ),
    .ZN(u_multiplier_pp1_38 [7]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_37_5__18_  (.A(u_multiplier_STAGE1_pp1_36_e42_5_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_5__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_5__19_  (.A1(u_multiplier_STAGE1__1035_ ),
    .A2(u_multiplier_STAGE1__1034_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_5__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_5__20_  (.A(u_multiplier_STAGE1__1035_ ),
    .B(u_multiplier_STAGE1__1034_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_37_5__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_5__21_  (.A1(u_multiplier_STAGE1__1036_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_5__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_5__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_5__22_  (.A(u_multiplier_STAGE1__1036_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_5__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_37_5__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_5__23_  (.A1(u_multiplier_STAGE1__1037_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_5__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_5__24_  (.A(u_multiplier_STAGE1__1037_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_5__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_5__25_  (.A(u_multiplier_STAGE1_pp1_36_e42_5_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_5__16_ ),
    .ZN(u_multiplier_pp1_37 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_5__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_37_5__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_5__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_37_e42_5_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_37_5__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_37_5__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_37_5__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_37_5__17_ ),
    .ZN(u_multiplier_pp1_38 [6]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_38_1__18_  (.A(u_multiplier_STAGE1_pp1_37_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_1__19_  (.A1(u_multiplier_STAGE1__1041_ ),
    .A2(u_multiplier_STAGE1__1040_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_1__20_  (.A(u_multiplier_STAGE1__1041_ ),
    .B(u_multiplier_STAGE1__1040_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_38_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_1__21_  (.A1(u_multiplier_STAGE1__1042_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_1__22_  (.A(u_multiplier_STAGE1__1042_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_38_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_1__23_  (.A1(u_multiplier_STAGE1__1043_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_1__24_  (.A(u_multiplier_STAGE1__1043_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_1__25_  (.A(u_multiplier_STAGE1_pp1_37_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_1__16_ ),
    .ZN(u_multiplier_pp1_38 [4]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_38_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_38_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_38_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_38_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_38_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_38_1__17_ ),
    .ZN(u_multiplier_pp1_39 [9]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_38_2__18_  (.A(u_multiplier_STAGE1_pp1_37_e42_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_2__19_  (.A1(u_multiplier_STAGE1__1045_ ),
    .A2(u_multiplier_STAGE1__1044_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_2__20_  (.A(u_multiplier_STAGE1__1045_ ),
    .B(u_multiplier_STAGE1__1044_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_38_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_2__21_  (.A1(u_multiplier_STAGE1__1046_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_2__22_  (.A(u_multiplier_STAGE1__1046_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_38_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_2__23_  (.A1(u_multiplier_STAGE1__1047_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_2__24_  (.A(u_multiplier_STAGE1__1047_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_2__25_  (.A(u_multiplier_STAGE1_pp1_37_e42_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_2__16_ ),
    .ZN(u_multiplier_pp1_38 [3]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_38_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_38_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_38_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_38_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_38_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_38_2__17_ ),
    .ZN(u_multiplier_pp1_39 [8]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_38_3__18_  (.A(u_multiplier_STAGE1_pp1_37_e42_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_3__19_  (.A1(u_multiplier_STAGE1__1049_ ),
    .A2(u_multiplier_STAGE1__1048_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_3__20_  (.A(u_multiplier_STAGE1__1049_ ),
    .B(u_multiplier_STAGE1__1048_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_38_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_3__21_  (.A1(u_multiplier_STAGE1__1050_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_3__22_  (.A(u_multiplier_STAGE1__1050_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_38_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_3__23_  (.A1(u_multiplier_STAGE1__1051_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_3__24_  (.A(u_multiplier_STAGE1__1051_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_3__25_  (.A(u_multiplier_STAGE1_pp1_37_e42_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_3__16_ ),
    .ZN(u_multiplier_pp1_38 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_38_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_38_e42_3_cout ));
 OAI21_X1 u_multiplier_STAGE1_E_4_2_pp_38_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_38_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_38_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_38_3__17_ ),
    .ZN(u_multiplier_pp1_39 [7]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_38_4__18_  (.A(u_multiplier_STAGE1_pp1_37_e42_4_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_4__19_  (.A1(u_multiplier_STAGE1__1053_ ),
    .A2(u_multiplier_STAGE1__1052_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_4__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_4__20_  (.A(u_multiplier_STAGE1__1053_ ),
    .B(u_multiplier_STAGE1__1052_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_38_4__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_4__21_  (.A1(u_multiplier_STAGE1__1054_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_4__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_4__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_4__22_  (.A(u_multiplier_STAGE1__1054_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_4__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_38_4__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_4__23_  (.A1(u_multiplier_STAGE1__1055_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_4__24_  (.A(u_multiplier_STAGE1__1055_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_4__25_  (.A(u_multiplier_STAGE1_pp1_37_e42_4_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_4__16_ ),
    .ZN(u_multiplier_pp1_38 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_4__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_38_4__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_4__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_38_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_38_4__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_38_4__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_38_4__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_38_4__17_ ),
    .ZN(u_multiplier_pp1_39 [6]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_38_5__18_  (.A(u_multiplier_STAGE1_pp1_37_e42_5_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_5__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_5__19_  (.A1(u_multiplier_STAGE1__1057_ ),
    .A2(u_multiplier_STAGE1__1056_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_5__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_5__20_  (.A(u_multiplier_STAGE1__1057_ ),
    .B(u_multiplier_STAGE1__1056_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_38_5__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_5__21_  (.A1(u_multiplier_STAGE1__1058_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_5__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_5__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_5__22_  (.A(u_multiplier_STAGE1__1058_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_5__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_38_5__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_5__23_  (.A1(u_multiplier_STAGE1__1059_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_5__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_5__24_  (.A(u_multiplier_STAGE1__1059_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_5__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_5__25_  (.A(u_multiplier_STAGE1_pp1_37_e42_5_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_5__16_ ),
    .ZN(u_multiplier_pp1_38 [0]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_5__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_38_5__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_5__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_38_e42_5_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_38_5__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_38_5__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_38_5__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_38_5__17_ ),
    .ZN(u_multiplier_pp1_39 [5]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_39_1__18_  (.A(u_multiplier_STAGE1_pp1_38_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_1__19_  (.A1(u_multiplier_STAGE1__1061_ ),
    .A2(u_multiplier_STAGE1__1060_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_1__20_  (.A(u_multiplier_STAGE1__1061_ ),
    .B(u_multiplier_STAGE1__1060_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_39_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_1__21_  (.A1(u_multiplier_STAGE1__1062_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_39_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_1__22_  (.A(u_multiplier_STAGE1__1062_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_39_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_39_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_1__23_  (.A1(u_multiplier_STAGE1__1063_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_39_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_1__24_  (.A(u_multiplier_STAGE1__1063_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_39_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_1__25_  (.A(u_multiplier_STAGE1_pp1_38_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_39_1__16_ ),
    .ZN(u_multiplier_pp1_39 [4]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_39_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_39_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_39_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_39_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_39_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_39_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_39_1__17_ ),
    .ZN(u_multiplier_pp1_40 [8]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_39_2__18_  (.A(u_multiplier_STAGE1_pp1_38_e42_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_2__19_  (.A1(u_multiplier_STAGE1__1065_ ),
    .A2(u_multiplier_STAGE1__1064_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_2__20_  (.A(u_multiplier_STAGE1__1065_ ),
    .B(u_multiplier_STAGE1__1064_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_39_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_2__21_  (.A1(u_multiplier_STAGE1__1066_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_39_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_2__22_  (.A(u_multiplier_STAGE1__1066_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_39_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_39_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_2__23_  (.A1(u_multiplier_STAGE1__1067_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_39_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_2__24_  (.A(u_multiplier_STAGE1__1067_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_39_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_2__25_  (.A(u_multiplier_STAGE1_pp1_38_e42_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_39_2__16_ ),
    .ZN(u_multiplier_pp1_39 [3]));
 NAND2_X2 u_multiplier_STAGE1_E_4_2_pp_39_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_39_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_39_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_39_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_39_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_39_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_39_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_39_2__17_ ),
    .ZN(u_multiplier_pp1_40 [7]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_39_3__18_  (.A(u_multiplier_STAGE1_pp1_38_e42_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_3__19_  (.A1(u_multiplier_STAGE1__1069_ ),
    .A2(u_multiplier_STAGE1__1068_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_3__20_  (.A(u_multiplier_STAGE1__1069_ ),
    .B(u_multiplier_STAGE1__1068_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_39_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_3__21_  (.A1(u_multiplier_STAGE1__1070_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_39_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_3__22_  (.A(u_multiplier_STAGE1__1070_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_39_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_39_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_3__23_  (.A1(u_multiplier_STAGE1__1071_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_39_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_3__24_  (.A(u_multiplier_STAGE1__1071_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_39_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_3__25_  (.A(u_multiplier_STAGE1_pp1_38_e42_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_39_3__16_ ),
    .ZN(u_multiplier_pp1_39 [2]));
 NAND2_X2 u_multiplier_STAGE1_E_4_2_pp_39_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_39_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_39_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_39_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_39_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_39_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_39_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_39_3__17_ ),
    .ZN(u_multiplier_pp1_40 [6]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_39_4__18_  (.A(u_multiplier_STAGE1_pp1_38_e42_4_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_4__19_  (.A1(u_multiplier_STAGE1__1073_ ),
    .A2(u_multiplier_STAGE1__1072_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_4__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_4__20_  (.A(u_multiplier_STAGE1__1073_ ),
    .B(u_multiplier_STAGE1__1072_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_39_4__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_4__21_  (.A1(u_multiplier_STAGE1__1074_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_39_4__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_4__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_4__22_  (.A(u_multiplier_STAGE1__1074_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_39_4__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_39_4__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_4__23_  (.A1(u_multiplier_STAGE1__1075_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_39_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_4__24_  (.A(u_multiplier_STAGE1__1075_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_39_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_4__25_  (.A(u_multiplier_STAGE1_pp1_38_e42_4_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_39_4__16_ ),
    .ZN(u_multiplier_pp1_39 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_4__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_39_4__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_39_4__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_39_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_39_4__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_39_4__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_39_4__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_39_4__17_ ),
    .ZN(u_multiplier_pp1_40 [5]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_40_1__18_  (.A(u_multiplier_STAGE1_pp1_39_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_1__19_  (.A1(u_multiplier_STAGE1__1079_ ),
    .A2(u_multiplier_STAGE1__1078_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_1__20_  (.A(u_multiplier_STAGE1__1079_ ),
    .B(u_multiplier_STAGE1__1078_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_40_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_1__21_  (.A1(u_multiplier_STAGE1__1080_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_40_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_1__22_  (.A(u_multiplier_STAGE1__1080_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_40_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_40_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_1__23_  (.A1(u_multiplier_STAGE1__1081_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_40_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_1__24_  (.A(u_multiplier_STAGE1__1081_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_40_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_1__25_  (.A(u_multiplier_STAGE1_pp1_39_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_40_1__16_ ),
    .ZN(u_multiplier_pp1_40 [3]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_40_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_40_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_40_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE1_E_4_2_pp_40_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_40_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_40_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_40_1__17_ ),
    .ZN(u_multiplier_pp1_41 [7]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_40_2__18_  (.A(u_multiplier_STAGE1_pp1_39_e42_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_2__19_  (.A1(u_multiplier_STAGE1__1083_ ),
    .A2(u_multiplier_STAGE1__1082_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_2__20_  (.A(u_multiplier_STAGE1__1083_ ),
    .B(u_multiplier_STAGE1__1082_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_40_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_2__21_  (.A1(u_multiplier_STAGE1__1084_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_40_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_2__22_  (.A(u_multiplier_STAGE1__1084_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_40_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_40_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_2__23_  (.A1(u_multiplier_STAGE1__1085_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_40_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_2__24_  (.A(u_multiplier_STAGE1__1085_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_40_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_2__25_  (.A(u_multiplier_STAGE1_pp1_39_e42_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_40_2__16_ ),
    .ZN(u_multiplier_pp1_40 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_40_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_40_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_40_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_40_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_40_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_40_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_40_2__17_ ),
    .ZN(u_multiplier_pp1_41 [6]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_40_3__18_  (.A(u_multiplier_STAGE1_pp1_39_e42_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_3__19_  (.A1(u_multiplier_STAGE1__1087_ ),
    .A2(u_multiplier_STAGE1__1086_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_3__20_  (.A(u_multiplier_STAGE1__1087_ ),
    .B(u_multiplier_STAGE1__1086_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_40_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_3__21_  (.A1(u_multiplier_STAGE1__1088_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_40_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_3__22_  (.A(u_multiplier_STAGE1__1088_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_40_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_40_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_3__23_  (.A1(u_multiplier_STAGE1__1089_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_40_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_3__24_  (.A(u_multiplier_STAGE1__1089_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_40_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_3__25_  (.A(u_multiplier_STAGE1_pp1_39_e42_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_40_3__16_ ),
    .ZN(u_multiplier_pp1_40 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_40_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_40_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_40_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_40_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_40_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_40_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_40_3__17_ ),
    .ZN(u_multiplier_pp1_41 [5]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_40_4__18_  (.A(u_multiplier_STAGE1_pp1_39_e42_4_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_4__19_  (.A1(u_multiplier_STAGE1__1091_ ),
    .A2(u_multiplier_STAGE1__1090_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_4__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_4__20_  (.A(u_multiplier_STAGE1__1091_ ),
    .B(u_multiplier_STAGE1__1090_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_40_4__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_4__21_  (.A1(u_multiplier_STAGE1__1092_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_40_4__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_4__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_4__22_  (.A(u_multiplier_STAGE1__1092_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_40_4__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_40_4__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_4__23_  (.A1(u_multiplier_STAGE1__1093_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_40_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_4__24_  (.A(u_multiplier_STAGE1__1093_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_40_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_4__25_  (.A(u_multiplier_STAGE1_pp1_39_e42_4_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_40_4__16_ ),
    .ZN(u_multiplier_pp1_40 [0]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_4__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_40_4__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_40_4__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_40_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_40_4__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_40_4__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_40_4__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_40_4__17_ ),
    .ZN(u_multiplier_pp1_41 [4]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_41_1__18_  (.A(u_multiplier_STAGE1_pp1_40_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_41_1__19_  (.A1(u_multiplier_STAGE1__1095_ ),
    .A2(u_multiplier_STAGE1__1094_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_41_1__20_  (.A(u_multiplier_STAGE1__1095_ ),
    .B(u_multiplier_STAGE1__1094_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_41_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_41_1__21_  (.A1(u_multiplier_STAGE1__1096_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_41_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_41_1__22_  (.A(u_multiplier_STAGE1__1096_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_41_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_41_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_41_1__23_  (.A1(u_multiplier_STAGE1__1097_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_41_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_41_1__24_  (.A(u_multiplier_STAGE1__1097_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_41_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_41_1__25_  (.A(u_multiplier_STAGE1_pp1_40_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_41_1__16_ ),
    .ZN(u_multiplier_pp1_41 [3]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_41_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_41_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_41_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_41_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_41_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_41_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_41_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_41_1__17_ ),
    .ZN(u_multiplier_pp1_42 [6]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_41_2__18_  (.A(u_multiplier_STAGE1_pp1_40_e42_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_41_2__19_  (.A1(u_multiplier_STAGE1__1099_ ),
    .A2(u_multiplier_STAGE1__1098_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_41_2__20_  (.A(u_multiplier_STAGE1__1099_ ),
    .B(u_multiplier_STAGE1__1098_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_41_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_41_2__21_  (.A1(u_multiplier_STAGE1__1100_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_41_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_41_2__22_  (.A(u_multiplier_STAGE1__1100_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_41_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_41_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_41_2__23_  (.A1(u_multiplier_STAGE1__1101_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_41_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_41_2__24_  (.A(u_multiplier_STAGE1__1101_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_41_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_41_2__25_  (.A(u_multiplier_STAGE1_pp1_40_e42_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_41_2__16_ ),
    .ZN(u_multiplier_pp1_41 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_41_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_41_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_41_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_41_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_41_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_41_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_41_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_41_2__17_ ),
    .ZN(u_multiplier_pp1_42 [5]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_41_3__18_  (.A(u_multiplier_STAGE1_pp1_40_e42_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_41_3__19_  (.A1(u_multiplier_STAGE1__1103_ ),
    .A2(u_multiplier_STAGE1__1102_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_41_3__20_  (.A(u_multiplier_STAGE1__1103_ ),
    .B(u_multiplier_STAGE1__1102_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_41_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_41_3__21_  (.A1(u_multiplier_STAGE1__1104_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_41_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_41_3__22_  (.A(u_multiplier_STAGE1__1104_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_41_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_41_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_41_3__23_  (.A1(u_multiplier_STAGE1__1105_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_41_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_41_3__24_  (.A(u_multiplier_STAGE1__1105_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_41_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_41_3__25_  (.A(u_multiplier_STAGE1_pp1_40_e42_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_41_3__16_ ),
    .ZN(u_multiplier_pp1_41 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_41_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_41_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_41_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_41_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_41_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_41_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_41_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_41_3__17_ ),
    .ZN(u_multiplier_pp1_42 [4]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_42_1__18_  (.A(u_multiplier_STAGE1_pp1_41_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_42_1__19_  (.A1(u_multiplier_STAGE1__1109_ ),
    .A2(u_multiplier_STAGE1__1108_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_42_1__20_  (.A(u_multiplier_STAGE1__1109_ ),
    .B(u_multiplier_STAGE1__1108_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_42_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_42_1__21_  (.A1(u_multiplier_STAGE1__1110_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_42_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_42_1__22_  (.A(u_multiplier_STAGE1__1110_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_42_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_42_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_42_1__23_  (.A1(u_multiplier_STAGE1__1111_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_42_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_42_1__24_  (.A(u_multiplier_STAGE1__1111_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_42_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_42_1__25_  (.A(u_multiplier_STAGE1_pp1_41_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_42_1__16_ ),
    .ZN(u_multiplier_pp1_42 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_42_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_42_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_42_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_42_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_42_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_42_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_42_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_42_1__17_ ),
    .ZN(u_multiplier_pp1_43 [5]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_42_2__18_  (.A(u_multiplier_STAGE1_pp1_41_e42_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_42_2__19_  (.A1(u_multiplier_STAGE1__1113_ ),
    .A2(u_multiplier_STAGE1__1112_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_42_2__20_  (.A(u_multiplier_STAGE1__1113_ ),
    .B(u_multiplier_STAGE1__1112_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_42_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_42_2__21_  (.A1(u_multiplier_STAGE1__1114_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_42_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_42_2__22_  (.A(u_multiplier_STAGE1__1114_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_42_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_42_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_42_2__23_  (.A1(u_multiplier_STAGE1__1115_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_42_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_42_2__24_  (.A(u_multiplier_STAGE1__1115_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_42_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_42_2__25_  (.A(u_multiplier_STAGE1_pp1_41_e42_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_42_2__16_ ),
    .ZN(u_multiplier_pp1_42 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_42_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_42_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_42_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_42_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_42_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_42_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_42_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_42_2__17_ ),
    .ZN(u_multiplier_pp1_43 [4]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_42_3__18_  (.A(u_multiplier_STAGE1_pp1_41_e42_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_42_3__19_  (.A1(u_multiplier_STAGE1__1117_ ),
    .A2(u_multiplier_STAGE1__1116_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_42_3__20_  (.A(u_multiplier_STAGE1__1117_ ),
    .B(u_multiplier_STAGE1__1116_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_42_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_42_3__21_  (.A1(u_multiplier_STAGE1__1118_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_42_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_42_3__22_  (.A(u_multiplier_STAGE1__1118_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_42_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_42_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_42_3__23_  (.A1(u_multiplier_STAGE1__1119_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_42_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_42_3__24_  (.A(u_multiplier_STAGE1__1119_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_42_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_42_3__25_  (.A(u_multiplier_STAGE1_pp1_41_e42_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_42_3__16_ ),
    .ZN(u_multiplier_pp1_42 [0]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_42_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_42_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_42_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_42_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_42_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_42_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_42_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_42_3__17_ ),
    .ZN(u_multiplier_pp1_43 [3]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_43_1__18_  (.A(u_multiplier_STAGE1_pp1_42_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_43_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_43_1__19_  (.A1(u_multiplier_STAGE1__1121_ ),
    .A2(u_multiplier_STAGE1__1120_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_43_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_43_1__20_  (.A(u_multiplier_STAGE1__1121_ ),
    .B(u_multiplier_STAGE1__1120_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_43_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_43_1__21_  (.A1(u_multiplier_STAGE1__1122_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_43_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_43_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_43_1__22_  (.A(u_multiplier_STAGE1__1122_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_43_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_43_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_43_1__23_  (.A1(u_multiplier_STAGE1__1123_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_43_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_43_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_43_1__24_  (.A(u_multiplier_STAGE1__1123_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_43_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_43_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_43_1__25_  (.A(u_multiplier_STAGE1_pp1_42_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_43_1__16_ ),
    .ZN(u_multiplier_pp1_43 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_43_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_43_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_43_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_43_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_43_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_43_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_43_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_43_1__17_ ),
    .ZN(u_multiplier_pp1_44 [4]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_43_2__18_  (.A(u_multiplier_STAGE1_pp1_42_e42_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_43_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_43_2__19_  (.A1(u_multiplier_STAGE1__1125_ ),
    .A2(u_multiplier_STAGE1__1124_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_43_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_43_2__20_  (.A(u_multiplier_STAGE1__1125_ ),
    .B(u_multiplier_STAGE1__1124_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_43_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_43_2__21_  (.A1(u_multiplier_STAGE1__1126_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_43_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_43_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_43_2__22_  (.A(u_multiplier_STAGE1__1126_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_43_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_43_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_43_2__23_  (.A1(u_multiplier_STAGE1__1127_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_43_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_43_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_43_2__24_  (.A(u_multiplier_STAGE1__1127_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_43_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_43_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_43_2__25_  (.A(u_multiplier_STAGE1_pp1_42_e42_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_43_2__16_ ),
    .ZN(u_multiplier_pp1_43 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_43_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_43_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_43_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_43_e42_2_cout ));
 OAI21_X1 u_multiplier_STAGE1_E_4_2_pp_43_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_43_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_43_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_43_2__17_ ),
    .ZN(u_multiplier_pp1_44 [3]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_44_1__18_  (.A(u_multiplier_STAGE1_pp1_43_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_44_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_44_1__19_  (.A1(u_multiplier_STAGE1__1131_ ),
    .A2(u_multiplier_STAGE1__1130_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_44_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_44_1__20_  (.A(u_multiplier_STAGE1__1131_ ),
    .B(u_multiplier_STAGE1__1130_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_44_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_44_1__21_  (.A1(u_multiplier_STAGE1__1132_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_44_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_44_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_44_1__22_  (.A(u_multiplier_STAGE1__1132_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_44_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_44_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_44_1__23_  (.A1(u_multiplier_STAGE1__1133_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_44_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_44_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_44_1__24_  (.A(u_multiplier_STAGE1__1133_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_44_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_44_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_44_1__25_  (.A(u_multiplier_STAGE1_pp1_43_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_44_1__16_ ),
    .ZN(u_multiplier_pp1_44 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_44_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_44_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_44_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_44_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_44_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_44_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_44_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_44_1__17_ ),
    .ZN(u_multiplier_pp1_45 [3]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_44_2__18_  (.A(u_multiplier_STAGE1_pp1_43_e42_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_44_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_44_2__19_  (.A1(u_multiplier_STAGE1__1135_ ),
    .A2(u_multiplier_STAGE1__1134_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_44_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_44_2__20_  (.A(u_multiplier_STAGE1__1135_ ),
    .B(u_multiplier_STAGE1__1134_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_44_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_44_2__21_  (.A1(u_multiplier_STAGE1__1136_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_44_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_44_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_44_2__22_  (.A(u_multiplier_STAGE1__1136_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_44_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_44_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_44_2__23_  (.A1(u_multiplier_STAGE1__1137_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_44_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_44_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_44_2__24_  (.A(u_multiplier_STAGE1__1137_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_44_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_44_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_44_2__25_  (.A(u_multiplier_STAGE1_pp1_43_e42_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_44_2__16_ ),
    .ZN(u_multiplier_pp1_44 [0]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_44_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_44_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_44_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_44_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_44_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_44_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_44_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_44_2__17_ ),
    .ZN(u_multiplier_pp1_45 [2]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_45_1__18_  (.A(u_multiplier_STAGE1_pp1_44_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_45_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_45_1__19_  (.A1(u_multiplier_STAGE1__1139_ ),
    .A2(u_multiplier_STAGE1__1138_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_45_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_45_1__20_  (.A(u_multiplier_STAGE1__1139_ ),
    .B(u_multiplier_STAGE1__1138_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_45_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_45_1__21_  (.A1(u_multiplier_STAGE1__1140_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_45_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_45_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_45_1__22_  (.A(u_multiplier_STAGE1__1140_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_45_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_45_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_45_1__23_  (.A1(u_multiplier_STAGE1__1141_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_45_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_45_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_45_1__24_  (.A(u_multiplier_STAGE1__1141_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_45_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_45_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_45_1__25_  (.A(u_multiplier_STAGE1_pp1_44_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_45_1__16_ ),
    .ZN(u_multiplier_pp1_45 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_45_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_45_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_45_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_45_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_45_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_45_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_45_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_45_1__17_ ),
    .ZN(u_multiplier_pp1_46 [2]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_46_1__18_  (.A(u_multiplier_STAGE1_pp1_45_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_46_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_46_1__19_  (.A1(u_multiplier_STAGE1__1145_ ),
    .A2(u_multiplier_STAGE1__1144_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_46_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_46_1__20_  (.A(u_multiplier_STAGE1__1145_ ),
    .B(u_multiplier_STAGE1__1144_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_46_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_46_1__21_  (.A1(u_multiplier_STAGE1__1146_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_46_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_46_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_46_1__22_  (.A(u_multiplier_STAGE1__1146_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_46_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_46_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_46_1__23_  (.A1(u_multiplier_STAGE1__1147_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_46_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_46_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_46_1__24_  (.A(u_multiplier_STAGE1__1147_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_46_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_46_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_46_1__25_  (.A(u_multiplier_STAGE1_pp1_45_e42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_46_1__16_ ),
    .ZN(u_multiplier_pp1_46 [0]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_46_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_46_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_46_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_46_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_46_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_46_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_46_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_46_1__17_ ),
    .ZN(u_multiplier_pp1_47 [1]));
 INV_X1 u_multiplier_STAGE1_Full_adder_pp_33_1__12_  (.A(u_multiplier_STAGE1_pp1_32_e42_8_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_33_1__08_ ));
 NAND3_X2 u_multiplier_STAGE1_Full_adder_pp_33_1__13_  (.A1(u_multiplier_STAGE1__0939_ ),
    .A2(u_multiplier_STAGE1__0938_ ),
    .A3(u_multiplier_STAGE1_pp1_32_e42_8_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_33_1__09_ ));
 NOR2_X4 u_multiplier_STAGE1_Full_adder_pp_33_1__14_  (.A1(u_multiplier_STAGE1__0939_ ),
    .A2(u_multiplier_STAGE1__0938_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_33_1__10_ ));
 AOI21_X2 u_multiplier_STAGE1_Full_adder_pp_33_1__15_  (.A(u_multiplier_STAGE1_pp1_32_e42_8_cout ),
    .B1(u_multiplier_STAGE1__0938_ ),
    .B2(u_multiplier_STAGE1__0939_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_33_1__11_ ));
 NOR2_X4 u_multiplier_STAGE1_Full_adder_pp_33_1__16_  (.A1(u_multiplier_STAGE1_Full_adder_pp_33_1__10_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_33_1__11_ ),
    .ZN(u_multiplier_pp1_34 [7]));
 AOI22_X4 u_multiplier_STAGE1_Full_adder_pp_33_1__17_  (.A1(u_multiplier_STAGE1_Full_adder_pp_33_1__08_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_33_1__10_ ),
    .B1(u_multiplier_pp1_34 [7]),
    .B2(u_multiplier_STAGE1_Full_adder_pp_33_1__09_ ),
    .ZN(u_multiplier_pp1_33 [0]));
 INV_X1 u_multiplier_STAGE1_Full_adder_pp_35_1__12_  (.A(u_multiplier_STAGE1_pp1_34_e42_7_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_35_1__08_ ));
 NAND3_X2 u_multiplier_STAGE1_Full_adder_pp_35_1__13_  (.A1(u_multiplier_STAGE1__0993_ ),
    .A2(u_multiplier_STAGE1__0992_ ),
    .A3(u_multiplier_STAGE1_pp1_34_e42_7_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_35_1__09_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_35_1__14_  (.A1(u_multiplier_STAGE1__0993_ ),
    .A2(u_multiplier_STAGE1__0992_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_35_1__10_ ));
 AOI21_X1 u_multiplier_STAGE1_Full_adder_pp_35_1__15_  (.A(u_multiplier_STAGE1_pp1_34_e42_7_cout ),
    .B1(u_multiplier_STAGE1__0992_ ),
    .B2(u_multiplier_STAGE1__0993_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_35_1__11_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_35_1__16_  (.A1(u_multiplier_STAGE1_Full_adder_pp_35_1__10_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_35_1__11_ ),
    .ZN(u_multiplier_pp1_36 [6]));
 AOI22_X4 u_multiplier_STAGE1_Full_adder_pp_35_1__17_  (.A1(u_multiplier_STAGE1_Full_adder_pp_35_1__08_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_35_1__10_ ),
    .B1(u_multiplier_pp1_36 [6]),
    .B2(u_multiplier_STAGE1_Full_adder_pp_35_1__09_ ),
    .ZN(u_multiplier_pp1_35 [0]));
 INV_X1 u_multiplier_STAGE1_Full_adder_pp_37_1__12_  (.A(u_multiplier_STAGE1_pp1_36_e42_6_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_37_1__08_ ));
 NAND3_X1 u_multiplier_STAGE1_Full_adder_pp_37_1__13_  (.A1(u_multiplier_STAGE1__1039_ ),
    .A2(u_multiplier_STAGE1__1038_ ),
    .A3(u_multiplier_STAGE1_pp1_36_e42_6_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_37_1__09_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_37_1__14_  (.A1(u_multiplier_STAGE1__1039_ ),
    .A2(u_multiplier_STAGE1__1038_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_37_1__10_ ));
 AOI21_X1 u_multiplier_STAGE1_Full_adder_pp_37_1__15_  (.A(u_multiplier_STAGE1_pp1_36_e42_6_cout ),
    .B1(u_multiplier_STAGE1__1038_ ),
    .B2(u_multiplier_STAGE1__1039_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_37_1__11_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_37_1__16_  (.A1(u_multiplier_STAGE1_Full_adder_pp_37_1__10_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_37_1__11_ ),
    .ZN(u_multiplier_pp1_38 [5]));
 AOI22_X2 u_multiplier_STAGE1_Full_adder_pp_37_1__17_  (.A1(u_multiplier_STAGE1_Full_adder_pp_37_1__08_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_37_1__10_ ),
    .B1(u_multiplier_pp1_38 [5]),
    .B2(u_multiplier_STAGE1_Full_adder_pp_37_1__09_ ),
    .ZN(u_multiplier_pp1_37 [0]));
 INV_X1 u_multiplier_STAGE1_Full_adder_pp_39_1__12_  (.A(u_multiplier_STAGE1_pp1_38_e42_5_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_39_1__08_ ));
 NAND3_X2 u_multiplier_STAGE1_Full_adder_pp_39_1__13_  (.A1(u_multiplier_STAGE1__1077_ ),
    .A2(u_multiplier_STAGE1__1076_ ),
    .A3(u_multiplier_STAGE1_pp1_38_e42_5_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_39_1__09_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_39_1__14_  (.A1(u_multiplier_STAGE1__1077_ ),
    .A2(u_multiplier_STAGE1__1076_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_39_1__10_ ));
 AOI21_X1 u_multiplier_STAGE1_Full_adder_pp_39_1__15_  (.A(u_multiplier_STAGE1_pp1_38_e42_5_cout ),
    .B1(u_multiplier_STAGE1__1076_ ),
    .B2(u_multiplier_STAGE1__1077_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_39_1__11_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_39_1__16_  (.A1(u_multiplier_STAGE1_Full_adder_pp_39_1__10_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_39_1__11_ ),
    .ZN(u_multiplier_pp1_40 [4]));
 AOI22_X4 u_multiplier_STAGE1_Full_adder_pp_39_1__17_  (.A1(u_multiplier_STAGE1_Full_adder_pp_39_1__08_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_39_1__10_ ),
    .B1(u_multiplier_pp1_40 [4]),
    .B2(u_multiplier_STAGE1_Full_adder_pp_39_1__09_ ),
    .ZN(u_multiplier_pp1_39 [0]));
 INV_X1 u_multiplier_STAGE1_Full_adder_pp_41_1__12_  (.A(u_multiplier_STAGE1_pp1_40_e42_4_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_41_1__08_ ));
 NAND3_X2 u_multiplier_STAGE1_Full_adder_pp_41_1__13_  (.A1(u_multiplier_STAGE1__1107_ ),
    .A2(u_multiplier_STAGE1__1106_ ),
    .A3(u_multiplier_STAGE1_pp1_40_e42_4_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_41_1__09_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_41_1__14_  (.A1(u_multiplier_STAGE1__1107_ ),
    .A2(u_multiplier_STAGE1__1106_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_41_1__10_ ));
 AOI21_X1 u_multiplier_STAGE1_Full_adder_pp_41_1__15_  (.A(u_multiplier_STAGE1_pp1_40_e42_4_cout ),
    .B1(u_multiplier_STAGE1__1106_ ),
    .B2(u_multiplier_STAGE1__1107_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_41_1__11_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_41_1__16_  (.A1(u_multiplier_STAGE1_Full_adder_pp_41_1__10_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_41_1__11_ ),
    .ZN(u_multiplier_pp1_42 [3]));
 AOI22_X4 u_multiplier_STAGE1_Full_adder_pp_41_1__17_  (.A1(u_multiplier_STAGE1_Full_adder_pp_41_1__08_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_41_1__10_ ),
    .B1(u_multiplier_pp1_42 [3]),
    .B2(u_multiplier_STAGE1_Full_adder_pp_41_1__09_ ),
    .ZN(u_multiplier_pp1_41 [0]));
 INV_X1 u_multiplier_STAGE1_Full_adder_pp_43_1__12_  (.A(u_multiplier_STAGE1_pp1_42_e42_3_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_43_1__08_ ));
 NAND3_X2 u_multiplier_STAGE1_Full_adder_pp_43_1__13_  (.A1(u_multiplier_STAGE1__1129_ ),
    .A2(u_multiplier_STAGE1__1128_ ),
    .A3(u_multiplier_STAGE1_pp1_42_e42_3_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_43_1__09_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_43_1__14_  (.A1(u_multiplier_STAGE1__1129_ ),
    .A2(u_multiplier_STAGE1__1128_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_43_1__10_ ));
 AOI21_X1 u_multiplier_STAGE1_Full_adder_pp_43_1__15_  (.A(u_multiplier_STAGE1_pp1_42_e42_3_cout ),
    .B1(u_multiplier_STAGE1__1128_ ),
    .B2(u_multiplier_STAGE1__1129_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_43_1__11_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_43_1__16_  (.A1(u_multiplier_STAGE1_Full_adder_pp_43_1__10_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_43_1__11_ ),
    .ZN(u_multiplier_pp1_44 [2]));
 AOI22_X4 u_multiplier_STAGE1_Full_adder_pp_43_1__17_  (.A1(u_multiplier_STAGE1_Full_adder_pp_43_1__08_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_43_1__10_ ),
    .B1(u_multiplier_pp1_44 [2]),
    .B2(u_multiplier_STAGE1_Full_adder_pp_43_1__09_ ),
    .ZN(u_multiplier_pp1_43 [0]));
 INV_X1 u_multiplier_STAGE1_Full_adder_pp_45_1__12_  (.A(u_multiplier_STAGE1_pp1_44_e42_2_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_45_1__08_ ));
 NAND3_X1 u_multiplier_STAGE1_Full_adder_pp_45_1__13_  (.A1(u_multiplier_STAGE1__1143_ ),
    .A2(u_multiplier_STAGE1__1142_ ),
    .A3(u_multiplier_STAGE1_pp1_44_e42_2_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_45_1__09_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_45_1__14_  (.A1(u_multiplier_STAGE1__1143_ ),
    .A2(u_multiplier_STAGE1__1142_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_45_1__10_ ));
 AOI21_X1 u_multiplier_STAGE1_Full_adder_pp_45_1__15_  (.A(u_multiplier_STAGE1_pp1_44_e42_2_cout ),
    .B1(u_multiplier_STAGE1__1142_ ),
    .B2(u_multiplier_STAGE1__1143_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_45_1__11_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_45_1__16_  (.A1(u_multiplier_STAGE1_Full_adder_pp_45_1__10_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_45_1__11_ ),
    .ZN(u_multiplier_pp1_46 [1]));
 AOI22_X2 u_multiplier_STAGE1_Full_adder_pp_45_1__17_  (.A1(u_multiplier_STAGE1_Full_adder_pp_45_1__08_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_45_1__10_ ),
    .B1(u_multiplier_pp1_46 [1]),
    .B2(u_multiplier_STAGE1_Full_adder_pp_45_1__09_ ),
    .ZN(u_multiplier_pp1_45 [0]));
 INV_X1 u_multiplier_STAGE1_Full_adder_pp_47_1__12_  (.A(u_multiplier_STAGE1_pp1_46_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_47_1__08_ ));
 NAND3_X2 u_multiplier_STAGE1_Full_adder_pp_47_1__13_  (.A1(u_multiplier_STAGE1__1149_ ),
    .A2(u_multiplier_STAGE1__1148_ ),
    .A3(u_multiplier_STAGE1_pp1_46_e42_1_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_47_1__09_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_47_1__14_  (.A1(u_multiplier_STAGE1__1149_ ),
    .A2(u_multiplier_STAGE1__1148_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_47_1__10_ ));
 AOI21_X1 u_multiplier_STAGE1_Full_adder_pp_47_1__15_  (.A(u_multiplier_STAGE1_pp1_46_e42_1_cout ),
    .B1(u_multiplier_STAGE1__1148_ ),
    .B2(u_multiplier_STAGE1__1149_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_47_1__11_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_47_1__16_  (.A1(u_multiplier_STAGE1_Full_adder_pp_47_1__10_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_47_1__11_ ),
    .ZN(u_multiplier_pp1_48 [0]));
 AOI22_X4 u_multiplier_STAGE1_Full_adder_pp_47_1__17_  (.A1(u_multiplier_STAGE1_Full_adder_pp_47_1__08_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_47_1__10_ ),
    .B1(u_multiplier_pp1_48 [0]),
    .B2(u_multiplier_STAGE1_Full_adder_pp_47_1__09_ ),
    .ZN(u_multiplier_pp1_47 [0]));
 AND2_X1 u_multiplier_STAGE1_Half_adder_pp_16_1__4_  (.A1(u_multiplier_STAGE1__0608_ ),
    .A2(u_multiplier_STAGE1__0607_ ),
    .ZN(u_multiplier_pp1_17 [1]));
 XOR2_X2 u_multiplier_STAGE1_Half_adder_pp_16_1__5_  (.A(u_multiplier_STAGE1__0608_ ),
    .B(u_multiplier_STAGE1__0607_ ),
    .Z(u_multiplier_pp1_16 [0]));
 AND2_X1 u_multiplier_STAGE1_Half_adder_pp_18_1__4_  (.A1(u_multiplier_STAGE1__0618_ ),
    .A2(u_multiplier_STAGE1__0617_ ),
    .ZN(u_multiplier_pp1_19 [2]));
 XOR2_X2 u_multiplier_STAGE1_Half_adder_pp_18_1__5_  (.A(u_multiplier_STAGE1__0618_ ),
    .B(u_multiplier_STAGE1__0617_ ),
    .Z(u_multiplier_pp1_18 [0]));
 AND2_X1 u_multiplier_STAGE1_Half_adder_pp_20_1__4_  (.A1(u_multiplier_STAGE1__0636_ ),
    .A2(u_multiplier_STAGE1__0635_ ),
    .ZN(u_multiplier_pp1_21 [3]));
 XOR2_X2 u_multiplier_STAGE1_Half_adder_pp_20_1__5_  (.A(u_multiplier_STAGE1__0636_ ),
    .B(u_multiplier_STAGE1__0635_ ),
    .Z(u_multiplier_pp1_20 [0]));
 AND2_X1 u_multiplier_STAGE1_Half_adder_pp_22_1__4_  (.A1(u_multiplier_STAGE1__0662_ ),
    .A2(u_multiplier_STAGE1__0661_ ),
    .ZN(u_multiplier_pp1_23 [4]));
 XOR2_X2 u_multiplier_STAGE1_Half_adder_pp_22_1__5_  (.A(u_multiplier_STAGE1__0662_ ),
    .B(u_multiplier_STAGE1__0661_ ),
    .Z(u_multiplier_pp1_22 [0]));
 AND2_X1 u_multiplier_STAGE1_Half_adder_pp_24_1__4_  (.A1(u_multiplier_STAGE1__0696_ ),
    .A2(u_multiplier_STAGE1__0695_ ),
    .ZN(u_multiplier_pp1_25 [5]));
 XOR2_X2 u_multiplier_STAGE1_Half_adder_pp_24_1__5_  (.A(u_multiplier_STAGE1__0696_ ),
    .B(u_multiplier_STAGE1__0695_ ),
    .Z(u_multiplier_pp1_24 [0]));
 AND2_X1 u_multiplier_STAGE1_Half_adder_pp_26_1__4_  (.A1(u_multiplier_STAGE1__0738_ ),
    .A2(u_multiplier_STAGE1__0737_ ),
    .ZN(u_multiplier_pp1_27 [6]));
 XOR2_X2 u_multiplier_STAGE1_Half_adder_pp_26_1__5_  (.A(u_multiplier_STAGE1__0738_ ),
    .B(u_multiplier_STAGE1__0737_ ),
    .Z(u_multiplier_pp1_26 [0]));
 AND2_X1 u_multiplier_STAGE1_Half_adder_pp_28_1__4_  (.A1(u_multiplier_STAGE1__0788_ ),
    .A2(u_multiplier_STAGE1__0787_ ),
    .ZN(u_multiplier_pp1_29 [7]));
 XOR2_X2 u_multiplier_STAGE1_Half_adder_pp_28_1__5_  (.A(u_multiplier_STAGE1__0788_ ),
    .B(u_multiplier_STAGE1__0787_ ),
    .Z(u_multiplier_pp1_28 [0]));
 AND2_X1 u_multiplier_STAGE1_Half_adder_pp_30_1__4_  (.A1(u_multiplier_STAGE1__0846_ ),
    .A2(u_multiplier_STAGE1__0845_ ),
    .ZN(u_multiplier_pp1_31 [8]));
 XOR2_X2 u_multiplier_STAGE1_Half_adder_pp_30_1__5_  (.A(u_multiplier_STAGE1__0846_ ),
    .B(u_multiplier_STAGE1__0845_ ),
    .Z(u_multiplier_pp1_30 [0]));
 AND2_X1 u_multiplier_STAGE1__1631_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[0]),
    .ZN(u_multiplier_pp3_0 ));
 AND2_X1 u_multiplier_STAGE1__1632_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[1]),
    .ZN(u_multiplier_pp3_1 [0]));
 AND2_X1 u_multiplier_STAGE1__1633_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[1]),
    .ZN(u_multiplier_pp3_1 [1]));
 AND2_X1 u_multiplier_STAGE1__1634_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[2]),
    .ZN(u_multiplier_pp3_2 [0]));
 AND2_X1 u_multiplier_STAGE1__1635_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[1]),
    .ZN(u_multiplier_pp3_2 [1]));
 AND2_X1 u_multiplier_STAGE1__1636_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[2]),
    .ZN(u_multiplier_pp3_2 [2]));
 AND2_X1 u_multiplier_STAGE1__1637_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[3]),
    .ZN(u_multiplier_pp3_3 [0]));
 AND2_X1 u_multiplier_STAGE1__1638_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[2]),
    .ZN(u_multiplier_pp3_3 [1]));
 AND2_X1 u_multiplier_STAGE1__1639_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[2]),
    .ZN(u_multiplier_pp3_3 [2]));
 AND2_X1 u_multiplier_STAGE1__1640_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[3]),
    .ZN(u_multiplier_pp3_3 [3]));
 AND2_X1 u_multiplier_STAGE1__1641_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[4]),
    .ZN(u_multiplier_pp3_4 [1]));
 AND2_X1 u_multiplier_STAGE1__1642_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[3]),
    .ZN(u_multiplier_pp3_4 [2]));
 AND2_X1 u_multiplier_STAGE1__1643_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[2]),
    .ZN(u_multiplier_pp3_4 [3]));
 AND2_X1 u_multiplier_STAGE1__1644_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[3]),
    .ZN(u_multiplier_pp2_4 [1]));
 AND2_X1 u_multiplier_STAGE1__1645_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[4]),
    .ZN(u_multiplier_pp2_4 [0]));
 AND2_X1 u_multiplier_STAGE1__1646_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[5]),
    .ZN(u_multiplier_pp3_5 [2]));
 AND2_X1 u_multiplier_STAGE1__1647_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[4]),
    .ZN(u_multiplier_pp3_5 [3]));
 AND2_X1 u_multiplier_STAGE1__1648_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[3]),
    .ZN(u_multiplier_pp2_5 [3]));
 AND2_X1 u_multiplier_STAGE1__1649_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[3]),
    .ZN(u_multiplier_pp2_5 [2]));
 AND2_X1 u_multiplier_STAGE1__1650_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[4]),
    .ZN(u_multiplier_pp2_5 [1]));
 AND2_X1 u_multiplier_STAGE1__1651_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[5]),
    .ZN(u_multiplier_pp2_5 [0]));
 AND2_X1 u_multiplier_STAGE1__1652_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[6]),
    .ZN(u_multiplier_pp3_6 [3]));
 AND2_X1 u_multiplier_STAGE1__1653_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[5]),
    .ZN(u_multiplier_pp2_6 [5]));
 AND2_X1 u_multiplier_STAGE1__1654_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[4]),
    .ZN(u_multiplier_pp2_6 [4]));
 AND2_X1 u_multiplier_STAGE1__1655_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[3]),
    .ZN(u_multiplier_pp2_6 [3]));
 AND2_X1 u_multiplier_STAGE1__1656_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[4]),
    .ZN(u_multiplier_pp2_6 [2]));
 AND2_X1 u_multiplier_STAGE1__1657_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[5]),
    .ZN(u_multiplier_pp2_6 [1]));
 AND2_X1 u_multiplier_STAGE1__1658_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[6]),
    .ZN(u_multiplier_pp2_6 [0]));
 AND2_X1 u_multiplier_STAGE1__1659_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[7]),
    .ZN(u_multiplier_pp2_7 [7]));
 AND2_X1 u_multiplier_STAGE1__1660_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[6]),
    .ZN(u_multiplier_pp2_7 [6]));
 AND2_X1 u_multiplier_STAGE1__1661_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[5]),
    .ZN(u_multiplier_pp2_7 [5]));
 AND2_X1 u_multiplier_STAGE1__1662_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[4]),
    .ZN(u_multiplier_pp2_7 [4]));
 AND2_X1 u_multiplier_STAGE1__1663_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[4]),
    .ZN(u_multiplier_pp2_7 [3]));
 AND2_X1 u_multiplier_STAGE1__1664_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[5]),
    .ZN(u_multiplier_pp2_7 [2]));
 AND2_X1 u_multiplier_STAGE1__1665_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[6]),
    .ZN(u_multiplier_pp2_7 [1]));
 AND2_X1 u_multiplier_STAGE1__1666_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[7]),
    .ZN(u_multiplier_pp2_7 [0]));
 AND2_X1 u_multiplier_STAGE1__1667_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[8]),
    .ZN(u_multiplier_pp1_8 [0]));
 AND2_X1 u_multiplier_STAGE1__1668_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[7]),
    .ZN(u_multiplier_pp1_8 [1]));
 AND2_X1 u_multiplier_STAGE1__1669_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[6]),
    .ZN(u_multiplier_pp2_8 [7]));
 AND2_X1 u_multiplier_STAGE1__1670_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[5]),
    .ZN(u_multiplier_pp2_8 [6]));
 AND2_X1 u_multiplier_STAGE1__1671_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[4]),
    .ZN(u_multiplier_pp2_8 [5]));
 AND2_X1 u_multiplier_STAGE1__1672_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[5]),
    .ZN(u_multiplier_pp2_8 [4]));
 AND2_X1 u_multiplier_STAGE1__1673_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[6]),
    .ZN(u_multiplier_pp2_8 [3]));
 AND2_X1 u_multiplier_STAGE1__1674_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[7]),
    .ZN(u_multiplier_pp2_8 [2]));
 AND2_X1 u_multiplier_STAGE1__1675_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[8]),
    .ZN(u_multiplier_pp2_8 [1]));
 AND2_X1 u_multiplier_STAGE1__1676_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[9]),
    .ZN(u_multiplier_pp1_9 [0]));
 AND2_X1 u_multiplier_STAGE1__1677_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[8]),
    .ZN(u_multiplier_pp1_9 [1]));
 AND2_X1 u_multiplier_STAGE1__1678_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[7]),
    .ZN(u_multiplier_pp1_9 [2]));
 AND2_X1 u_multiplier_STAGE1__1679_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[6]),
    .ZN(u_multiplier_pp1_9 [3]));
 AND2_X1 u_multiplier_STAGE1__1680_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[5]),
    .ZN(u_multiplier_pp2_9 [7]));
 AND2_X1 u_multiplier_STAGE1__1681_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[5]),
    .ZN(u_multiplier_pp2_9 [6]));
 AND2_X1 u_multiplier_STAGE1__1682_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[6]),
    .ZN(u_multiplier_pp2_9 [5]));
 AND2_X1 u_multiplier_STAGE1__1683_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[7]),
    .ZN(u_multiplier_pp2_9 [4]));
 AND2_X1 u_multiplier_STAGE1__1684_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[8]),
    .ZN(u_multiplier_pp2_9 [3]));
 AND2_X1 u_multiplier_STAGE1__1685_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[9]),
    .ZN(u_multiplier_pp2_9 [2]));
 AND2_X1 u_multiplier_STAGE1__1686_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[10]),
    .ZN(u_multiplier_pp1_10 [0]));
 AND2_X1 u_multiplier_STAGE1__1687_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[9]),
    .ZN(u_multiplier_pp1_10 [1]));
 AND2_X1 u_multiplier_STAGE1__1688_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[8]),
    .ZN(u_multiplier_pp1_10 [2]));
 AND2_X1 u_multiplier_STAGE1__1689_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[7]),
    .ZN(u_multiplier_pp1_10 [3]));
 AND2_X1 u_multiplier_STAGE1__1690_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[6]),
    .ZN(u_multiplier_pp1_10 [4]));
 AND2_X1 u_multiplier_STAGE1__1691_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[5]),
    .ZN(u_multiplier_pp1_10 [5]));
 AND2_X1 u_multiplier_STAGE1__1692_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[6]),
    .ZN(u_multiplier_pp2_10 [7]));
 AND2_X1 u_multiplier_STAGE1__1693_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[7]),
    .ZN(u_multiplier_pp2_10 [6]));
 AND2_X1 u_multiplier_STAGE1__1694_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[8]),
    .ZN(u_multiplier_pp2_10 [5]));
 AND2_X1 u_multiplier_STAGE1__1695_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[9]),
    .ZN(u_multiplier_pp2_10 [4]));
 AND2_X1 u_multiplier_STAGE1__1696_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[10]),
    .ZN(u_multiplier_pp2_10 [3]));
 AND2_X1 u_multiplier_STAGE1__1697_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[11]),
    .ZN(u_multiplier_pp1_11 [0]));
 AND2_X1 u_multiplier_STAGE1__1698_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[10]),
    .ZN(u_multiplier_pp1_11 [1]));
 AND2_X1 u_multiplier_STAGE1__1699_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[9]),
    .ZN(u_multiplier_pp1_11 [2]));
 AND2_X1 u_multiplier_STAGE1__1700_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[8]),
    .ZN(u_multiplier_pp1_11 [3]));
 AND2_X1 u_multiplier_STAGE1__1701_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[7]),
    .ZN(u_multiplier_pp1_11 [4]));
 AND2_X1 u_multiplier_STAGE1__1702_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[6]),
    .ZN(u_multiplier_pp1_11 [5]));
 AND2_X1 u_multiplier_STAGE1__1703_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[6]),
    .ZN(u_multiplier_pp1_11 [6]));
 AND2_X1 u_multiplier_STAGE1__1704_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[7]),
    .ZN(u_multiplier_pp1_11 [7]));
 AND2_X1 u_multiplier_STAGE1__1705_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[8]),
    .ZN(u_multiplier_pp2_11 [7]));
 AND2_X1 u_multiplier_STAGE1__1706_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[9]),
    .ZN(u_multiplier_pp2_11 [6]));
 AND2_X1 u_multiplier_STAGE1__1707_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[10]),
    .ZN(u_multiplier_pp2_11 [5]));
 AND2_X1 u_multiplier_STAGE1__1708_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[11]),
    .ZN(u_multiplier_pp2_11 [4]));
 AND2_X1 u_multiplier_STAGE1__1709_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[12]),
    .ZN(u_multiplier_pp1_12 [0]));
 AND2_X1 u_multiplier_STAGE1__1710_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[11]),
    .ZN(u_multiplier_pp1_12 [1]));
 AND2_X1 u_multiplier_STAGE1__1711_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[10]),
    .ZN(u_multiplier_pp1_12 [2]));
 AND2_X1 u_multiplier_STAGE1__1712_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[9]),
    .ZN(u_multiplier_pp1_12 [3]));
 AND2_X1 u_multiplier_STAGE1__1713_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[8]),
    .ZN(u_multiplier_pp1_12 [4]));
 AND2_X1 u_multiplier_STAGE1__1714_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[7]),
    .ZN(u_multiplier_pp1_12 [5]));
 AND2_X1 u_multiplier_STAGE1__1715_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[6]),
    .ZN(u_multiplier_pp1_12 [6]));
 AND2_X1 u_multiplier_STAGE1__1716_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[7]),
    .ZN(u_multiplier_pp1_12 [7]));
 AND2_X1 u_multiplier_STAGE1__1717_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[8]),
    .ZN(u_multiplier_pp1_12 [8]));
 AND2_X1 u_multiplier_STAGE1__1718_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[9]),
    .ZN(u_multiplier_pp1_12 [9]));
 AND2_X1 u_multiplier_STAGE1__1719_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[10]),
    .ZN(u_multiplier_pp2_12 [7]));
 AND2_X1 u_multiplier_STAGE1__1720_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[11]),
    .ZN(u_multiplier_pp2_12 [6]));
 AND2_X1 u_multiplier_STAGE1__1721_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[12]),
    .ZN(u_multiplier_pp2_12 [5]));
 AND2_X1 u_multiplier_STAGE1__1722_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[13]),
    .ZN(u_multiplier_pp1_13 [0]));
 AND2_X1 u_multiplier_STAGE1__1723_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[12]),
    .ZN(u_multiplier_pp1_13 [1]));
 AND2_X1 u_multiplier_STAGE1__1724_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[11]),
    .ZN(u_multiplier_pp1_13 [2]));
 AND2_X1 u_multiplier_STAGE1__1725_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[10]),
    .ZN(u_multiplier_pp1_13 [3]));
 AND2_X1 u_multiplier_STAGE1__1726_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[9]),
    .ZN(u_multiplier_pp1_13 [4]));
 AND2_X1 u_multiplier_STAGE1__1727_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[8]),
    .ZN(u_multiplier_pp1_13 [5]));
 AND2_X1 u_multiplier_STAGE1__1728_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[7]),
    .ZN(u_multiplier_pp1_13 [6]));
 AND2_X1 u_multiplier_STAGE1__1729_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[7]),
    .ZN(u_multiplier_pp1_13 [7]));
 AND2_X1 u_multiplier_STAGE1__1730_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[8]),
    .ZN(u_multiplier_pp1_13 [8]));
 AND2_X1 u_multiplier_STAGE1__1731_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[9]),
    .ZN(u_multiplier_pp1_13 [9]));
 AND2_X1 u_multiplier_STAGE1__1732_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[10]),
    .ZN(u_multiplier_pp1_13 [10]));
 AND2_X1 u_multiplier_STAGE1__1733_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[11]),
    .ZN(u_multiplier_pp1_13 [11]));
 AND2_X1 u_multiplier_STAGE1__1734_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[12]),
    .ZN(u_multiplier_pp2_13 [7]));
 AND2_X1 u_multiplier_STAGE1__1735_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_pp2_13 [6]));
 AND2_X1 u_multiplier_STAGE1__1736_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_pp1_14 [0]));
 AND2_X1 u_multiplier_STAGE1__1737_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[13]),
    .ZN(u_multiplier_pp1_14 [1]));
 AND2_X1 u_multiplier_STAGE1__1738_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[12]),
    .ZN(u_multiplier_pp1_14 [2]));
 AND2_X1 u_multiplier_STAGE1__1739_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[11]),
    .ZN(u_multiplier_pp1_14 [3]));
 AND2_X1 u_multiplier_STAGE1__1740_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[10]),
    .ZN(u_multiplier_pp1_14 [4]));
 AND2_X1 u_multiplier_STAGE1__1741_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[9]),
    .ZN(u_multiplier_pp1_14 [5]));
 AND2_X1 u_multiplier_STAGE1__1742_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[8]),
    .ZN(u_multiplier_pp1_14 [6]));
 AND2_X1 u_multiplier_STAGE1__1743_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[7]),
    .ZN(u_multiplier_pp1_14 [7]));
 AND2_X1 u_multiplier_STAGE1__1744_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[8]),
    .ZN(u_multiplier_pp1_14 [8]));
 AND2_X1 u_multiplier_STAGE1__1745_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[9]),
    .ZN(u_multiplier_pp1_14 [9]));
 AND2_X1 u_multiplier_STAGE1__1746_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[10]),
    .ZN(u_multiplier_pp1_14 [10]));
 AND2_X1 u_multiplier_STAGE1__1747_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[11]),
    .ZN(u_multiplier_pp1_14 [11]));
 AND2_X1 u_multiplier_STAGE1__1748_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[12]),
    .ZN(u_multiplier_pp1_14 [12]));
 AND2_X1 u_multiplier_STAGE1__1749_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_pp1_14 [13]));
 AND2_X1 u_multiplier_STAGE1__1750_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_pp2_14 [7]));
 AND2_X1 u_multiplier_STAGE1__1751_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_pp1_15 [0]));
 AND2_X1 u_multiplier_STAGE1__1752_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_pp1_15 [1]));
 AND2_X1 u_multiplier_STAGE1__1753_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[13]),
    .ZN(u_multiplier_pp1_15 [2]));
 AND2_X1 u_multiplier_STAGE1__1754_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[12]),
    .ZN(u_multiplier_pp1_15 [3]));
 AND2_X1 u_multiplier_STAGE1__1755_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[11]),
    .ZN(u_multiplier_pp1_15 [4]));
 AND2_X1 u_multiplier_STAGE1__1756_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[10]),
    .ZN(u_multiplier_pp1_15 [5]));
 AND2_X1 u_multiplier_STAGE1__1757_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[9]),
    .ZN(u_multiplier_pp1_15 [6]));
 AND2_X1 u_multiplier_STAGE1__1758_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[8]),
    .ZN(u_multiplier_pp1_15 [7]));
 AND2_X1 u_multiplier_STAGE1__1759_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[8]),
    .ZN(u_multiplier_pp1_15 [8]));
 AND2_X1 u_multiplier_STAGE1__1760_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[9]),
    .ZN(u_multiplier_pp1_15 [9]));
 AND2_X1 u_multiplier_STAGE1__1761_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[10]),
    .ZN(u_multiplier_pp1_15 [10]));
 AND2_X1 u_multiplier_STAGE1__1762_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[11]),
    .ZN(u_multiplier_pp1_15 [11]));
 AND2_X1 u_multiplier_STAGE1__1763_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[12]),
    .ZN(u_multiplier_pp1_15 [12]));
 AND2_X1 u_multiplier_STAGE1__1764_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_pp1_15 [13]));
 AND2_X1 u_multiplier_STAGE1__1765_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_pp1_15 [14]));
 AND2_X1 u_multiplier_STAGE1__1766_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_pp1_15 [15]));
 AND2_X1 u_multiplier_STAGE1__1767_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_STAGE1__0607_ ));
 AND2_X1 u_multiplier_STAGE1__1768_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_STAGE1__0608_ ));
 AND2_X1 u_multiplier_STAGE1__1769_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_pp1_16 [1]));
 AND2_X1 u_multiplier_STAGE1__1770_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_pp1_16 [2]));
 AND2_X1 u_multiplier_STAGE1__1771_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_pp1_16 [3]));
 AND2_X1 u_multiplier_STAGE1__1772_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[13]),
    .ZN(u_multiplier_pp1_16 [4]));
 AND2_X1 u_multiplier_STAGE1__1773_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[12]),
    .ZN(u_multiplier_pp1_16 [5]));
 AND2_X1 u_multiplier_STAGE1__1774_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[11]),
    .ZN(u_multiplier_pp1_16 [6]));
 AND2_X1 u_multiplier_STAGE1__1775_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[10]),
    .ZN(u_multiplier_pp1_16 [7]));
 AND2_X1 u_multiplier_STAGE1__1776_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[9]),
    .ZN(u_multiplier_pp1_16 [8]));
 AND2_X1 u_multiplier_STAGE1__1777_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[8]),
    .ZN(u_multiplier_pp1_16 [9]));
 AND2_X1 u_multiplier_STAGE1__1778_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[9]),
    .ZN(u_multiplier_pp1_16 [10]));
 AND2_X1 u_multiplier_STAGE1__1779_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[10]),
    .ZN(u_multiplier_pp1_16 [11]));
 AND2_X1 u_multiplier_STAGE1__1780_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[11]),
    .ZN(u_multiplier_pp1_16 [12]));
 AND2_X1 u_multiplier_STAGE1__1781_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[12]),
    .ZN(u_multiplier_pp1_16 [13]));
 AND2_X1 u_multiplier_STAGE1__1782_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_pp1_16 [14]));
 AND2_X1 u_multiplier_STAGE1__1783_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_pp1_16 [15]));
 AND2_X1 u_multiplier_STAGE1__1784_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0609_ ));
 AND2_X1 u_multiplier_STAGE1__1785_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_STAGE1__0610_ ));
 AND2_X1 u_multiplier_STAGE1__1786_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_STAGE1__0611_ ));
 AND2_X1 u_multiplier_STAGE1__1787_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_STAGE1__0612_ ));
 AND2_X1 u_multiplier_STAGE1__1788_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_pp1_17 [2]));
 AND2_X1 u_multiplier_STAGE1__1789_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_pp1_17 [3]));
 AND2_X1 u_multiplier_STAGE1__1790_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_pp1_17 [4]));
 AND2_X1 u_multiplier_STAGE1__1791_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_pp1_17 [5]));
 AND2_X1 u_multiplier_STAGE1__1792_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[13]),
    .ZN(u_multiplier_pp1_17 [6]));
 AND2_X1 u_multiplier_STAGE1__1793_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[12]),
    .ZN(u_multiplier_pp1_17 [7]));
 AND2_X1 u_multiplier_STAGE1__1794_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[11]),
    .ZN(u_multiplier_pp1_17 [8]));
 AND2_X1 u_multiplier_STAGE1__1795_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[10]),
    .ZN(u_multiplier_pp1_17 [9]));
 AND2_X1 u_multiplier_STAGE1__1796_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[9]),
    .ZN(u_multiplier_pp1_17 [10]));
 AND2_X1 u_multiplier_STAGE1__1797_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[9]),
    .ZN(u_multiplier_pp1_17 [11]));
 AND2_X1 u_multiplier_STAGE1__1798_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[10]),
    .ZN(u_multiplier_pp1_17 [12]));
 AND2_X1 u_multiplier_STAGE1__1799_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[11]),
    .ZN(u_multiplier_pp1_17 [13]));
 AND2_X1 u_multiplier_STAGE1__1800_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[12]),
    .ZN(u_multiplier_pp1_17 [14]));
 AND2_X1 u_multiplier_STAGE1__1801_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_pp1_17 [15]));
 AND2_X1 u_multiplier_STAGE1__1802_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0613_ ));
 AND2_X1 u_multiplier_STAGE1__1803_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0614_ ));
 AND2_X1 u_multiplier_STAGE1__1804_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_STAGE1__0615_ ));
 AND2_X1 u_multiplier_STAGE1__1805_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_STAGE1__0616_ ));
 AND2_X1 u_multiplier_STAGE1__1806_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_STAGE1__0617_ ));
 AND2_X1 u_multiplier_STAGE1__1807_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_STAGE1__0618_ ));
 AND2_X1 u_multiplier_STAGE1__1808_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_pp1_18 [3]));
 AND2_X1 u_multiplier_STAGE1__1809_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_pp1_18 [4]));
 AND2_X1 u_multiplier_STAGE1__1810_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_pp1_18 [5]));
 AND2_X1 u_multiplier_STAGE1__1811_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_pp1_18 [6]));
 AND2_X1 u_multiplier_STAGE1__1812_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_pp1_18 [7]));
 AND2_X1 u_multiplier_STAGE1__1813_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[13]),
    .ZN(u_multiplier_pp1_18 [8]));
 AND2_X1 u_multiplier_STAGE1__1814_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[12]),
    .ZN(u_multiplier_pp1_18 [9]));
 AND2_X1 u_multiplier_STAGE1__1815_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[11]),
    .ZN(u_multiplier_pp1_18 [10]));
 AND2_X1 u_multiplier_STAGE1__1816_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[10]),
    .ZN(u_multiplier_pp1_18 [11]));
 AND2_X1 u_multiplier_STAGE1__1817_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[9]),
    .ZN(u_multiplier_pp1_18 [12]));
 AND2_X1 u_multiplier_STAGE1__1818_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[10]),
    .ZN(u_multiplier_pp1_18 [13]));
 AND2_X1 u_multiplier_STAGE1__1819_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[11]),
    .ZN(u_multiplier_pp1_18 [14]));
 AND2_X1 u_multiplier_STAGE1__1820_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[12]),
    .ZN(u_multiplier_pp1_18 [15]));
 AND2_X1 u_multiplier_STAGE1__1821_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0619_ ));
 AND2_X1 u_multiplier_STAGE1__1822_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0620_ ));
 AND2_X1 u_multiplier_STAGE1__1823_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0621_ ));
 AND2_X1 u_multiplier_STAGE1__1824_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_STAGE1__0622_ ));
 AND2_X1 u_multiplier_STAGE1__1825_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_STAGE1__0623_ ));
 AND2_X1 u_multiplier_STAGE1__1826_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_STAGE1__0624_ ));
 AND2_X1 u_multiplier_STAGE1__1827_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_STAGE1__0625_ ));
 AND2_X1 u_multiplier_STAGE1__1828_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[12]),
    .ZN(u_multiplier_STAGE1__0626_ ));
 AND2_X1 u_multiplier_STAGE1__1829_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_pp1_19 [4]));
 AND2_X1 u_multiplier_STAGE1__1830_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_pp1_19 [5]));
 AND2_X1 u_multiplier_STAGE1__1831_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_pp1_19 [6]));
 AND2_X1 u_multiplier_STAGE1__1832_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_pp1_19 [7]));
 AND2_X1 u_multiplier_STAGE1__1833_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_pp1_19 [8]));
 AND2_X1 u_multiplier_STAGE1__1834_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_pp1_19 [9]));
 AND2_X1 u_multiplier_STAGE1__1835_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[13]),
    .ZN(u_multiplier_pp1_19 [10]));
 AND2_X1 u_multiplier_STAGE1__1836_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[12]),
    .ZN(u_multiplier_pp1_19 [11]));
 AND2_X1 u_multiplier_STAGE1__1837_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[11]),
    .ZN(u_multiplier_pp1_19 [12]));
 AND2_X1 u_multiplier_STAGE1__1838_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[10]),
    .ZN(u_multiplier_pp1_19 [13]));
 AND2_X1 u_multiplier_STAGE1__1839_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[10]),
    .ZN(u_multiplier_pp1_19 [14]));
 AND2_X1 u_multiplier_STAGE1__1840_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[11]),
    .ZN(u_multiplier_pp1_19 [15]));
 AND2_X1 u_multiplier_STAGE1__1841_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__0627_ ));
 AND2_X1 u_multiplier_STAGE1__1842_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0628_ ));
 AND2_X1 u_multiplier_STAGE1__1843_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0629_ ));
 AND2_X1 u_multiplier_STAGE1__1844_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0630_ ));
 AND2_X1 u_multiplier_STAGE1__1845_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_STAGE1__0631_ ));
 AND2_X1 u_multiplier_STAGE1__1846_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_STAGE1__0632_ ));
 AND2_X1 u_multiplier_STAGE1__1847_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_STAGE1__0633_ ));
 AND2_X1 u_multiplier_STAGE1__1848_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_STAGE1__0634_ ));
 AND2_X1 u_multiplier_STAGE1__1849_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[12]),
    .ZN(u_multiplier_STAGE1__0635_ ));
 AND2_X1 u_multiplier_STAGE1__1850_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[11]),
    .ZN(u_multiplier_STAGE1__0636_ ));
 AND2_X1 u_multiplier_STAGE1__1851_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_pp1_20 [5]));
 AND2_X1 u_multiplier_STAGE1__1852_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_pp1_20 [6]));
 AND2_X1 u_multiplier_STAGE1__1853_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_pp1_20 [7]));
 AND2_X1 u_multiplier_STAGE1__1854_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_pp1_20 [8]));
 AND2_X1 u_multiplier_STAGE1__1855_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_pp1_20 [9]));
 AND2_X1 u_multiplier_STAGE1__1856_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_pp1_20 [10]));
 AND2_X1 u_multiplier_STAGE1__1857_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_pp1_20 [11]));
 AND2_X1 u_multiplier_STAGE1__1858_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[13]),
    .ZN(u_multiplier_pp1_20 [12]));
 AND2_X1 u_multiplier_STAGE1__1859_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[12]),
    .ZN(u_multiplier_pp1_20 [13]));
 AND2_X1 u_multiplier_STAGE1__1860_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[11]),
    .ZN(u_multiplier_pp1_20 [14]));
 AND2_X1 u_multiplier_STAGE1__1861_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[10]),
    .ZN(u_multiplier_pp1_20 [15]));
 AND2_X1 u_multiplier_STAGE1__1862_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__0637_ ));
 AND2_X1 u_multiplier_STAGE1__1863_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__0638_ ));
 AND2_X1 u_multiplier_STAGE1__1864_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0639_ ));
 AND2_X1 u_multiplier_STAGE1__1865_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0640_ ));
 AND2_X1 u_multiplier_STAGE1__1866_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0641_ ));
 AND2_X1 u_multiplier_STAGE1__1867_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_STAGE1__0642_ ));
 AND2_X1 u_multiplier_STAGE1__1868_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_STAGE1__0643_ ));
 AND2_X1 u_multiplier_STAGE1__1869_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_STAGE1__0644_ ));
 AND2_X1 u_multiplier_STAGE1__1870_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_STAGE1__0645_ ));
 AND2_X1 u_multiplier_STAGE1__1871_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[12]),
    .ZN(u_multiplier_STAGE1__0646_ ));
 AND2_X1 u_multiplier_STAGE1__1872_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[11]),
    .ZN(u_multiplier_STAGE1__0647_ ));
 AND2_X1 u_multiplier_STAGE1__1873_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[11]),
    .ZN(u_multiplier_STAGE1__0648_ ));
 AND2_X1 u_multiplier_STAGE1__1874_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_pp1_21 [6]));
 AND2_X1 u_multiplier_STAGE1__1875_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_pp1_21 [7]));
 AND2_X1 u_multiplier_STAGE1__1876_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_pp1_21 [8]));
 AND2_X1 u_multiplier_STAGE1__1877_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_pp1_21 [9]));
 AND2_X1 u_multiplier_STAGE1__1878_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_pp1_21 [10]));
 AND2_X1 u_multiplier_STAGE1__1879_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_pp1_21 [11]));
 AND2_X1 u_multiplier_STAGE1__1880_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_pp1_21 [12]));
 AND2_X1 u_multiplier_STAGE1__1881_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_pp1_21 [13]));
 AND2_X1 u_multiplier_STAGE1__1882_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[13]),
    .ZN(u_multiplier_pp1_21 [14]));
 AND2_X1 u_multiplier_STAGE1__1883_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[12]),
    .ZN(u_multiplier_pp1_21 [15]));
 AND2_X1 u_multiplier_STAGE1__1884_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__0649_ ));
 AND2_X1 u_multiplier_STAGE1__1885_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__0650_ ));
 AND2_X1 u_multiplier_STAGE1__1886_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__0651_ ));
 AND2_X1 u_multiplier_STAGE1__1887_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0652_ ));
 AND2_X1 u_multiplier_STAGE1__1888_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0653_ ));
 AND2_X1 u_multiplier_STAGE1__1889_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0654_ ));
 AND2_X1 u_multiplier_STAGE1__1890_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_STAGE1__0655_ ));
 AND2_X1 u_multiplier_STAGE1__1891_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_STAGE1__0656_ ));
 AND2_X1 u_multiplier_STAGE1__1892_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_STAGE1__0657_ ));
 AND2_X1 u_multiplier_STAGE1__1893_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_STAGE1__0658_ ));
 AND2_X1 u_multiplier_STAGE1__1894_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[12]),
    .ZN(u_multiplier_STAGE1__0659_ ));
 AND2_X1 u_multiplier_STAGE1__1895_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[11]),
    .ZN(u_multiplier_STAGE1__0660_ ));
 AND2_X1 u_multiplier_STAGE1__1896_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[12]),
    .ZN(u_multiplier_STAGE1__0661_ ));
 AND2_X1 u_multiplier_STAGE1__1897_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[13]),
    .ZN(u_multiplier_STAGE1__0662_ ));
 AND2_X1 u_multiplier_STAGE1__1898_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_pp1_22 [7]));
 AND2_X1 u_multiplier_STAGE1__1899_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_pp1_22 [8]));
 AND2_X1 u_multiplier_STAGE1__1900_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_pp1_22 [9]));
 AND2_X1 u_multiplier_STAGE1__1901_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_pp1_22 [10]));
 AND2_X1 u_multiplier_STAGE1__1902_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_pp1_22 [11]));
 AND2_X1 u_multiplier_STAGE1__1903_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_pp1_22 [12]));
 AND2_X1 u_multiplier_STAGE1__1904_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_pp1_22 [13]));
 AND2_X1 u_multiplier_STAGE1__1905_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_pp1_22 [14]));
 AND2_X1 u_multiplier_STAGE1__1906_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_pp1_22 [15]));
 AND2_X1 u_multiplier_STAGE1__1907_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__0663_ ));
 AND2_X1 u_multiplier_STAGE1__1908_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__0664_ ));
 AND2_X1 u_multiplier_STAGE1__1909_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__0665_ ));
 AND2_X1 u_multiplier_STAGE1__1910_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__0666_ ));
 AND2_X1 u_multiplier_STAGE1__1911_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0667_ ));
 AND2_X1 u_multiplier_STAGE1__1912_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0668_ ));
 AND2_X1 u_multiplier_STAGE1__1913_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0669_ ));
 AND2_X1 u_multiplier_STAGE1__1914_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_STAGE1__0670_ ));
 AND2_X1 u_multiplier_STAGE1__1915_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_STAGE1__0671_ ));
 AND2_X1 u_multiplier_STAGE1__1916_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_STAGE1__0672_ ));
 AND2_X1 u_multiplier_STAGE1__1917_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_STAGE1__0673_ ));
 AND2_X1 u_multiplier_STAGE1__1918_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[12]),
    .ZN(u_multiplier_STAGE1__0674_ ));
 AND2_X1 u_multiplier_STAGE1__1919_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[12]),
    .ZN(u_multiplier_STAGE1__0675_ ));
 AND2_X1 u_multiplier_STAGE1__1920_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[13]),
    .ZN(u_multiplier_STAGE1__0676_ ));
 AND2_X1 u_multiplier_STAGE1__1921_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_STAGE1__0677_ ));
 AND2_X1 u_multiplier_STAGE1__1922_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_STAGE1__0678_ ));
 AND2_X1 u_multiplier_STAGE1__1923_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_pp1_23 [8]));
 AND2_X1 u_multiplier_STAGE1__1924_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_pp1_23 [9]));
 AND2_X1 u_multiplier_STAGE1__1925_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_pp1_23 [10]));
 AND2_X1 u_multiplier_STAGE1__1926_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_pp1_23 [11]));
 AND2_X1 u_multiplier_STAGE1__1927_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_pp1_23 [12]));
 AND2_X1 u_multiplier_STAGE1__1928_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_pp1_23 [13]));
 AND2_X1 u_multiplier_STAGE1__1929_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_pp1_23 [14]));
 AND2_X1 u_multiplier_STAGE1__1930_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_pp1_23 [15]));
 AND2_X1 u_multiplier_STAGE1__1931_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__0679_ ));
 AND2_X1 u_multiplier_STAGE1__1932_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__0680_ ));
 AND2_X1 u_multiplier_STAGE1__1933_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__0681_ ));
 AND2_X1 u_multiplier_STAGE1__1934_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__0682_ ));
 AND2_X1 u_multiplier_STAGE1__1935_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__0683_ ));
 AND2_X1 u_multiplier_STAGE1__1936_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0684_ ));
 AND2_X1 u_multiplier_STAGE1__1937_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0685_ ));
 AND2_X1 u_multiplier_STAGE1__1938_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0686_ ));
 AND2_X1 u_multiplier_STAGE1__1939_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_STAGE1__0687_ ));
 AND2_X1 u_multiplier_STAGE1__1940_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_STAGE1__0688_ ));
 AND2_X1 u_multiplier_STAGE1__1941_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_STAGE1__0689_ ));
 AND2_X1 u_multiplier_STAGE1__1942_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_STAGE1__0690_ ));
 AND2_X1 u_multiplier_STAGE1__1943_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[12]),
    .ZN(u_multiplier_STAGE1__0691_ ));
 AND2_X1 u_multiplier_STAGE1__1944_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[13]),
    .ZN(u_multiplier_STAGE1__0692_ ));
 AND2_X1 u_multiplier_STAGE1__1945_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_STAGE1__0693_ ));
 AND2_X1 u_multiplier_STAGE1__1946_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_STAGE1__0694_ ));
 AND2_X1 u_multiplier_STAGE1__1947_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_STAGE1__0695_ ));
 AND2_X1 u_multiplier_STAGE1__1948_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0696_ ));
 AND2_X1 u_multiplier_STAGE1__1949_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_pp1_24 [9]));
 AND2_X1 u_multiplier_STAGE1__1950_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_pp1_24 [10]));
 AND2_X1 u_multiplier_STAGE1__1951_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_pp1_24 [11]));
 AND2_X1 u_multiplier_STAGE1__1952_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_pp1_24 [12]));
 AND2_X1 u_multiplier_STAGE1__1953_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_pp1_24 [13]));
 AND2_X1 u_multiplier_STAGE1__1954_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_pp1_24 [14]));
 AND2_X1 u_multiplier_STAGE1__1955_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_pp1_24 [15]));
 AND2_X1 u_multiplier_STAGE1__1956_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__0697_ ));
 AND2_X1 u_multiplier_STAGE1__1957_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__0698_ ));
 AND2_X1 u_multiplier_STAGE1__1958_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__0699_ ));
 AND2_X1 u_multiplier_STAGE1__1959_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__0700_ ));
 AND2_X1 u_multiplier_STAGE1__1960_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__0701_ ));
 AND2_X1 u_multiplier_STAGE1__1961_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__0702_ ));
 AND2_X1 u_multiplier_STAGE1__1962_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0703_ ));
 AND2_X1 u_multiplier_STAGE1__1963_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0704_ ));
 AND2_X1 u_multiplier_STAGE1__1964_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0705_ ));
 AND2_X1 u_multiplier_STAGE1__1965_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_STAGE1__0706_ ));
 AND2_X1 u_multiplier_STAGE1__1966_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_STAGE1__0707_ ));
 AND2_X1 u_multiplier_STAGE1__1967_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_STAGE1__0708_ ));
 AND2_X1 u_multiplier_STAGE1__1968_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_STAGE1__0709_ ));
 AND2_X1 u_multiplier_STAGE1__1969_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[13]),
    .ZN(u_multiplier_STAGE1__0710_ ));
 AND2_X1 u_multiplier_STAGE1__1970_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_STAGE1__0711_ ));
 AND2_X1 u_multiplier_STAGE1__1971_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_STAGE1__0712_ ));
 AND2_X1 u_multiplier_STAGE1__1972_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_STAGE1__0713_ ));
 AND2_X1 u_multiplier_STAGE1__1973_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0714_ ));
 AND2_X1 u_multiplier_STAGE1__1974_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0715_ ));
 AND2_X1 u_multiplier_STAGE1__1975_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0716_ ));
 AND2_X1 u_multiplier_STAGE1__1976_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_pp1_25 [10]));
 AND2_X1 u_multiplier_STAGE1__1977_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_pp1_25 [11]));
 AND2_X1 u_multiplier_STAGE1__1978_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_pp1_25 [12]));
 AND2_X1 u_multiplier_STAGE1__1979_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_pp1_25 [13]));
 AND2_X1 u_multiplier_STAGE1__1980_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_pp1_25 [14]));
 AND2_X1 u_multiplier_STAGE1__1981_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_pp1_25 [15]));
 AND2_X1 u_multiplier_STAGE1__1982_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__0717_ ));
 AND2_X1 u_multiplier_STAGE1__1983_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__0718_ ));
 AND2_X1 u_multiplier_STAGE1__1984_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__0719_ ));
 AND2_X1 u_multiplier_STAGE1__1985_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__0720_ ));
 AND2_X1 u_multiplier_STAGE1__1986_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__0721_ ));
 AND2_X1 u_multiplier_STAGE1__1987_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__0722_ ));
 AND2_X1 u_multiplier_STAGE1__1988_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__0723_ ));
 AND2_X1 u_multiplier_STAGE1__1989_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0724_ ));
 AND2_X1 u_multiplier_STAGE1__1990_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0725_ ));
 AND2_X1 u_multiplier_STAGE1__1991_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0726_ ));
 AND2_X1 u_multiplier_STAGE1__1992_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_STAGE1__0727_ ));
 AND2_X1 u_multiplier_STAGE1__1993_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_STAGE1__0728_ ));
 AND2_X1 u_multiplier_STAGE1__1994_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_STAGE1__0729_ ));
 AND2_X1 u_multiplier_STAGE1__1995_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_STAGE1__0730_ ));
 AND2_X1 u_multiplier_STAGE1__1996_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_STAGE1__0731_ ));
 AND2_X1 u_multiplier_STAGE1__1997_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_STAGE1__0732_ ));
 AND2_X1 u_multiplier_STAGE1__1998_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_STAGE1__0733_ ));
 AND2_X1 u_multiplier_STAGE1__1999_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0734_ ));
 AND2_X1 u_multiplier_STAGE1__2000_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0735_ ));
 AND2_X1 u_multiplier_STAGE1__2001_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0736_ ));
 AND2_X1 u_multiplier_STAGE1__2002_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__0737_ ));
 AND2_X1 u_multiplier_STAGE1__2003_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__0738_ ));
 AND2_X1 u_multiplier_STAGE1__2004_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_pp1_26 [11]));
 AND2_X1 u_multiplier_STAGE1__2005_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_pp1_26 [12]));
 AND2_X1 u_multiplier_STAGE1__2006_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_pp1_26 [13]));
 AND2_X1 u_multiplier_STAGE1__2007_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_pp1_26 [14]));
 AND2_X1 u_multiplier_STAGE1__2008_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_pp1_26 [15]));
 AND2_X1 u_multiplier_STAGE1__2009_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__0739_ ));
 AND2_X1 u_multiplier_STAGE1__2010_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__0740_ ));
 AND2_X1 u_multiplier_STAGE1__2011_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__0741_ ));
 AND2_X1 u_multiplier_STAGE1__2012_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__0742_ ));
 AND2_X1 u_multiplier_STAGE1__2013_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__0743_ ));
 AND2_X1 u_multiplier_STAGE1__2014_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__0744_ ));
 AND2_X1 u_multiplier_STAGE1__2015_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__0745_ ));
 AND2_X1 u_multiplier_STAGE1__2016_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__0746_ ));
 AND2_X1 u_multiplier_STAGE1__2017_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0747_ ));
 AND2_X1 u_multiplier_STAGE1__2018_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0748_ ));
 AND2_X1 u_multiplier_STAGE1__2019_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0749_ ));
 AND2_X1 u_multiplier_STAGE1__2020_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_STAGE1__0750_ ));
 AND2_X1 u_multiplier_STAGE1__2021_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_STAGE1__0751_ ));
 AND2_X1 u_multiplier_STAGE1__2022_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_STAGE1__0752_ ));
 AND2_X1 u_multiplier_STAGE1__2023_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_STAGE1__0753_ ));
 AND2_X1 u_multiplier_STAGE1__2024_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_STAGE1__0754_ ));
 AND2_X1 u_multiplier_STAGE1__2025_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_STAGE1__0755_ ));
 AND2_X1 u_multiplier_STAGE1__2026_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0756_ ));
 AND2_X1 u_multiplier_STAGE1__2027_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0757_ ));
 AND2_X1 u_multiplier_STAGE1__2028_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0758_ ));
 AND2_X1 u_multiplier_STAGE1__2029_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__0759_ ));
 AND2_X1 u_multiplier_STAGE1__2030_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__0760_ ));
 AND2_X1 u_multiplier_STAGE1__2031_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__0761_ ));
 AND2_X1 u_multiplier_STAGE1__2032_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__0762_ ));
 AND2_X1 u_multiplier_STAGE1__2033_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_pp1_27 [12]));
 AND2_X1 u_multiplier_STAGE1__2034_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_pp1_27 [13]));
 AND2_X1 u_multiplier_STAGE1__2035_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_pp1_27 [14]));
 AND2_X1 u_multiplier_STAGE1__2036_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_pp1_27 [15]));
 AND2_X1 u_multiplier_STAGE1__2037_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_STAGE1__0763_ ));
 AND2_X1 u_multiplier_STAGE1__2038_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__0764_ ));
 AND2_X1 u_multiplier_STAGE1__2039_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__0765_ ));
 AND2_X1 u_multiplier_STAGE1__2040_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__0766_ ));
 AND2_X1 u_multiplier_STAGE1__2041_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__0767_ ));
 AND2_X1 u_multiplier_STAGE1__2042_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__0768_ ));
 AND2_X1 u_multiplier_STAGE1__2043_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__0769_ ));
 AND2_X1 u_multiplier_STAGE1__2044_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__0770_ ));
 AND2_X1 u_multiplier_STAGE1__2045_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__0771_ ));
 AND2_X1 u_multiplier_STAGE1__2046_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0772_ ));
 AND2_X1 u_multiplier_STAGE1__2047_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0773_ ));
 AND2_X1 u_multiplier_STAGE1__2048_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0774_ ));
 AND2_X1 u_multiplier_STAGE1__2049_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_STAGE1__0775_ ));
 AND2_X1 u_multiplier_STAGE1__2050_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_STAGE1__0776_ ));
 AND2_X1 u_multiplier_STAGE1__2051_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_STAGE1__0777_ ));
 AND2_X1 u_multiplier_STAGE1__2052_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_STAGE1__0778_ ));
 AND2_X1 u_multiplier_STAGE1__2053_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_STAGE1__0779_ ));
 AND2_X1 u_multiplier_STAGE1__2054_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0780_ ));
 AND2_X1 u_multiplier_STAGE1__2055_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0781_ ));
 AND2_X1 u_multiplier_STAGE1__2056_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0782_ ));
 AND2_X1 u_multiplier_STAGE1__2057_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__0783_ ));
 AND2_X1 u_multiplier_STAGE1__2058_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__0784_ ));
 AND2_X1 u_multiplier_STAGE1__2059_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__0785_ ));
 AND2_X1 u_multiplier_STAGE1__2060_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__0786_ ));
 AND2_X1 u_multiplier_STAGE1__2061_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__0787_ ));
 AND2_X1 u_multiplier_STAGE1__2062_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__0788_ ));
 AND2_X1 u_multiplier_STAGE1__2063_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_28 [13]));
 AND2_X1 u_multiplier_STAGE1__2064_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_pp1_28 [14]));
 AND2_X1 u_multiplier_STAGE1__2065_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_pp1_28 [15]));
 AND2_X1 u_multiplier_STAGE1__2066_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_STAGE1__0789_ ));
 AND2_X1 u_multiplier_STAGE1__2067_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_STAGE1__0790_ ));
 AND2_X1 u_multiplier_STAGE1__2068_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__0791_ ));
 AND2_X1 u_multiplier_STAGE1__2069_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__0792_ ));
 AND2_X1 u_multiplier_STAGE1__2070_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__0793_ ));
 AND2_X1 u_multiplier_STAGE1__2071_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__0794_ ));
 AND2_X1 u_multiplier_STAGE1__2072_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__0795_ ));
 AND2_X1 u_multiplier_STAGE1__2073_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__0796_ ));
 AND2_X1 u_multiplier_STAGE1__2074_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__0797_ ));
 AND2_X1 u_multiplier_STAGE1__2075_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__0798_ ));
 AND2_X1 u_multiplier_STAGE1__2076_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0799_ ));
 AND2_X1 u_multiplier_STAGE1__2077_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0800_ ));
 AND2_X1 u_multiplier_STAGE1__2078_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0801_ ));
 AND2_X1 u_multiplier_STAGE1__2079_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_STAGE1__0802_ ));
 AND2_X1 u_multiplier_STAGE1__2080_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_STAGE1__0803_ ));
 AND2_X1 u_multiplier_STAGE1__2081_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_STAGE1__0804_ ));
 AND2_X1 u_multiplier_STAGE1__2082_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_STAGE1__0805_ ));
 AND2_X1 u_multiplier_STAGE1__2083_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0806_ ));
 AND2_X1 u_multiplier_STAGE1__2084_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0807_ ));
 AND2_X1 u_multiplier_STAGE1__2085_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0808_ ));
 AND2_X1 u_multiplier_STAGE1__2086_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__0809_ ));
 AND2_X1 u_multiplier_STAGE1__2087_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__0810_ ));
 AND2_X1 u_multiplier_STAGE1__2088_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__0811_ ));
 AND2_X1 u_multiplier_STAGE1__2089_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__0812_ ));
 AND2_X1 u_multiplier_STAGE1__2090_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__0813_ ));
 AND2_X1 u_multiplier_STAGE1__2091_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__0814_ ));
 AND2_X1 u_multiplier_STAGE1__2092_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__0815_ ));
 AND2_X1 u_multiplier_STAGE1__2093_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__0816_ ));
 AND2_X1 u_multiplier_STAGE1__2094_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_29 [14]));
 AND2_X1 u_multiplier_STAGE1__2095_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_29 [15]));
 AND2_X1 u_multiplier_STAGE1__2096_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_STAGE1__0817_ ));
 AND2_X1 u_multiplier_STAGE1__2097_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_STAGE1__0818_ ));
 AND2_X1 u_multiplier_STAGE1__2098_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_STAGE1__0819_ ));
 AND2_X1 u_multiplier_STAGE1__2099_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__0820_ ));
 AND2_X1 u_multiplier_STAGE1__2100_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__0821_ ));
 AND2_X1 u_multiplier_STAGE1__2101_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__0822_ ));
 AND2_X1 u_multiplier_STAGE1__2102_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__0823_ ));
 AND2_X1 u_multiplier_STAGE1__2103_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__0824_ ));
 AND2_X1 u_multiplier_STAGE1__2104_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__0825_ ));
 AND2_X1 u_multiplier_STAGE1__2105_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__0826_ ));
 AND2_X1 u_multiplier_STAGE1__2106_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__0827_ ));
 AND2_X1 u_multiplier_STAGE1__2107_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0828_ ));
 AND2_X1 u_multiplier_STAGE1__2108_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0829_ ));
 AND2_X1 u_multiplier_STAGE1__2109_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0830_ ));
 AND2_X1 u_multiplier_STAGE1__2110_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_STAGE1__0831_ ));
 AND2_X1 u_multiplier_STAGE1__2111_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_STAGE1__0832_ ));
 AND2_X1 u_multiplier_STAGE1__2112_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_STAGE1__0833_ ));
 AND2_X1 u_multiplier_STAGE1__2113_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0834_ ));
 AND2_X1 u_multiplier_STAGE1__2114_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0835_ ));
 AND2_X1 u_multiplier_STAGE1__2115_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0836_ ));
 AND2_X1 u_multiplier_STAGE1__2116_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__0837_ ));
 AND2_X1 u_multiplier_STAGE1__2117_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__0838_ ));
 AND2_X1 u_multiplier_STAGE1__2118_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__0839_ ));
 AND2_X1 u_multiplier_STAGE1__2119_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__0840_ ));
 AND2_X1 u_multiplier_STAGE1__2120_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__0841_ ));
 AND2_X1 u_multiplier_STAGE1__2121_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__0842_ ));
 AND2_X1 u_multiplier_STAGE1__2122_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__0843_ ));
 AND2_X1 u_multiplier_STAGE1__2123_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__0844_ ));
 AND2_X1 u_multiplier_STAGE1__2124_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_STAGE1__0845_ ));
 AND2_X1 u_multiplier_STAGE1__2125_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_STAGE1__0846_ ));
 AND2_X1 u_multiplier_STAGE1__2126_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_30 [15]));
 AND2_X1 u_multiplier_STAGE1__2127_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_STAGE1__0847_ ));
 AND2_X1 u_multiplier_STAGE1__2128_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_STAGE1__0848_ ));
 AND2_X1 u_multiplier_STAGE1__2129_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_STAGE1__0849_ ));
 AND2_X1 u_multiplier_STAGE1__2130_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_STAGE1__0850_ ));
 AND2_X1 u_multiplier_STAGE1__2131_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__0851_ ));
 AND2_X1 u_multiplier_STAGE1__2132_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__0852_ ));
 AND2_X1 u_multiplier_STAGE1__2133_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__0853_ ));
 AND2_X1 u_multiplier_STAGE1__2134_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__0854_ ));
 AND2_X1 u_multiplier_STAGE1__2135_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__0855_ ));
 AND2_X1 u_multiplier_STAGE1__2136_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__0856_ ));
 AND2_X1 u_multiplier_STAGE1__2137_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__0857_ ));
 AND2_X1 u_multiplier_STAGE1__2138_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__0858_ ));
 AND2_X1 u_multiplier_STAGE1__2139_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0859_ ));
 AND2_X1 u_multiplier_STAGE1__2140_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0860_ ));
 AND2_X1 u_multiplier_STAGE1__2141_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0861_ ));
 AND2_X1 u_multiplier_STAGE1__2142_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_STAGE1__0862_ ));
 AND2_X1 u_multiplier_STAGE1__2143_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_STAGE1__0863_ ));
 AND2_X1 u_multiplier_STAGE1__2144_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0864_ ));
 AND2_X1 u_multiplier_STAGE1__2145_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0865_ ));
 AND2_X1 u_multiplier_STAGE1__2146_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0866_ ));
 AND2_X1 u_multiplier_STAGE1__2147_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__0867_ ));
 AND2_X1 u_multiplier_STAGE1__2148_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__0868_ ));
 AND2_X1 u_multiplier_STAGE1__2149_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__0869_ ));
 AND2_X1 u_multiplier_STAGE1__2150_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__0870_ ));
 AND2_X1 u_multiplier_STAGE1__2151_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__0871_ ));
 AND2_X1 u_multiplier_STAGE1__2152_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__0872_ ));
 AND2_X1 u_multiplier_STAGE1__2153_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__0873_ ));
 AND2_X1 u_multiplier_STAGE1__2154_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__0874_ ));
 AND2_X1 u_multiplier_STAGE1__2155_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_STAGE1__0875_ ));
 AND2_X1 u_multiplier_STAGE1__2156_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_STAGE1__0876_ ));
 AND2_X1 u_multiplier_STAGE1__2157_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_STAGE1__0877_ ));
 AND2_X1 u_multiplier_STAGE1__2158_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_STAGE1__0878_ ));
 AND2_X1 u_multiplier_STAGE1__2159_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_STAGE1__0879_ ));
 AND2_X1 u_multiplier_STAGE1__2160_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_STAGE1__0880_ ));
 AND2_X1 u_multiplier_STAGE1__2161_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_STAGE1__0881_ ));
 AND2_X1 u_multiplier_STAGE1__2162_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_STAGE1__0882_ ));
 AND2_X1 u_multiplier_STAGE1__2163_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__0883_ ));
 AND2_X1 u_multiplier_STAGE1__2164_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__0884_ ));
 AND2_X1 u_multiplier_STAGE1__2165_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__0885_ ));
 AND2_X1 u_multiplier_STAGE1__2166_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__0886_ ));
 AND2_X1 u_multiplier_STAGE1__2167_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__0887_ ));
 AND2_X1 u_multiplier_STAGE1__2168_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__0888_ ));
 AND2_X1 u_multiplier_STAGE1__2169_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__0889_ ));
 AND2_X1 u_multiplier_STAGE1__2170_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__0890_ ));
 AND2_X1 u_multiplier_STAGE1__2171_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0891_ ));
 AND2_X1 u_multiplier_STAGE1__2172_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0892_ ));
 AND2_X1 u_multiplier_STAGE1__2173_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0893_ ));
 AND2_X1 u_multiplier_STAGE1__2174_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_STAGE1__0894_ ));
 AND2_X1 u_multiplier_STAGE1__2175_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0895_ ));
 AND2_X1 u_multiplier_STAGE1__2176_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0896_ ));
 AND2_X1 u_multiplier_STAGE1__2177_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0897_ ));
 AND2_X1 u_multiplier_STAGE1__2178_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__0898_ ));
 AND2_X1 u_multiplier_STAGE1__2179_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__0899_ ));
 AND2_X1 u_multiplier_STAGE1__2180_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__0900_ ));
 AND2_X1 u_multiplier_STAGE1__2181_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__0901_ ));
 AND2_X1 u_multiplier_STAGE1__2182_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__0902_ ));
 AND2_X1 u_multiplier_STAGE1__2183_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__0903_ ));
 AND2_X1 u_multiplier_STAGE1__2184_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__0904_ ));
 AND2_X1 u_multiplier_STAGE1__2185_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__0905_ ));
 AND2_X1 u_multiplier_STAGE1__2186_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_STAGE1__0906_ ));
 AND2_X1 u_multiplier_STAGE1__2187_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_STAGE1__0907_ ));
 AND2_X1 u_multiplier_STAGE1__2188_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_STAGE1__0908_ ));
 AND2_X1 u_multiplier_STAGE1__2189_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_STAGE1__0909_ ));
 AND2_X1 u_multiplier_STAGE1__2190_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_STAGE1__0910_ ));
 AND2_X1 u_multiplier_STAGE1__2191_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_STAGE1__0911_ ));
 AND2_X1 u_multiplier_STAGE1__2192_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_STAGE1__0912_ ));
 AND2_X1 u_multiplier_STAGE1__2193_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_STAGE1__0913_ ));
 AND2_X1 u_multiplier_STAGE1__2194_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__0914_ ));
 AND2_X1 u_multiplier_STAGE1__2195_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__0915_ ));
 AND2_X1 u_multiplier_STAGE1__2196_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__0916_ ));
 AND2_X1 u_multiplier_STAGE1__2197_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__0917_ ));
 AND2_X1 u_multiplier_STAGE1__2198_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__0918_ ));
 AND2_X1 u_multiplier_STAGE1__2199_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__0919_ ));
 AND2_X1 u_multiplier_STAGE1__2200_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__0920_ ));
 AND2_X1 u_multiplier_STAGE1__2201_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__0921_ ));
 AND2_X1 u_multiplier_STAGE1__2202_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0922_ ));
 AND2_X1 u_multiplier_STAGE1__2203_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0923_ ));
 AND2_X1 u_multiplier_STAGE1__2204_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0924_ ));
 AND2_X1 u_multiplier_STAGE1__2205_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0925_ ));
 AND2_X1 u_multiplier_STAGE1__2206_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0926_ ));
 AND2_X1 u_multiplier_STAGE1__2207_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0927_ ));
 AND2_X1 u_multiplier_STAGE1__2208_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__0928_ ));
 AND2_X1 u_multiplier_STAGE1__2209_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__0929_ ));
 AND2_X1 u_multiplier_STAGE1__2210_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__0930_ ));
 AND2_X1 u_multiplier_STAGE1__2211_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__0931_ ));
 AND2_X1 u_multiplier_STAGE1__2212_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__0932_ ));
 AND2_X1 u_multiplier_STAGE1__2213_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__0933_ ));
 AND2_X1 u_multiplier_STAGE1__2214_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__0934_ ));
 AND2_X1 u_multiplier_STAGE1__2215_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__0935_ ));
 AND2_X1 u_multiplier_STAGE1__2216_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_STAGE1__0936_ ));
 AND2_X1 u_multiplier_STAGE1__2217_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_STAGE1__0937_ ));
 AND2_X2 u_multiplier_STAGE1__2218_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_STAGE1__0938_ ));
 AND2_X2 u_multiplier_STAGE1__2219_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_STAGE1__0939_ ));
 AND2_X1 u_multiplier_STAGE1__2220_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_STAGE1__0940_ ));
 AND2_X1 u_multiplier_STAGE1__2221_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_STAGE1__0941_ ));
 AND2_X1 u_multiplier_STAGE1__2222_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_STAGE1__0942_ ));
 AND2_X1 u_multiplier_STAGE1__2223_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_STAGE1__0943_ ));
 AND2_X1 u_multiplier_STAGE1__2224_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__0944_ ));
 AND2_X1 u_multiplier_STAGE1__2225_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__0945_ ));
 AND2_X1 u_multiplier_STAGE1__2226_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__0946_ ));
 AND2_X1 u_multiplier_STAGE1__2227_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__0947_ ));
 AND2_X1 u_multiplier_STAGE1__2228_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__0948_ ));
 AND2_X1 u_multiplier_STAGE1__2229_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__0949_ ));
 AND2_X1 u_multiplier_STAGE1__2230_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__0950_ ));
 AND2_X1 u_multiplier_STAGE1__2231_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__0951_ ));
 AND2_X1 u_multiplier_STAGE1__2232_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0952_ ));
 AND2_X1 u_multiplier_STAGE1__2233_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0953_ ));
 AND2_X1 u_multiplier_STAGE1__2234_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0954_ ));
 AND2_X1 u_multiplier_STAGE1__2235_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0955_ ));
 AND2_X1 u_multiplier_STAGE1__2236_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0956_ ));
 AND2_X1 u_multiplier_STAGE1__2237_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__0957_ ));
 AND2_X1 u_multiplier_STAGE1__2238_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__0958_ ));
 AND2_X1 u_multiplier_STAGE1__2239_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__0959_ ));
 AND2_X1 u_multiplier_STAGE1__2240_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__0960_ ));
 AND2_X1 u_multiplier_STAGE1__2241_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__0961_ ));
 AND2_X1 u_multiplier_STAGE1__2242_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__0962_ ));
 AND2_X1 u_multiplier_STAGE1__2243_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__0963_ ));
 AND2_X1 u_multiplier_STAGE1__2244_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__0964_ ));
 AND2_X1 u_multiplier_STAGE1__2245_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_STAGE1__0965_ ));
 AND2_X1 u_multiplier_STAGE1__2246_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_STAGE1__0966_ ));
 AND2_X1 u_multiplier_STAGE1__2247_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_STAGE1__0967_ ));
 AND2_X1 u_multiplier_STAGE1__2248_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_34 [15]));
 AND2_X1 u_multiplier_STAGE1__2249_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_STAGE1__0968_ ));
 AND2_X1 u_multiplier_STAGE1__2250_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_STAGE1__0969_ ));
 AND2_X1 u_multiplier_STAGE1__2251_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_STAGE1__0970_ ));
 AND2_X1 u_multiplier_STAGE1__2252_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_STAGE1__0971_ ));
 AND2_X1 u_multiplier_STAGE1__2253_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__0972_ ));
 AND2_X1 u_multiplier_STAGE1__2254_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__0973_ ));
 AND2_X1 u_multiplier_STAGE1__2255_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__0974_ ));
 AND2_X1 u_multiplier_STAGE1__2256_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__0975_ ));
 AND2_X1 u_multiplier_STAGE1__2257_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__0976_ ));
 AND2_X1 u_multiplier_STAGE1__2258_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__0977_ ));
 AND2_X1 u_multiplier_STAGE1__2259_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__0978_ ));
 AND2_X1 u_multiplier_STAGE1__2260_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__0979_ ));
 AND2_X1 u_multiplier_STAGE1__2261_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0980_ ));
 AND2_X1 u_multiplier_STAGE1__2262_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0981_ ));
 AND2_X1 u_multiplier_STAGE1__2263_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0982_ ));
 AND2_X1 u_multiplier_STAGE1__2264_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0983_ ));
 AND2_X1 u_multiplier_STAGE1__2265_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__0984_ ));
 AND2_X1 u_multiplier_STAGE1__2266_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__0985_ ));
 AND2_X1 u_multiplier_STAGE1__2267_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__0986_ ));
 AND2_X1 u_multiplier_STAGE1__2268_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__0987_ ));
 AND2_X1 u_multiplier_STAGE1__2269_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__0988_ ));
 AND2_X1 u_multiplier_STAGE1__2270_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__0989_ ));
 AND2_X1 u_multiplier_STAGE1__2271_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__0990_ ));
 AND2_X1 u_multiplier_STAGE1__2272_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__0991_ ));
 AND2_X1 u_multiplier_STAGE1__2273_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_STAGE1__0992_ ));
 AND2_X1 u_multiplier_STAGE1__2274_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_STAGE1__0993_ ));
 AND2_X1 u_multiplier_STAGE1__2275_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_35 [14]));
 AND2_X1 u_multiplier_STAGE1__2276_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_35 [15]));
 AND2_X1 u_multiplier_STAGE1__2277_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_STAGE1__0994_ ));
 AND2_X1 u_multiplier_STAGE1__2278_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_STAGE1__0995_ ));
 AND2_X1 u_multiplier_STAGE1__2279_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_STAGE1__0996_ ));
 AND2_X1 u_multiplier_STAGE1__2280_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_STAGE1__0997_ ));
 AND2_X1 u_multiplier_STAGE1__2281_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__0998_ ));
 AND2_X1 u_multiplier_STAGE1__2282_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__0999_ ));
 AND2_X1 u_multiplier_STAGE1__2283_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__1000_ ));
 AND2_X1 u_multiplier_STAGE1__2284_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__1001_ ));
 AND2_X1 u_multiplier_STAGE1__2285_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__1002_ ));
 AND2_X1 u_multiplier_STAGE1__2286_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__1003_ ));
 AND2_X1 u_multiplier_STAGE1__2287_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__1004_ ));
 AND2_X1 u_multiplier_STAGE1__2288_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__1005_ ));
 AND2_X1 u_multiplier_STAGE1__2289_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__1006_ ));
 AND2_X1 u_multiplier_STAGE1__2290_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__1007_ ));
 AND2_X1 u_multiplier_STAGE1__2291_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__1008_ ));
 AND2_X1 u_multiplier_STAGE1__2292_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__1009_ ));
 AND2_X1 u_multiplier_STAGE1__2293_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__1010_ ));
 AND2_X1 u_multiplier_STAGE1__2294_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__1011_ ));
 AND2_X1 u_multiplier_STAGE1__2295_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__1012_ ));
 AND2_X1 u_multiplier_STAGE1__2296_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__1013_ ));
 AND2_X1 u_multiplier_STAGE1__2297_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__1014_ ));
 AND2_X1 u_multiplier_STAGE1__2298_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__1015_ ));
 AND2_X1 u_multiplier_STAGE1__2299_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__1016_ ));
 AND2_X1 u_multiplier_STAGE1__2300_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_STAGE1__1017_ ));
 AND2_X1 u_multiplier_STAGE1__2301_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_36 [13]));
 AND2_X1 u_multiplier_STAGE1__2302_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_36 [14]));
 AND2_X1 u_multiplier_STAGE1__2303_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_36 [15]));
 AND2_X1 u_multiplier_STAGE1__2304_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_STAGE1__1018_ ));
 AND2_X1 u_multiplier_STAGE1__2305_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_STAGE1__1019_ ));
 AND2_X1 u_multiplier_STAGE1__2306_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_STAGE1__1020_ ));
 AND2_X1 u_multiplier_STAGE1__2307_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_STAGE1__1021_ ));
 AND2_X1 u_multiplier_STAGE1__2308_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__1022_ ));
 AND2_X1 u_multiplier_STAGE1__2309_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__1023_ ));
 AND2_X1 u_multiplier_STAGE1__2310_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__1024_ ));
 AND2_X1 u_multiplier_STAGE1__2311_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__1025_ ));
 AND2_X1 u_multiplier_STAGE1__2312_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__1026_ ));
 AND2_X1 u_multiplier_STAGE1__2313_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__1027_ ));
 AND2_X1 u_multiplier_STAGE1__2314_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__1028_ ));
 AND2_X1 u_multiplier_STAGE1__2315_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__1029_ ));
 AND2_X1 u_multiplier_STAGE1__2316_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__1030_ ));
 AND2_X1 u_multiplier_STAGE1__2317_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__1031_ ));
 AND2_X1 u_multiplier_STAGE1__2318_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__1032_ ));
 AND2_X1 u_multiplier_STAGE1__2319_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__1033_ ));
 AND2_X1 u_multiplier_STAGE1__2320_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__1034_ ));
 AND2_X1 u_multiplier_STAGE1__2321_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__1035_ ));
 AND2_X1 u_multiplier_STAGE1__2322_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__1036_ ));
 AND2_X1 u_multiplier_STAGE1__2323_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__1037_ ));
 AND2_X1 u_multiplier_STAGE1__2324_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__1038_ ));
 AND2_X1 u_multiplier_STAGE1__2325_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__1039_ ));
 AND2_X1 u_multiplier_STAGE1__2326_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_37 [12]));
 AND2_X1 u_multiplier_STAGE1__2327_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_37 [13]));
 AND2_X1 u_multiplier_STAGE1__2328_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_37 [14]));
 AND2_X1 u_multiplier_STAGE1__2329_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_37 [15]));
 AND2_X1 u_multiplier_STAGE1__2330_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_STAGE1__1040_ ));
 AND2_X1 u_multiplier_STAGE1__2331_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_STAGE1__1041_ ));
 AND2_X1 u_multiplier_STAGE1__2332_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_STAGE1__1042_ ));
 AND2_X1 u_multiplier_STAGE1__2333_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_STAGE1__1043_ ));
 AND2_X1 u_multiplier_STAGE1__2334_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__1044_ ));
 AND2_X1 u_multiplier_STAGE1__2335_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__1045_ ));
 AND2_X1 u_multiplier_STAGE1__2336_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__1046_ ));
 AND2_X1 u_multiplier_STAGE1__2337_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__1047_ ));
 AND2_X1 u_multiplier_STAGE1__2338_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__1048_ ));
 AND2_X1 u_multiplier_STAGE1__2339_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__1049_ ));
 AND2_X1 u_multiplier_STAGE1__2340_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__1050_ ));
 AND2_X1 u_multiplier_STAGE1__2341_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__1051_ ));
 AND2_X1 u_multiplier_STAGE1__2342_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__1052_ ));
 AND2_X1 u_multiplier_STAGE1__2343_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__1053_ ));
 AND2_X1 u_multiplier_STAGE1__2344_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__1054_ ));
 AND2_X1 u_multiplier_STAGE1__2345_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__1055_ ));
 AND2_X1 u_multiplier_STAGE1__2346_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__1056_ ));
 AND2_X1 u_multiplier_STAGE1__2347_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__1057_ ));
 AND2_X1 u_multiplier_STAGE1__2348_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__1058_ ));
 AND2_X1 u_multiplier_STAGE1__2349_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__1059_ ));
 AND2_X1 u_multiplier_STAGE1__2350_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_38 [11]));
 AND2_X1 u_multiplier_STAGE1__2351_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_38 [12]));
 AND2_X1 u_multiplier_STAGE1__2352_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_38 [13]));
 AND2_X1 u_multiplier_STAGE1__2353_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_38 [14]));
 AND2_X1 u_multiplier_STAGE1__2354_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_pp1_38 [15]));
 AND2_X1 u_multiplier_STAGE1__2355_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_STAGE1__1060_ ));
 AND2_X1 u_multiplier_STAGE1__2356_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_STAGE1__1061_ ));
 AND2_X1 u_multiplier_STAGE1__2357_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_STAGE1__1062_ ));
 AND2_X1 u_multiplier_STAGE1__2358_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_STAGE1__1063_ ));
 AND2_X1 u_multiplier_STAGE1__2359_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__1064_ ));
 AND2_X1 u_multiplier_STAGE1__2360_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__1065_ ));
 AND2_X1 u_multiplier_STAGE1__2361_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__1066_ ));
 AND2_X1 u_multiplier_STAGE1__2362_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__1067_ ));
 AND2_X1 u_multiplier_STAGE1__2363_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__1068_ ));
 AND2_X1 u_multiplier_STAGE1__2364_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__1069_ ));
 AND2_X1 u_multiplier_STAGE1__2365_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__1070_ ));
 AND2_X1 u_multiplier_STAGE1__2366_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__1071_ ));
 AND2_X1 u_multiplier_STAGE1__2367_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__1072_ ));
 AND2_X1 u_multiplier_STAGE1__2368_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__1073_ ));
 AND2_X1 u_multiplier_STAGE1__2369_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__1074_ ));
 AND2_X1 u_multiplier_STAGE1__2370_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__1075_ ));
 AND2_X1 u_multiplier_STAGE1__2371_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__1076_ ));
 AND2_X1 u_multiplier_STAGE1__2372_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__1077_ ));
 AND2_X1 u_multiplier_STAGE1__2373_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_39 [10]));
 AND2_X1 u_multiplier_STAGE1__2374_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_39 [11]));
 AND2_X1 u_multiplier_STAGE1__2375_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_39 [12]));
 AND2_X1 u_multiplier_STAGE1__2376_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_39 [13]));
 AND2_X1 u_multiplier_STAGE1__2377_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_pp1_39 [14]));
 AND2_X1 u_multiplier_STAGE1__2378_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_pp1_39 [15]));
 AND2_X1 u_multiplier_STAGE1__2379_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_STAGE1__1078_ ));
 AND2_X1 u_multiplier_STAGE1__2380_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_STAGE1__1079_ ));
 AND2_X1 u_multiplier_STAGE1__2381_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_STAGE1__1080_ ));
 AND2_X1 u_multiplier_STAGE1__2382_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_STAGE1__1081_ ));
 AND2_X1 u_multiplier_STAGE1__2383_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__1082_ ));
 AND2_X1 u_multiplier_STAGE1__2384_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__1083_ ));
 AND2_X1 u_multiplier_STAGE1__2385_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__1084_ ));
 AND2_X1 u_multiplier_STAGE1__2386_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__1085_ ));
 AND2_X1 u_multiplier_STAGE1__2387_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__1086_ ));
 AND2_X1 u_multiplier_STAGE1__2388_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__1087_ ));
 AND2_X1 u_multiplier_STAGE1__2389_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__1088_ ));
 AND2_X1 u_multiplier_STAGE1__2390_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__1089_ ));
 AND2_X1 u_multiplier_STAGE1__2391_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__1090_ ));
 AND2_X1 u_multiplier_STAGE1__2392_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__1091_ ));
 AND2_X1 u_multiplier_STAGE1__2393_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__1092_ ));
 AND2_X1 u_multiplier_STAGE1__2394_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__1093_ ));
 AND2_X1 u_multiplier_STAGE1__2395_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_40 [9]));
 AND2_X1 u_multiplier_STAGE1__2396_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_40 [10]));
 AND2_X1 u_multiplier_STAGE1__2397_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_40 [11]));
 AND2_X1 u_multiplier_STAGE1__2398_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_40 [12]));
 AND2_X1 u_multiplier_STAGE1__2399_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_pp1_40 [13]));
 AND2_X1 u_multiplier_STAGE1__2400_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_pp1_40 [14]));
 AND2_X1 u_multiplier_STAGE1__2401_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_pp1_40 [15]));
 AND2_X1 u_multiplier_STAGE1__2402_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_STAGE1__1094_ ));
 AND2_X1 u_multiplier_STAGE1__2403_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_STAGE1__1095_ ));
 AND2_X1 u_multiplier_STAGE1__2404_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_STAGE1__1096_ ));
 AND2_X1 u_multiplier_STAGE1__2405_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_STAGE1__1097_ ));
 AND2_X1 u_multiplier_STAGE1__2406_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__1098_ ));
 AND2_X1 u_multiplier_STAGE1__2407_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__1099_ ));
 AND2_X1 u_multiplier_STAGE1__2408_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__1100_ ));
 AND2_X1 u_multiplier_STAGE1__2409_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__1101_ ));
 AND2_X1 u_multiplier_STAGE1__2410_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__1102_ ));
 AND2_X1 u_multiplier_STAGE1__2411_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__1103_ ));
 AND2_X1 u_multiplier_STAGE1__2412_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__1104_ ));
 AND2_X1 u_multiplier_STAGE1__2413_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__1105_ ));
 AND2_X1 u_multiplier_STAGE1__2414_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__1106_ ));
 AND2_X1 u_multiplier_STAGE1__2415_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__1107_ ));
 AND2_X1 u_multiplier_STAGE1__2416_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_41 [8]));
 AND2_X1 u_multiplier_STAGE1__2417_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_41 [9]));
 AND2_X1 u_multiplier_STAGE1__2418_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_41 [10]));
 AND2_X1 u_multiplier_STAGE1__2419_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_41 [11]));
 AND2_X1 u_multiplier_STAGE1__2420_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_pp1_41 [12]));
 AND2_X1 u_multiplier_STAGE1__2421_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_pp1_41 [13]));
 AND2_X1 u_multiplier_STAGE1__2422_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_pp1_41 [14]));
 AND2_X1 u_multiplier_STAGE1__2423_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_pp1_41 [15]));
 AND2_X1 u_multiplier_STAGE1__2424_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_STAGE1__1108_ ));
 AND2_X1 u_multiplier_STAGE1__2425_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_STAGE1__1109_ ));
 AND2_X1 u_multiplier_STAGE1__2426_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_STAGE1__1110_ ));
 AND2_X1 u_multiplier_STAGE1__2427_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_STAGE1__1111_ ));
 AND2_X1 u_multiplier_STAGE1__2428_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__1112_ ));
 AND2_X1 u_multiplier_STAGE1__2429_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__1113_ ));
 AND2_X1 u_multiplier_STAGE1__2430_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__1114_ ));
 AND2_X1 u_multiplier_STAGE1__2431_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__1115_ ));
 AND2_X1 u_multiplier_STAGE1__2432_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__1116_ ));
 AND2_X1 u_multiplier_STAGE1__2433_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__1117_ ));
 AND2_X1 u_multiplier_STAGE1__2434_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__1118_ ));
 AND2_X1 u_multiplier_STAGE1__2435_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__1119_ ));
 AND2_X1 u_multiplier_STAGE1__2436_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_42 [7]));
 AND2_X1 u_multiplier_STAGE1__2437_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_42 [8]));
 AND2_X1 u_multiplier_STAGE1__2438_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_42 [9]));
 AND2_X1 u_multiplier_STAGE1__2439_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_42 [10]));
 AND2_X1 u_multiplier_STAGE1__2440_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_pp1_42 [11]));
 AND2_X1 u_multiplier_STAGE1__2441_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_pp1_42 [12]));
 AND2_X1 u_multiplier_STAGE1__2442_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_pp1_42 [13]));
 AND2_X1 u_multiplier_STAGE1__2443_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_pp1_42 [14]));
 AND2_X1 u_multiplier_STAGE1__2444_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_pp1_42 [15]));
 AND2_X1 u_multiplier_STAGE1__2445_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_STAGE1__1120_ ));
 AND2_X1 u_multiplier_STAGE1__2446_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_STAGE1__1121_ ));
 AND2_X1 u_multiplier_STAGE1__2447_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_STAGE1__1122_ ));
 AND2_X1 u_multiplier_STAGE1__2448_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_STAGE1__1123_ ));
 AND2_X1 u_multiplier_STAGE1__2449_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__1124_ ));
 AND2_X1 u_multiplier_STAGE1__2450_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__1125_ ));
 AND2_X1 u_multiplier_STAGE1__2451_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__1126_ ));
 AND2_X1 u_multiplier_STAGE1__2452_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__1127_ ));
 AND2_X1 u_multiplier_STAGE1__2453_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__1128_ ));
 AND2_X1 u_multiplier_STAGE1__2454_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__1129_ ));
 AND2_X1 u_multiplier_STAGE1__2455_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_43 [6]));
 AND2_X1 u_multiplier_STAGE1__2456_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_43 [7]));
 AND2_X1 u_multiplier_STAGE1__2457_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_43 [8]));
 AND2_X1 u_multiplier_STAGE1__2458_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_43 [9]));
 AND2_X1 u_multiplier_STAGE1__2459_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_pp1_43 [10]));
 AND2_X1 u_multiplier_STAGE1__2460_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_pp1_43 [11]));
 AND2_X1 u_multiplier_STAGE1__2461_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_pp1_43 [12]));
 AND2_X1 u_multiplier_STAGE1__2462_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_pp1_43 [13]));
 AND2_X1 u_multiplier_STAGE1__2463_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_pp1_43 [14]));
 AND2_X1 u_multiplier_STAGE1__2464_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_pp1_43 [15]));
 AND2_X1 u_multiplier_STAGE1__2465_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_STAGE1__1130_ ));
 AND2_X1 u_multiplier_STAGE1__2466_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_STAGE1__1131_ ));
 AND2_X1 u_multiplier_STAGE1__2467_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_STAGE1__1132_ ));
 AND2_X1 u_multiplier_STAGE1__2468_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_STAGE1__1133_ ));
 AND2_X1 u_multiplier_STAGE1__2469_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__1134_ ));
 AND2_X1 u_multiplier_STAGE1__2470_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__1135_ ));
 AND2_X1 u_multiplier_STAGE1__2471_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__1136_ ));
 AND2_X1 u_multiplier_STAGE1__2472_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__1137_ ));
 AND2_X1 u_multiplier_STAGE1__2473_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_44 [5]));
 AND2_X1 u_multiplier_STAGE1__2474_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_44 [6]));
 AND2_X1 u_multiplier_STAGE1__2475_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_44 [7]));
 AND2_X1 u_multiplier_STAGE1__2476_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_44 [8]));
 AND2_X1 u_multiplier_STAGE1__2477_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_pp1_44 [9]));
 AND2_X1 u_multiplier_STAGE1__2478_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_pp1_44 [10]));
 AND2_X1 u_multiplier_STAGE1__2479_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_pp1_44 [11]));
 AND2_X1 u_multiplier_STAGE1__2480_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_pp1_44 [12]));
 AND2_X1 u_multiplier_STAGE1__2481_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_pp1_44 [13]));
 AND2_X1 u_multiplier_STAGE1__2482_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_pp1_44 [14]));
 AND2_X1 u_multiplier_STAGE1__2483_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_pp1_44 [15]));
 AND2_X1 u_multiplier_STAGE1__2484_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_STAGE1__1138_ ));
 AND2_X1 u_multiplier_STAGE1__2485_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_STAGE1__1139_ ));
 AND2_X1 u_multiplier_STAGE1__2486_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_STAGE1__1140_ ));
 AND2_X1 u_multiplier_STAGE1__2487_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_STAGE1__1141_ ));
 AND2_X1 u_multiplier_STAGE1__2488_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__1142_ ));
 AND2_X1 u_multiplier_STAGE1__2489_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__1143_ ));
 AND2_X1 u_multiplier_STAGE1__2490_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_45 [4]));
 AND2_X1 u_multiplier_STAGE1__2491_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_45 [5]));
 AND2_X1 u_multiplier_STAGE1__2492_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_45 [6]));
 AND2_X1 u_multiplier_STAGE1__2493_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_45 [7]));
 AND2_X1 u_multiplier_STAGE1__2494_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_pp1_45 [8]));
 AND2_X1 u_multiplier_STAGE1__2495_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_pp1_45 [9]));
 AND2_X1 u_multiplier_STAGE1__2496_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_pp1_45 [10]));
 AND2_X1 u_multiplier_STAGE1__2497_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_pp1_45 [11]));
 AND2_X1 u_multiplier_STAGE1__2498_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_pp1_45 [12]));
 AND2_X1 u_multiplier_STAGE1__2499_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_pp1_45 [13]));
 AND2_X1 u_multiplier_STAGE1__2500_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_pp1_45 [14]));
 AND2_X1 u_multiplier_STAGE1__2501_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_pp1_45 [15]));
 AND2_X1 u_multiplier_STAGE1__2502_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_STAGE1__1144_ ));
 AND2_X1 u_multiplier_STAGE1__2503_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_STAGE1__1145_ ));
 AND2_X1 u_multiplier_STAGE1__2504_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_STAGE1__1146_ ));
 AND2_X1 u_multiplier_STAGE1__2505_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_STAGE1__1147_ ));
 AND2_X1 u_multiplier_STAGE1__2506_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_46 [3]));
 AND2_X1 u_multiplier_STAGE1__2507_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_46 [4]));
 AND2_X1 u_multiplier_STAGE1__2508_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_46 [5]));
 AND2_X1 u_multiplier_STAGE1__2509_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_46 [6]));
 AND2_X1 u_multiplier_STAGE1__2510_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_pp1_46 [7]));
 AND2_X1 u_multiplier_STAGE1__2511_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_pp1_46 [8]));
 AND2_X1 u_multiplier_STAGE1__2512_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_pp1_46 [9]));
 AND2_X1 u_multiplier_STAGE1__2513_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_pp1_46 [10]));
 AND2_X1 u_multiplier_STAGE1__2514_  (.A1(sram_rdata_reg[23]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_pp1_46 [11]));
 AND2_X1 u_multiplier_STAGE1__2515_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_pp1_46 [12]));
 AND2_X1 u_multiplier_STAGE1__2516_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_pp1_46 [13]));
 AND2_X1 u_multiplier_STAGE1__2517_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_pp1_46 [14]));
 AND2_X1 u_multiplier_STAGE1__2518_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_pp1_46 [15]));
 AND2_X1 u_multiplier_STAGE1__2519_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_STAGE1__1148_ ));
 AND2_X1 u_multiplier_STAGE1__2520_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_STAGE1__1149_ ));
 AND2_X1 u_multiplier_STAGE1__2521_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_47 [2]));
 AND2_X1 u_multiplier_STAGE1__2522_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_47 [3]));
 AND2_X1 u_multiplier_STAGE1__2523_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_47 [4]));
 AND2_X1 u_multiplier_STAGE1__2524_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_47 [5]));
 AND2_X1 u_multiplier_STAGE1__2525_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_pp1_47 [6]));
 AND2_X1 u_multiplier_STAGE1__2526_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_pp1_47 [7]));
 AND2_X1 u_multiplier_STAGE1__2527_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_pp1_47 [8]));
 AND2_X1 u_multiplier_STAGE1__2528_  (.A1(sram_rdata_reg[23]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_pp1_47 [9]));
 AND2_X1 u_multiplier_STAGE1__2529_  (.A1(data_in_reg[23]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_pp1_47 [10]));
 AND2_X1 u_multiplier_STAGE1__2530_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_pp1_47 [11]));
 AND2_X1 u_multiplier_STAGE1__2531_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_pp1_47 [12]));
 AND2_X1 u_multiplier_STAGE1__2532_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_pp1_47 [13]));
 AND2_X1 u_multiplier_STAGE1__2533_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp1_47 [14]));
 AND2_X1 u_multiplier_STAGE1__2534_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp1_47 [15]));
 AND2_X1 u_multiplier_STAGE1__2535_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_48 [1]));
 AND2_X1 u_multiplier_STAGE1__2536_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_48 [2]));
 AND2_X1 u_multiplier_STAGE1__2537_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_48 [3]));
 AND2_X1 u_multiplier_STAGE1__2538_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_48 [4]));
 AND2_X1 u_multiplier_STAGE1__2539_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_pp1_48 [5]));
 AND2_X1 u_multiplier_STAGE1__2540_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_pp1_48 [6]));
 AND2_X1 u_multiplier_STAGE1__2541_  (.A1(sram_rdata_reg[23]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_pp1_48 [7]));
 AND2_X1 u_multiplier_STAGE1__2542_  (.A1(sram_rdata_reg[24]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_pp1_48 [8]));
 AND2_X1 u_multiplier_STAGE1__2543_  (.A1(data_in_reg[23]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_pp1_48 [9]));
 AND2_X1 u_multiplier_STAGE1__2544_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_pp1_48 [10]));
 AND2_X1 u_multiplier_STAGE1__2545_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_pp1_48 [11]));
 AND2_X1 u_multiplier_STAGE1__2546_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp1_48 [12]));
 AND2_X1 u_multiplier_STAGE1__2547_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp1_48 [13]));
 AND2_X1 u_multiplier_STAGE1__2548_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp1_48 [14]));
 AND2_X1 u_multiplier_STAGE1__2549_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp1_48 [15]));
 AND2_X1 u_multiplier_STAGE1__2550_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_49 [0]));
 AND2_X1 u_multiplier_STAGE1__2551_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_49 [1]));
 AND2_X1 u_multiplier_STAGE1__2552_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_49 [2]));
 AND2_X1 u_multiplier_STAGE1__2553_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_49 [3]));
 AND2_X1 u_multiplier_STAGE1__2554_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_pp1_49 [4]));
 AND2_X1 u_multiplier_STAGE1__2555_  (.A1(sram_rdata_reg[23]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_pp1_49 [5]));
 AND2_X1 u_multiplier_STAGE1__2556_  (.A1(sram_rdata_reg[24]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_pp1_49 [6]));
 AND2_X1 u_multiplier_STAGE1__2557_  (.A1(data_in_reg[24]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_pp1_49 [7]));
 AND2_X1 u_multiplier_STAGE1__2558_  (.A1(data_in_reg[23]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_pp1_49 [8]));
 AND2_X1 u_multiplier_STAGE1__2559_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_pp1_49 [9]));
 AND2_X1 u_multiplier_STAGE1__2560_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp1_49 [10]));
 AND2_X1 u_multiplier_STAGE1__2561_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp1_49 [11]));
 AND2_X1 u_multiplier_STAGE1__2562_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp1_49 [12]));
 AND2_X1 u_multiplier_STAGE1__2563_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp1_49 [13]));
 AND2_X1 u_multiplier_STAGE1__2564_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_50 [0]));
 AND2_X1 u_multiplier_STAGE1__2565_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_50 [1]));
 AND2_X1 u_multiplier_STAGE1__2566_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_50 [2]));
 AND2_X1 u_multiplier_STAGE1__2567_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_50 [3]));
 AND2_X1 u_multiplier_STAGE1__2568_  (.A1(sram_rdata_reg[23]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_pp1_50 [4]));
 AND2_X1 u_multiplier_STAGE1__2569_  (.A1(sram_rdata_reg[24]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_pp1_50 [5]));
 AND2_X1 u_multiplier_STAGE1__2570_  (.A1(sram_rdata_reg[25]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_pp1_50 [6]));
 AND2_X1 u_multiplier_STAGE1__2571_  (.A1(data_in_reg[24]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_pp1_50 [7]));
 AND2_X1 u_multiplier_STAGE1__2572_  (.A1(data_in_reg[23]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_pp1_50 [8]));
 AND2_X1 u_multiplier_STAGE1__2573_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp1_50 [9]));
 AND2_X1 u_multiplier_STAGE1__2574_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp1_50 [10]));
 AND2_X1 u_multiplier_STAGE1__2575_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp1_50 [11]));
 AND2_X1 u_multiplier_STAGE1__2576_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp2_50 [7]));
 AND2_X1 u_multiplier_STAGE1__2577_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_51 [0]));
 AND2_X1 u_multiplier_STAGE1__2578_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_51 [1]));
 AND2_X1 u_multiplier_STAGE1__2579_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_51 [2]));
 AND2_X1 u_multiplier_STAGE1__2580_  (.A1(sram_rdata_reg[23]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_51 [3]));
 AND2_X1 u_multiplier_STAGE1__2581_  (.A1(sram_rdata_reg[24]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_pp1_51 [4]));
 AND2_X1 u_multiplier_STAGE1__2582_  (.A1(sram_rdata_reg[25]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_pp1_51 [5]));
 AND2_X1 u_multiplier_STAGE1__2583_  (.A1(data_in_reg[25]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_pp1_51 [6]));
 AND2_X1 u_multiplier_STAGE1__2584_  (.A1(data_in_reg[24]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_pp1_51 [7]));
 AND2_X2 u_multiplier_STAGE1__2585_  (.A1(data_in_reg[23]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp1_51 [8]));
 AND2_X2 u_multiplier_STAGE1__2586_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp1_51 [9]));
 AND2_X1 u_multiplier_STAGE1__2587_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp2_51 [7]));
 AND2_X1 u_multiplier_STAGE1__2588_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp2_51 [6]));
 AND2_X1 u_multiplier_STAGE1__2589_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_52 [0]));
 AND2_X1 u_multiplier_STAGE1__2590_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_52 [1]));
 AND2_X1 u_multiplier_STAGE1__2591_  (.A1(sram_rdata_reg[23]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_52 [2]));
 AND2_X1 u_multiplier_STAGE1__2592_  (.A1(sram_rdata_reg[24]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_52 [3]));
 AND2_X1 u_multiplier_STAGE1__2593_  (.A1(sram_rdata_reg[25]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_pp1_52 [4]));
 AND2_X1 u_multiplier_STAGE1__2594_  (.A1(sram_rdata_reg[26]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_pp1_52 [5]));
 AND2_X1 u_multiplier_STAGE1__2595_  (.A1(data_in_reg[25]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_pp1_52 [6]));
 AND2_X1 u_multiplier_STAGE1__2596_  (.A1(data_in_reg[24]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp1_52 [7]));
 AND2_X1 u_multiplier_STAGE1__2597_  (.A1(data_in_reg[23]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp2_52 [7]));
 AND2_X1 u_multiplier_STAGE1__2598_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp2_52 [6]));
 AND2_X1 u_multiplier_STAGE1__2599_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp2_52 [5]));
 AND2_X1 u_multiplier_STAGE1__2600_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_53 [0]));
 AND2_X1 u_multiplier_STAGE1__2601_  (.A1(sram_rdata_reg[23]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_53 [1]));
 AND2_X1 u_multiplier_STAGE1__2602_  (.A1(sram_rdata_reg[24]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_53 [2]));
 AND2_X1 u_multiplier_STAGE1__2603_  (.A1(sram_rdata_reg[25]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_53 [3]));
 AND2_X1 u_multiplier_STAGE1__2604_  (.A1(sram_rdata_reg[26]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_pp1_53 [4]));
 AND2_X1 u_multiplier_STAGE1__2605_  (.A1(data_in_reg[26]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_pp1_53 [5]));
 AND2_X1 u_multiplier_STAGE1__2606_  (.A1(data_in_reg[25]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp2_53 [7]));
 AND2_X1 u_multiplier_STAGE1__2607_  (.A1(data_in_reg[24]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp2_53 [6]));
 AND2_X1 u_multiplier_STAGE1__2608_  (.A1(data_in_reg[23]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp2_53 [5]));
 AND2_X1 u_multiplier_STAGE1__2609_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp2_53 [4]));
 AND2_X1 u_multiplier_STAGE1__2610_  (.A1(sram_rdata_reg[23]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_54 [0]));
 AND2_X1 u_multiplier_STAGE1__2611_  (.A1(sram_rdata_reg[24]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_54 [1]));
 AND2_X1 u_multiplier_STAGE1__2612_  (.A1(sram_rdata_reg[25]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_54 [2]));
 AND2_X1 u_multiplier_STAGE1__2613_  (.A1(sram_rdata_reg[26]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_54 [3]));
 AND2_X1 u_multiplier_STAGE1__2614_  (.A1(sram_rdata_reg[27]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_pp2_54 [7]));
 AND2_X1 u_multiplier_STAGE1__2615_  (.A1(data_in_reg[26]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp2_54 [6]));
 AND2_X1 u_multiplier_STAGE1__2616_  (.A1(data_in_reg[25]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp2_54 [5]));
 AND2_X1 u_multiplier_STAGE1__2617_  (.A1(data_in_reg[24]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp2_54 [4]));
 AND2_X1 u_multiplier_STAGE1__2618_  (.A1(data_in_reg[23]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp2_54 [3]));
 AND2_X1 u_multiplier_STAGE1__2619_  (.A1(sram_rdata_reg[24]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_55 [0]));
 AND2_X1 u_multiplier_STAGE1__2620_  (.A1(sram_rdata_reg[25]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_55 [1]));
 AND2_X1 u_multiplier_STAGE1__2621_  (.A1(sram_rdata_reg[26]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp2_55 [7]));
 AND2_X1 u_multiplier_STAGE1__2622_  (.A1(sram_rdata_reg[27]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp2_55 [6]));
 AND2_X1 u_multiplier_STAGE1__2623_  (.A1(data_in_reg[27]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp2_55 [5]));
 AND2_X1 u_multiplier_STAGE1__2624_  (.A1(data_in_reg[26]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp2_55 [4]));
 AND2_X1 u_multiplier_STAGE1__2625_  (.A1(data_in_reg[25]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp2_55 [3]));
 AND2_X1 u_multiplier_STAGE1__2626_  (.A1(data_in_reg[24]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp2_55 [2]));
 AND2_X1 u_multiplier_STAGE1__2627_  (.A1(sram_rdata_reg[25]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp2_56 [7]));
 AND2_X1 u_multiplier_STAGE1__2628_  (.A1(sram_rdata_reg[26]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp2_56 [6]));
 AND2_X1 u_multiplier_STAGE1__2629_  (.A1(sram_rdata_reg[27]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp2_56 [5]));
 AND2_X1 u_multiplier_STAGE1__2630_  (.A1(sram_rdata_reg[28]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp2_56 [4]));
 AND2_X1 u_multiplier_STAGE1__2631_  (.A1(data_in_reg[27]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp2_56 [3]));
 AND2_X1 u_multiplier_STAGE1__2632_  (.A1(data_in_reg[26]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp2_56 [2]));
 AND2_X1 u_multiplier_STAGE1__2633_  (.A1(data_in_reg[25]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp2_56 [1]));
 AND2_X1 u_multiplier_STAGE1__2634_  (.A1(sram_rdata_reg[26]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp2_57 [5]));
 AND2_X1 u_multiplier_STAGE1__2635_  (.A1(sram_rdata_reg[27]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp2_57 [4]));
 AND2_X1 u_multiplier_STAGE1__2636_  (.A1(sram_rdata_reg[28]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp2_57 [3]));
 AND2_X1 u_multiplier_STAGE1__2637_  (.A1(data_in_reg[28]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp2_57 [2]));
 AND2_X1 u_multiplier_STAGE1__2638_  (.A1(data_in_reg[27]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp2_57 [1]));
 AND2_X1 u_multiplier_STAGE1__2639_  (.A1(data_in_reg[26]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp2_57 [0]));
 AND2_X1 u_multiplier_STAGE1__2640_  (.A1(sram_rdata_reg[27]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp3_58 [3]));
 AND2_X1 u_multiplier_STAGE1__2641_  (.A1(sram_rdata_reg[28]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp2_58 [3]));
 AND2_X1 u_multiplier_STAGE1__2642_  (.A1(sram_rdata_reg[29]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp2_58 [2]));
 AND2_X1 u_multiplier_STAGE1__2643_  (.A1(data_in_reg[28]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp2_58 [1]));
 AND2_X1 u_multiplier_STAGE1__2644_  (.A1(data_in_reg[27]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp2_58 [0]));
 AND2_X1 u_multiplier_STAGE1__2645_  (.A1(sram_rdata_reg[28]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp3_59 [2]));
 AND2_X1 u_multiplier_STAGE1__2646_  (.A1(sram_rdata_reg[29]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp3_59 [3]));
 AND2_X1 u_multiplier_STAGE1__2647_  (.A1(data_in_reg[29]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp2_59 [1]));
 AND2_X1 u_multiplier_STAGE1__2648_  (.A1(data_in_reg[28]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp2_59 [0]));
 AND2_X1 u_multiplier_STAGE1__2649_  (.A1(sram_rdata_reg[29]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp3_60 [1]));
 AND2_X1 u_multiplier_STAGE1__2650_  (.A1(sram_rdata_reg[30]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp3_60 [2]));
 AND2_X1 u_multiplier_STAGE1__2651_  (.A1(data_in_reg[29]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp3_60 [3]));
 AND2_X1 u_multiplier_STAGE1__2652_  (.A1(sram_rdata_reg[30]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp3_61 [0]));
 AND2_X1 u_multiplier_STAGE1__2653_  (.A1(data_in_reg[30]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp3_61 [1]));
 AND2_X1 u_multiplier_STAGE1__2654_  (.A1(sram_rdata_reg[31]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp3_62 ));
 LOGIC0_X1 u_multiplier_STAGE2_E_4_2_pp2_11_2__25__133  (.Z(net133));
 LOGIC0_X1 u_multiplier_STAGE2_E_4_2_pp2_11_2__18__132  (.Z(net132));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_10_1__18_  (.A(u_multiplier_STAGE2_pp2_9_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_10_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_10_1__19_  (.A1(u_multiplier_pp1_10 [1]),
    .A2(u_multiplier_pp1_10 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_10_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_10_1__20_  (.A(u_multiplier_pp1_10 [1]),
    .B(u_multiplier_pp1_10 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_10_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_10_1__21_  (.A1(u_multiplier_pp1_10 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_10_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_10_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_10_1__22_  (.A(u_multiplier_pp1_10 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_10_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_10_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_10_1__23_  (.A1(u_multiplier_pp1_10 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_10_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_10_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_10_1__24_  (.A(u_multiplier_pp1_10 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_10_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_10_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_10_1__25_  (.A(u_multiplier_STAGE2_pp2_9_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_10_1__16_ ),
    .ZN(u_multiplier_pp2_10 [1]));
 NAND2_X2 u_multiplier_STAGE2_E_4_2_pp2_10_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_10_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_10_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_10_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_10_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_10_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_10_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_10_1__17_ ),
    .ZN(u_multiplier_pp2_11 [3]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_11_1__18_  (.A(u_multiplier_STAGE2_pp2_10_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_11_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_11_1__19_  (.A1(u_multiplier_pp1_11 [1]),
    .A2(u_multiplier_pp1_11 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_11_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_11_1__20_  (.A(u_multiplier_pp1_11 [1]),
    .B(u_multiplier_pp1_11 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_11_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_11_1__21_  (.A1(u_multiplier_pp1_11 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_11_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_11_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_11_1__22_  (.A(u_multiplier_pp1_11 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_11_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_11_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_11_1__23_  (.A1(u_multiplier_pp1_11 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_11_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_11_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_11_1__24_  (.A(u_multiplier_pp1_11 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_11_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_11_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_11_1__25_  (.A(u_multiplier_STAGE2_pp2_10_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_11_1__16_ ),
    .ZN(u_multiplier_pp2_11 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_11_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_11_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_11_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_11_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_11_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_11_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_11_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_11_1__17_ ),
    .ZN(u_multiplier_pp2_12 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_11_2__18_  (.A(net132),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_11_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_11_2__19_  (.A1(u_multiplier_pp1_11 [5]),
    .A2(u_multiplier_pp1_11 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_11_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_11_2__20_  (.A(u_multiplier_pp1_11 [5]),
    .B(u_multiplier_pp1_11 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_11_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_11_2__21_  (.A1(u_multiplier_pp1_11 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_11_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_11_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_11_2__22_  (.A(u_multiplier_pp1_11 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_11_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_11_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_11_2__23_  (.A1(u_multiplier_pp1_11 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_11_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_11_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_11_2__24_  (.A(u_multiplier_pp1_11 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_11_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_11_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_11_2__25_  (.A(net133),
    .B(u_multiplier_STAGE2_E_4_2_pp2_11_2__16_ ),
    .ZN(u_multiplier_pp2_11 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_11_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_11_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_11_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_11_e42_2_cout ));
 OAI21_X1 u_multiplier_STAGE2_E_4_2_pp2_11_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_11_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_11_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_11_2__17_ ),
    .ZN(u_multiplier_pp2_12 [3]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_12_1__18_  (.A(u_multiplier_STAGE2_pp2_11_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_12_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_12_1__19_  (.A1(u_multiplier_pp1_12 [1]),
    .A2(u_multiplier_pp1_12 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_12_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_12_1__20_  (.A(u_multiplier_pp1_12 [1]),
    .B(u_multiplier_pp1_12 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_12_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_12_1__21_  (.A1(u_multiplier_pp1_12 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_12_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_12_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_12_1__22_  (.A(u_multiplier_pp1_12 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_12_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_12_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_12_1__23_  (.A1(u_multiplier_pp1_12 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_12_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_12_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_12_1__24_  (.A(u_multiplier_pp1_12 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_12_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_12_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_12_1__25_  (.A(u_multiplier_STAGE2_pp2_11_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_12_1__16_ ),
    .ZN(u_multiplier_pp2_12 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_12_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_12_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_12_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_12_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_12_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_12_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_12_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_12_1__17_ ),
    .ZN(u_multiplier_pp2_13 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_12_2__18_  (.A(u_multiplier_STAGE2_pp2_11_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_12_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_12_2__19_  (.A1(u_multiplier_pp1_12 [5]),
    .A2(u_multiplier_pp1_12 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_12_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_12_2__20_  (.A(u_multiplier_pp1_12 [5]),
    .B(u_multiplier_pp1_12 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_12_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_12_2__21_  (.A1(u_multiplier_pp1_12 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_12_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_12_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_12_2__22_  (.A(u_multiplier_pp1_12 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_12_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_12_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_12_2__23_  (.A1(u_multiplier_pp1_12 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_12_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_12_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_12_2__24_  (.A(u_multiplier_pp1_12 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_12_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_12_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_12_2__25_  (.A(u_multiplier_STAGE2_pp2_11_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_12_2__16_ ),
    .ZN(u_multiplier_pp2_12 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_12_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_12_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_12_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_12_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_12_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_12_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_12_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_12_2__17_ ),
    .ZN(u_multiplier_pp2_13 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_13_1__18_  (.A(u_multiplier_STAGE2_pp2_12_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_13_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_13_1__19_  (.A1(u_multiplier_pp1_13 [1]),
    .A2(u_multiplier_pp1_13 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_13_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_13_1__20_  (.A(u_multiplier_pp1_13 [1]),
    .B(u_multiplier_pp1_13 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_13_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_13_1__21_  (.A1(u_multiplier_pp1_13 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_13_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_13_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_13_1__22_  (.A(u_multiplier_pp1_13 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_13_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_13_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_13_1__23_  (.A1(u_multiplier_pp1_13 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_13_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_13_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_13_1__24_  (.A(u_multiplier_pp1_13 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_13_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_13_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_13_1__25_  (.A(u_multiplier_STAGE2_pp2_12_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_13_1__16_ ),
    .ZN(u_multiplier_pp2_13 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_13_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_13_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_13_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_13_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_13_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_13_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_13_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_13_1__17_ ),
    .ZN(u_multiplier_pp2_14 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_13_2__18_  (.A(u_multiplier_STAGE2_pp2_12_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_13_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_13_2__19_  (.A1(u_multiplier_pp1_13 [5]),
    .A2(u_multiplier_pp1_13 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_13_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_13_2__20_  (.A(u_multiplier_pp1_13 [5]),
    .B(u_multiplier_pp1_13 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_13_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_13_2__21_  (.A1(u_multiplier_pp1_13 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_13_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_13_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_13_2__22_  (.A(u_multiplier_pp1_13 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_13_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_13_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_13_2__23_  (.A1(u_multiplier_pp1_13 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_13_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_13_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_13_2__24_  (.A(u_multiplier_pp1_13 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_13_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_13_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_13_2__25_  (.A(u_multiplier_STAGE2_pp2_12_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_13_2__16_ ),
    .ZN(u_multiplier_pp2_13 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_13_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_13_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_13_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_13_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_13_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_13_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_13_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_13_2__17_ ),
    .ZN(u_multiplier_pp2_14 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_13_3__18_  (.A(net134),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_13_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_13_3__19_  (.A1(u_multiplier_pp1_13 [9]),
    .A2(u_multiplier_pp1_13 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_13_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_13_3__20_  (.A(u_multiplier_pp1_13 [9]),
    .B(u_multiplier_pp1_13 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_13_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_13_3__21_  (.A1(u_multiplier_pp1_13 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_13_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_13_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_13_3__22_  (.A(u_multiplier_pp1_13 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_13_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_13_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_13_3__23_  (.A1(u_multiplier_pp1_13 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_13_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_13_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_13_3__24_  (.A(u_multiplier_pp1_13 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_13_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_13_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_13_3__25_  (.A(net135),
    .B(u_multiplier_STAGE2_E_4_2_pp2_13_3__16_ ),
    .ZN(u_multiplier_pp2_13 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_13_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_13_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_13_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_13_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_13_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_13_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_13_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_13_3__17_ ),
    .ZN(u_multiplier_pp2_14 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_14_1__18_  (.A(u_multiplier_STAGE2_pp2_13_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_14_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_14_1__19_  (.A1(u_multiplier_pp1_14 [1]),
    .A2(u_multiplier_pp1_14 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_14_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_14_1__20_  (.A(u_multiplier_pp1_14 [1]),
    .B(u_multiplier_pp1_14 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_14_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_14_1__21_  (.A1(u_multiplier_pp1_14 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_14_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_14_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_14_1__22_  (.A(u_multiplier_pp1_14 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_14_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_14_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_14_1__23_  (.A1(u_multiplier_pp1_14 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_14_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_14_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_14_1__24_  (.A(u_multiplier_pp1_14 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_14_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_14_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_14_1__25_  (.A(u_multiplier_STAGE2_pp2_13_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_14_1__16_ ),
    .ZN(u_multiplier_pp2_14 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_14_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_14_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_14_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_14_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE2_E_4_2_pp2_14_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_14_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_14_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_14_1__17_ ),
    .ZN(u_multiplier_pp2_15 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_14_2__18_  (.A(u_multiplier_STAGE2_pp2_13_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_14_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_14_2__19_  (.A1(u_multiplier_pp1_14 [5]),
    .A2(u_multiplier_pp1_14 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_14_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_14_2__20_  (.A(u_multiplier_pp1_14 [5]),
    .B(u_multiplier_pp1_14 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_14_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_14_2__21_  (.A1(u_multiplier_pp1_14 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_14_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_14_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_14_2__22_  (.A(u_multiplier_pp1_14 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_14_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_14_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_14_2__23_  (.A1(u_multiplier_pp1_14 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_14_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_14_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_14_2__24_  (.A(u_multiplier_pp1_14 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_14_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_14_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_14_2__25_  (.A(u_multiplier_STAGE2_pp2_13_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_14_2__16_ ),
    .ZN(u_multiplier_pp2_14 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_14_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_14_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_14_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_14_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_14_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_14_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_14_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_14_2__17_ ),
    .ZN(u_multiplier_pp2_15 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_14_3__18_  (.A(u_multiplier_STAGE2_pp2_13_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_14_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_14_3__19_  (.A1(u_multiplier_pp1_14 [9]),
    .A2(u_multiplier_pp1_14 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_14_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_14_3__20_  (.A(u_multiplier_pp1_14 [9]),
    .B(u_multiplier_pp1_14 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_14_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_14_3__21_  (.A1(u_multiplier_pp1_14 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_14_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_14_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_14_3__22_  (.A(u_multiplier_pp1_14 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_14_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_14_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_14_3__23_  (.A1(u_multiplier_pp1_14 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_14_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_14_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_14_3__24_  (.A(u_multiplier_pp1_14 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_14_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_14_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_14_3__25_  (.A(u_multiplier_STAGE2_pp2_13_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_14_3__16_ ),
    .ZN(u_multiplier_pp2_14 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_14_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_14_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_14_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_14_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_14_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_14_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_14_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_14_3__17_ ),
    .ZN(u_multiplier_pp2_15 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_15_1__18_  (.A(u_multiplier_STAGE2_pp2_14_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_15_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_15_1__19_  (.A1(u_multiplier_pp1_15 [1]),
    .A2(u_multiplier_pp1_15 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_15_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_15_1__20_  (.A(u_multiplier_pp1_15 [1]),
    .B(u_multiplier_pp1_15 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_15_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_15_1__21_  (.A1(u_multiplier_pp1_15 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_15_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_15_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_15_1__22_  (.A(u_multiplier_pp1_15 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_15_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_15_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_15_1__23_  (.A1(u_multiplier_pp1_15 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_15_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_15_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_15_1__24_  (.A(u_multiplier_pp1_15 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_15_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_15_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_15_1__25_  (.A(u_multiplier_STAGE2_pp2_14_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_15_1__16_ ),
    .ZN(u_multiplier_pp2_15 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_15_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_15_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_15_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_15_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_15_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_15_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_15_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_15_1__17_ ),
    .ZN(u_multiplier_pp2_16 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_15_2__18_  (.A(u_multiplier_STAGE2_pp2_14_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_15_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_15_2__19_  (.A1(u_multiplier_pp1_15 [5]),
    .A2(u_multiplier_pp1_15 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_15_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_15_2__20_  (.A(u_multiplier_pp1_15 [5]),
    .B(u_multiplier_pp1_15 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_15_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_15_2__21_  (.A1(u_multiplier_pp1_15 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_15_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_15_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_15_2__22_  (.A(u_multiplier_pp1_15 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_15_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_15_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_15_2__23_  (.A1(u_multiplier_pp1_15 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_15_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_15_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_15_2__24_  (.A(u_multiplier_pp1_15 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_15_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_15_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_15_2__25_  (.A(u_multiplier_STAGE2_pp2_14_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_15_2__16_ ),
    .ZN(u_multiplier_pp2_15 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_15_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_15_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_15_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_15_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_15_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_15_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_15_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_15_2__17_ ),
    .ZN(u_multiplier_pp2_16 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_15_3__18_  (.A(u_multiplier_STAGE2_pp2_14_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_15_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_15_3__19_  (.A1(u_multiplier_pp1_15 [9]),
    .A2(u_multiplier_pp1_15 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_15_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_15_3__20_  (.A(u_multiplier_pp1_15 [9]),
    .B(u_multiplier_pp1_15 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_15_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_15_3__21_  (.A1(u_multiplier_pp1_15 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_15_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_15_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_15_3__22_  (.A(u_multiplier_pp1_15 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_15_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_15_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_15_3__23_  (.A1(u_multiplier_pp1_15 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_15_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_15_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_15_3__24_  (.A(u_multiplier_pp1_15 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_15_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_15_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_15_3__25_  (.A(u_multiplier_STAGE2_pp2_14_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_15_3__16_ ),
    .ZN(u_multiplier_pp2_15 [1]));
 NAND2_X2 u_multiplier_STAGE2_E_4_2_pp2_15_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_15_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_15_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_15_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_15_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_15_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_15_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_15_3__17_ ),
    .ZN(u_multiplier_pp2_16 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_15_4__18_  (.A(net136),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_15_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_15_4__19_  (.A1(u_multiplier_pp1_15 [13]),
    .A2(u_multiplier_pp1_15 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_15_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_15_4__20_  (.A(u_multiplier_pp1_15 [13]),
    .B(u_multiplier_pp1_15 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_15_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_15_4__21_  (.A1(u_multiplier_pp1_15 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_15_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_15_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_15_4__22_  (.A(u_multiplier_pp1_15 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_15_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_15_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_15_4__23_  (.A1(u_multiplier_pp1_15 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_15_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_15_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_15_4__24_  (.A(u_multiplier_pp1_15 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_15_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_15_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_15_4__25_  (.A(net137),
    .B(u_multiplier_STAGE2_E_4_2_pp2_15_4__16_ ),
    .ZN(u_multiplier_pp2_15 [0]));
 NAND2_X2 u_multiplier_STAGE2_E_4_2_pp2_15_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_15_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_15_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_15_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_15_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_15_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_15_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_15_4__17_ ),
    .ZN(u_multiplier_pp2_16 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_16_1__18_  (.A(u_multiplier_STAGE2_pp2_15_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_16_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_16_1__19_  (.A1(u_multiplier_pp1_16 [1]),
    .A2(u_multiplier_pp1_16 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_16_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_16_1__20_  (.A(u_multiplier_pp1_16 [1]),
    .B(u_multiplier_pp1_16 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_16_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_16_1__21_  (.A1(u_multiplier_pp1_16 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_16_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_16_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_16_1__22_  (.A(u_multiplier_pp1_16 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_16_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_16_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_16_1__23_  (.A1(u_multiplier_pp1_16 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_16_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_16_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_16_1__24_  (.A(u_multiplier_pp1_16 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_16_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_16_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_16_1__25_  (.A(u_multiplier_STAGE2_pp2_15_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_16_1__16_ ),
    .ZN(u_multiplier_pp2_16 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_16_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_16_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_16_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_16_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE2_E_4_2_pp2_16_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_16_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_16_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_16_1__17_ ),
    .ZN(u_multiplier_pp2_17 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_16_2__18_  (.A(u_multiplier_STAGE2_pp2_15_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_16_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_16_2__19_  (.A1(u_multiplier_pp1_16 [5]),
    .A2(u_multiplier_pp1_16 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_16_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_16_2__20_  (.A(u_multiplier_pp1_16 [5]),
    .B(u_multiplier_pp1_16 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_16_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_16_2__21_  (.A1(u_multiplier_pp1_16 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_16_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_16_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_16_2__22_  (.A(u_multiplier_pp1_16 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_16_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_16_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_16_2__23_  (.A1(u_multiplier_pp1_16 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_16_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_16_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_16_2__24_  (.A(u_multiplier_pp1_16 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_16_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_16_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_16_2__25_  (.A(u_multiplier_STAGE2_pp2_15_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_16_2__16_ ),
    .ZN(u_multiplier_pp2_16 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_16_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_16_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_16_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_16_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_16_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_16_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_16_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_16_2__17_ ),
    .ZN(u_multiplier_pp2_17 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_16_3__18_  (.A(u_multiplier_STAGE2_pp2_15_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_16_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_16_3__19_  (.A1(u_multiplier_pp1_16 [9]),
    .A2(u_multiplier_pp1_16 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_16_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_16_3__20_  (.A(u_multiplier_pp1_16 [9]),
    .B(u_multiplier_pp1_16 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_16_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_16_3__21_  (.A1(u_multiplier_pp1_16 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_16_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_16_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_16_3__22_  (.A(u_multiplier_pp1_16 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_16_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_16_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_16_3__23_  (.A1(u_multiplier_pp1_16 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_16_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_16_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_16_3__24_  (.A(u_multiplier_pp1_16 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_16_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_16_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_16_3__25_  (.A(u_multiplier_STAGE2_pp2_15_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_16_3__16_ ),
    .ZN(u_multiplier_pp2_16 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_16_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_16_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_16_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_16_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_16_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_16_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_16_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_16_3__17_ ),
    .ZN(u_multiplier_pp2_17 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_16_4__18_  (.A(u_multiplier_STAGE2_pp2_15_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_16_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_16_4__19_  (.A1(u_multiplier_pp1_16 [13]),
    .A2(u_multiplier_pp1_16 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_16_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_16_4__20_  (.A(u_multiplier_pp1_16 [13]),
    .B(u_multiplier_pp1_16 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_16_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_16_4__21_  (.A1(u_multiplier_pp1_16 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_16_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_16_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_16_4__22_  (.A(u_multiplier_pp1_16 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_16_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_16_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_16_4__23_  (.A1(u_multiplier_pp1_16 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_16_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_16_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_16_4__24_  (.A(u_multiplier_pp1_16 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_16_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_16_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_16_4__25_  (.A(u_multiplier_STAGE2_pp2_15_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_16_4__16_ ),
    .ZN(u_multiplier_pp2_16 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_16_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_16_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_16_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_16_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_16_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_16_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_16_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_16_4__17_ ),
    .ZN(u_multiplier_pp2_17 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_17_1__18_  (.A(u_multiplier_STAGE2_pp2_16_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_17_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_17_1__19_  (.A1(u_multiplier_pp1_17 [1]),
    .A2(u_multiplier_pp1_17 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_17_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_17_1__20_  (.A(u_multiplier_pp1_17 [1]),
    .B(u_multiplier_pp1_17 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_17_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_17_1__21_  (.A1(u_multiplier_pp1_17 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_17_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_17_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_17_1__22_  (.A(u_multiplier_pp1_17 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_17_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_17_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_17_1__23_  (.A1(u_multiplier_pp1_17 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_17_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_17_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_17_1__24_  (.A(u_multiplier_pp1_17 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_17_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_17_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_17_1__25_  (.A(u_multiplier_STAGE2_pp2_16_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_17_1__16_ ),
    .ZN(u_multiplier_pp2_17 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_17_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_17_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_17_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_17_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE2_E_4_2_pp2_17_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_17_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_17_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_17_1__17_ ),
    .ZN(u_multiplier_pp2_18 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_17_2__18_  (.A(u_multiplier_STAGE2_pp2_16_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_17_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_17_2__19_  (.A1(u_multiplier_pp1_17 [5]),
    .A2(u_multiplier_pp1_17 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_17_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_17_2__20_  (.A(u_multiplier_pp1_17 [5]),
    .B(u_multiplier_pp1_17 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_17_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_17_2__21_  (.A1(u_multiplier_pp1_17 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_17_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_17_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_17_2__22_  (.A(u_multiplier_pp1_17 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_17_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_17_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_17_2__23_  (.A1(u_multiplier_pp1_17 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_17_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_17_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_17_2__24_  (.A(u_multiplier_pp1_17 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_17_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_17_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_17_2__25_  (.A(u_multiplier_STAGE2_pp2_16_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_17_2__16_ ),
    .ZN(u_multiplier_pp2_17 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_17_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_17_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_17_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_17_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_17_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_17_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_17_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_17_2__17_ ),
    .ZN(u_multiplier_pp2_18 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_17_3__18_  (.A(u_multiplier_STAGE2_pp2_16_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_17_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_17_3__19_  (.A1(u_multiplier_pp1_17 [9]),
    .A2(u_multiplier_pp1_17 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_17_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_17_3__20_  (.A(u_multiplier_pp1_17 [9]),
    .B(u_multiplier_pp1_17 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_17_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_17_3__21_  (.A1(u_multiplier_pp1_17 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_17_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_17_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_17_3__22_  (.A(u_multiplier_pp1_17 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_17_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_17_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_17_3__23_  (.A1(u_multiplier_pp1_17 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_17_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_17_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_17_3__24_  (.A(u_multiplier_pp1_17 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_17_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_17_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_17_3__25_  (.A(u_multiplier_STAGE2_pp2_16_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_17_3__16_ ),
    .ZN(u_multiplier_pp2_17 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_17_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_17_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_17_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_17_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_17_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_17_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_17_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_17_3__17_ ),
    .ZN(u_multiplier_pp2_18 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_17_4__18_  (.A(u_multiplier_STAGE2_pp2_16_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_17_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_17_4__19_  (.A1(u_multiplier_pp1_17 [13]),
    .A2(u_multiplier_pp1_17 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_17_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_17_4__20_  (.A(u_multiplier_pp1_17 [13]),
    .B(u_multiplier_pp1_17 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_17_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_17_4__21_  (.A1(u_multiplier_pp1_17 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_17_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_17_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_17_4__22_  (.A(u_multiplier_pp1_17 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_17_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_17_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_17_4__23_  (.A1(u_multiplier_pp1_17 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_17_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_17_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_17_4__24_  (.A(u_multiplier_pp1_17 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_17_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_17_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_17_4__25_  (.A(u_multiplier_STAGE2_pp2_16_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_17_4__16_ ),
    .ZN(u_multiplier_pp2_17 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_17_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_17_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_17_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_17_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_17_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_17_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_17_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_17_4__17_ ),
    .ZN(u_multiplier_pp2_18 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_18_1__18_  (.A(u_multiplier_STAGE2_pp2_17_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_18_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_18_1__19_  (.A1(u_multiplier_pp1_18 [1]),
    .A2(u_multiplier_pp1_18 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_18_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_18_1__20_  (.A(u_multiplier_pp1_18 [1]),
    .B(u_multiplier_pp1_18 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_18_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_18_1__21_  (.A1(u_multiplier_pp1_18 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_18_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_18_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_18_1__22_  (.A(u_multiplier_pp1_18 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_18_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_18_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_18_1__23_  (.A1(u_multiplier_pp1_18 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_18_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_18_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_18_1__24_  (.A(u_multiplier_pp1_18 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_18_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_18_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_18_1__25_  (.A(u_multiplier_STAGE2_pp2_17_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_18_1__16_ ),
    .ZN(u_multiplier_pp2_18 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_18_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_18_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_18_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_18_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE2_E_4_2_pp2_18_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_18_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_18_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_18_1__17_ ),
    .ZN(u_multiplier_pp2_19 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_18_2__18_  (.A(u_multiplier_STAGE2_pp2_17_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_18_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_18_2__19_  (.A1(u_multiplier_pp1_18 [5]),
    .A2(u_multiplier_pp1_18 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_18_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_18_2__20_  (.A(u_multiplier_pp1_18 [5]),
    .B(u_multiplier_pp1_18 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_18_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_18_2__21_  (.A1(u_multiplier_pp1_18 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_18_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_18_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_18_2__22_  (.A(u_multiplier_pp1_18 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_18_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_18_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_18_2__23_  (.A1(u_multiplier_pp1_18 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_18_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_18_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_18_2__24_  (.A(u_multiplier_pp1_18 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_18_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_18_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_18_2__25_  (.A(u_multiplier_STAGE2_pp2_17_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_18_2__16_ ),
    .ZN(u_multiplier_pp2_18 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_18_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_18_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_18_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_18_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_18_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_18_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_18_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_18_2__17_ ),
    .ZN(u_multiplier_pp2_19 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_18_3__18_  (.A(u_multiplier_STAGE2_pp2_17_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_18_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_18_3__19_  (.A1(u_multiplier_pp1_18 [9]),
    .A2(u_multiplier_pp1_18 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_18_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_18_3__20_  (.A(u_multiplier_pp1_18 [9]),
    .B(u_multiplier_pp1_18 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_18_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_18_3__21_  (.A1(u_multiplier_pp1_18 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_18_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_18_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_18_3__22_  (.A(u_multiplier_pp1_18 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_18_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_18_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_18_3__23_  (.A1(u_multiplier_pp1_18 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_18_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_18_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_18_3__24_  (.A(u_multiplier_pp1_18 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_18_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_18_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_18_3__25_  (.A(u_multiplier_STAGE2_pp2_17_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_18_3__16_ ),
    .ZN(u_multiplier_pp2_18 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_18_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_18_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_18_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_18_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_18_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_18_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_18_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_18_3__17_ ),
    .ZN(u_multiplier_pp2_19 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_18_4__18_  (.A(u_multiplier_STAGE2_pp2_17_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_18_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_18_4__19_  (.A1(u_multiplier_pp1_18 [13]),
    .A2(u_multiplier_pp1_18 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_18_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_18_4__20_  (.A(u_multiplier_pp1_18 [13]),
    .B(u_multiplier_pp1_18 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_18_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_18_4__21_  (.A1(u_multiplier_pp1_18 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_18_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_18_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_18_4__22_  (.A(u_multiplier_pp1_18 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_18_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_18_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_18_4__23_  (.A1(u_multiplier_pp1_18 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_18_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_18_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_18_4__24_  (.A(u_multiplier_pp1_18 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_18_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_18_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_18_4__25_  (.A(u_multiplier_STAGE2_pp2_17_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_18_4__16_ ),
    .ZN(u_multiplier_pp2_18 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_18_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_18_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_18_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_18_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_18_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_18_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_18_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_18_4__17_ ),
    .ZN(u_multiplier_pp2_19 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_19_1__18_  (.A(u_multiplier_STAGE2_pp2_18_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_19_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_19_1__19_  (.A1(u_multiplier_pp1_19 [1]),
    .A2(u_multiplier_pp1_19 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_19_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_19_1__20_  (.A(u_multiplier_pp1_19 [1]),
    .B(u_multiplier_pp1_19 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_19_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_19_1__21_  (.A1(u_multiplier_pp1_19 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_19_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_19_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_19_1__22_  (.A(u_multiplier_pp1_19 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_19_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_19_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_19_1__23_  (.A1(u_multiplier_pp1_19 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_19_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_19_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_19_1__24_  (.A(u_multiplier_pp1_19 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_19_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_19_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_19_1__25_  (.A(u_multiplier_STAGE2_pp2_18_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_19_1__16_ ),
    .ZN(u_multiplier_pp2_19 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_19_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_19_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_19_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_19_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_19_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_19_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_19_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_19_1__17_ ),
    .ZN(u_multiplier_pp2_20 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_19_2__18_  (.A(u_multiplier_STAGE2_pp2_18_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_19_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_19_2__19_  (.A1(u_multiplier_pp1_19 [5]),
    .A2(u_multiplier_pp1_19 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_19_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_19_2__20_  (.A(u_multiplier_pp1_19 [5]),
    .B(u_multiplier_pp1_19 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_19_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_19_2__21_  (.A1(u_multiplier_pp1_19 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_19_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_19_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_19_2__22_  (.A(u_multiplier_pp1_19 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_19_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_19_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_19_2__23_  (.A1(u_multiplier_pp1_19 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_19_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_19_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_19_2__24_  (.A(u_multiplier_pp1_19 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_19_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_19_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_19_2__25_  (.A(u_multiplier_STAGE2_pp2_18_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_19_2__16_ ),
    .ZN(u_multiplier_pp2_19 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_19_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_19_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_19_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_19_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_19_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_19_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_19_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_19_2__17_ ),
    .ZN(u_multiplier_pp2_20 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_19_3__18_  (.A(u_multiplier_STAGE2_pp2_18_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_19_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_19_3__19_  (.A1(u_multiplier_pp1_19 [9]),
    .A2(u_multiplier_pp1_19 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_19_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_19_3__20_  (.A(u_multiplier_pp1_19 [9]),
    .B(u_multiplier_pp1_19 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_19_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_19_3__21_  (.A1(u_multiplier_pp1_19 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_19_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_19_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_19_3__22_  (.A(u_multiplier_pp1_19 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_19_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_19_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_19_3__23_  (.A1(u_multiplier_pp1_19 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_19_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_19_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_19_3__24_  (.A(u_multiplier_pp1_19 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_19_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_19_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_19_3__25_  (.A(u_multiplier_STAGE2_pp2_18_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_19_3__16_ ),
    .ZN(u_multiplier_pp2_19 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_19_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_19_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_19_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_19_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_19_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_19_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_19_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_19_3__17_ ),
    .ZN(u_multiplier_pp2_20 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_19_4__18_  (.A(u_multiplier_STAGE2_pp2_18_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_19_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_19_4__19_  (.A1(u_multiplier_pp1_19 [13]),
    .A2(u_multiplier_pp1_19 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_19_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_19_4__20_  (.A(u_multiplier_pp1_19 [13]),
    .B(u_multiplier_pp1_19 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_19_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_19_4__21_  (.A1(u_multiplier_pp1_19 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_19_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_19_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_19_4__22_  (.A(u_multiplier_pp1_19 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_19_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_19_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_19_4__23_  (.A1(u_multiplier_pp1_19 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_19_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_19_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_19_4__24_  (.A(u_multiplier_pp1_19 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_19_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_19_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_19_4__25_  (.A(u_multiplier_STAGE2_pp2_18_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_19_4__16_ ),
    .ZN(u_multiplier_pp2_19 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_19_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_19_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_19_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_19_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_19_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_19_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_19_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_19_4__17_ ),
    .ZN(u_multiplier_pp2_20 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_20_1__18_  (.A(u_multiplier_STAGE2_pp2_19_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_20_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_20_1__19_  (.A1(u_multiplier_pp1_20 [1]),
    .A2(u_multiplier_pp1_20 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_20_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_20_1__20_  (.A(u_multiplier_pp1_20 [1]),
    .B(u_multiplier_pp1_20 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_20_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_20_1__21_  (.A1(u_multiplier_pp1_20 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_20_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_20_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_20_1__22_  (.A(u_multiplier_pp1_20 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_20_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_20_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_20_1__23_  (.A1(u_multiplier_pp1_20 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_20_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_20_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_20_1__24_  (.A(u_multiplier_pp1_20 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_20_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_20_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_20_1__25_  (.A(u_multiplier_STAGE2_pp2_19_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_20_1__16_ ),
    .ZN(u_multiplier_pp2_20 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_20_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_20_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_20_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_20_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_20_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_20_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_20_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_20_1__17_ ),
    .ZN(u_multiplier_pp2_21 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_20_2__18_  (.A(u_multiplier_STAGE2_pp2_19_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_20_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_20_2__19_  (.A1(u_multiplier_pp1_20 [5]),
    .A2(u_multiplier_pp1_20 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_20_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_20_2__20_  (.A(u_multiplier_pp1_20 [5]),
    .B(u_multiplier_pp1_20 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_20_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_20_2__21_  (.A1(u_multiplier_pp1_20 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_20_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_20_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_20_2__22_  (.A(u_multiplier_pp1_20 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_20_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_20_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_20_2__23_  (.A1(u_multiplier_pp1_20 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_20_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_20_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_20_2__24_  (.A(u_multiplier_pp1_20 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_20_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_20_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_20_2__25_  (.A(u_multiplier_STAGE2_pp2_19_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_20_2__16_ ),
    .ZN(u_multiplier_pp2_20 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_20_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_20_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_20_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_20_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_20_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_20_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_20_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_20_2__17_ ),
    .ZN(u_multiplier_pp2_21 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_20_3__18_  (.A(u_multiplier_STAGE2_pp2_19_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_20_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_20_3__19_  (.A1(u_multiplier_pp1_20 [9]),
    .A2(u_multiplier_pp1_20 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_20_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_20_3__20_  (.A(u_multiplier_pp1_20 [9]),
    .B(u_multiplier_pp1_20 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_20_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_20_3__21_  (.A1(u_multiplier_pp1_20 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_20_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_20_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_20_3__22_  (.A(u_multiplier_pp1_20 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_20_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_20_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_20_3__23_  (.A1(u_multiplier_pp1_20 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_20_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_20_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_20_3__24_  (.A(u_multiplier_pp1_20 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_20_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_20_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_20_3__25_  (.A(u_multiplier_STAGE2_pp2_19_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_20_3__16_ ),
    .ZN(u_multiplier_pp2_20 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_20_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_20_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_20_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_20_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_20_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_20_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_20_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_20_3__17_ ),
    .ZN(u_multiplier_pp2_21 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_20_4__18_  (.A(u_multiplier_STAGE2_pp2_19_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_20_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_20_4__19_  (.A1(u_multiplier_pp1_20 [13]),
    .A2(u_multiplier_pp1_20 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_20_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_20_4__20_  (.A(u_multiplier_pp1_20 [13]),
    .B(u_multiplier_pp1_20 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_20_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_20_4__21_  (.A1(u_multiplier_pp1_20 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_20_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_20_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_20_4__22_  (.A(u_multiplier_pp1_20 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_20_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_20_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_20_4__23_  (.A1(u_multiplier_pp1_20 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_20_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_20_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_20_4__24_  (.A(u_multiplier_pp1_20 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_20_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_20_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_20_4__25_  (.A(u_multiplier_STAGE2_pp2_19_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_20_4__16_ ),
    .ZN(u_multiplier_pp2_20 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_20_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_20_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_20_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_20_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_20_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_20_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_20_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_20_4__17_ ),
    .ZN(u_multiplier_pp2_21 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_21_1__18_  (.A(u_multiplier_STAGE2_pp2_20_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_21_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_21_1__19_  (.A1(u_multiplier_pp1_21 [1]),
    .A2(u_multiplier_pp1_21 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_21_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_21_1__20_  (.A(u_multiplier_pp1_21 [1]),
    .B(u_multiplier_pp1_21 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_21_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_21_1__21_  (.A1(u_multiplier_pp1_21 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_21_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_21_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_21_1__22_  (.A(u_multiplier_pp1_21 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_21_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_21_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_21_1__23_  (.A1(u_multiplier_pp1_21 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_21_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_21_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_21_1__24_  (.A(u_multiplier_pp1_21 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_21_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_21_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_21_1__25_  (.A(u_multiplier_STAGE2_pp2_20_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_21_1__16_ ),
    .ZN(u_multiplier_pp2_21 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_21_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_21_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_21_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_21_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_21_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_21_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_21_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_21_1__17_ ),
    .ZN(u_multiplier_pp2_22 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_21_2__18_  (.A(u_multiplier_STAGE2_pp2_20_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_21_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_21_2__19_  (.A1(u_multiplier_pp1_21 [5]),
    .A2(u_multiplier_pp1_21 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_21_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_21_2__20_  (.A(u_multiplier_pp1_21 [5]),
    .B(u_multiplier_pp1_21 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_21_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_21_2__21_  (.A1(u_multiplier_pp1_21 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_21_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_21_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_21_2__22_  (.A(u_multiplier_pp1_21 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_21_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_21_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_21_2__23_  (.A1(u_multiplier_pp1_21 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_21_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_21_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_21_2__24_  (.A(u_multiplier_pp1_21 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_21_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_21_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_21_2__25_  (.A(u_multiplier_STAGE2_pp2_20_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_21_2__16_ ),
    .ZN(u_multiplier_pp2_21 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_21_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_21_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_21_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_21_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_21_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_21_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_21_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_21_2__17_ ),
    .ZN(u_multiplier_pp2_22 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_21_3__18_  (.A(u_multiplier_STAGE2_pp2_20_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_21_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_21_3__19_  (.A1(u_multiplier_pp1_21 [9]),
    .A2(u_multiplier_pp1_21 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_21_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_21_3__20_  (.A(u_multiplier_pp1_21 [9]),
    .B(u_multiplier_pp1_21 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_21_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_21_3__21_  (.A1(u_multiplier_pp1_21 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_21_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_21_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_21_3__22_  (.A(u_multiplier_pp1_21 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_21_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_21_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_21_3__23_  (.A1(u_multiplier_pp1_21 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_21_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_21_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_21_3__24_  (.A(u_multiplier_pp1_21 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_21_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_21_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_21_3__25_  (.A(u_multiplier_STAGE2_pp2_20_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_21_3__16_ ),
    .ZN(u_multiplier_pp2_21 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_21_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_21_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_21_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_21_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_21_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_21_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_21_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_21_3__17_ ),
    .ZN(u_multiplier_pp2_22 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_21_4__18_  (.A(u_multiplier_STAGE2_pp2_20_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_21_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_21_4__19_  (.A1(u_multiplier_pp1_21 [13]),
    .A2(u_multiplier_pp1_21 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_21_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_21_4__20_  (.A(u_multiplier_pp1_21 [13]),
    .B(u_multiplier_pp1_21 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_21_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_21_4__21_  (.A1(u_multiplier_pp1_21 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_21_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_21_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_21_4__22_  (.A(u_multiplier_pp1_21 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_21_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_21_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_21_4__23_  (.A1(u_multiplier_pp1_21 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_21_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_21_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_21_4__24_  (.A(u_multiplier_pp1_21 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_21_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_21_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_21_4__25_  (.A(u_multiplier_STAGE2_pp2_20_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_21_4__16_ ),
    .ZN(u_multiplier_pp2_21 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_21_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_21_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_21_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_21_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_21_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_21_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_21_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_21_4__17_ ),
    .ZN(u_multiplier_pp2_22 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_22_1__18_  (.A(u_multiplier_STAGE2_pp2_21_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_22_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_22_1__19_  (.A1(u_multiplier_pp1_22 [1]),
    .A2(u_multiplier_pp1_22 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_22_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_22_1__20_  (.A(u_multiplier_pp1_22 [1]),
    .B(u_multiplier_pp1_22 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_22_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_22_1__21_  (.A1(u_multiplier_pp1_22 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_22_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_22_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_22_1__22_  (.A(u_multiplier_pp1_22 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_22_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_22_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_22_1__23_  (.A1(u_multiplier_pp1_22 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_22_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_22_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_22_1__24_  (.A(u_multiplier_pp1_22 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_22_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_22_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_22_1__25_  (.A(u_multiplier_STAGE2_pp2_21_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_22_1__16_ ),
    .ZN(u_multiplier_pp2_22 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_22_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_22_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_22_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_22_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_22_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_22_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_22_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_22_1__17_ ),
    .ZN(u_multiplier_pp2_23 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_22_2__18_  (.A(u_multiplier_STAGE2_pp2_21_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_22_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_22_2__19_  (.A1(u_multiplier_pp1_22 [5]),
    .A2(u_multiplier_pp1_22 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_22_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_22_2__20_  (.A(u_multiplier_pp1_22 [5]),
    .B(u_multiplier_pp1_22 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_22_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_22_2__21_  (.A1(u_multiplier_pp1_22 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_22_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_22_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_22_2__22_  (.A(u_multiplier_pp1_22 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_22_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_22_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_22_2__23_  (.A1(u_multiplier_pp1_22 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_22_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_22_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_22_2__24_  (.A(u_multiplier_pp1_22 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_22_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_22_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_22_2__25_  (.A(u_multiplier_STAGE2_pp2_21_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_22_2__16_ ),
    .ZN(u_multiplier_pp2_22 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_22_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_22_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_22_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_22_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_22_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_22_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_22_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_22_2__17_ ),
    .ZN(u_multiplier_pp2_23 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_22_3__18_  (.A(u_multiplier_STAGE2_pp2_21_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_22_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_22_3__19_  (.A1(u_multiplier_pp1_22 [9]),
    .A2(u_multiplier_pp1_22 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_22_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_22_3__20_  (.A(u_multiplier_pp1_22 [9]),
    .B(u_multiplier_pp1_22 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_22_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_22_3__21_  (.A1(u_multiplier_pp1_22 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_22_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_22_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_22_3__22_  (.A(u_multiplier_pp1_22 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_22_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_22_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_22_3__23_  (.A1(u_multiplier_pp1_22 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_22_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_22_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_22_3__24_  (.A(u_multiplier_pp1_22 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_22_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_22_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_22_3__25_  (.A(u_multiplier_STAGE2_pp2_21_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_22_3__16_ ),
    .ZN(u_multiplier_pp2_22 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_22_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_22_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_22_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_22_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_22_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_22_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_22_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_22_3__17_ ),
    .ZN(u_multiplier_pp2_23 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_22_4__18_  (.A(u_multiplier_STAGE2_pp2_21_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_22_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_22_4__19_  (.A1(u_multiplier_pp1_22 [13]),
    .A2(u_multiplier_pp1_22 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_22_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_22_4__20_  (.A(u_multiplier_pp1_22 [13]),
    .B(u_multiplier_pp1_22 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_22_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_22_4__21_  (.A1(u_multiplier_pp1_22 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_22_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_22_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_22_4__22_  (.A(u_multiplier_pp1_22 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_22_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_22_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_22_4__23_  (.A1(u_multiplier_pp1_22 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_22_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_22_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_22_4__24_  (.A(u_multiplier_pp1_22 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_22_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_22_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_22_4__25_  (.A(u_multiplier_STAGE2_pp2_21_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_22_4__16_ ),
    .ZN(u_multiplier_pp2_22 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_22_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_22_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_22_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_22_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_22_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_22_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_22_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_22_4__17_ ),
    .ZN(u_multiplier_pp2_23 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_23_1__18_  (.A(u_multiplier_STAGE2_pp2_22_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_23_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_23_1__19_  (.A1(u_multiplier_pp1_23 [1]),
    .A2(u_multiplier_pp1_23 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_23_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_23_1__20_  (.A(u_multiplier_pp1_23 [1]),
    .B(u_multiplier_pp1_23 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_23_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_23_1__21_  (.A1(u_multiplier_pp1_23 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_23_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_23_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_23_1__22_  (.A(u_multiplier_pp1_23 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_23_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_23_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_23_1__23_  (.A1(u_multiplier_pp1_23 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_23_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_23_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_23_1__24_  (.A(u_multiplier_pp1_23 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_23_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_23_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_23_1__25_  (.A(u_multiplier_STAGE2_pp2_22_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_23_1__16_ ),
    .ZN(u_multiplier_pp2_23 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_23_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_23_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_23_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_23_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_23_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_23_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_23_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_23_1__17_ ),
    .ZN(u_multiplier_pp2_24 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_23_2__18_  (.A(u_multiplier_STAGE2_pp2_22_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_23_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_23_2__19_  (.A1(u_multiplier_pp1_23 [5]),
    .A2(u_multiplier_pp1_23 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_23_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_23_2__20_  (.A(u_multiplier_pp1_23 [5]),
    .B(u_multiplier_pp1_23 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_23_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_23_2__21_  (.A1(u_multiplier_pp1_23 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_23_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_23_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_23_2__22_  (.A(u_multiplier_pp1_23 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_23_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_23_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_23_2__23_  (.A1(u_multiplier_pp1_23 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_23_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_23_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_23_2__24_  (.A(u_multiplier_pp1_23 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_23_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_23_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_23_2__25_  (.A(u_multiplier_STAGE2_pp2_22_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_23_2__16_ ),
    .ZN(u_multiplier_pp2_23 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_23_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_23_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_23_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_23_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_23_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_23_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_23_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_23_2__17_ ),
    .ZN(u_multiplier_pp2_24 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_23_3__18_  (.A(u_multiplier_STAGE2_pp2_22_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_23_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_23_3__19_  (.A1(u_multiplier_pp1_23 [9]),
    .A2(u_multiplier_pp1_23 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_23_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_23_3__20_  (.A(u_multiplier_pp1_23 [9]),
    .B(u_multiplier_pp1_23 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_23_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_23_3__21_  (.A1(u_multiplier_pp1_23 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_23_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_23_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_23_3__22_  (.A(u_multiplier_pp1_23 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_23_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_23_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_23_3__23_  (.A1(u_multiplier_pp1_23 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_23_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_23_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_23_3__24_  (.A(u_multiplier_pp1_23 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_23_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_23_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_23_3__25_  (.A(u_multiplier_STAGE2_pp2_22_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_23_3__16_ ),
    .ZN(u_multiplier_pp2_23 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_23_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_23_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_23_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_23_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_23_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_23_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_23_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_23_3__17_ ),
    .ZN(u_multiplier_pp2_24 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_23_4__18_  (.A(u_multiplier_STAGE2_pp2_22_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_23_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_23_4__19_  (.A1(u_multiplier_pp1_23 [13]),
    .A2(u_multiplier_pp1_23 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_23_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_23_4__20_  (.A(u_multiplier_pp1_23 [13]),
    .B(u_multiplier_pp1_23 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_23_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_23_4__21_  (.A1(u_multiplier_pp1_23 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_23_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_23_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_23_4__22_  (.A(u_multiplier_pp1_23 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_23_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_23_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_23_4__23_  (.A1(u_multiplier_pp1_23 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_23_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_23_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_23_4__24_  (.A(u_multiplier_pp1_23 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_23_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_23_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_23_4__25_  (.A(u_multiplier_STAGE2_pp2_22_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_23_4__16_ ),
    .ZN(u_multiplier_pp2_23 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_23_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_23_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_23_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_23_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_23_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_23_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_23_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_23_4__17_ ),
    .ZN(u_multiplier_pp2_24 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_24_1__18_  (.A(u_multiplier_STAGE2_pp2_23_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_24_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_24_1__19_  (.A1(u_multiplier_pp1_24 [1]),
    .A2(u_multiplier_pp1_24 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_24_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_24_1__20_  (.A(u_multiplier_pp1_24 [1]),
    .B(u_multiplier_pp1_24 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_24_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_24_1__21_  (.A1(u_multiplier_pp1_24 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_24_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_24_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_24_1__22_  (.A(u_multiplier_pp1_24 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_24_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_24_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_24_1__23_  (.A1(u_multiplier_pp1_24 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_24_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_24_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_24_1__24_  (.A(u_multiplier_pp1_24 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_24_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_24_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_24_1__25_  (.A(u_multiplier_STAGE2_pp2_23_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_24_1__16_ ),
    .ZN(u_multiplier_pp2_24 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_24_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_24_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_24_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_24_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_24_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_24_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_24_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_24_1__17_ ),
    .ZN(u_multiplier_pp2_25 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_24_2__18_  (.A(u_multiplier_STAGE2_pp2_23_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_24_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_24_2__19_  (.A1(u_multiplier_pp1_24 [5]),
    .A2(u_multiplier_pp1_24 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_24_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_24_2__20_  (.A(u_multiplier_pp1_24 [5]),
    .B(u_multiplier_pp1_24 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_24_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_24_2__21_  (.A1(u_multiplier_pp1_24 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_24_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_24_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_24_2__22_  (.A(u_multiplier_pp1_24 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_24_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_24_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_24_2__23_  (.A1(u_multiplier_pp1_24 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_24_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_24_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_24_2__24_  (.A(u_multiplier_pp1_24 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_24_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_24_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_24_2__25_  (.A(u_multiplier_STAGE2_pp2_23_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_24_2__16_ ),
    .ZN(u_multiplier_pp2_24 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_24_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_24_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_24_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_24_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_24_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_24_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_24_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_24_2__17_ ),
    .ZN(u_multiplier_pp2_25 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_24_3__18_  (.A(u_multiplier_STAGE2_pp2_23_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_24_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_24_3__19_  (.A1(u_multiplier_pp1_24 [9]),
    .A2(u_multiplier_pp1_24 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_24_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_24_3__20_  (.A(u_multiplier_pp1_24 [9]),
    .B(u_multiplier_pp1_24 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_24_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_24_3__21_  (.A1(u_multiplier_pp1_24 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_24_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_24_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_24_3__22_  (.A(u_multiplier_pp1_24 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_24_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_24_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_24_3__23_  (.A1(u_multiplier_pp1_24 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_24_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_24_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_24_3__24_  (.A(u_multiplier_pp1_24 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_24_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_24_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_24_3__25_  (.A(u_multiplier_STAGE2_pp2_23_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_24_3__16_ ),
    .ZN(u_multiplier_pp2_24 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_24_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_24_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_24_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_24_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_24_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_24_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_24_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_24_3__17_ ),
    .ZN(u_multiplier_pp2_25 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_24_4__18_  (.A(u_multiplier_STAGE2_pp2_23_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_24_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_24_4__19_  (.A1(u_multiplier_pp1_24 [13]),
    .A2(u_multiplier_pp1_24 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_24_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_24_4__20_  (.A(u_multiplier_pp1_24 [13]),
    .B(u_multiplier_pp1_24 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_24_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_24_4__21_  (.A1(u_multiplier_pp1_24 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_24_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_24_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_24_4__22_  (.A(u_multiplier_pp1_24 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_24_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_24_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_24_4__23_  (.A1(u_multiplier_pp1_24 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_24_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_24_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_24_4__24_  (.A(u_multiplier_pp1_24 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_24_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_24_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_24_4__25_  (.A(u_multiplier_STAGE2_pp2_23_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_24_4__16_ ),
    .ZN(u_multiplier_pp2_24 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_24_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_24_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_24_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_24_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_24_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_24_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_24_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_24_4__17_ ),
    .ZN(u_multiplier_pp2_25 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_25_1__18_  (.A(u_multiplier_STAGE2_pp2_24_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_25_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_25_1__19_  (.A1(u_multiplier_pp1_25 [1]),
    .A2(u_multiplier_pp1_25 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_25_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_25_1__20_  (.A(u_multiplier_pp1_25 [1]),
    .B(u_multiplier_pp1_25 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_25_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_25_1__21_  (.A1(u_multiplier_pp1_25 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_25_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_25_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_25_1__22_  (.A(u_multiplier_pp1_25 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_25_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_25_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_25_1__23_  (.A1(u_multiplier_pp1_25 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_25_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_25_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_25_1__24_  (.A(u_multiplier_pp1_25 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_25_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_25_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_25_1__25_  (.A(u_multiplier_STAGE2_pp2_24_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_25_1__16_ ),
    .ZN(u_multiplier_pp2_25 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_25_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_25_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_25_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_25_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_25_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_25_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_25_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_25_1__17_ ),
    .ZN(u_multiplier_pp2_26 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_25_2__18_  (.A(u_multiplier_STAGE2_pp2_24_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_25_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_25_2__19_  (.A1(u_multiplier_pp1_25 [5]),
    .A2(u_multiplier_pp1_25 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_25_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_25_2__20_  (.A(u_multiplier_pp1_25 [5]),
    .B(u_multiplier_pp1_25 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_25_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_25_2__21_  (.A1(u_multiplier_pp1_25 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_25_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_25_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_25_2__22_  (.A(u_multiplier_pp1_25 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_25_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_25_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_25_2__23_  (.A1(u_multiplier_pp1_25 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_25_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_25_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_25_2__24_  (.A(u_multiplier_pp1_25 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_25_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_25_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_25_2__25_  (.A(u_multiplier_STAGE2_pp2_24_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_25_2__16_ ),
    .ZN(u_multiplier_pp2_25 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_25_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_25_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_25_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_25_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_25_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_25_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_25_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_25_2__17_ ),
    .ZN(u_multiplier_pp2_26 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_25_3__18_  (.A(u_multiplier_STAGE2_pp2_24_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_25_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_25_3__19_  (.A1(u_multiplier_pp1_25 [9]),
    .A2(u_multiplier_pp1_25 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_25_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_25_3__20_  (.A(u_multiplier_pp1_25 [9]),
    .B(u_multiplier_pp1_25 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_25_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_25_3__21_  (.A1(u_multiplier_pp1_25 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_25_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_25_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_25_3__22_  (.A(u_multiplier_pp1_25 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_25_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_25_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_25_3__23_  (.A1(u_multiplier_pp1_25 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_25_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_25_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_25_3__24_  (.A(u_multiplier_pp1_25 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_25_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_25_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_25_3__25_  (.A(u_multiplier_STAGE2_pp2_24_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_25_3__16_ ),
    .ZN(u_multiplier_pp2_25 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_25_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_25_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_25_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_25_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_25_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_25_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_25_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_25_3__17_ ),
    .ZN(u_multiplier_pp2_26 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_25_4__18_  (.A(u_multiplier_STAGE2_pp2_24_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_25_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_25_4__19_  (.A1(u_multiplier_pp1_25 [13]),
    .A2(u_multiplier_pp1_25 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_25_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_25_4__20_  (.A(u_multiplier_pp1_25 [13]),
    .B(u_multiplier_pp1_25 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_25_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_25_4__21_  (.A1(u_multiplier_pp1_25 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_25_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_25_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_25_4__22_  (.A(u_multiplier_pp1_25 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_25_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_25_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_25_4__23_  (.A1(u_multiplier_pp1_25 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_25_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_25_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_25_4__24_  (.A(u_multiplier_pp1_25 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_25_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_25_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_25_4__25_  (.A(u_multiplier_STAGE2_pp2_24_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_25_4__16_ ),
    .ZN(u_multiplier_pp2_25 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_25_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_25_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_25_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_25_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_25_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_25_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_25_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_25_4__17_ ),
    .ZN(u_multiplier_pp2_26 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_26_1__18_  (.A(u_multiplier_STAGE2_pp2_25_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_26_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_26_1__19_  (.A1(u_multiplier_pp1_26 [1]),
    .A2(u_multiplier_pp1_26 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_26_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_26_1__20_  (.A(u_multiplier_pp1_26 [1]),
    .B(u_multiplier_pp1_26 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_26_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_26_1__21_  (.A1(u_multiplier_pp1_26 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_26_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_26_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_26_1__22_  (.A(u_multiplier_pp1_26 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_26_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_26_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_26_1__23_  (.A1(u_multiplier_pp1_26 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_26_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_26_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_26_1__24_  (.A(u_multiplier_pp1_26 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_26_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_26_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_26_1__25_  (.A(u_multiplier_STAGE2_pp2_25_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_26_1__16_ ),
    .ZN(u_multiplier_pp2_26 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_26_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_26_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_26_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_26_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_26_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_26_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_26_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_26_1__17_ ),
    .ZN(u_multiplier_pp2_27 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_26_2__18_  (.A(u_multiplier_STAGE2_pp2_25_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_26_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_26_2__19_  (.A1(u_multiplier_pp1_26 [5]),
    .A2(u_multiplier_pp1_26 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_26_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_26_2__20_  (.A(u_multiplier_pp1_26 [5]),
    .B(u_multiplier_pp1_26 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_26_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_26_2__21_  (.A1(u_multiplier_pp1_26 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_26_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_26_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_26_2__22_  (.A(u_multiplier_pp1_26 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_26_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_26_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_26_2__23_  (.A1(u_multiplier_pp1_26 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_26_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_26_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_26_2__24_  (.A(u_multiplier_pp1_26 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_26_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_26_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_26_2__25_  (.A(u_multiplier_STAGE2_pp2_25_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_26_2__16_ ),
    .ZN(u_multiplier_pp2_26 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_26_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_26_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_26_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_26_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_26_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_26_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_26_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_26_2__17_ ),
    .ZN(u_multiplier_pp2_27 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_26_3__18_  (.A(u_multiplier_STAGE2_pp2_25_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_26_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_26_3__19_  (.A1(u_multiplier_pp1_26 [9]),
    .A2(u_multiplier_pp1_26 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_26_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_26_3__20_  (.A(u_multiplier_pp1_26 [9]),
    .B(u_multiplier_pp1_26 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_26_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_26_3__21_  (.A1(u_multiplier_pp1_26 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_26_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_26_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_26_3__22_  (.A(u_multiplier_pp1_26 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_26_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_26_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_26_3__23_  (.A1(u_multiplier_pp1_26 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_26_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_26_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_26_3__24_  (.A(u_multiplier_pp1_26 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_26_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_26_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_26_3__25_  (.A(u_multiplier_STAGE2_pp2_25_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_26_3__16_ ),
    .ZN(u_multiplier_pp2_26 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_26_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_26_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_26_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_26_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_26_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_26_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_26_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_26_3__17_ ),
    .ZN(u_multiplier_pp2_27 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_26_4__18_  (.A(u_multiplier_STAGE2_pp2_25_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_26_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_26_4__19_  (.A1(u_multiplier_pp1_26 [13]),
    .A2(u_multiplier_pp1_26 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_26_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_26_4__20_  (.A(u_multiplier_pp1_26 [13]),
    .B(u_multiplier_pp1_26 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_26_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_26_4__21_  (.A1(u_multiplier_pp1_26 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_26_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_26_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_26_4__22_  (.A(u_multiplier_pp1_26 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_26_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_26_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_26_4__23_  (.A1(u_multiplier_pp1_26 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_26_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_26_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_26_4__24_  (.A(u_multiplier_pp1_26 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_26_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_26_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_26_4__25_  (.A(u_multiplier_STAGE2_pp2_25_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_26_4__16_ ),
    .ZN(u_multiplier_pp2_26 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_26_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_26_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_26_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_26_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_26_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_26_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_26_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_26_4__17_ ),
    .ZN(u_multiplier_pp2_27 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_27_1__18_  (.A(u_multiplier_STAGE2_pp2_26_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_27_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_27_1__19_  (.A1(u_multiplier_pp1_27 [1]),
    .A2(u_multiplier_pp1_27 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_27_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_27_1__20_  (.A(u_multiplier_pp1_27 [1]),
    .B(u_multiplier_pp1_27 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_27_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_27_1__21_  (.A1(u_multiplier_pp1_27 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_27_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_27_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_27_1__22_  (.A(u_multiplier_pp1_27 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_27_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_27_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_27_1__23_  (.A1(u_multiplier_pp1_27 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_27_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_27_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_27_1__24_  (.A(u_multiplier_pp1_27 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_27_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_27_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_27_1__25_  (.A(u_multiplier_STAGE2_pp2_26_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_27_1__16_ ),
    .ZN(u_multiplier_pp2_27 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_27_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_27_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_27_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_27_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_27_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_27_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_27_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_27_1__17_ ),
    .ZN(u_multiplier_pp2_28 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_27_2__18_  (.A(u_multiplier_STAGE2_pp2_26_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_27_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_27_2__19_  (.A1(u_multiplier_pp1_27 [5]),
    .A2(u_multiplier_pp1_27 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_27_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_27_2__20_  (.A(u_multiplier_pp1_27 [5]),
    .B(u_multiplier_pp1_27 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_27_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_27_2__21_  (.A1(u_multiplier_pp1_27 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_27_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_27_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_27_2__22_  (.A(u_multiplier_pp1_27 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_27_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_27_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_27_2__23_  (.A1(u_multiplier_pp1_27 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_27_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_27_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_27_2__24_  (.A(u_multiplier_pp1_27 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_27_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_27_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_27_2__25_  (.A(u_multiplier_STAGE2_pp2_26_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_27_2__16_ ),
    .ZN(u_multiplier_pp2_27 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_27_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_27_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_27_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_27_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_27_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_27_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_27_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_27_2__17_ ),
    .ZN(u_multiplier_pp2_28 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_27_3__18_  (.A(u_multiplier_STAGE2_pp2_26_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_27_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_27_3__19_  (.A1(u_multiplier_pp1_27 [9]),
    .A2(u_multiplier_pp1_27 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_27_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_27_3__20_  (.A(u_multiplier_pp1_27 [9]),
    .B(u_multiplier_pp1_27 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_27_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_27_3__21_  (.A1(u_multiplier_pp1_27 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_27_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_27_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_27_3__22_  (.A(u_multiplier_pp1_27 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_27_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_27_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_27_3__23_  (.A1(u_multiplier_pp1_27 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_27_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_27_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_27_3__24_  (.A(u_multiplier_pp1_27 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_27_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_27_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_27_3__25_  (.A(u_multiplier_STAGE2_pp2_26_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_27_3__16_ ),
    .ZN(u_multiplier_pp2_27 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_27_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_27_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_27_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_27_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_27_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_27_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_27_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_27_3__17_ ),
    .ZN(u_multiplier_pp2_28 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_27_4__18_  (.A(u_multiplier_STAGE2_pp2_26_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_27_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_27_4__19_  (.A1(u_multiplier_pp1_27 [13]),
    .A2(u_multiplier_pp1_27 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_27_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_27_4__20_  (.A(u_multiplier_pp1_27 [13]),
    .B(u_multiplier_pp1_27 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_27_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_27_4__21_  (.A1(u_multiplier_pp1_27 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_27_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_27_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_27_4__22_  (.A(u_multiplier_pp1_27 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_27_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_27_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_27_4__23_  (.A1(u_multiplier_pp1_27 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_27_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_27_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_27_4__24_  (.A(u_multiplier_pp1_27 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_27_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_27_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_27_4__25_  (.A(u_multiplier_STAGE2_pp2_26_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_27_4__16_ ),
    .ZN(u_multiplier_pp2_27 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_27_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_27_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_27_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_27_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_27_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_27_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_27_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_27_4__17_ ),
    .ZN(u_multiplier_pp2_28 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_28_1__18_  (.A(u_multiplier_STAGE2_pp2_27_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_28_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_28_1__19_  (.A1(u_multiplier_pp1_28 [1]),
    .A2(u_multiplier_pp1_28 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_28_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_28_1__20_  (.A(u_multiplier_pp1_28 [1]),
    .B(u_multiplier_pp1_28 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_28_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_28_1__21_  (.A1(u_multiplier_pp1_28 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_28_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_28_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_28_1__22_  (.A(u_multiplier_pp1_28 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_28_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_28_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_28_1__23_  (.A1(u_multiplier_pp1_28 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_28_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_28_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_28_1__24_  (.A(u_multiplier_pp1_28 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_28_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_28_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_28_1__25_  (.A(u_multiplier_STAGE2_pp2_27_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_28_1__16_ ),
    .ZN(u_multiplier_pp2_28 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_28_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_28_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_28_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_28_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_28_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_28_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_28_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_28_1__17_ ),
    .ZN(u_multiplier_pp2_29 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_28_2__18_  (.A(u_multiplier_STAGE2_pp2_27_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_28_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_28_2__19_  (.A1(u_multiplier_pp1_28 [5]),
    .A2(u_multiplier_pp1_28 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_28_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_28_2__20_  (.A(u_multiplier_pp1_28 [5]),
    .B(u_multiplier_pp1_28 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_28_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_28_2__21_  (.A1(u_multiplier_pp1_28 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_28_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_28_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_28_2__22_  (.A(u_multiplier_pp1_28 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_28_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_28_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_28_2__23_  (.A1(u_multiplier_pp1_28 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_28_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_28_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_28_2__24_  (.A(u_multiplier_pp1_28 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_28_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_28_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_28_2__25_  (.A(u_multiplier_STAGE2_pp2_27_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_28_2__16_ ),
    .ZN(u_multiplier_pp2_28 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_28_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_28_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_28_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_28_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_28_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_28_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_28_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_28_2__17_ ),
    .ZN(u_multiplier_pp2_29 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_28_3__18_  (.A(u_multiplier_STAGE2_pp2_27_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_28_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_28_3__19_  (.A1(u_multiplier_pp1_28 [9]),
    .A2(u_multiplier_pp1_28 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_28_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_28_3__20_  (.A(u_multiplier_pp1_28 [9]),
    .B(u_multiplier_pp1_28 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_28_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_28_3__21_  (.A1(u_multiplier_pp1_28 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_28_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_28_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_28_3__22_  (.A(u_multiplier_pp1_28 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_28_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_28_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_28_3__23_  (.A1(u_multiplier_pp1_28 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_28_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_28_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_28_3__24_  (.A(u_multiplier_pp1_28 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_28_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_28_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_28_3__25_  (.A(u_multiplier_STAGE2_pp2_27_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_28_3__16_ ),
    .ZN(u_multiplier_pp2_28 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_28_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_28_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_28_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_28_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_28_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_28_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_28_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_28_3__17_ ),
    .ZN(u_multiplier_pp2_29 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_28_4__18_  (.A(u_multiplier_STAGE2_pp2_27_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_28_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_28_4__19_  (.A1(u_multiplier_pp1_28 [13]),
    .A2(u_multiplier_pp1_28 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_28_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_28_4__20_  (.A(u_multiplier_pp1_28 [13]),
    .B(u_multiplier_pp1_28 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_28_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_28_4__21_  (.A1(u_multiplier_pp1_28 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_28_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_28_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_28_4__22_  (.A(u_multiplier_pp1_28 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_28_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_28_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_28_4__23_  (.A1(u_multiplier_pp1_28 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_28_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_28_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_28_4__24_  (.A(u_multiplier_pp1_28 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_28_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_28_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_28_4__25_  (.A(u_multiplier_STAGE2_pp2_27_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_28_4__16_ ),
    .ZN(u_multiplier_pp2_28 [0]));
 NAND2_X2 u_multiplier_STAGE2_E_4_2_pp2_28_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_28_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_28_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_28_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_28_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_28_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_28_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_28_4__17_ ),
    .ZN(u_multiplier_pp2_29 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_29_1__18_  (.A(u_multiplier_STAGE2_pp2_28_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_29_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_29_1__19_  (.A1(u_multiplier_pp1_29 [1]),
    .A2(u_multiplier_pp1_29 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_29_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_29_1__20_  (.A(u_multiplier_pp1_29 [1]),
    .B(u_multiplier_pp1_29 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_29_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_29_1__21_  (.A1(u_multiplier_pp1_29 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_29_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_29_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_29_1__22_  (.A(u_multiplier_pp1_29 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_29_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_29_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_29_1__23_  (.A1(u_multiplier_pp1_29 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_29_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_29_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_29_1__24_  (.A(u_multiplier_pp1_29 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_29_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_29_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_29_1__25_  (.A(u_multiplier_STAGE2_pp2_28_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_29_1__16_ ),
    .ZN(u_multiplier_pp2_29 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_29_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_29_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_29_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_29_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_29_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_29_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_29_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_29_1__17_ ),
    .ZN(u_multiplier_pp2_30 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_29_2__18_  (.A(u_multiplier_STAGE2_pp2_28_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_29_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_29_2__19_  (.A1(u_multiplier_pp1_29 [5]),
    .A2(u_multiplier_pp1_29 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_29_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_29_2__20_  (.A(u_multiplier_pp1_29 [5]),
    .B(u_multiplier_pp1_29 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_29_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_29_2__21_  (.A1(u_multiplier_pp1_29 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_29_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_29_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_29_2__22_  (.A(u_multiplier_pp1_29 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_29_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_29_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_29_2__23_  (.A1(u_multiplier_pp1_29 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_29_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_29_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_29_2__24_  (.A(u_multiplier_pp1_29 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_29_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_29_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_29_2__25_  (.A(u_multiplier_STAGE2_pp2_28_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_29_2__16_ ),
    .ZN(u_multiplier_pp2_29 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_29_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_29_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_29_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_29_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_29_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_29_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_29_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_29_2__17_ ),
    .ZN(u_multiplier_pp2_30 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_29_3__18_  (.A(u_multiplier_STAGE2_pp2_28_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_29_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_29_3__19_  (.A1(u_multiplier_pp1_29 [9]),
    .A2(u_multiplier_pp1_29 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_29_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_29_3__20_  (.A(u_multiplier_pp1_29 [9]),
    .B(u_multiplier_pp1_29 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_29_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_29_3__21_  (.A1(u_multiplier_pp1_29 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_29_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_29_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_29_3__22_  (.A(u_multiplier_pp1_29 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_29_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_29_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_29_3__23_  (.A1(u_multiplier_pp1_29 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_29_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_29_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_29_3__24_  (.A(u_multiplier_pp1_29 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_29_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_29_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_29_3__25_  (.A(u_multiplier_STAGE2_pp2_28_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_29_3__16_ ),
    .ZN(u_multiplier_pp2_29 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_29_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_29_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_29_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_29_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_29_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_29_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_29_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_29_3__17_ ),
    .ZN(u_multiplier_pp2_30 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_29_4__18_  (.A(u_multiplier_STAGE2_pp2_28_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_29_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_29_4__19_  (.A1(u_multiplier_pp1_29 [13]),
    .A2(u_multiplier_pp1_29 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_29_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_29_4__20_  (.A(u_multiplier_pp1_29 [13]),
    .B(u_multiplier_pp1_29 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_29_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_29_4__21_  (.A1(u_multiplier_pp1_29 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_29_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_29_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_29_4__22_  (.A(u_multiplier_pp1_29 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_29_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_29_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_29_4__23_  (.A1(u_multiplier_pp1_29 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_29_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_29_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_29_4__24_  (.A(u_multiplier_pp1_29 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_29_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_29_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_29_4__25_  (.A(u_multiplier_STAGE2_pp2_28_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_29_4__16_ ),
    .ZN(u_multiplier_pp2_29 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_29_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_29_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_29_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_29_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_29_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_29_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_29_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_29_4__17_ ),
    .ZN(u_multiplier_pp2_30 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_30_1__18_  (.A(u_multiplier_STAGE2_pp2_29_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_30_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_30_1__19_  (.A1(u_multiplier_pp1_30 [1]),
    .A2(u_multiplier_pp1_30 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_30_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_30_1__20_  (.A(u_multiplier_pp1_30 [1]),
    .B(u_multiplier_pp1_30 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_30_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_30_1__21_  (.A1(u_multiplier_pp1_30 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_30_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_30_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_30_1__22_  (.A(u_multiplier_pp1_30 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_30_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_30_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_30_1__23_  (.A1(u_multiplier_pp1_30 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_30_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_30_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_30_1__24_  (.A(u_multiplier_pp1_30 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_30_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_30_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_30_1__25_  (.A(u_multiplier_STAGE2_pp2_29_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_30_1__16_ ),
    .ZN(u_multiplier_pp2_30 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_30_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_30_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_30_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_30_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE2_E_4_2_pp2_30_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_30_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_30_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_30_1__17_ ),
    .ZN(u_multiplier_pp2_31 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_30_2__18_  (.A(u_multiplier_STAGE2_pp2_29_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_30_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_30_2__19_  (.A1(u_multiplier_pp1_30 [5]),
    .A2(u_multiplier_pp1_30 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_30_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_30_2__20_  (.A(u_multiplier_pp1_30 [5]),
    .B(u_multiplier_pp1_30 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_30_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_30_2__21_  (.A1(u_multiplier_pp1_30 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_30_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_30_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_30_2__22_  (.A(u_multiplier_pp1_30 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_30_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_30_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_30_2__23_  (.A1(u_multiplier_pp1_30 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_30_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_30_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_30_2__24_  (.A(u_multiplier_pp1_30 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_30_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_30_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_30_2__25_  (.A(u_multiplier_STAGE2_pp2_29_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_30_2__16_ ),
    .ZN(u_multiplier_pp2_30 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_30_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_30_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_30_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_30_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_30_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_30_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_30_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_30_2__17_ ),
    .ZN(u_multiplier_pp2_31 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_30_3__18_  (.A(u_multiplier_STAGE2_pp2_29_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_30_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_30_3__19_  (.A1(u_multiplier_pp1_30 [9]),
    .A2(u_multiplier_pp1_30 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_30_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_30_3__20_  (.A(u_multiplier_pp1_30 [9]),
    .B(u_multiplier_pp1_30 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_30_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_30_3__21_  (.A1(u_multiplier_pp1_30 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_30_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_30_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_30_3__22_  (.A(u_multiplier_pp1_30 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_30_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_30_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_30_3__23_  (.A1(u_multiplier_pp1_30 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_30_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_30_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_30_3__24_  (.A(u_multiplier_pp1_30 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_30_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_30_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_30_3__25_  (.A(u_multiplier_STAGE2_pp2_29_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_30_3__16_ ),
    .ZN(u_multiplier_pp2_30 [1]));
 NAND2_X2 u_multiplier_STAGE2_E_4_2_pp2_30_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_30_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_30_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_30_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_30_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_30_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_30_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_30_3__17_ ),
    .ZN(u_multiplier_pp2_31 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_30_4__18_  (.A(u_multiplier_STAGE2_pp2_29_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_30_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_30_4__19_  (.A1(u_multiplier_pp1_30 [13]),
    .A2(u_multiplier_pp1_30 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_30_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_30_4__20_  (.A(u_multiplier_pp1_30 [13]),
    .B(u_multiplier_pp1_30 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_30_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_30_4__21_  (.A1(u_multiplier_pp1_30 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_30_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_30_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_30_4__22_  (.A(u_multiplier_pp1_30 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_30_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_30_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_30_4__23_  (.A1(u_multiplier_pp1_30 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_30_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_30_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_30_4__24_  (.A(u_multiplier_pp1_30 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_30_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_30_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_30_4__25_  (.A(u_multiplier_STAGE2_pp2_29_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_30_4__16_ ),
    .ZN(u_multiplier_pp2_30 [0]));
 NAND2_X2 u_multiplier_STAGE2_E_4_2_pp2_30_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_30_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_30_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_30_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_30_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_30_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_30_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_30_4__17_ ),
    .ZN(u_multiplier_pp2_31 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_31_1__18_  (.A(u_multiplier_STAGE2_pp2_30_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_31_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_31_1__19_  (.A1(u_multiplier_pp1_31 [1]),
    .A2(u_multiplier_pp1_31 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_31_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_31_1__20_  (.A(u_multiplier_pp1_31 [1]),
    .B(u_multiplier_pp1_31 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_31_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_31_1__21_  (.A1(u_multiplier_pp1_31 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_31_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_31_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_31_1__22_  (.A(u_multiplier_pp1_31 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_31_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_31_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_31_1__23_  (.A1(u_multiplier_pp1_31 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_31_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_31_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_31_1__24_  (.A(u_multiplier_pp1_31 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_31_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_31_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_31_1__25_  (.A(u_multiplier_STAGE2_pp2_30_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_31_1__16_ ),
    .ZN(u_multiplier_pp2_31 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_31_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_31_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_31_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_31_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE2_E_4_2_pp2_31_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_31_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_31_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_31_1__17_ ),
    .ZN(u_multiplier_pp2_32 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_31_2__18_  (.A(u_multiplier_STAGE2_pp2_30_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_31_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_31_2__19_  (.A1(u_multiplier_pp1_31 [5]),
    .A2(u_multiplier_pp1_31 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_31_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_31_2__20_  (.A(u_multiplier_pp1_31 [5]),
    .B(u_multiplier_pp1_31 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_31_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_31_2__21_  (.A1(u_multiplier_pp1_31 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_31_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_31_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_31_2__22_  (.A(u_multiplier_pp1_31 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_31_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_31_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_31_2__23_  (.A1(u_multiplier_pp1_31 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_31_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_31_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_31_2__24_  (.A(u_multiplier_pp1_31 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_31_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_31_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_31_2__25_  (.A(u_multiplier_STAGE2_pp2_30_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_31_2__16_ ),
    .ZN(u_multiplier_pp2_31 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_31_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_31_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_31_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_31_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_31_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_31_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_31_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_31_2__17_ ),
    .ZN(u_multiplier_pp2_32 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_31_3__18_  (.A(u_multiplier_STAGE2_pp2_30_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_31_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_31_3__19_  (.A1(u_multiplier_pp1_31 [9]),
    .A2(u_multiplier_pp1_31 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_31_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_31_3__20_  (.A(u_multiplier_pp1_31 [9]),
    .B(u_multiplier_pp1_31 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_31_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_31_3__21_  (.A1(u_multiplier_pp1_31 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_31_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_31_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_31_3__22_  (.A(u_multiplier_pp1_31 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_31_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_31_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_31_3__23_  (.A1(u_multiplier_pp1_31 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_31_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_31_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_31_3__24_  (.A(u_multiplier_pp1_31 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_31_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_31_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_31_3__25_  (.A(u_multiplier_STAGE2_pp2_30_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_31_3__16_ ),
    .ZN(u_multiplier_pp2_31 [1]));
 NAND2_X2 u_multiplier_STAGE2_E_4_2_pp2_31_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_31_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_31_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_31_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_31_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_31_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_31_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_31_3__17_ ),
    .ZN(u_multiplier_pp2_32 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_31_4__18_  (.A(u_multiplier_STAGE2_pp2_30_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_31_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_31_4__19_  (.A1(u_multiplier_pp1_31 [13]),
    .A2(u_multiplier_pp1_31 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_31_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_31_4__20_  (.A(u_multiplier_pp1_31 [13]),
    .B(u_multiplier_pp1_31 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_31_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_31_4__21_  (.A1(u_multiplier_pp1_31 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_31_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_31_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_31_4__22_  (.A(u_multiplier_pp1_31 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_31_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_31_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_31_4__23_  (.A1(u_multiplier_pp1_31 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_31_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_31_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_31_4__24_  (.A(u_multiplier_pp1_31 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_31_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_31_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_31_4__25_  (.A(u_multiplier_STAGE2_pp2_30_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_31_4__16_ ),
    .ZN(u_multiplier_pp2_31 [0]));
 NAND2_X2 u_multiplier_STAGE2_E_4_2_pp2_31_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_31_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_31_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_31_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_31_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_31_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_31_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_31_4__17_ ),
    .ZN(u_multiplier_pp2_32 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_32_1__18_  (.A(u_multiplier_STAGE2_pp2_31_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_1__19_  (.A1(u_multiplier_pp1_32 [1]),
    .A2(u_multiplier_pp1_32 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_1__20_  (.A(u_multiplier_pp1_32 [1]),
    .B(u_multiplier_pp1_32 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_32_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_1__21_  (.A1(u_multiplier_pp1_32 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_32_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_1__22_  (.A(u_multiplier_pp1_32 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_32_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_32_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_1__23_  (.A1(u_multiplier_pp1_32 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_32_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_1__24_  (.A(u_multiplier_pp1_32 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_32_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_1__25_  (.A(u_multiplier_STAGE2_pp2_31_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_32_1__16_ ),
    .ZN(u_multiplier_pp2_32 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_32_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_32_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_32_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_32_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_32_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_32_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_32_1__17_ ),
    .ZN(u_multiplier_pp2_33 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_32_2__18_  (.A(u_multiplier_STAGE2_pp2_31_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_2__19_  (.A1(u_multiplier_pp1_32 [5]),
    .A2(u_multiplier_pp1_32 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_2__20_  (.A(u_multiplier_pp1_32 [5]),
    .B(u_multiplier_pp1_32 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_32_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_2__21_  (.A1(u_multiplier_pp1_32 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_32_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_2__22_  (.A(u_multiplier_pp1_32 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_32_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_32_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_2__23_  (.A1(u_multiplier_pp1_32 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_32_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_2__24_  (.A(u_multiplier_pp1_32 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_32_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_2__25_  (.A(u_multiplier_STAGE2_pp2_31_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_32_2__16_ ),
    .ZN(u_multiplier_pp2_32 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_32_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_32_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_32_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_32_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_32_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_32_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_32_2__17_ ),
    .ZN(u_multiplier_pp2_33 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_32_3__18_  (.A(u_multiplier_STAGE2_pp2_31_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_3__19_  (.A1(u_multiplier_pp1_32 [9]),
    .A2(u_multiplier_pp1_32 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_3__20_  (.A(u_multiplier_pp1_32 [9]),
    .B(u_multiplier_pp1_32 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_32_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_3__21_  (.A1(u_multiplier_pp1_32 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_32_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_3__22_  (.A(u_multiplier_pp1_32 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_32_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_32_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_3__23_  (.A1(u_multiplier_pp1_32 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_32_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_3__24_  (.A(u_multiplier_pp1_32 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_32_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_3__25_  (.A(u_multiplier_STAGE2_pp2_31_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_32_3__16_ ),
    .ZN(u_multiplier_pp2_32 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_32_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_32_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_32_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_32_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_32_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_32_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_32_3__17_ ),
    .ZN(u_multiplier_pp2_33 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_32_4__18_  (.A(u_multiplier_STAGE2_pp2_31_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_4__19_  (.A1(u_multiplier_pp1_32 [13]),
    .A2(u_multiplier_pp1_32 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_4__20_  (.A(u_multiplier_pp1_32 [13]),
    .B(u_multiplier_pp1_32 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_32_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_4__21_  (.A1(u_multiplier_pp1_32 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_32_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_4__22_  (.A(u_multiplier_pp1_32 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_32_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_32_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_4__23_  (.A1(u_multiplier_pp1_32 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_32_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_4__24_  (.A(u_multiplier_pp1_32 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_32_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_4__25_  (.A(u_multiplier_STAGE2_pp2_31_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_32_4__16_ ),
    .ZN(u_multiplier_pp2_32 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_32_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_32_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_32_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_32_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_32_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_32_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_32_4__17_ ),
    .ZN(u_multiplier_pp2_33 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_33_1__18_  (.A(u_multiplier_STAGE2_pp2_32_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_1__19_  (.A1(u_multiplier_pp1_33 [1]),
    .A2(u_multiplier_pp1_33 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_1__20_  (.A(u_multiplier_pp1_33 [1]),
    .B(u_multiplier_pp1_33 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_33_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_1__21_  (.A1(u_multiplier_pp1_33 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_33_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_1__22_  (.A(u_multiplier_pp1_33 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_33_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_33_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_1__23_  (.A1(u_multiplier_pp1_33 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_33_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_1__24_  (.A(u_multiplier_pp1_33 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_33_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_1__25_  (.A(u_multiplier_STAGE2_pp2_32_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_33_1__16_ ),
    .ZN(u_multiplier_pp2_33 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_33_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_33_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_33_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_33_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_33_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_33_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_33_1__17_ ),
    .ZN(u_multiplier_pp2_34 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_33_2__18_  (.A(u_multiplier_STAGE2_pp2_32_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_2__19_  (.A1(u_multiplier_pp1_33 [5]),
    .A2(u_multiplier_pp1_33 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_2__20_  (.A(u_multiplier_pp1_33 [5]),
    .B(u_multiplier_pp1_33 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_33_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_2__21_  (.A1(u_multiplier_pp1_33 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_33_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_2__22_  (.A(u_multiplier_pp1_33 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_33_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_33_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_2__23_  (.A1(u_multiplier_pp1_33 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_33_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_2__24_  (.A(u_multiplier_pp1_33 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_33_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_2__25_  (.A(u_multiplier_STAGE2_pp2_32_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_33_2__16_ ),
    .ZN(u_multiplier_pp2_33 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_33_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_33_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_33_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_33_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_33_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_33_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_33_2__17_ ),
    .ZN(u_multiplier_pp2_34 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_33_3__18_  (.A(u_multiplier_STAGE2_pp2_32_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_3__19_  (.A1(u_multiplier_pp1_33 [9]),
    .A2(u_multiplier_pp1_33 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_3__20_  (.A(u_multiplier_pp1_33 [9]),
    .B(u_multiplier_pp1_33 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_33_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_3__21_  (.A1(u_multiplier_pp1_33 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_33_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_3__22_  (.A(u_multiplier_pp1_33 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_33_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_33_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_3__23_  (.A1(u_multiplier_pp1_33 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_33_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_3__24_  (.A(u_multiplier_pp1_33 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_33_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_3__25_  (.A(u_multiplier_STAGE2_pp2_32_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_33_3__16_ ),
    .ZN(u_multiplier_pp2_33 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_33_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_33_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_33_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_33_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_33_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_33_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_33_3__17_ ),
    .ZN(u_multiplier_pp2_34 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_33_4__18_  (.A(u_multiplier_STAGE2_pp2_32_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_4__19_  (.A1(u_multiplier_pp1_33 [13]),
    .A2(u_multiplier_pp1_33 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_4__20_  (.A(u_multiplier_pp1_33 [13]),
    .B(u_multiplier_pp1_33 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_33_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_4__21_  (.A1(u_multiplier_pp1_33 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_33_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_4__22_  (.A(u_multiplier_pp1_33 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_33_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_33_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_4__23_  (.A1(u_multiplier_pp1_33 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_33_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_4__24_  (.A(u_multiplier_pp1_33 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_33_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_4__25_  (.A(u_multiplier_STAGE2_pp2_32_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_33_4__16_ ),
    .ZN(u_multiplier_pp2_33 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_33_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_33_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_33_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_33_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_33_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_33_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_33_4__17_ ),
    .ZN(u_multiplier_pp2_34 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_34_1__18_  (.A(u_multiplier_STAGE2_pp2_33_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_1__19_  (.A1(u_multiplier_pp1_34 [1]),
    .A2(u_multiplier_pp1_34 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_1__20_  (.A(u_multiplier_pp1_34 [1]),
    .B(u_multiplier_pp1_34 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_34_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_1__21_  (.A1(u_multiplier_pp1_34 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_34_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_1__22_  (.A(u_multiplier_pp1_34 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_34_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_34_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_1__23_  (.A1(u_multiplier_pp1_34 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_34_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_1__24_  (.A(u_multiplier_pp1_34 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_34_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_1__25_  (.A(u_multiplier_STAGE2_pp2_33_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_34_1__16_ ),
    .ZN(u_multiplier_pp2_34 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_34_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_34_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_34_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_34_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_34_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_34_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_34_1__17_ ),
    .ZN(u_multiplier_pp2_35 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_34_2__18_  (.A(u_multiplier_STAGE2_pp2_33_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_2__19_  (.A1(u_multiplier_pp1_34 [5]),
    .A2(u_multiplier_pp1_34 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_2__20_  (.A(u_multiplier_pp1_34 [5]),
    .B(u_multiplier_pp1_34 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_34_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_2__21_  (.A1(u_multiplier_pp1_34 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_34_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_2__22_  (.A(u_multiplier_pp1_34 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_34_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_34_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_2__23_  (.A1(u_multiplier_pp1_34 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_34_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_2__24_  (.A(u_multiplier_pp1_34 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_34_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_2__25_  (.A(u_multiplier_STAGE2_pp2_33_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_34_2__16_ ),
    .ZN(u_multiplier_pp2_34 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_34_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_34_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_34_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_34_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_34_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_34_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_34_2__17_ ),
    .ZN(u_multiplier_pp2_35 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_34_3__18_  (.A(u_multiplier_STAGE2_pp2_33_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_3__19_  (.A1(u_multiplier_pp1_34 [9]),
    .A2(u_multiplier_pp1_34 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_3__20_  (.A(u_multiplier_pp1_34 [9]),
    .B(u_multiplier_pp1_34 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_34_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_3__21_  (.A1(u_multiplier_pp1_34 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_34_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_3__22_  (.A(u_multiplier_pp1_34 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_34_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_34_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_3__23_  (.A1(u_multiplier_pp1_34 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_34_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_3__24_  (.A(u_multiplier_pp1_34 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_34_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_3__25_  (.A(u_multiplier_STAGE2_pp2_33_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_34_3__16_ ),
    .ZN(u_multiplier_pp2_34 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_34_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_34_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_34_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_34_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_34_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_34_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_34_3__17_ ),
    .ZN(u_multiplier_pp2_35 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_34_4__18_  (.A(u_multiplier_STAGE2_pp2_33_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_4__19_  (.A1(u_multiplier_pp1_34 [13]),
    .A2(u_multiplier_pp1_34 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_4__20_  (.A(u_multiplier_pp1_34 [13]),
    .B(u_multiplier_pp1_34 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_34_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_4__21_  (.A1(u_multiplier_pp1_34 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_34_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_4__22_  (.A(u_multiplier_pp1_34 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_34_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_34_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_4__23_  (.A1(u_multiplier_pp1_34 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_34_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_4__24_  (.A(u_multiplier_pp1_34 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_34_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_4__25_  (.A(u_multiplier_STAGE2_pp2_33_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_34_4__16_ ),
    .ZN(u_multiplier_pp2_34 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_34_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_34_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_34_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_34_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_34_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_34_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_34_4__17_ ),
    .ZN(u_multiplier_pp2_35 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_35_1__18_  (.A(u_multiplier_STAGE2_pp2_34_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_1__19_  (.A1(u_multiplier_pp1_35 [1]),
    .A2(u_multiplier_pp1_35 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_1__20_  (.A(u_multiplier_pp1_35 [1]),
    .B(u_multiplier_pp1_35 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_35_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_1__21_  (.A1(u_multiplier_pp1_35 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_35_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_1__22_  (.A(u_multiplier_pp1_35 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_35_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_35_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_1__23_  (.A1(u_multiplier_pp1_35 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_35_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_1__24_  (.A(u_multiplier_pp1_35 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_35_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_1__25_  (.A(u_multiplier_STAGE2_pp2_34_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_35_1__16_ ),
    .ZN(u_multiplier_pp2_35 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_35_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_35_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_35_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_35_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_35_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_35_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_35_1__17_ ),
    .ZN(u_multiplier_pp2_36 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_35_2__18_  (.A(u_multiplier_STAGE2_pp2_34_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_2__19_  (.A1(u_multiplier_pp1_35 [5]),
    .A2(u_multiplier_pp1_35 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_2__20_  (.A(u_multiplier_pp1_35 [5]),
    .B(u_multiplier_pp1_35 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_35_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_2__21_  (.A1(u_multiplier_pp1_35 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_35_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_2__22_  (.A(u_multiplier_pp1_35 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_35_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_35_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_2__23_  (.A1(u_multiplier_pp1_35 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_35_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_2__24_  (.A(u_multiplier_pp1_35 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_35_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_2__25_  (.A(u_multiplier_STAGE2_pp2_34_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_35_2__16_ ),
    .ZN(u_multiplier_pp2_35 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_35_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_35_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_35_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_35_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_35_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_35_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_35_2__17_ ),
    .ZN(u_multiplier_pp2_36 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_35_3__18_  (.A(u_multiplier_STAGE2_pp2_34_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_3__19_  (.A1(u_multiplier_pp1_35 [9]),
    .A2(u_multiplier_pp1_35 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_3__20_  (.A(u_multiplier_pp1_35 [9]),
    .B(u_multiplier_pp1_35 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_35_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_3__21_  (.A1(u_multiplier_pp1_35 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_35_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_3__22_  (.A(u_multiplier_pp1_35 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_35_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_35_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_3__23_  (.A1(u_multiplier_pp1_35 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_35_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_3__24_  (.A(u_multiplier_pp1_35 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_35_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_3__25_  (.A(u_multiplier_STAGE2_pp2_34_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_35_3__16_ ),
    .ZN(u_multiplier_pp2_35 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_35_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_35_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_35_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_35_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_35_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_35_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_35_3__17_ ),
    .ZN(u_multiplier_pp2_36 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_35_4__18_  (.A(u_multiplier_STAGE2_pp2_34_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_4__19_  (.A1(u_multiplier_pp1_35 [13]),
    .A2(u_multiplier_pp1_35 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_4__20_  (.A(u_multiplier_pp1_35 [13]),
    .B(u_multiplier_pp1_35 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_35_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_4__21_  (.A1(u_multiplier_pp1_35 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_35_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_4__22_  (.A(u_multiplier_pp1_35 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_35_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_35_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_4__23_  (.A1(u_multiplier_pp1_35 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_35_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_4__24_  (.A(u_multiplier_pp1_35 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_35_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_4__25_  (.A(u_multiplier_STAGE2_pp2_34_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_35_4__16_ ),
    .ZN(u_multiplier_pp2_35 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_35_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_35_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_35_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_35_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_35_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_35_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_35_4__17_ ),
    .ZN(u_multiplier_pp2_36 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_36_1__18_  (.A(u_multiplier_STAGE2_pp2_35_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_1__19_  (.A1(u_multiplier_pp1_36 [1]),
    .A2(u_multiplier_pp1_36 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_1__20_  (.A(u_multiplier_pp1_36 [1]),
    .B(u_multiplier_pp1_36 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_36_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_1__21_  (.A1(u_multiplier_pp1_36 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_36_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_1__22_  (.A(u_multiplier_pp1_36 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_36_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_36_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_1__23_  (.A1(u_multiplier_pp1_36 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_36_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_1__24_  (.A(u_multiplier_pp1_36 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_36_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_1__25_  (.A(u_multiplier_STAGE2_pp2_35_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_36_1__16_ ),
    .ZN(u_multiplier_pp2_36 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_36_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_36_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_36_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_36_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_36_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_36_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_36_1__17_ ),
    .ZN(u_multiplier_pp2_37 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_36_2__18_  (.A(u_multiplier_STAGE2_pp2_35_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_2__19_  (.A1(u_multiplier_pp1_36 [5]),
    .A2(u_multiplier_pp1_36 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_2__20_  (.A(u_multiplier_pp1_36 [5]),
    .B(u_multiplier_pp1_36 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_36_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_2__21_  (.A1(u_multiplier_pp1_36 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_36_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_2__22_  (.A(u_multiplier_pp1_36 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_36_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_36_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_2__23_  (.A1(u_multiplier_pp1_36 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_36_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_2__24_  (.A(u_multiplier_pp1_36 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_36_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_2__25_  (.A(u_multiplier_STAGE2_pp2_35_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_36_2__16_ ),
    .ZN(u_multiplier_pp2_36 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_36_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_36_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_36_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_36_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_36_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_36_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_36_2__17_ ),
    .ZN(u_multiplier_pp2_37 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_36_3__18_  (.A(u_multiplier_STAGE2_pp2_35_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_3__19_  (.A1(u_multiplier_pp1_36 [9]),
    .A2(u_multiplier_pp1_36 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_3__20_  (.A(u_multiplier_pp1_36 [9]),
    .B(u_multiplier_pp1_36 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_36_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_3__21_  (.A1(u_multiplier_pp1_36 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_36_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_3__22_  (.A(u_multiplier_pp1_36 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_36_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_36_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_3__23_  (.A1(u_multiplier_pp1_36 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_36_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_3__24_  (.A(u_multiplier_pp1_36 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_36_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_3__25_  (.A(u_multiplier_STAGE2_pp2_35_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_36_3__16_ ),
    .ZN(u_multiplier_pp2_36 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_36_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_36_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_36_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_36_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_36_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_36_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_36_3__17_ ),
    .ZN(u_multiplier_pp2_37 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_36_4__18_  (.A(u_multiplier_STAGE2_pp2_35_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_4__19_  (.A1(u_multiplier_pp1_36 [13]),
    .A2(u_multiplier_pp1_36 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_4__20_  (.A(u_multiplier_pp1_36 [13]),
    .B(u_multiplier_pp1_36 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_36_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_4__21_  (.A1(u_multiplier_pp1_36 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_36_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_4__22_  (.A(u_multiplier_pp1_36 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_36_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_36_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_4__23_  (.A1(u_multiplier_pp1_36 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_36_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_4__24_  (.A(u_multiplier_pp1_36 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_36_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_4__25_  (.A(u_multiplier_STAGE2_pp2_35_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_36_4__16_ ),
    .ZN(u_multiplier_pp2_36 [0]));
 NAND2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_36_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_36_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_36_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_36_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_36_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_36_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_36_4__17_ ),
    .ZN(u_multiplier_pp2_37 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_37_1__18_  (.A(u_multiplier_STAGE2_pp2_36_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_1__19_  (.A1(u_multiplier_pp1_37 [1]),
    .A2(u_multiplier_pp1_37 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_1__20_  (.A(u_multiplier_pp1_37 [1]),
    .B(u_multiplier_pp1_37 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_37_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_1__21_  (.A1(u_multiplier_pp1_37 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_37_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_1__22_  (.A(u_multiplier_pp1_37 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_37_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_37_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_1__23_  (.A1(u_multiplier_pp1_37 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_37_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_1__24_  (.A(u_multiplier_pp1_37 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_37_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_1__25_  (.A(u_multiplier_STAGE2_pp2_36_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_37_1__16_ ),
    .ZN(u_multiplier_pp2_37 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_37_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_37_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_37_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_37_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_37_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_37_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_37_1__17_ ),
    .ZN(u_multiplier_pp2_38 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_37_2__18_  (.A(u_multiplier_STAGE2_pp2_36_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_2__19_  (.A1(u_multiplier_pp1_37 [5]),
    .A2(u_multiplier_pp1_37 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_2__20_  (.A(u_multiplier_pp1_37 [5]),
    .B(u_multiplier_pp1_37 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_37_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_2__21_  (.A1(u_multiplier_pp1_37 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_37_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_2__22_  (.A(u_multiplier_pp1_37 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_37_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_37_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_2__23_  (.A1(u_multiplier_pp1_37 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_37_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_2__24_  (.A(u_multiplier_pp1_37 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_37_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_2__25_  (.A(u_multiplier_STAGE2_pp2_36_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_37_2__16_ ),
    .ZN(u_multiplier_pp2_37 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_37_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_37_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_37_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_37_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_37_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_37_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_37_2__17_ ),
    .ZN(u_multiplier_pp2_38 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_37_3__18_  (.A(u_multiplier_STAGE2_pp2_36_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_3__19_  (.A1(u_multiplier_pp1_37 [9]),
    .A2(u_multiplier_pp1_37 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_3__20_  (.A(u_multiplier_pp1_37 [9]),
    .B(u_multiplier_pp1_37 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_37_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_3__21_  (.A1(u_multiplier_pp1_37 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_37_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_3__22_  (.A(u_multiplier_pp1_37 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_37_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_37_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_3__23_  (.A1(u_multiplier_pp1_37 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_37_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_3__24_  (.A(u_multiplier_pp1_37 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_37_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_3__25_  (.A(u_multiplier_STAGE2_pp2_36_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_37_3__16_ ),
    .ZN(u_multiplier_pp2_37 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_37_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_37_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_37_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_37_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_37_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_37_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_37_3__17_ ),
    .ZN(u_multiplier_pp2_38 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_37_4__18_  (.A(u_multiplier_STAGE2_pp2_36_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_4__19_  (.A1(u_multiplier_pp1_37 [13]),
    .A2(u_multiplier_pp1_37 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_4__20_  (.A(u_multiplier_pp1_37 [13]),
    .B(u_multiplier_pp1_37 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_37_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_4__21_  (.A1(u_multiplier_pp1_37 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_37_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_4__22_  (.A(u_multiplier_pp1_37 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_37_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_37_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_4__23_  (.A1(u_multiplier_pp1_37 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_37_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_4__24_  (.A(u_multiplier_pp1_37 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_37_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_4__25_  (.A(u_multiplier_STAGE2_pp2_36_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_37_4__16_ ),
    .ZN(u_multiplier_pp2_37 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_37_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_37_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_37_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_37_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_37_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_37_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_37_4__17_ ),
    .ZN(u_multiplier_pp2_38 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_38_1__18_  (.A(u_multiplier_STAGE2_pp2_37_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_1__19_  (.A1(u_multiplier_pp1_38 [1]),
    .A2(u_multiplier_pp1_38 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_1__20_  (.A(u_multiplier_pp1_38 [1]),
    .B(u_multiplier_pp1_38 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_38_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_1__21_  (.A1(u_multiplier_pp1_38 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_38_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_1__22_  (.A(u_multiplier_pp1_38 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_38_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_38_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_1__23_  (.A1(u_multiplier_pp1_38 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_38_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_1__24_  (.A(u_multiplier_pp1_38 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_38_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_1__25_  (.A(u_multiplier_STAGE2_pp2_37_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_38_1__16_ ),
    .ZN(u_multiplier_pp2_38 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_38_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_38_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_38_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE2_E_4_2_pp2_38_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_38_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_38_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_38_1__17_ ),
    .ZN(u_multiplier_pp2_39 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_38_2__18_  (.A(u_multiplier_STAGE2_pp2_37_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_2__19_  (.A1(u_multiplier_pp1_38 [5]),
    .A2(u_multiplier_pp1_38 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_2__20_  (.A(u_multiplier_pp1_38 [5]),
    .B(u_multiplier_pp1_38 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_38_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_2__21_  (.A1(u_multiplier_pp1_38 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_38_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_2__22_  (.A(u_multiplier_pp1_38 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_38_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_38_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_2__23_  (.A1(u_multiplier_pp1_38 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_38_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_2__24_  (.A(u_multiplier_pp1_38 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_38_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_2__25_  (.A(u_multiplier_STAGE2_pp2_37_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_38_2__16_ ),
    .ZN(u_multiplier_pp2_38 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_38_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_38_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_38_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_38_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_38_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_38_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_38_2__17_ ),
    .ZN(u_multiplier_pp2_39 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_38_3__18_  (.A(u_multiplier_STAGE2_pp2_37_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_3__19_  (.A1(u_multiplier_pp1_38 [9]),
    .A2(u_multiplier_pp1_38 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_3__20_  (.A(u_multiplier_pp1_38 [9]),
    .B(u_multiplier_pp1_38 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_38_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_3__21_  (.A1(u_multiplier_pp1_38 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_38_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_3__22_  (.A(u_multiplier_pp1_38 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_38_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_38_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_3__23_  (.A1(u_multiplier_pp1_38 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_38_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_3__24_  (.A(u_multiplier_pp1_38 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_38_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_3__25_  (.A(u_multiplier_STAGE2_pp2_37_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_38_3__16_ ),
    .ZN(u_multiplier_pp2_38 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_38_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_38_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_38_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_38_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_38_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_38_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_38_3__17_ ),
    .ZN(u_multiplier_pp2_39 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_38_4__18_  (.A(u_multiplier_STAGE2_pp2_37_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_4__19_  (.A1(u_multiplier_pp1_38 [13]),
    .A2(u_multiplier_pp1_38 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_4__20_  (.A(u_multiplier_pp1_38 [13]),
    .B(u_multiplier_pp1_38 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_38_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_4__21_  (.A1(u_multiplier_pp1_38 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_38_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_4__22_  (.A(u_multiplier_pp1_38 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_38_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_38_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_4__23_  (.A1(u_multiplier_pp1_38 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_38_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_4__24_  (.A(u_multiplier_pp1_38 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_38_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_4__25_  (.A(u_multiplier_STAGE2_pp2_37_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_38_4__16_ ),
    .ZN(u_multiplier_pp2_38 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_38_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_38_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_38_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_38_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_38_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_38_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_38_4__17_ ),
    .ZN(u_multiplier_pp2_39 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_39_1__18_  (.A(u_multiplier_STAGE2_pp2_38_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_1__19_  (.A1(u_multiplier_pp1_39 [1]),
    .A2(u_multiplier_pp1_39 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_1__20_  (.A(u_multiplier_pp1_39 [1]),
    .B(u_multiplier_pp1_39 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_39_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_1__21_  (.A1(u_multiplier_pp1_39 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_39_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_1__22_  (.A(u_multiplier_pp1_39 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_39_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_39_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_1__23_  (.A1(u_multiplier_pp1_39 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_39_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_1__24_  (.A(u_multiplier_pp1_39 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_39_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_1__25_  (.A(u_multiplier_STAGE2_pp2_38_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_39_1__16_ ),
    .ZN(u_multiplier_pp2_39 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_39_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_39_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_39_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_39_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_39_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_39_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_39_1__17_ ),
    .ZN(u_multiplier_pp2_40 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_39_2__18_  (.A(u_multiplier_STAGE2_pp2_38_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_2__19_  (.A1(u_multiplier_pp1_39 [5]),
    .A2(u_multiplier_pp1_39 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_2__20_  (.A(u_multiplier_pp1_39 [5]),
    .B(u_multiplier_pp1_39 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_39_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_2__21_  (.A1(u_multiplier_pp1_39 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_39_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_2__22_  (.A(u_multiplier_pp1_39 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_39_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_39_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_2__23_  (.A1(u_multiplier_pp1_39 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_39_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_2__24_  (.A(u_multiplier_pp1_39 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_39_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_2__25_  (.A(u_multiplier_STAGE2_pp2_38_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_39_2__16_ ),
    .ZN(u_multiplier_pp2_39 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_39_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_39_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_39_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_39_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_39_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_39_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_39_2__17_ ),
    .ZN(u_multiplier_pp2_40 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_39_3__18_  (.A(u_multiplier_STAGE2_pp2_38_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_3__19_  (.A1(u_multiplier_pp1_39 [9]),
    .A2(u_multiplier_pp1_39 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_3__20_  (.A(u_multiplier_pp1_39 [9]),
    .B(u_multiplier_pp1_39 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_39_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_3__21_  (.A1(u_multiplier_pp1_39 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_39_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_3__22_  (.A(u_multiplier_pp1_39 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_39_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_39_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_3__23_  (.A1(u_multiplier_pp1_39 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_39_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_3__24_  (.A(u_multiplier_pp1_39 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_39_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_3__25_  (.A(u_multiplier_STAGE2_pp2_38_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_39_3__16_ ),
    .ZN(u_multiplier_pp2_39 [1]));
 NAND2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_39_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_39_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_39_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_39_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_39_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_39_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_39_3__17_ ),
    .ZN(u_multiplier_pp2_40 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_39_4__18_  (.A(u_multiplier_STAGE2_pp2_38_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_4__19_  (.A1(u_multiplier_pp1_39 [13]),
    .A2(u_multiplier_pp1_39 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_4__20_  (.A(u_multiplier_pp1_39 [13]),
    .B(u_multiplier_pp1_39 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_39_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_4__21_  (.A1(u_multiplier_pp1_39 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_39_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_4__22_  (.A(u_multiplier_pp1_39 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_39_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_39_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_4__23_  (.A1(u_multiplier_pp1_39 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_39_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_4__24_  (.A(u_multiplier_pp1_39 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_39_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_4__25_  (.A(u_multiplier_STAGE2_pp2_38_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_39_4__16_ ),
    .ZN(u_multiplier_pp2_39 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_39_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_39_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_39_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_39_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_39_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_39_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_39_4__17_ ),
    .ZN(u_multiplier_pp2_40 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_40_1__18_  (.A(u_multiplier_STAGE2_pp2_39_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_1__19_  (.A1(u_multiplier_pp1_40 [1]),
    .A2(u_multiplier_pp1_40 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_1__20_  (.A(u_multiplier_pp1_40 [1]),
    .B(u_multiplier_pp1_40 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_40_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_1__21_  (.A1(u_multiplier_pp1_40 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_40_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_1__22_  (.A(u_multiplier_pp1_40 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_40_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_40_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_1__23_  (.A1(u_multiplier_pp1_40 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_40_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_1__24_  (.A(u_multiplier_pp1_40 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_40_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_1__25_  (.A(u_multiplier_STAGE2_pp2_39_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_40_1__16_ ),
    .ZN(u_multiplier_pp2_40 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_40_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_40_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_40_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE2_E_4_2_pp2_40_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_40_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_40_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_40_1__17_ ),
    .ZN(u_multiplier_pp2_41 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_40_2__18_  (.A(u_multiplier_STAGE2_pp2_39_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_2__19_  (.A1(u_multiplier_pp1_40 [5]),
    .A2(u_multiplier_pp1_40 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_2__20_  (.A(u_multiplier_pp1_40 [5]),
    .B(u_multiplier_pp1_40 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_40_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_2__21_  (.A1(u_multiplier_pp1_40 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_40_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_2__22_  (.A(u_multiplier_pp1_40 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_40_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_40_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_2__23_  (.A1(u_multiplier_pp1_40 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_40_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_2__24_  (.A(u_multiplier_pp1_40 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_40_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_2__25_  (.A(u_multiplier_STAGE2_pp2_39_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_40_2__16_ ),
    .ZN(u_multiplier_pp2_40 [2]));
 NAND2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_40_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_40_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_40_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_40_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_40_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_40_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_40_2__17_ ),
    .ZN(u_multiplier_pp2_41 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_40_3__18_  (.A(u_multiplier_STAGE2_pp2_39_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_3__19_  (.A1(u_multiplier_pp1_40 [9]),
    .A2(u_multiplier_pp1_40 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_3__20_  (.A(u_multiplier_pp1_40 [9]),
    .B(u_multiplier_pp1_40 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_40_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_3__21_  (.A1(u_multiplier_pp1_40 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_40_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_3__22_  (.A(u_multiplier_pp1_40 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_40_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_40_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_3__23_  (.A1(u_multiplier_pp1_40 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_40_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_3__24_  (.A(u_multiplier_pp1_40 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_40_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_3__25_  (.A(u_multiplier_STAGE2_pp2_39_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_40_3__16_ ),
    .ZN(u_multiplier_pp2_40 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_40_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_40_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_40_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_40_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_40_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_40_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_40_3__17_ ),
    .ZN(u_multiplier_pp2_41 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_40_4__18_  (.A(u_multiplier_STAGE2_pp2_39_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_4__19_  (.A1(u_multiplier_pp1_40 [13]),
    .A2(u_multiplier_pp1_40 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_4__20_  (.A(u_multiplier_pp1_40 [13]),
    .B(u_multiplier_pp1_40 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_40_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_4__21_  (.A1(u_multiplier_pp1_40 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_40_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_4__22_  (.A(u_multiplier_pp1_40 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_40_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_40_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_4__23_  (.A1(u_multiplier_pp1_40 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_40_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_4__24_  (.A(u_multiplier_pp1_40 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_40_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_4__25_  (.A(u_multiplier_STAGE2_pp2_39_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_40_4__16_ ),
    .ZN(u_multiplier_pp2_40 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_40_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_40_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_40_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_40_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_40_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_40_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_40_4__17_ ),
    .ZN(u_multiplier_pp2_41 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_41_1__18_  (.A(u_multiplier_STAGE2_pp2_40_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_1__19_  (.A1(u_multiplier_pp1_41 [1]),
    .A2(u_multiplier_pp1_41 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_1__20_  (.A(u_multiplier_pp1_41 [1]),
    .B(u_multiplier_pp1_41 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_41_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_1__21_  (.A1(u_multiplier_pp1_41 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_41_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_1__22_  (.A(u_multiplier_pp1_41 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_41_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_41_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_1__23_  (.A1(u_multiplier_pp1_41 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_41_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_1__24_  (.A(u_multiplier_pp1_41 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_41_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_1__25_  (.A(u_multiplier_STAGE2_pp2_40_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_41_1__16_ ),
    .ZN(u_multiplier_pp2_41 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_41_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_41_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_41_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_41_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_41_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_41_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_41_1__17_ ),
    .ZN(u_multiplier_pp2_42 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_41_2__18_  (.A(u_multiplier_STAGE2_pp2_40_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_2__19_  (.A1(u_multiplier_pp1_41 [5]),
    .A2(u_multiplier_pp1_41 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_2__20_  (.A(u_multiplier_pp1_41 [5]),
    .B(u_multiplier_pp1_41 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_41_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_2__21_  (.A1(u_multiplier_pp1_41 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_41_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_2__22_  (.A(u_multiplier_pp1_41 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_41_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_41_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_2__23_  (.A1(u_multiplier_pp1_41 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_41_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_2__24_  (.A(u_multiplier_pp1_41 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_41_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_2__25_  (.A(u_multiplier_STAGE2_pp2_40_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_41_2__16_ ),
    .ZN(u_multiplier_pp2_41 [2]));
 NAND2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_41_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_41_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_41_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_41_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_41_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_41_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_41_2__17_ ),
    .ZN(u_multiplier_pp2_42 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_41_3__18_  (.A(u_multiplier_STAGE2_pp2_40_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_3__19_  (.A1(u_multiplier_pp1_41 [9]),
    .A2(u_multiplier_pp1_41 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_3__20_  (.A(u_multiplier_pp1_41 [9]),
    .B(u_multiplier_pp1_41 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_41_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_3__21_  (.A1(u_multiplier_pp1_41 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_41_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_3__22_  (.A(u_multiplier_pp1_41 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_41_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_41_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_3__23_  (.A1(u_multiplier_pp1_41 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_41_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_3__24_  (.A(u_multiplier_pp1_41 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_41_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_3__25_  (.A(u_multiplier_STAGE2_pp2_40_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_41_3__16_ ),
    .ZN(u_multiplier_pp2_41 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_41_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_41_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_41_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_41_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_41_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_41_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_41_3__17_ ),
    .ZN(u_multiplier_pp2_42 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_41_4__18_  (.A(u_multiplier_STAGE2_pp2_40_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_4__19_  (.A1(u_multiplier_pp1_41 [13]),
    .A2(u_multiplier_pp1_41 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_4__20_  (.A(u_multiplier_pp1_41 [13]),
    .B(u_multiplier_pp1_41 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_41_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_4__21_  (.A1(u_multiplier_pp1_41 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_41_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_4__22_  (.A(u_multiplier_pp1_41 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_41_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_41_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_4__23_  (.A1(u_multiplier_pp1_41 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_41_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_4__24_  (.A(u_multiplier_pp1_41 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_41_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_4__25_  (.A(u_multiplier_STAGE2_pp2_40_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_41_4__16_ ),
    .ZN(u_multiplier_pp2_41 [0]));
 NAND2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_41_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_41_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_41_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_41_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_41_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_41_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_41_4__17_ ),
    .ZN(u_multiplier_pp2_42 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_42_1__18_  (.A(u_multiplier_STAGE2_pp2_41_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_1__19_  (.A1(u_multiplier_pp1_42 [1]),
    .A2(u_multiplier_pp1_42 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_1__20_  (.A(u_multiplier_pp1_42 [1]),
    .B(u_multiplier_pp1_42 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_42_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_1__21_  (.A1(u_multiplier_pp1_42 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_42_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_1__22_  (.A(u_multiplier_pp1_42 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_42_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_42_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_1__23_  (.A1(u_multiplier_pp1_42 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_42_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_1__24_  (.A(u_multiplier_pp1_42 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_42_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_1__25_  (.A(u_multiplier_STAGE2_pp2_41_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_42_1__16_ ),
    .ZN(u_multiplier_pp2_42 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_42_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_42_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_42_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE2_E_4_2_pp2_42_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_42_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_42_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_42_1__17_ ),
    .ZN(u_multiplier_pp2_43 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_42_2__18_  (.A(u_multiplier_STAGE2_pp2_41_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_2__19_  (.A1(u_multiplier_pp1_42 [5]),
    .A2(u_multiplier_pp1_42 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_2__20_  (.A(u_multiplier_pp1_42 [5]),
    .B(u_multiplier_pp1_42 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_42_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_2__21_  (.A1(u_multiplier_pp1_42 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_42_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_2__22_  (.A(u_multiplier_pp1_42 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_42_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_42_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_2__23_  (.A1(u_multiplier_pp1_42 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_42_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_2__24_  (.A(u_multiplier_pp1_42 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_42_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_2__25_  (.A(u_multiplier_STAGE2_pp2_41_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_42_2__16_ ),
    .ZN(u_multiplier_pp2_42 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_42_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_42_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_42_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_42_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_42_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_42_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_42_2__17_ ),
    .ZN(u_multiplier_pp2_43 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_42_3__18_  (.A(u_multiplier_STAGE2_pp2_41_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_3__19_  (.A1(u_multiplier_pp1_42 [9]),
    .A2(u_multiplier_pp1_42 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_3__20_  (.A(u_multiplier_pp1_42 [9]),
    .B(u_multiplier_pp1_42 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_42_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_3__21_  (.A1(u_multiplier_pp1_42 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_42_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_3__22_  (.A(u_multiplier_pp1_42 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_42_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_42_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_3__23_  (.A1(u_multiplier_pp1_42 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_42_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_3__24_  (.A(u_multiplier_pp1_42 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_42_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_3__25_  (.A(u_multiplier_STAGE2_pp2_41_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_42_3__16_ ),
    .ZN(u_multiplier_pp2_42 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_42_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_42_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_42_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_42_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_42_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_42_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_42_3__17_ ),
    .ZN(u_multiplier_pp2_43 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_42_4__18_  (.A(u_multiplier_STAGE2_pp2_41_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_4__19_  (.A1(u_multiplier_pp1_42 [13]),
    .A2(u_multiplier_pp1_42 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_4__20_  (.A(u_multiplier_pp1_42 [13]),
    .B(u_multiplier_pp1_42 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_42_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_4__21_  (.A1(u_multiplier_pp1_42 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_42_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_4__22_  (.A(u_multiplier_pp1_42 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_42_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_42_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_4__23_  (.A1(u_multiplier_pp1_42 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_42_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_4__24_  (.A(u_multiplier_pp1_42 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_42_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_4__25_  (.A(u_multiplier_STAGE2_pp2_41_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_42_4__16_ ),
    .ZN(u_multiplier_pp2_42 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_42_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_42_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_42_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_42_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_42_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_42_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_42_4__17_ ),
    .ZN(u_multiplier_pp2_43 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_43_1__18_  (.A(u_multiplier_STAGE2_pp2_42_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_1__19_  (.A1(u_multiplier_pp1_43 [1]),
    .A2(u_multiplier_pp1_43 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_1__20_  (.A(u_multiplier_pp1_43 [1]),
    .B(u_multiplier_pp1_43 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_43_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_1__21_  (.A1(u_multiplier_pp1_43 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_43_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_1__22_  (.A(u_multiplier_pp1_43 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_43_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_43_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_1__23_  (.A1(u_multiplier_pp1_43 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_43_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_1__24_  (.A(u_multiplier_pp1_43 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_43_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_1__25_  (.A(u_multiplier_STAGE2_pp2_42_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_43_1__16_ ),
    .ZN(u_multiplier_pp2_43 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_43_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_43_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_43_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE2_E_4_2_pp2_43_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_43_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_43_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_43_1__17_ ),
    .ZN(u_multiplier_pp2_44 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_43_2__18_  (.A(u_multiplier_STAGE2_pp2_42_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_2__19_  (.A1(u_multiplier_pp1_43 [5]),
    .A2(u_multiplier_pp1_43 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_2__20_  (.A(u_multiplier_pp1_43 [5]),
    .B(u_multiplier_pp1_43 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_43_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_2__21_  (.A1(u_multiplier_pp1_43 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_43_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_2__22_  (.A(u_multiplier_pp1_43 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_43_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_43_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_2__23_  (.A1(u_multiplier_pp1_43 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_43_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_2__24_  (.A(u_multiplier_pp1_43 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_43_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_2__25_  (.A(u_multiplier_STAGE2_pp2_42_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_43_2__16_ ),
    .ZN(u_multiplier_pp2_43 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_43_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_43_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_43_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_43_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_43_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_43_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_43_2__17_ ),
    .ZN(u_multiplier_pp2_44 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_43_3__18_  (.A(u_multiplier_STAGE2_pp2_42_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_3__19_  (.A1(u_multiplier_pp1_43 [9]),
    .A2(u_multiplier_pp1_43 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_3__20_  (.A(u_multiplier_pp1_43 [9]),
    .B(u_multiplier_pp1_43 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_43_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_3__21_  (.A1(u_multiplier_pp1_43 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_43_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_3__22_  (.A(u_multiplier_pp1_43 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_43_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_43_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_3__23_  (.A1(u_multiplier_pp1_43 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_43_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_3__24_  (.A(u_multiplier_pp1_43 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_43_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_3__25_  (.A(u_multiplier_STAGE2_pp2_42_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_43_3__16_ ),
    .ZN(u_multiplier_pp2_43 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_43_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_43_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_43_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_43_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_43_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_43_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_43_3__17_ ),
    .ZN(u_multiplier_pp2_44 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_43_4__18_  (.A(u_multiplier_STAGE2_pp2_42_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_4__19_  (.A1(u_multiplier_pp1_43 [13]),
    .A2(u_multiplier_pp1_43 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_4__20_  (.A(u_multiplier_pp1_43 [13]),
    .B(u_multiplier_pp1_43 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_43_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_4__21_  (.A1(u_multiplier_pp1_43 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_43_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_4__22_  (.A(u_multiplier_pp1_43 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_43_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_43_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_4__23_  (.A1(u_multiplier_pp1_43 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_43_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_4__24_  (.A(u_multiplier_pp1_43 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_43_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_4__25_  (.A(u_multiplier_STAGE2_pp2_42_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_43_4__16_ ),
    .ZN(u_multiplier_pp2_43 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_43_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_43_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_43_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_43_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_43_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_43_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_43_4__17_ ),
    .ZN(u_multiplier_pp2_44 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_44_1__18_  (.A(u_multiplier_STAGE2_pp2_43_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_1__19_  (.A1(u_multiplier_pp1_44 [1]),
    .A2(u_multiplier_pp1_44 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_1__20_  (.A(u_multiplier_pp1_44 [1]),
    .B(u_multiplier_pp1_44 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_44_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_1__21_  (.A1(u_multiplier_pp1_44 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_44_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_1__22_  (.A(u_multiplier_pp1_44 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_44_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_44_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_1__23_  (.A1(u_multiplier_pp1_44 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_44_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_1__24_  (.A(u_multiplier_pp1_44 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_44_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_1__25_  (.A(u_multiplier_STAGE2_pp2_43_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_44_1__16_ ),
    .ZN(u_multiplier_pp2_44 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_44_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_44_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_44_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE2_E_4_2_pp2_44_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_44_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_44_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_44_1__17_ ),
    .ZN(u_multiplier_pp2_45 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_44_2__18_  (.A(u_multiplier_STAGE2_pp2_43_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_2__19_  (.A1(u_multiplier_pp1_44 [5]),
    .A2(u_multiplier_pp1_44 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_2__20_  (.A(u_multiplier_pp1_44 [5]),
    .B(u_multiplier_pp1_44 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_44_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_2__21_  (.A1(u_multiplier_pp1_44 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_44_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_2__22_  (.A(u_multiplier_pp1_44 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_44_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_44_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_2__23_  (.A1(u_multiplier_pp1_44 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_44_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_2__24_  (.A(u_multiplier_pp1_44 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_44_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_2__25_  (.A(u_multiplier_STAGE2_pp2_43_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_44_2__16_ ),
    .ZN(u_multiplier_pp2_44 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_44_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_44_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_44_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_44_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_44_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_44_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_44_2__17_ ),
    .ZN(u_multiplier_pp2_45 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_44_3__18_  (.A(u_multiplier_STAGE2_pp2_43_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_3__19_  (.A1(u_multiplier_pp1_44 [9]),
    .A2(u_multiplier_pp1_44 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_3__20_  (.A(u_multiplier_pp1_44 [9]),
    .B(u_multiplier_pp1_44 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_44_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_3__21_  (.A1(u_multiplier_pp1_44 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_44_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_3__22_  (.A(u_multiplier_pp1_44 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_44_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_44_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_3__23_  (.A1(u_multiplier_pp1_44 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_44_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_3__24_  (.A(u_multiplier_pp1_44 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_44_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_3__25_  (.A(u_multiplier_STAGE2_pp2_43_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_44_3__16_ ),
    .ZN(u_multiplier_pp2_44 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_44_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_44_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_44_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_44_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_44_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_44_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_44_3__17_ ),
    .ZN(u_multiplier_pp2_45 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_44_4__18_  (.A(u_multiplier_STAGE2_pp2_43_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_4__19_  (.A1(u_multiplier_pp1_44 [13]),
    .A2(u_multiplier_pp1_44 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_4__20_  (.A(u_multiplier_pp1_44 [13]),
    .B(u_multiplier_pp1_44 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_44_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_4__21_  (.A1(u_multiplier_pp1_44 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_44_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_4__22_  (.A(u_multiplier_pp1_44 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_44_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_44_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_4__23_  (.A1(u_multiplier_pp1_44 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_44_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_4__24_  (.A(u_multiplier_pp1_44 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_44_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_4__25_  (.A(u_multiplier_STAGE2_pp2_43_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_44_4__16_ ),
    .ZN(u_multiplier_pp2_44 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_44_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_44_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_44_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_44_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_44_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_44_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_44_4__17_ ),
    .ZN(u_multiplier_pp2_45 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_45_1__18_  (.A(u_multiplier_STAGE2_pp2_44_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_1__19_  (.A1(u_multiplier_pp1_45 [1]),
    .A2(u_multiplier_pp1_45 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_1__20_  (.A(u_multiplier_pp1_45 [1]),
    .B(u_multiplier_pp1_45 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_45_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_1__21_  (.A1(u_multiplier_pp1_45 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_45_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_1__22_  (.A(u_multiplier_pp1_45 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_45_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_45_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_1__23_  (.A1(u_multiplier_pp1_45 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_45_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_1__24_  (.A(u_multiplier_pp1_45 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_45_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_1__25_  (.A(u_multiplier_STAGE2_pp2_44_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_45_1__16_ ),
    .ZN(u_multiplier_pp2_45 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_45_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_45_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_45_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_45_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_45_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_45_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_45_1__17_ ),
    .ZN(u_multiplier_pp2_46 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_45_2__18_  (.A(u_multiplier_STAGE2_pp2_44_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_2__19_  (.A1(u_multiplier_pp1_45 [5]),
    .A2(u_multiplier_pp1_45 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_2__20_  (.A(u_multiplier_pp1_45 [5]),
    .B(u_multiplier_pp1_45 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_45_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_2__21_  (.A1(u_multiplier_pp1_45 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_45_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_2__22_  (.A(u_multiplier_pp1_45 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_45_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_45_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_2__23_  (.A1(u_multiplier_pp1_45 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_45_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_2__24_  (.A(u_multiplier_pp1_45 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_45_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_2__25_  (.A(u_multiplier_STAGE2_pp2_44_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_45_2__16_ ),
    .ZN(u_multiplier_pp2_45 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_45_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_45_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_45_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_45_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_45_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_45_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_45_2__17_ ),
    .ZN(u_multiplier_pp2_46 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_45_3__18_  (.A(u_multiplier_STAGE2_pp2_44_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_3__19_  (.A1(u_multiplier_pp1_45 [9]),
    .A2(u_multiplier_pp1_45 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_3__20_  (.A(u_multiplier_pp1_45 [9]),
    .B(u_multiplier_pp1_45 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_45_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_3__21_  (.A1(u_multiplier_pp1_45 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_45_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_3__22_  (.A(u_multiplier_pp1_45 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_45_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_45_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_3__23_  (.A1(u_multiplier_pp1_45 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_45_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_3__24_  (.A(u_multiplier_pp1_45 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_45_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_3__25_  (.A(u_multiplier_STAGE2_pp2_44_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_45_3__16_ ),
    .ZN(u_multiplier_pp2_45 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_45_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_45_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_45_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_45_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_45_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_45_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_45_3__17_ ),
    .ZN(u_multiplier_pp2_46 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_45_4__18_  (.A(u_multiplier_STAGE2_pp2_44_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_4__19_  (.A1(u_multiplier_pp1_45 [13]),
    .A2(u_multiplier_pp1_45 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_4__20_  (.A(u_multiplier_pp1_45 [13]),
    .B(u_multiplier_pp1_45 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_45_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_4__21_  (.A1(u_multiplier_pp1_45 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_45_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_4__22_  (.A(u_multiplier_pp1_45 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_45_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_45_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_4__23_  (.A1(u_multiplier_pp1_45 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_45_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_4__24_  (.A(u_multiplier_pp1_45 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_45_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_4__25_  (.A(u_multiplier_STAGE2_pp2_44_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_45_4__16_ ),
    .ZN(u_multiplier_pp2_45 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_45_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_45_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_45_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_45_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_45_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_45_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_45_4__17_ ),
    .ZN(u_multiplier_pp2_46 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_46_1__18_  (.A(u_multiplier_STAGE2_pp2_45_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_1__19_  (.A1(u_multiplier_pp1_46 [1]),
    .A2(u_multiplier_pp1_46 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_1__20_  (.A(u_multiplier_pp1_46 [1]),
    .B(u_multiplier_pp1_46 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_46_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_1__21_  (.A1(u_multiplier_pp1_46 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_46_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_1__22_  (.A(u_multiplier_pp1_46 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_46_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_46_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_1__23_  (.A1(u_multiplier_pp1_46 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_46_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_1__24_  (.A(u_multiplier_pp1_46 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_46_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_1__25_  (.A(u_multiplier_STAGE2_pp2_45_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_46_1__16_ ),
    .ZN(u_multiplier_pp2_46 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_46_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_46_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_46_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_46_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_46_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_46_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_46_1__17_ ),
    .ZN(u_multiplier_pp2_47 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_46_2__18_  (.A(u_multiplier_STAGE2_pp2_45_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_2__19_  (.A1(u_multiplier_pp1_46 [5]),
    .A2(u_multiplier_pp1_46 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_2__20_  (.A(u_multiplier_pp1_46 [5]),
    .B(u_multiplier_pp1_46 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_46_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_2__21_  (.A1(u_multiplier_pp1_46 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_46_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_2__22_  (.A(u_multiplier_pp1_46 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_46_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_46_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_2__23_  (.A1(u_multiplier_pp1_46 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_46_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_2__24_  (.A(u_multiplier_pp1_46 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_46_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_2__25_  (.A(u_multiplier_STAGE2_pp2_45_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_46_2__16_ ),
    .ZN(u_multiplier_pp2_46 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_46_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_46_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_46_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_46_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_46_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_46_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_46_2__17_ ),
    .ZN(u_multiplier_pp2_47 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_46_3__18_  (.A(u_multiplier_STAGE2_pp2_45_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_3__19_  (.A1(u_multiplier_pp1_46 [9]),
    .A2(u_multiplier_pp1_46 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_3__20_  (.A(u_multiplier_pp1_46 [9]),
    .B(u_multiplier_pp1_46 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_46_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_3__21_  (.A1(u_multiplier_pp1_46 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_46_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_3__22_  (.A(u_multiplier_pp1_46 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_46_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_46_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_3__23_  (.A1(u_multiplier_pp1_46 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_46_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_3__24_  (.A(u_multiplier_pp1_46 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_46_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_3__25_  (.A(u_multiplier_STAGE2_pp2_45_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_46_3__16_ ),
    .ZN(u_multiplier_pp2_46 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_46_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_46_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_46_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_46_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_46_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_46_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_46_3__17_ ),
    .ZN(u_multiplier_pp2_47 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_46_4__18_  (.A(u_multiplier_STAGE2_pp2_45_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_4__19_  (.A1(u_multiplier_pp1_46 [13]),
    .A2(u_multiplier_pp1_46 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_4__20_  (.A(u_multiplier_pp1_46 [13]),
    .B(u_multiplier_pp1_46 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_46_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_4__21_  (.A1(u_multiplier_pp1_46 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_46_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_4__22_  (.A(u_multiplier_pp1_46 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_46_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_46_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_4__23_  (.A1(u_multiplier_pp1_46 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_46_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_4__24_  (.A(u_multiplier_pp1_46 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_46_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_4__25_  (.A(u_multiplier_STAGE2_pp2_45_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_46_4__16_ ),
    .ZN(u_multiplier_pp2_46 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_46_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_46_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_46_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_46_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_46_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_46_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_46_4__17_ ),
    .ZN(u_multiplier_pp2_47 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_47_1__18_  (.A(u_multiplier_STAGE2_pp2_46_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_1__19_  (.A1(u_multiplier_pp1_47 [1]),
    .A2(u_multiplier_pp1_47 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_1__20_  (.A(u_multiplier_pp1_47 [1]),
    .B(u_multiplier_pp1_47 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_47_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_1__21_  (.A1(u_multiplier_pp1_47 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_47_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_1__22_  (.A(u_multiplier_pp1_47 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_47_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_47_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_1__23_  (.A1(u_multiplier_pp1_47 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_47_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_1__24_  (.A(u_multiplier_pp1_47 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_47_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_1__25_  (.A(u_multiplier_STAGE2_pp2_46_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_47_1__16_ ),
    .ZN(u_multiplier_pp2_47 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_47_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_47_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_47_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_47_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_47_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_47_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_47_1__17_ ),
    .ZN(u_multiplier_pp2_48 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_47_2__18_  (.A(u_multiplier_STAGE2_pp2_46_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_2__19_  (.A1(u_multiplier_pp1_47 [5]),
    .A2(u_multiplier_pp1_47 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_2__20_  (.A(u_multiplier_pp1_47 [5]),
    .B(u_multiplier_pp1_47 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_47_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_2__21_  (.A1(u_multiplier_pp1_47 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_47_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_2__22_  (.A(u_multiplier_pp1_47 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_47_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_47_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_2__23_  (.A1(u_multiplier_pp1_47 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_47_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_2__24_  (.A(u_multiplier_pp1_47 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_47_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_2__25_  (.A(u_multiplier_STAGE2_pp2_46_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_47_2__16_ ),
    .ZN(u_multiplier_pp2_47 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_47_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_47_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_47_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_47_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_47_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_47_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_47_2__17_ ),
    .ZN(u_multiplier_pp2_48 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_47_3__18_  (.A(u_multiplier_STAGE2_pp2_46_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_3__19_  (.A1(u_multiplier_pp1_47 [9]),
    .A2(u_multiplier_pp1_47 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_3__20_  (.A(u_multiplier_pp1_47 [9]),
    .B(u_multiplier_pp1_47 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_47_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_3__21_  (.A1(u_multiplier_pp1_47 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_47_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_3__22_  (.A(u_multiplier_pp1_47 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_47_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_47_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_3__23_  (.A1(u_multiplier_pp1_47 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_47_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_3__24_  (.A(u_multiplier_pp1_47 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_47_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_3__25_  (.A(u_multiplier_STAGE2_pp2_46_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_47_3__16_ ),
    .ZN(u_multiplier_pp2_47 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_47_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_47_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_47_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_47_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_47_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_47_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_47_3__17_ ),
    .ZN(u_multiplier_pp2_48 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_47_4__18_  (.A(u_multiplier_STAGE2_pp2_46_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_4__19_  (.A1(u_multiplier_pp1_47 [13]),
    .A2(u_multiplier_pp1_47 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_4__20_  (.A(u_multiplier_pp1_47 [13]),
    .B(u_multiplier_pp1_47 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_47_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_4__21_  (.A1(u_multiplier_pp1_47 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_47_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_4__22_  (.A(u_multiplier_pp1_47 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_47_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_47_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_4__23_  (.A1(u_multiplier_pp1_47 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_47_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_4__24_  (.A(u_multiplier_pp1_47 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_47_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_4__25_  (.A(u_multiplier_STAGE2_pp2_46_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_47_4__16_ ),
    .ZN(u_multiplier_pp2_47 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_47_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_47_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_47_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_47_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_47_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_47_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_47_4__17_ ),
    .ZN(u_multiplier_pp2_48 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_48_1__18_  (.A(u_multiplier_STAGE2_pp2_47_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_1__19_  (.A1(u_multiplier_pp1_48 [1]),
    .A2(u_multiplier_pp1_48 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_1__20_  (.A(u_multiplier_pp1_48 [1]),
    .B(u_multiplier_pp1_48 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_48_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_1__21_  (.A1(u_multiplier_pp1_48 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_48_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_1__22_  (.A(u_multiplier_pp1_48 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_48_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_48_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_1__23_  (.A1(u_multiplier_pp1_48 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_48_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_1__24_  (.A(u_multiplier_pp1_48 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_48_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_1__25_  (.A(u_multiplier_STAGE2_pp2_47_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_48_1__16_ ),
    .ZN(u_multiplier_pp2_48 [3]));
 NAND2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_48_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_48_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_48_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_48_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_48_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_48_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_48_1__17_ ),
    .ZN(u_multiplier_pp2_49 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_48_2__18_  (.A(u_multiplier_STAGE2_pp2_47_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_2__19_  (.A1(u_multiplier_pp1_48 [5]),
    .A2(u_multiplier_pp1_48 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_2__20_  (.A(u_multiplier_pp1_48 [5]),
    .B(u_multiplier_pp1_48 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_48_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_2__21_  (.A1(u_multiplier_pp1_48 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_48_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_2__22_  (.A(u_multiplier_pp1_48 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_48_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_48_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_2__23_  (.A1(u_multiplier_pp1_48 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_48_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_2__24_  (.A(u_multiplier_pp1_48 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_48_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_2__25_  (.A(u_multiplier_STAGE2_pp2_47_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_48_2__16_ ),
    .ZN(u_multiplier_pp2_48 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_48_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_48_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_48_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_48_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_48_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_48_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_48_2__17_ ),
    .ZN(u_multiplier_pp2_49 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_48_3__18_  (.A(u_multiplier_STAGE2_pp2_47_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_3__19_  (.A1(u_multiplier_pp1_48 [9]),
    .A2(u_multiplier_pp1_48 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_3__20_  (.A(u_multiplier_pp1_48 [9]),
    .B(u_multiplier_pp1_48 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_48_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_3__21_  (.A1(u_multiplier_pp1_48 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_48_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_3__22_  (.A(u_multiplier_pp1_48 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_48_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_48_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_3__23_  (.A1(u_multiplier_pp1_48 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_48_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_3__24_  (.A(u_multiplier_pp1_48 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_48_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_3__25_  (.A(u_multiplier_STAGE2_pp2_47_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_48_3__16_ ),
    .ZN(u_multiplier_pp2_48 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_48_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_48_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_48_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_48_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_48_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_48_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_48_3__17_ ),
    .ZN(u_multiplier_pp2_49 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_48_4__18_  (.A(u_multiplier_STAGE2_pp2_47_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_4__19_  (.A1(u_multiplier_pp1_48 [13]),
    .A2(u_multiplier_pp1_48 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_4__20_  (.A(u_multiplier_pp1_48 [13]),
    .B(u_multiplier_pp1_48 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_48_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_4__21_  (.A1(u_multiplier_pp1_48 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_48_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_4__22_  (.A(u_multiplier_pp1_48 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_48_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_48_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_4__23_  (.A1(u_multiplier_pp1_48 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_48_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_4__24_  (.A(u_multiplier_pp1_48 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_48_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_4__25_  (.A(u_multiplier_STAGE2_pp2_47_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_48_4__16_ ),
    .ZN(u_multiplier_pp2_48 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_48_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_48_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_48_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_48_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_48_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_48_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_48_4__17_ ),
    .ZN(u_multiplier_pp2_49 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_49_1__18_  (.A(u_multiplier_STAGE2_pp2_48_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_49_1__19_  (.A1(u_multiplier_pp1_49 [1]),
    .A2(u_multiplier_pp1_49 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_49_1__20_  (.A(u_multiplier_pp1_49 [1]),
    .B(u_multiplier_pp1_49 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_49_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_49_1__21_  (.A1(u_multiplier_pp1_49 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_49_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_49_1__22_  (.A(u_multiplier_pp1_49 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_49_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_49_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_49_1__23_  (.A1(u_multiplier_pp1_49 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_49_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_49_1__24_  (.A(u_multiplier_pp1_49 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_49_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_49_1__25_  (.A(u_multiplier_STAGE2_pp2_48_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_49_1__16_ ),
    .ZN(u_multiplier_pp2_49 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_49_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_49_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_49_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_49_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_49_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_49_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_49_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_49_1__17_ ),
    .ZN(u_multiplier_pp2_50 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_49_2__18_  (.A(u_multiplier_STAGE2_pp2_48_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_49_2__19_  (.A1(u_multiplier_pp1_49 [5]),
    .A2(u_multiplier_pp1_49 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_49_2__20_  (.A(u_multiplier_pp1_49 [5]),
    .B(u_multiplier_pp1_49 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_49_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_49_2__21_  (.A1(u_multiplier_pp1_49 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_49_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_49_2__22_  (.A(u_multiplier_pp1_49 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_49_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_49_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_49_2__23_  (.A1(u_multiplier_pp1_49 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_49_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_49_2__24_  (.A(u_multiplier_pp1_49 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_49_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_49_2__25_  (.A(u_multiplier_STAGE2_pp2_48_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_49_2__16_ ),
    .ZN(u_multiplier_pp2_49 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_49_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_49_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_49_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_49_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_49_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_49_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_49_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_49_2__17_ ),
    .ZN(u_multiplier_pp2_50 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_49_3__18_  (.A(u_multiplier_STAGE2_pp2_48_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_49_3__19_  (.A1(u_multiplier_pp1_49 [9]),
    .A2(u_multiplier_pp1_49 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_49_3__20_  (.A(u_multiplier_pp1_49 [9]),
    .B(u_multiplier_pp1_49 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_49_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_49_3__21_  (.A1(u_multiplier_pp1_49 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_49_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_49_3__22_  (.A(u_multiplier_pp1_49 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_49_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_49_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_49_3__23_  (.A1(u_multiplier_pp1_49 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_49_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_49_3__24_  (.A(u_multiplier_pp1_49 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_49_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_49_3__25_  (.A(u_multiplier_STAGE2_pp2_48_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_49_3__16_ ),
    .ZN(u_multiplier_pp2_49 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_49_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_49_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_49_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_49_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_49_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_49_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_49_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_49_3__17_ ),
    .ZN(u_multiplier_pp2_50 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_50_1__18_  (.A(u_multiplier_STAGE2_pp2_49_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_50_1__19_  (.A1(u_multiplier_pp1_50 [1]),
    .A2(u_multiplier_pp1_50 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_50_1__20_  (.A(u_multiplier_pp1_50 [1]),
    .B(u_multiplier_pp1_50 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_50_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_50_1__21_  (.A1(u_multiplier_pp1_50 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_50_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_50_1__22_  (.A(u_multiplier_pp1_50 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_50_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_50_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_50_1__23_  (.A1(u_multiplier_pp1_50 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_50_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_50_1__24_  (.A(u_multiplier_pp1_50 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_50_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_50_1__25_  (.A(u_multiplier_STAGE2_pp2_49_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_50_1__16_ ),
    .ZN(u_multiplier_pp2_50 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_50_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_50_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_50_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_50_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_50_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_50_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_50_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_50_1__17_ ),
    .ZN(u_multiplier_pp2_51 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_50_2__18_  (.A(u_multiplier_STAGE2_pp2_49_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_50_2__19_  (.A1(u_multiplier_pp1_50 [5]),
    .A2(u_multiplier_pp1_50 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_50_2__20_  (.A(u_multiplier_pp1_50 [5]),
    .B(u_multiplier_pp1_50 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_50_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_50_2__21_  (.A1(u_multiplier_pp1_50 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_50_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_50_2__22_  (.A(u_multiplier_pp1_50 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_50_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_50_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_50_2__23_  (.A1(u_multiplier_pp1_50 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_50_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_50_2__24_  (.A(u_multiplier_pp1_50 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_50_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_50_2__25_  (.A(u_multiplier_STAGE2_pp2_49_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_50_2__16_ ),
    .ZN(u_multiplier_pp2_50 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_50_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_50_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_50_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_50_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_50_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_50_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_50_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_50_2__17_ ),
    .ZN(u_multiplier_pp2_51 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_50_3__18_  (.A(u_multiplier_STAGE2_pp2_49_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_50_3__19_  (.A1(u_multiplier_pp1_50 [9]),
    .A2(u_multiplier_pp1_50 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_50_3__20_  (.A(u_multiplier_pp1_50 [9]),
    .B(u_multiplier_pp1_50 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_50_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_50_3__21_  (.A1(u_multiplier_pp1_50 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_50_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_50_3__22_  (.A(u_multiplier_pp1_50 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_50_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_50_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_50_3__23_  (.A1(u_multiplier_pp1_50 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_50_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_50_3__24_  (.A(u_multiplier_pp1_50 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_50_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_50_3__25_  (.A(u_multiplier_STAGE2_pp2_49_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_50_3__16_ ),
    .ZN(u_multiplier_pp2_50 [0]));
 NAND2_X2 u_multiplier_STAGE2_E_4_2_pp2_50_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_50_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_50_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_50_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_50_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_50_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_50_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_50_3__17_ ),
    .ZN(u_multiplier_pp2_51 [3]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_51_1__18_  (.A(u_multiplier_STAGE2_pp2_50_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_51_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_51_1__19_  (.A1(u_multiplier_pp1_51 [1]),
    .A2(u_multiplier_pp1_51 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_51_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_51_1__20_  (.A(u_multiplier_pp1_51 [1]),
    .B(u_multiplier_pp1_51 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_51_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_51_1__21_  (.A1(u_multiplier_pp1_51 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_51_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_51_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_51_1__22_  (.A(u_multiplier_pp1_51 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_51_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_51_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_51_1__23_  (.A1(u_multiplier_pp1_51 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_51_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_51_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_51_1__24_  (.A(u_multiplier_pp1_51 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_51_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_51_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_51_1__25_  (.A(u_multiplier_STAGE2_pp2_50_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_51_1__16_ ),
    .ZN(u_multiplier_pp2_51 [2]));
 NAND2_X2 u_multiplier_STAGE2_E_4_2_pp2_51_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_51_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_51_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_51_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_51_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_51_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_51_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_51_1__17_ ),
    .ZN(u_multiplier_pp2_52 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_51_2__18_  (.A(u_multiplier_STAGE2_pp2_50_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_51_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_51_2__19_  (.A1(u_multiplier_pp1_51 [5]),
    .A2(u_multiplier_pp1_51 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_51_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_51_2__20_  (.A(u_multiplier_pp1_51 [5]),
    .B(u_multiplier_pp1_51 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_51_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_51_2__21_  (.A1(u_multiplier_pp1_51 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_51_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_51_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_51_2__22_  (.A(u_multiplier_pp1_51 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_51_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_51_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_51_2__23_  (.A1(u_multiplier_pp1_51 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_51_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_51_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_51_2__24_  (.A(u_multiplier_pp1_51 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_51_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_51_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_51_2__25_  (.A(u_multiplier_STAGE2_pp2_50_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_51_2__16_ ),
    .ZN(u_multiplier_pp2_51 [1]));
 NAND2_X2 u_multiplier_STAGE2_E_4_2_pp2_51_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_51_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_51_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_51_e42_2_cout ));
 OAI21_X1 u_multiplier_STAGE2_E_4_2_pp2_51_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_51_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_51_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_51_2__17_ ),
    .ZN(u_multiplier_pp2_52 [3]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_52_1__18_  (.A(u_multiplier_STAGE2_pp2_51_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_52_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_52_1__19_  (.A1(u_multiplier_pp1_52 [1]),
    .A2(u_multiplier_pp1_52 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_52_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_52_1__20_  (.A(u_multiplier_pp1_52 [1]),
    .B(u_multiplier_pp1_52 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_52_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_52_1__21_  (.A1(u_multiplier_pp1_52 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_52_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_52_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_52_1__22_  (.A(u_multiplier_pp1_52 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_52_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_52_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_52_1__23_  (.A1(u_multiplier_pp1_52 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_52_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_52_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_52_1__24_  (.A(u_multiplier_pp1_52 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_52_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_52_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_52_1__25_  (.A(u_multiplier_STAGE2_pp2_51_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_52_1__16_ ),
    .ZN(u_multiplier_pp2_52 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_52_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_52_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_52_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_52_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE2_E_4_2_pp2_52_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_52_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_52_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_52_1__17_ ),
    .ZN(u_multiplier_pp2_53 [3]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_52_2__18_  (.A(u_multiplier_STAGE2_pp2_51_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_52_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_52_2__19_  (.A1(u_multiplier_pp1_52 [5]),
    .A2(u_multiplier_pp1_52 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_52_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_52_2__20_  (.A(u_multiplier_pp1_52 [5]),
    .B(u_multiplier_pp1_52 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_52_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_52_2__21_  (.A1(u_multiplier_pp1_52 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_52_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_52_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_52_2__22_  (.A(u_multiplier_pp1_52 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_52_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_52_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_52_2__23_  (.A1(u_multiplier_pp1_52 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_52_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_52_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_52_2__24_  (.A(u_multiplier_pp1_52 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_52_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_52_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_52_2__25_  (.A(u_multiplier_STAGE2_pp2_51_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_52_2__16_ ),
    .ZN(u_multiplier_pp2_52 [0]));
 NAND2_X2 u_multiplier_STAGE2_E_4_2_pp2_52_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_52_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_52_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_52_e42_2_cout ));
 OAI21_X4 u_multiplier_STAGE2_E_4_2_pp2_52_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_52_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_52_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_52_2__17_ ),
    .ZN(u_multiplier_pp2_53 [2]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_53_1__18_  (.A(u_multiplier_STAGE2_pp2_52_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_53_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_53_1__19_  (.A1(u_multiplier_pp1_53 [1]),
    .A2(u_multiplier_pp1_53 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_53_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_53_1__20_  (.A(u_multiplier_pp1_53 [1]),
    .B(u_multiplier_pp1_53 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_53_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_53_1__21_  (.A1(u_multiplier_pp1_53 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_53_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_53_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_53_1__22_  (.A(u_multiplier_pp1_53 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_53_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_53_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_53_1__23_  (.A1(u_multiplier_pp1_53 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_53_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_53_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_53_1__24_  (.A(u_multiplier_pp1_53 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_53_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_53_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_53_1__25_  (.A(u_multiplier_STAGE2_pp2_52_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_53_1__16_ ),
    .ZN(u_multiplier_pp2_53 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_53_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_53_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_53_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_53_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_53_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_53_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_53_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_53_1__17_ ),
    .ZN(u_multiplier_pp2_54 [2]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_54_1__18_  (.A(u_multiplier_STAGE2_pp2_53_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_54_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_54_1__19_  (.A1(u_multiplier_pp1_54 [1]),
    .A2(u_multiplier_pp1_54 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_54_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_54_1__20_  (.A(u_multiplier_pp1_54 [1]),
    .B(u_multiplier_pp1_54 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_54_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_54_1__21_  (.A1(u_multiplier_pp1_54 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_54_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_54_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_54_1__22_  (.A(u_multiplier_pp1_54 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_54_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_54_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_54_1__23_  (.A1(u_multiplier_pp1_54 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_54_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_54_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_54_1__24_  (.A(u_multiplier_pp1_54 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_54_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_54_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_54_1__25_  (.A(u_multiplier_STAGE2_pp2_53_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_54_1__16_ ),
    .ZN(u_multiplier_pp2_54 [0]));
 NAND2_X2 u_multiplier_STAGE2_E_4_2_pp2_54_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_54_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_54_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_54_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_54_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_54_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_54_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_54_1__17_ ),
    .ZN(u_multiplier_pp2_55 [1]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_9_1__18_  (.A(net138),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_9_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_9_1__19_  (.A1(u_multiplier_pp1_9 [1]),
    .A2(u_multiplier_pp1_9 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_9_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_9_1__20_  (.A(u_multiplier_pp1_9 [1]),
    .B(u_multiplier_pp1_9 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_9_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_9_1__21_  (.A1(u_multiplier_pp1_9 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_9_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_9_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_9_1__22_  (.A(u_multiplier_pp1_9 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_9_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_9_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_9_1__23_  (.A1(u_multiplier_pp1_9 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_9_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_9_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_9_1__24_  (.A(u_multiplier_pp1_9 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_9_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_9_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_9_1__25_  (.A(net139),
    .B(u_multiplier_STAGE2_E_4_2_pp2_9_1__16_ ),
    .ZN(u_multiplier_pp2_9 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_9_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_9_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_9_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_9_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_9_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_9_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_9_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_9_1__17_ ),
    .ZN(u_multiplier_pp2_10 [2]));
 INV_X1 u_multiplier_STAGE2_Full_adder_pp2_49_1__12_  (.A(u_multiplier_STAGE2_pp2_48_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_49_1__08_ ));
 NAND3_X2 u_multiplier_STAGE2_Full_adder_pp2_49_1__13_  (.A1(u_multiplier_pp1_49 [13]),
    .A2(u_multiplier_pp1_49 [12]),
    .A3(u_multiplier_STAGE2_pp2_48_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_49_1__09_ ));
 NOR2_X2 u_multiplier_STAGE2_Full_adder_pp2_49_1__14_  (.A1(u_multiplier_pp1_49 [13]),
    .A2(u_multiplier_pp1_49 [12]),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_49_1__10_ ));
 AOI21_X1 u_multiplier_STAGE2_Full_adder_pp2_49_1__15_  (.A(u_multiplier_STAGE2_pp2_48_e42_4_cout ),
    .B1(u_multiplier_pp1_49 [12]),
    .B2(u_multiplier_pp1_49 [13]),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_49_1__11_ ));
 NOR2_X2 u_multiplier_STAGE2_Full_adder_pp2_49_1__16_  (.A1(u_multiplier_STAGE2_Full_adder_pp2_49_1__10_ ),
    .A2(u_multiplier_STAGE2_Full_adder_pp2_49_1__11_ ),
    .ZN(u_multiplier_pp2_50 [3]));
 AOI22_X4 u_multiplier_STAGE2_Full_adder_pp2_49_1__17_  (.A1(u_multiplier_STAGE2_Full_adder_pp2_49_1__08_ ),
    .A2(u_multiplier_STAGE2_Full_adder_pp2_49_1__10_ ),
    .B1(u_multiplier_pp2_50 [3]),
    .B2(u_multiplier_STAGE2_Full_adder_pp2_49_1__09_ ),
    .ZN(u_multiplier_pp2_49 [0]));
 INV_X1 u_multiplier_STAGE2_Full_adder_pp2_51_1__12_  (.A(u_multiplier_STAGE2_pp2_50_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_51_1__08_ ));
 NAND3_X2 u_multiplier_STAGE2_Full_adder_pp2_51_1__13_  (.A1(u_multiplier_pp1_51 [9]),
    .A2(u_multiplier_pp1_51 [8]),
    .A3(u_multiplier_STAGE2_pp2_50_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_51_1__09_ ));
 NOR2_X4 u_multiplier_STAGE2_Full_adder_pp2_51_1__14_  (.A1(u_multiplier_pp1_51 [9]),
    .A2(u_multiplier_pp1_51 [8]),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_51_1__10_ ));
 AOI21_X2 u_multiplier_STAGE2_Full_adder_pp2_51_1__15_  (.A(u_multiplier_STAGE2_pp2_50_e42_3_cout ),
    .B1(u_multiplier_pp1_51 [8]),
    .B2(u_multiplier_pp1_51 [9]),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_51_1__11_ ));
 NOR2_X4 u_multiplier_STAGE2_Full_adder_pp2_51_1__16_  (.A1(u_multiplier_STAGE2_Full_adder_pp2_51_1__10_ ),
    .A2(u_multiplier_STAGE2_Full_adder_pp2_51_1__11_ ),
    .ZN(u_multiplier_pp2_52 [2]));
 AOI22_X4 u_multiplier_STAGE2_Full_adder_pp2_51_1__17_  (.A1(u_multiplier_STAGE2_Full_adder_pp2_51_1__08_ ),
    .A2(u_multiplier_STAGE2_Full_adder_pp2_51_1__10_ ),
    .B1(u_multiplier_pp2_52 [2]),
    .B2(u_multiplier_STAGE2_Full_adder_pp2_51_1__09_ ),
    .ZN(u_multiplier_pp2_51 [0]));
 INV_X1 u_multiplier_STAGE2_Full_adder_pp2_53_1__12_  (.A(u_multiplier_STAGE2_pp2_52_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_53_1__08_ ));
 NAND3_X2 u_multiplier_STAGE2_Full_adder_pp2_53_1__13_  (.A1(u_multiplier_pp1_53 [5]),
    .A2(u_multiplier_pp1_53 [4]),
    .A3(u_multiplier_STAGE2_pp2_52_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_53_1__09_ ));
 NOR2_X2 u_multiplier_STAGE2_Full_adder_pp2_53_1__14_  (.A1(u_multiplier_pp1_53 [5]),
    .A2(u_multiplier_pp1_53 [4]),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_53_1__10_ ));
 AOI21_X1 u_multiplier_STAGE2_Full_adder_pp2_53_1__15_  (.A(u_multiplier_STAGE2_pp2_52_e42_2_cout ),
    .B1(u_multiplier_pp1_53 [4]),
    .B2(u_multiplier_pp1_53 [5]),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_53_1__11_ ));
 NOR2_X2 u_multiplier_STAGE2_Full_adder_pp2_53_1__16_  (.A1(u_multiplier_STAGE2_Full_adder_pp2_53_1__10_ ),
    .A2(u_multiplier_STAGE2_Full_adder_pp2_53_1__11_ ),
    .ZN(u_multiplier_pp2_54 [1]));
 AOI22_X4 u_multiplier_STAGE2_Full_adder_pp2_53_1__17_  (.A1(u_multiplier_STAGE2_Full_adder_pp2_53_1__08_ ),
    .A2(u_multiplier_STAGE2_Full_adder_pp2_53_1__10_ ),
    .B1(u_multiplier_pp2_54 [1]),
    .B2(u_multiplier_STAGE2_Full_adder_pp2_53_1__09_ ),
    .ZN(u_multiplier_pp2_53 [0]));
 INV_X1 u_multiplier_STAGE2_Full_adder_pp2_55_1__12_  (.A(u_multiplier_STAGE2_pp2_54_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_55_1__08_ ));
 NAND3_X2 u_multiplier_STAGE2_Full_adder_pp2_55_1__13_  (.A1(u_multiplier_pp1_55 [1]),
    .A2(u_multiplier_pp1_55 [0]),
    .A3(u_multiplier_STAGE2_pp2_54_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_55_1__09_ ));
 NOR2_X2 u_multiplier_STAGE2_Full_adder_pp2_55_1__14_  (.A1(u_multiplier_pp1_55 [1]),
    .A2(u_multiplier_pp1_55 [0]),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_55_1__10_ ));
 AOI21_X1 u_multiplier_STAGE2_Full_adder_pp2_55_1__15_  (.A(u_multiplier_STAGE2_pp2_54_e42_1_cout ),
    .B1(u_multiplier_pp1_55 [0]),
    .B2(u_multiplier_pp1_55 [1]),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_55_1__11_ ));
 NOR2_X2 u_multiplier_STAGE2_Full_adder_pp2_55_1__16_  (.A1(u_multiplier_STAGE2_Full_adder_pp2_55_1__10_ ),
    .A2(u_multiplier_STAGE2_Full_adder_pp2_55_1__11_ ),
    .ZN(u_multiplier_pp2_56 [0]));
 AOI22_X4 u_multiplier_STAGE2_Full_adder_pp2_55_1__17_  (.A1(u_multiplier_STAGE2_Full_adder_pp2_55_1__08_ ),
    .A2(u_multiplier_STAGE2_Full_adder_pp2_55_1__10_ ),
    .B1(u_multiplier_pp2_56 [0]),
    .B2(u_multiplier_STAGE2_Full_adder_pp2_55_1__09_ ),
    .ZN(u_multiplier_pp2_55 [0]));
 AND2_X1 u_multiplier_STAGE2_Half_adder_pp2_10_1__4_  (.A1(u_multiplier_pp1_10 [5]),
    .A2(u_multiplier_pp1_10 [4]),
    .ZN(u_multiplier_pp2_11 [2]));
 XOR2_X2 u_multiplier_STAGE2_Half_adder_pp2_10_1__5_  (.A(u_multiplier_pp1_10 [5]),
    .B(u_multiplier_pp1_10 [4]),
    .Z(u_multiplier_pp2_10 [0]));
 AND2_X1 u_multiplier_STAGE2_Half_adder_pp2_12_1__4_  (.A1(u_multiplier_pp1_12 [9]),
    .A2(u_multiplier_pp1_12 [8]),
    .ZN(u_multiplier_pp2_13 [3]));
 XOR2_X2 u_multiplier_STAGE2_Half_adder_pp2_12_1__5_  (.A(u_multiplier_pp1_12 [9]),
    .B(u_multiplier_pp1_12 [8]),
    .Z(u_multiplier_pp2_12 [0]));
 AND2_X1 u_multiplier_STAGE2_Half_adder_pp2_14_1__4_  (.A1(u_multiplier_pp1_14 [13]),
    .A2(u_multiplier_pp1_14 [12]),
    .ZN(u_multiplier_pp2_15 [4]));
 XOR2_X2 u_multiplier_STAGE2_Half_adder_pp2_14_1__5_  (.A(u_multiplier_pp1_14 [13]),
    .B(u_multiplier_pp1_14 [12]),
    .Z(u_multiplier_pp2_14 [0]));
 AND2_X1 u_multiplier_STAGE2_Half_adder_pp2_8_1__4_  (.A1(u_multiplier_pp1_8 [1]),
    .A2(u_multiplier_pp1_8 [0]),
    .ZN(u_multiplier_pp2_9 [1]));
 XOR2_X2 u_multiplier_STAGE2_Half_adder_pp2_8_1__5_  (.A(u_multiplier_pp1_8 [1]),
    .B(u_multiplier_pp1_8 [0]),
    .Z(u_multiplier_pp2_8 [0]));
 LOGIC0_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__55__140  (.Z(net140));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_10_1__18_  (.A(u_multiplier_STAGE3_pp3_9_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_10_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_10_1__19_  (.A1(u_multiplier_pp2_10 [1]),
    .A2(u_multiplier_pp2_10 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_10_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_10_1__20_  (.A(u_multiplier_pp2_10 [1]),
    .B(u_multiplier_pp2_10 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_10_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_10_1__21_  (.A1(u_multiplier_pp2_10 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_10_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_10_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_10_1__22_  (.A(u_multiplier_pp2_10 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_10_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_10_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_10_1__23_  (.A1(u_multiplier_pp2_10 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_10_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_10_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_10_1__24_  (.A(u_multiplier_pp2_10 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_10_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_10_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_10_1__25_  (.A(u_multiplier_STAGE3_pp3_9_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_10_1__16_ ),
    .ZN(u_multiplier_pp3_10 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_10_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_10_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_10_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_10_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_10_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_10_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_10_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_10_1__17_ ),
    .ZN(u_multiplier_pp3_11 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_10_2__18_  (.A(u_multiplier_STAGE3_pp3_9_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_10_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_10_2__19_  (.A1(u_multiplier_pp2_10 [5]),
    .A2(u_multiplier_pp2_10 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_10_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_10_2__20_  (.A(u_multiplier_pp2_10 [5]),
    .B(u_multiplier_pp2_10 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_10_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_10_2__21_  (.A1(u_multiplier_pp2_10 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_10_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_10_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_10_2__22_  (.A(u_multiplier_pp2_10 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_10_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_10_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_10_2__23_  (.A1(u_multiplier_pp2_10 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_10_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_10_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_10_2__24_  (.A(u_multiplier_pp2_10 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_10_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_10_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_10_2__25_  (.A(u_multiplier_STAGE3_pp3_9_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_10_2__16_ ),
    .ZN(u_multiplier_pp3_10 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_10_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_10_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_10_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_10_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_10_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_10_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_10_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_10_2__17_ ),
    .ZN(u_multiplier_pp3_11 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_11_1__18_  (.A(u_multiplier_STAGE3_pp3_10_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_11_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_11_1__19_  (.A1(u_multiplier_pp2_11 [1]),
    .A2(u_multiplier_pp2_11 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_11_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_11_1__20_  (.A(u_multiplier_pp2_11 [1]),
    .B(u_multiplier_pp2_11 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_11_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_11_1__21_  (.A1(u_multiplier_pp2_11 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_11_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_11_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_11_1__22_  (.A(u_multiplier_pp2_11 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_11_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_11_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_11_1__23_  (.A1(u_multiplier_pp2_11 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_11_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_11_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_11_1__24_  (.A(u_multiplier_pp2_11 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_11_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_11_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_11_1__25_  (.A(u_multiplier_STAGE3_pp3_10_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_11_1__16_ ),
    .ZN(u_multiplier_pp3_11 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_11_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_11_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_11_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_11_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_11_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_11_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_11_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_11_1__17_ ),
    .ZN(u_multiplier_pp3_12 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_11_2__18_  (.A(u_multiplier_STAGE3_pp3_10_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_11_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_11_2__19_  (.A1(u_multiplier_pp2_11 [5]),
    .A2(u_multiplier_pp2_11 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_11_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_11_2__20_  (.A(u_multiplier_pp2_11 [5]),
    .B(u_multiplier_pp2_11 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_11_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_11_2__21_  (.A1(u_multiplier_pp2_11 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_11_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_11_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_11_2__22_  (.A(u_multiplier_pp2_11 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_11_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_11_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_11_2__23_  (.A1(u_multiplier_pp2_11 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_11_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_11_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_11_2__24_  (.A(u_multiplier_pp2_11 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_11_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_11_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_11_2__25_  (.A(u_multiplier_STAGE3_pp3_10_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_11_2__16_ ),
    .ZN(u_multiplier_pp3_11 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_11_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_11_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_11_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_11_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_11_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_11_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_11_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_11_2__17_ ),
    .ZN(u_multiplier_pp3_12 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_12_1__18_  (.A(u_multiplier_STAGE3_pp3_11_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_12_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_12_1__19_  (.A1(u_multiplier_pp2_12 [1]),
    .A2(u_multiplier_pp2_12 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_12_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_12_1__20_  (.A(u_multiplier_pp2_12 [1]),
    .B(u_multiplier_pp2_12 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_12_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_12_1__21_  (.A1(u_multiplier_pp2_12 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_12_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_12_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_12_1__22_  (.A(u_multiplier_pp2_12 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_12_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_12_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_12_1__23_  (.A1(u_multiplier_pp2_12 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_12_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_12_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_12_1__24_  (.A(u_multiplier_pp2_12 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_12_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_12_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_12_1__25_  (.A(u_multiplier_STAGE3_pp3_11_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_12_1__16_ ),
    .ZN(u_multiplier_pp3_12 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_12_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_12_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_12_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_12_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_12_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_12_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_12_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_12_1__17_ ),
    .ZN(u_multiplier_pp3_13 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_12_2__18_  (.A(u_multiplier_STAGE3_pp3_11_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_12_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_12_2__19_  (.A1(u_multiplier_pp2_12 [5]),
    .A2(u_multiplier_pp2_12 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_12_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_12_2__20_  (.A(u_multiplier_pp2_12 [5]),
    .B(u_multiplier_pp2_12 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_12_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_12_2__21_  (.A1(u_multiplier_pp2_12 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_12_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_12_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_12_2__22_  (.A(u_multiplier_pp2_12 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_12_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_12_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_12_2__23_  (.A1(u_multiplier_pp2_12 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_12_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_12_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_12_2__24_  (.A(u_multiplier_pp2_12 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_12_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_12_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_12_2__25_  (.A(u_multiplier_STAGE3_pp3_11_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_12_2__16_ ),
    .ZN(u_multiplier_pp3_12 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_12_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_12_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_12_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_12_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_12_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_12_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_12_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_12_2__17_ ),
    .ZN(u_multiplier_pp3_13 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_13_1__18_  (.A(u_multiplier_STAGE3_pp3_12_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_13_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_13_1__19_  (.A1(u_multiplier_pp2_13 [1]),
    .A2(u_multiplier_pp2_13 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_13_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_13_1__20_  (.A(u_multiplier_pp2_13 [1]),
    .B(u_multiplier_pp2_13 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_13_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_13_1__21_  (.A1(u_multiplier_pp2_13 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_13_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_13_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_13_1__22_  (.A(u_multiplier_pp2_13 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_13_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_13_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_13_1__23_  (.A1(u_multiplier_pp2_13 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_13_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_13_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_13_1__24_  (.A(u_multiplier_pp2_13 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_13_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_13_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_13_1__25_  (.A(u_multiplier_STAGE3_pp3_12_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_13_1__16_ ),
    .ZN(u_multiplier_pp3_13 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_13_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_13_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_13_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_13_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_13_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_13_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_13_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_13_1__17_ ),
    .ZN(u_multiplier_pp3_14 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_13_2__18_  (.A(u_multiplier_STAGE3_pp3_12_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_13_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_13_2__19_  (.A1(u_multiplier_pp2_13 [5]),
    .A2(u_multiplier_pp2_13 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_13_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_13_2__20_  (.A(u_multiplier_pp2_13 [5]),
    .B(u_multiplier_pp2_13 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_13_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_13_2__21_  (.A1(u_multiplier_pp2_13 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_13_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_13_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_13_2__22_  (.A(u_multiplier_pp2_13 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_13_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_13_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_13_2__23_  (.A1(u_multiplier_pp2_13 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_13_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_13_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_13_2__24_  (.A(u_multiplier_pp2_13 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_13_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_13_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_13_2__25_  (.A(u_multiplier_STAGE3_pp3_12_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_13_2__16_ ),
    .ZN(u_multiplier_pp3_13 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_13_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_13_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_13_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_13_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_13_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_13_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_13_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_13_2__17_ ),
    .ZN(u_multiplier_pp3_14 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_14_1__18_  (.A(u_multiplier_STAGE3_pp3_13_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_14_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_14_1__19_  (.A1(u_multiplier_pp2_14 [1]),
    .A2(u_multiplier_pp2_14 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_14_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_14_1__20_  (.A(u_multiplier_pp2_14 [1]),
    .B(u_multiplier_pp2_14 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_14_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_14_1__21_  (.A1(u_multiplier_pp2_14 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_14_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_14_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_14_1__22_  (.A(u_multiplier_pp2_14 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_14_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_14_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_14_1__23_  (.A1(u_multiplier_pp2_14 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_14_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_14_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_14_1__24_  (.A(u_multiplier_pp2_14 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_14_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_14_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_14_1__25_  (.A(u_multiplier_STAGE3_pp3_13_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_14_1__16_ ),
    .ZN(u_multiplier_pp3_14 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_14_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_14_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_14_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_14_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_14_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_14_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_14_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_14_1__17_ ),
    .ZN(u_multiplier_pp3_15 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_14_2__18_  (.A(u_multiplier_STAGE3_pp3_13_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_14_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_14_2__19_  (.A1(u_multiplier_pp2_14 [5]),
    .A2(u_multiplier_pp2_14 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_14_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_14_2__20_  (.A(u_multiplier_pp2_14 [5]),
    .B(u_multiplier_pp2_14 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_14_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_14_2__21_  (.A1(u_multiplier_pp2_14 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_14_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_14_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_14_2__22_  (.A(u_multiplier_pp2_14 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_14_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_14_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_14_2__23_  (.A1(u_multiplier_pp2_14 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_14_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_14_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_14_2__24_  (.A(u_multiplier_pp2_14 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_14_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_14_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_14_2__25_  (.A(u_multiplier_STAGE3_pp3_13_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_14_2__16_ ),
    .ZN(u_multiplier_pp3_14 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_14_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_14_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_14_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_14_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_14_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_14_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_14_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_14_2__17_ ),
    .ZN(u_multiplier_pp3_15 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_15_1__18_  (.A(u_multiplier_STAGE3_pp3_14_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_15_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_15_1__19_  (.A1(u_multiplier_pp2_15 [1]),
    .A2(u_multiplier_pp2_15 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_15_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_15_1__20_  (.A(u_multiplier_pp2_15 [1]),
    .B(u_multiplier_pp2_15 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_15_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_15_1__21_  (.A1(u_multiplier_pp2_15 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_15_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_15_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_15_1__22_  (.A(u_multiplier_pp2_15 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_15_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_15_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_15_1__23_  (.A1(u_multiplier_pp2_15 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_15_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_15_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_15_1__24_  (.A(u_multiplier_pp2_15 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_15_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_15_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_15_1__25_  (.A(u_multiplier_STAGE3_pp3_14_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_15_1__16_ ),
    .ZN(u_multiplier_pp3_15 [1]));
 NAND2_X2 u_multiplier_STAGE3_E_4_2_pp3_15_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_15_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_15_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_15_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_15_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_15_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_15_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_15_1__17_ ),
    .ZN(u_multiplier_pp3_16 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_15_2__18_  (.A(u_multiplier_STAGE3_pp3_14_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_15_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_15_2__19_  (.A1(u_multiplier_pp2_15 [5]),
    .A2(u_multiplier_pp2_15 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_15_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_15_2__20_  (.A(u_multiplier_pp2_15 [5]),
    .B(u_multiplier_pp2_15 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_15_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_15_2__21_  (.A1(u_multiplier_pp2_15 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_15_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_15_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_15_2__22_  (.A(u_multiplier_pp2_15 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_15_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_15_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_15_2__23_  (.A1(u_multiplier_pp2_15 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_15_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_15_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_15_2__24_  (.A(u_multiplier_pp2_15 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_15_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_15_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_15_2__25_  (.A(u_multiplier_STAGE3_pp3_14_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_15_2__16_ ),
    .ZN(u_multiplier_pp3_15 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_15_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_15_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_15_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_15_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_15_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_15_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_15_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_15_2__17_ ),
    .ZN(u_multiplier_pp3_16 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_16_1__18_  (.A(u_multiplier_STAGE3_pp3_15_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_16_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_16_1__19_  (.A1(u_multiplier_pp2_16 [1]),
    .A2(u_multiplier_pp2_16 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_16_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_16_1__20_  (.A(u_multiplier_pp2_16 [1]),
    .B(u_multiplier_pp2_16 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_16_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_16_1__21_  (.A1(u_multiplier_pp2_16 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_16_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_16_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_16_1__22_  (.A(u_multiplier_pp2_16 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_16_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_16_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_16_1__23_  (.A1(u_multiplier_pp2_16 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_16_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_16_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_16_1__24_  (.A(u_multiplier_pp2_16 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_16_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_16_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_16_1__25_  (.A(u_multiplier_STAGE3_pp3_15_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_16_1__16_ ),
    .ZN(u_multiplier_pp3_16 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_16_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_16_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_16_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_16_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_16_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_16_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_16_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_16_1__17_ ),
    .ZN(u_multiplier_pp3_17 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_16_2__18_  (.A(u_multiplier_STAGE3_pp3_15_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_16_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_16_2__19_  (.A1(u_multiplier_pp2_16 [5]),
    .A2(u_multiplier_pp2_16 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_16_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_16_2__20_  (.A(u_multiplier_pp2_16 [5]),
    .B(u_multiplier_pp2_16 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_16_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_16_2__21_  (.A1(u_multiplier_pp2_16 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_16_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_16_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_16_2__22_  (.A(u_multiplier_pp2_16 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_16_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_16_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_16_2__23_  (.A1(u_multiplier_pp2_16 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_16_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_16_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_16_2__24_  (.A(u_multiplier_pp2_16 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_16_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_16_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_16_2__25_  (.A(u_multiplier_STAGE3_pp3_15_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_16_2__16_ ),
    .ZN(u_multiplier_pp3_16 [0]));
 NAND2_X2 u_multiplier_STAGE3_E_4_2_pp3_16_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_16_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_16_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_16_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_16_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_16_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_16_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_16_2__17_ ),
    .ZN(u_multiplier_pp3_17 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_17_1__18_  (.A(u_multiplier_STAGE3_pp3_16_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_17_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_17_1__19_  (.A1(u_multiplier_pp2_17 [1]),
    .A2(u_multiplier_pp2_17 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_17_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_17_1__20_  (.A(u_multiplier_pp2_17 [1]),
    .B(u_multiplier_pp2_17 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_17_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_17_1__21_  (.A1(u_multiplier_pp2_17 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_17_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_17_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_17_1__22_  (.A(u_multiplier_pp2_17 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_17_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_17_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_17_1__23_  (.A1(u_multiplier_pp2_17 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_17_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_17_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_17_1__24_  (.A(u_multiplier_pp2_17 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_17_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_17_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_17_1__25_  (.A(u_multiplier_STAGE3_pp3_16_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_17_1__16_ ),
    .ZN(u_multiplier_pp3_17 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_17_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_17_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_17_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_17_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_17_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_17_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_17_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_17_1__17_ ),
    .ZN(u_multiplier_pp3_18 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_17_2__18_  (.A(u_multiplier_STAGE3_pp3_16_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_17_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_17_2__19_  (.A1(u_multiplier_pp2_17 [5]),
    .A2(u_multiplier_pp2_17 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_17_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_17_2__20_  (.A(u_multiplier_pp2_17 [5]),
    .B(u_multiplier_pp2_17 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_17_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_17_2__21_  (.A1(u_multiplier_pp2_17 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_17_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_17_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_17_2__22_  (.A(u_multiplier_pp2_17 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_17_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_17_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_17_2__23_  (.A1(u_multiplier_pp2_17 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_17_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_17_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_17_2__24_  (.A(u_multiplier_pp2_17 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_17_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_17_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_17_2__25_  (.A(u_multiplier_STAGE3_pp3_16_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_17_2__16_ ),
    .ZN(u_multiplier_pp3_17 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_17_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_17_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_17_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_17_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_17_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_17_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_17_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_17_2__17_ ),
    .ZN(u_multiplier_pp3_18 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_18_1__18_  (.A(u_multiplier_STAGE3_pp3_17_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_18_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_18_1__19_  (.A1(u_multiplier_pp2_18 [1]),
    .A2(u_multiplier_pp2_18 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_18_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_18_1__20_  (.A(u_multiplier_pp2_18 [1]),
    .B(u_multiplier_pp2_18 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_18_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_18_1__21_  (.A1(u_multiplier_pp2_18 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_18_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_18_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_18_1__22_  (.A(u_multiplier_pp2_18 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_18_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_18_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_18_1__23_  (.A1(u_multiplier_pp2_18 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_18_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_18_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_18_1__24_  (.A(u_multiplier_pp2_18 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_18_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_18_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_18_1__25_  (.A(u_multiplier_STAGE3_pp3_17_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_18_1__16_ ),
    .ZN(u_multiplier_pp3_18 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_18_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_18_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_18_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_18_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_18_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_18_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_18_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_18_1__17_ ),
    .ZN(u_multiplier_pp3_19 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_18_2__18_  (.A(u_multiplier_STAGE3_pp3_17_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_18_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_18_2__19_  (.A1(u_multiplier_pp2_18 [5]),
    .A2(u_multiplier_pp2_18 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_18_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_18_2__20_  (.A(u_multiplier_pp2_18 [5]),
    .B(u_multiplier_pp2_18 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_18_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_18_2__21_  (.A1(u_multiplier_pp2_18 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_18_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_18_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_18_2__22_  (.A(u_multiplier_pp2_18 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_18_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_18_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_18_2__23_  (.A1(u_multiplier_pp2_18 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_18_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_18_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_18_2__24_  (.A(u_multiplier_pp2_18 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_18_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_18_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_18_2__25_  (.A(u_multiplier_STAGE3_pp3_17_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_18_2__16_ ),
    .ZN(u_multiplier_pp3_18 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_18_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_18_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_18_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_18_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_18_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_18_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_18_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_18_2__17_ ),
    .ZN(u_multiplier_pp3_19 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_19_1__18_  (.A(u_multiplier_STAGE3_pp3_18_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_19_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_19_1__19_  (.A1(u_multiplier_pp2_19 [1]),
    .A2(u_multiplier_pp2_19 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_19_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_19_1__20_  (.A(u_multiplier_pp2_19 [1]),
    .B(u_multiplier_pp2_19 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_19_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_19_1__21_  (.A1(u_multiplier_pp2_19 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_19_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_19_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_19_1__22_  (.A(u_multiplier_pp2_19 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_19_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_19_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_19_1__23_  (.A1(u_multiplier_pp2_19 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_19_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_19_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_19_1__24_  (.A(u_multiplier_pp2_19 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_19_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_19_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_19_1__25_  (.A(u_multiplier_STAGE3_pp3_18_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_19_1__16_ ),
    .ZN(u_multiplier_pp3_19 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_19_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_19_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_19_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_19_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_19_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_19_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_19_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_19_1__17_ ),
    .ZN(u_multiplier_pp3_20 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_19_2__18_  (.A(u_multiplier_STAGE3_pp3_18_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_19_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_19_2__19_  (.A1(u_multiplier_pp2_19 [5]),
    .A2(u_multiplier_pp2_19 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_19_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_19_2__20_  (.A(u_multiplier_pp2_19 [5]),
    .B(u_multiplier_pp2_19 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_19_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_19_2__21_  (.A1(u_multiplier_pp2_19 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_19_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_19_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_19_2__22_  (.A(u_multiplier_pp2_19 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_19_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_19_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_19_2__23_  (.A1(u_multiplier_pp2_19 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_19_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_19_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_19_2__24_  (.A(u_multiplier_pp2_19 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_19_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_19_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_19_2__25_  (.A(u_multiplier_STAGE3_pp3_18_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_19_2__16_ ),
    .ZN(u_multiplier_pp3_19 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_19_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_19_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_19_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_19_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_19_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_19_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_19_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_19_2__17_ ),
    .ZN(u_multiplier_pp3_20 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_20_1__18_  (.A(u_multiplier_STAGE3_pp3_19_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_20_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_20_1__19_  (.A1(u_multiplier_pp2_20 [1]),
    .A2(u_multiplier_pp2_20 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_20_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_20_1__20_  (.A(u_multiplier_pp2_20 [1]),
    .B(u_multiplier_pp2_20 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_20_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_20_1__21_  (.A1(u_multiplier_pp2_20 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_20_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_20_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_20_1__22_  (.A(u_multiplier_pp2_20 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_20_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_20_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_20_1__23_  (.A1(u_multiplier_pp2_20 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_20_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_20_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_20_1__24_  (.A(u_multiplier_pp2_20 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_20_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_20_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_20_1__25_  (.A(u_multiplier_STAGE3_pp3_19_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_20_1__16_ ),
    .ZN(u_multiplier_pp3_20 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_20_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_20_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_20_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_20_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_20_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_20_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_20_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_20_1__17_ ),
    .ZN(u_multiplier_pp3_21 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_20_2__18_  (.A(u_multiplier_STAGE3_pp3_19_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_20_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_20_2__19_  (.A1(u_multiplier_pp2_20 [5]),
    .A2(u_multiplier_pp2_20 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_20_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_20_2__20_  (.A(u_multiplier_pp2_20 [5]),
    .B(u_multiplier_pp2_20 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_20_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_20_2__21_  (.A1(u_multiplier_pp2_20 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_20_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_20_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_20_2__22_  (.A(u_multiplier_pp2_20 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_20_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_20_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_20_2__23_  (.A1(u_multiplier_pp2_20 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_20_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_20_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_20_2__24_  (.A(u_multiplier_pp2_20 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_20_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_20_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_20_2__25_  (.A(u_multiplier_STAGE3_pp3_19_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_20_2__16_ ),
    .ZN(u_multiplier_pp3_20 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_20_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_20_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_20_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_20_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_20_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_20_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_20_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_20_2__17_ ),
    .ZN(u_multiplier_pp3_21 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_21_1__18_  (.A(u_multiplier_STAGE3_pp3_20_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_21_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_21_1__19_  (.A1(u_multiplier_pp2_21 [1]),
    .A2(u_multiplier_pp2_21 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_21_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_21_1__20_  (.A(u_multiplier_pp2_21 [1]),
    .B(u_multiplier_pp2_21 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_21_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_21_1__21_  (.A1(u_multiplier_pp2_21 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_21_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_21_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_21_1__22_  (.A(u_multiplier_pp2_21 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_21_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_21_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_21_1__23_  (.A1(u_multiplier_pp2_21 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_21_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_21_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_21_1__24_  (.A(u_multiplier_pp2_21 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_21_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_21_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_21_1__25_  (.A(u_multiplier_STAGE3_pp3_20_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_21_1__16_ ),
    .ZN(u_multiplier_pp3_21 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_21_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_21_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_21_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_21_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_21_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_21_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_21_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_21_1__17_ ),
    .ZN(u_multiplier_pp3_22 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_21_2__18_  (.A(u_multiplier_STAGE3_pp3_20_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_21_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_21_2__19_  (.A1(u_multiplier_pp2_21 [5]),
    .A2(u_multiplier_pp2_21 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_21_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_21_2__20_  (.A(u_multiplier_pp2_21 [5]),
    .B(u_multiplier_pp2_21 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_21_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_21_2__21_  (.A1(u_multiplier_pp2_21 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_21_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_21_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_21_2__22_  (.A(u_multiplier_pp2_21 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_21_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_21_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_21_2__23_  (.A1(u_multiplier_pp2_21 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_21_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_21_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_21_2__24_  (.A(u_multiplier_pp2_21 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_21_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_21_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_21_2__25_  (.A(u_multiplier_STAGE3_pp3_20_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_21_2__16_ ),
    .ZN(u_multiplier_pp3_21 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_21_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_21_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_21_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_21_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_21_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_21_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_21_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_21_2__17_ ),
    .ZN(u_multiplier_pp3_22 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_22_1__18_  (.A(u_multiplier_STAGE3_pp3_21_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_22_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_22_1__19_  (.A1(u_multiplier_pp2_22 [1]),
    .A2(u_multiplier_pp2_22 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_22_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_22_1__20_  (.A(u_multiplier_pp2_22 [1]),
    .B(u_multiplier_pp2_22 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_22_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_22_1__21_  (.A1(u_multiplier_pp2_22 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_22_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_22_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_22_1__22_  (.A(u_multiplier_pp2_22 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_22_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_22_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_22_1__23_  (.A1(u_multiplier_pp2_22 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_22_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_22_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_22_1__24_  (.A(u_multiplier_pp2_22 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_22_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_22_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_22_1__25_  (.A(u_multiplier_STAGE3_pp3_21_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_22_1__16_ ),
    .ZN(u_multiplier_pp3_22 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_22_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_22_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_22_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_22_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_22_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_22_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_22_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_22_1__17_ ),
    .ZN(u_multiplier_pp3_23 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_22_2__18_  (.A(u_multiplier_STAGE3_pp3_21_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_22_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_22_2__19_  (.A1(u_multiplier_pp2_22 [5]),
    .A2(u_multiplier_pp2_22 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_22_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_22_2__20_  (.A(u_multiplier_pp2_22 [5]),
    .B(u_multiplier_pp2_22 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_22_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_22_2__21_  (.A1(u_multiplier_pp2_22 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_22_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_22_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_22_2__22_  (.A(u_multiplier_pp2_22 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_22_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_22_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_22_2__23_  (.A1(u_multiplier_pp2_22 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_22_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_22_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_22_2__24_  (.A(u_multiplier_pp2_22 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_22_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_22_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_22_2__25_  (.A(u_multiplier_STAGE3_pp3_21_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_22_2__16_ ),
    .ZN(u_multiplier_pp3_22 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_22_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_22_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_22_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_22_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_22_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_22_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_22_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_22_2__17_ ),
    .ZN(u_multiplier_pp3_23 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_23_1__18_  (.A(u_multiplier_STAGE3_pp3_22_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_23_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_23_1__19_  (.A1(u_multiplier_pp2_23 [1]),
    .A2(u_multiplier_pp2_23 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_23_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_23_1__20_  (.A(u_multiplier_pp2_23 [1]),
    .B(u_multiplier_pp2_23 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_23_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_23_1__21_  (.A1(u_multiplier_pp2_23 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_23_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_23_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_23_1__22_  (.A(u_multiplier_pp2_23 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_23_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_23_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_23_1__23_  (.A1(u_multiplier_pp2_23 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_23_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_23_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_23_1__24_  (.A(u_multiplier_pp2_23 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_23_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_23_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_23_1__25_  (.A(u_multiplier_STAGE3_pp3_22_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_23_1__16_ ),
    .ZN(u_multiplier_pp3_23 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_23_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_23_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_23_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_23_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_23_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_23_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_23_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_23_1__17_ ),
    .ZN(u_multiplier_pp3_24 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_23_2__18_  (.A(u_multiplier_STAGE3_pp3_22_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_23_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_23_2__19_  (.A1(u_multiplier_pp2_23 [5]),
    .A2(u_multiplier_pp2_23 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_23_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_23_2__20_  (.A(u_multiplier_pp2_23 [5]),
    .B(u_multiplier_pp2_23 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_23_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_23_2__21_  (.A1(u_multiplier_pp2_23 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_23_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_23_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_23_2__22_  (.A(u_multiplier_pp2_23 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_23_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_23_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_23_2__23_  (.A1(u_multiplier_pp2_23 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_23_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_23_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_23_2__24_  (.A(u_multiplier_pp2_23 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_23_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_23_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_23_2__25_  (.A(u_multiplier_STAGE3_pp3_22_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_23_2__16_ ),
    .ZN(u_multiplier_pp3_23 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_23_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_23_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_23_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_23_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_23_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_23_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_23_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_23_2__17_ ),
    .ZN(u_multiplier_pp3_24 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_24_1__18_  (.A(u_multiplier_STAGE3_pp3_23_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_24_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_24_1__19_  (.A1(u_multiplier_pp2_24 [1]),
    .A2(u_multiplier_pp2_24 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_24_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_24_1__20_  (.A(u_multiplier_pp2_24 [1]),
    .B(u_multiplier_pp2_24 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_24_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_24_1__21_  (.A1(u_multiplier_pp2_24 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_24_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_24_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_24_1__22_  (.A(u_multiplier_pp2_24 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_24_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_24_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_24_1__23_  (.A1(u_multiplier_pp2_24 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_24_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_24_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_24_1__24_  (.A(u_multiplier_pp2_24 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_24_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_24_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_24_1__25_  (.A(u_multiplier_STAGE3_pp3_23_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_24_1__16_ ),
    .ZN(u_multiplier_pp3_24 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_24_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_24_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_24_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_24_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_24_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_24_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_24_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_24_1__17_ ),
    .ZN(u_multiplier_pp3_25 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_24_2__18_  (.A(u_multiplier_STAGE3_pp3_23_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_24_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_24_2__19_  (.A1(u_multiplier_pp2_24 [5]),
    .A2(u_multiplier_pp2_24 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_24_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_24_2__20_  (.A(u_multiplier_pp2_24 [5]),
    .B(u_multiplier_pp2_24 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_24_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_24_2__21_  (.A1(u_multiplier_pp2_24 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_24_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_24_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_24_2__22_  (.A(u_multiplier_pp2_24 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_24_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_24_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_24_2__23_  (.A1(u_multiplier_pp2_24 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_24_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_24_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_24_2__24_  (.A(u_multiplier_pp2_24 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_24_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_24_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_24_2__25_  (.A(u_multiplier_STAGE3_pp3_23_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_24_2__16_ ),
    .ZN(u_multiplier_pp3_24 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_24_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_24_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_24_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_24_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_24_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_24_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_24_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_24_2__17_ ),
    .ZN(u_multiplier_pp3_25 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_25_1__18_  (.A(u_multiplier_STAGE3_pp3_24_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_25_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_25_1__19_  (.A1(u_multiplier_pp2_25 [1]),
    .A2(u_multiplier_pp2_25 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_25_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_25_1__20_  (.A(u_multiplier_pp2_25 [1]),
    .B(u_multiplier_pp2_25 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_25_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_25_1__21_  (.A1(u_multiplier_pp2_25 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_25_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_25_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_25_1__22_  (.A(u_multiplier_pp2_25 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_25_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_25_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_25_1__23_  (.A1(u_multiplier_pp2_25 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_25_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_25_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_25_1__24_  (.A(u_multiplier_pp2_25 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_25_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_25_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_25_1__25_  (.A(u_multiplier_STAGE3_pp3_24_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_25_1__16_ ),
    .ZN(u_multiplier_pp3_25 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_25_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_25_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_25_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_25_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_25_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_25_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_25_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_25_1__17_ ),
    .ZN(u_multiplier_pp3_26 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_25_2__18_  (.A(u_multiplier_STAGE3_pp3_24_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_25_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_25_2__19_  (.A1(u_multiplier_pp2_25 [5]),
    .A2(u_multiplier_pp2_25 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_25_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_25_2__20_  (.A(u_multiplier_pp2_25 [5]),
    .B(u_multiplier_pp2_25 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_25_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_25_2__21_  (.A1(u_multiplier_pp2_25 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_25_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_25_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_25_2__22_  (.A(u_multiplier_pp2_25 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_25_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_25_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_25_2__23_  (.A1(u_multiplier_pp2_25 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_25_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_25_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_25_2__24_  (.A(u_multiplier_pp2_25 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_25_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_25_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_25_2__25_  (.A(u_multiplier_STAGE3_pp3_24_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_25_2__16_ ),
    .ZN(u_multiplier_pp3_25 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_25_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_25_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_25_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_25_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_25_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_25_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_25_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_25_2__17_ ),
    .ZN(u_multiplier_pp3_26 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_26_1__18_  (.A(u_multiplier_STAGE3_pp3_25_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_26_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_26_1__19_  (.A1(u_multiplier_pp2_26 [1]),
    .A2(u_multiplier_pp2_26 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_26_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_26_1__20_  (.A(u_multiplier_pp2_26 [1]),
    .B(u_multiplier_pp2_26 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_26_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_26_1__21_  (.A1(u_multiplier_pp2_26 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_26_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_26_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_26_1__22_  (.A(u_multiplier_pp2_26 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_26_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_26_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_26_1__23_  (.A1(u_multiplier_pp2_26 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_26_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_26_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_26_1__24_  (.A(u_multiplier_pp2_26 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_26_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_26_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_26_1__25_  (.A(u_multiplier_STAGE3_pp3_25_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_26_1__16_ ),
    .ZN(u_multiplier_pp3_26 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_26_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_26_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_26_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_26_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_26_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_26_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_26_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_26_1__17_ ),
    .ZN(u_multiplier_pp3_27 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_26_2__18_  (.A(u_multiplier_STAGE3_pp3_25_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_26_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_26_2__19_  (.A1(u_multiplier_pp2_26 [5]),
    .A2(u_multiplier_pp2_26 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_26_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_26_2__20_  (.A(u_multiplier_pp2_26 [5]),
    .B(u_multiplier_pp2_26 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_26_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_26_2__21_  (.A1(u_multiplier_pp2_26 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_26_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_26_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_26_2__22_  (.A(u_multiplier_pp2_26 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_26_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_26_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_26_2__23_  (.A1(u_multiplier_pp2_26 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_26_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_26_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_26_2__24_  (.A(u_multiplier_pp2_26 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_26_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_26_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_26_2__25_  (.A(u_multiplier_STAGE3_pp3_25_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_26_2__16_ ),
    .ZN(u_multiplier_pp3_26 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_26_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_26_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_26_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_26_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_26_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_26_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_26_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_26_2__17_ ),
    .ZN(u_multiplier_pp3_27 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_27_1__18_  (.A(u_multiplier_STAGE3_pp3_26_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_27_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_27_1__19_  (.A1(u_multiplier_pp2_27 [1]),
    .A2(u_multiplier_pp2_27 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_27_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_27_1__20_  (.A(u_multiplier_pp2_27 [1]),
    .B(u_multiplier_pp2_27 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_27_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_27_1__21_  (.A1(u_multiplier_pp2_27 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_27_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_27_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_27_1__22_  (.A(u_multiplier_pp2_27 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_27_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_27_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_27_1__23_  (.A1(u_multiplier_pp2_27 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_27_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_27_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_27_1__24_  (.A(u_multiplier_pp2_27 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_27_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_27_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_27_1__25_  (.A(u_multiplier_STAGE3_pp3_26_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_27_1__16_ ),
    .ZN(u_multiplier_pp3_27 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_27_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_27_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_27_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_27_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_27_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_27_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_27_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_27_1__17_ ),
    .ZN(u_multiplier_pp3_28 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_27_2__18_  (.A(u_multiplier_STAGE3_pp3_26_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_27_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_27_2__19_  (.A1(u_multiplier_pp2_27 [5]),
    .A2(u_multiplier_pp2_27 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_27_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_27_2__20_  (.A(u_multiplier_pp2_27 [5]),
    .B(u_multiplier_pp2_27 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_27_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_27_2__21_  (.A1(u_multiplier_pp2_27 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_27_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_27_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_27_2__22_  (.A(u_multiplier_pp2_27 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_27_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_27_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_27_2__23_  (.A1(u_multiplier_pp2_27 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_27_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_27_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_27_2__24_  (.A(u_multiplier_pp2_27 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_27_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_27_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_27_2__25_  (.A(u_multiplier_STAGE3_pp3_26_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_27_2__16_ ),
    .ZN(u_multiplier_pp3_27 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_27_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_27_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_27_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_27_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_27_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_27_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_27_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_27_2__17_ ),
    .ZN(u_multiplier_pp3_28 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_28_1__18_  (.A(u_multiplier_STAGE3_pp3_27_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_28_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_28_1__19_  (.A1(u_multiplier_pp2_28 [1]),
    .A2(u_multiplier_pp2_28 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_28_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_28_1__20_  (.A(u_multiplier_pp2_28 [1]),
    .B(u_multiplier_pp2_28 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_28_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_28_1__21_  (.A1(u_multiplier_pp2_28 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_28_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_28_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_28_1__22_  (.A(u_multiplier_pp2_28 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_28_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_28_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_28_1__23_  (.A1(u_multiplier_pp2_28 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_28_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_28_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_28_1__24_  (.A(u_multiplier_pp2_28 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_28_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_28_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_28_1__25_  (.A(u_multiplier_STAGE3_pp3_27_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_28_1__16_ ),
    .ZN(u_multiplier_pp3_28 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_28_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_28_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_28_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_28_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_28_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_28_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_28_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_28_1__17_ ),
    .ZN(u_multiplier_pp3_29 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_28_2__18_  (.A(u_multiplier_STAGE3_pp3_27_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_28_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_28_2__19_  (.A1(u_multiplier_pp2_28 [5]),
    .A2(u_multiplier_pp2_28 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_28_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_28_2__20_  (.A(u_multiplier_pp2_28 [5]),
    .B(u_multiplier_pp2_28 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_28_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_28_2__21_  (.A1(u_multiplier_pp2_28 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_28_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_28_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_28_2__22_  (.A(u_multiplier_pp2_28 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_28_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_28_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_28_2__23_  (.A1(u_multiplier_pp2_28 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_28_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_28_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_28_2__24_  (.A(u_multiplier_pp2_28 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_28_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_28_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_28_2__25_  (.A(u_multiplier_STAGE3_pp3_27_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_28_2__16_ ),
    .ZN(u_multiplier_pp3_28 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_28_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_28_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_28_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_28_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_28_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_28_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_28_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_28_2__17_ ),
    .ZN(u_multiplier_pp3_29 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_29_1__18_  (.A(u_multiplier_STAGE3_pp3_28_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_29_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_29_1__19_  (.A1(u_multiplier_pp2_29 [1]),
    .A2(u_multiplier_pp2_29 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_29_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_29_1__20_  (.A(u_multiplier_pp2_29 [1]),
    .B(u_multiplier_pp2_29 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_29_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_29_1__21_  (.A1(u_multiplier_pp2_29 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_29_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_29_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_29_1__22_  (.A(u_multiplier_pp2_29 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_29_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_29_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_29_1__23_  (.A1(u_multiplier_pp2_29 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_29_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_29_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_29_1__24_  (.A(u_multiplier_pp2_29 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_29_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_29_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_29_1__25_  (.A(u_multiplier_STAGE3_pp3_28_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_29_1__16_ ),
    .ZN(u_multiplier_pp3_29 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_29_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_29_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_29_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_29_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_29_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_29_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_29_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_29_1__17_ ),
    .ZN(u_multiplier_pp3_30 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_29_2__18_  (.A(u_multiplier_STAGE3_pp3_28_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_29_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_29_2__19_  (.A1(u_multiplier_pp2_29 [5]),
    .A2(u_multiplier_pp2_29 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_29_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_29_2__20_  (.A(u_multiplier_pp2_29 [5]),
    .B(u_multiplier_pp2_29 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_29_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_29_2__21_  (.A1(u_multiplier_pp2_29 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_29_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_29_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_29_2__22_  (.A(u_multiplier_pp2_29 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_29_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_29_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_29_2__23_  (.A1(u_multiplier_pp2_29 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_29_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_29_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_29_2__24_  (.A(u_multiplier_pp2_29 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_29_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_29_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_29_2__25_  (.A(u_multiplier_STAGE3_pp3_28_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_29_2__16_ ),
    .ZN(u_multiplier_pp3_29 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_29_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_29_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_29_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_29_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_29_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_29_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_29_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_29_2__17_ ),
    .ZN(u_multiplier_pp3_30 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_30_1__18_  (.A(u_multiplier_STAGE3_pp3_29_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_30_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_30_1__19_  (.A1(u_multiplier_pp2_30 [1]),
    .A2(u_multiplier_pp2_30 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_30_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_30_1__20_  (.A(u_multiplier_pp2_30 [1]),
    .B(u_multiplier_pp2_30 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_30_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_30_1__21_  (.A1(u_multiplier_pp2_30 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_30_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_30_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_30_1__22_  (.A(u_multiplier_pp2_30 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_30_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_30_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_30_1__23_  (.A1(u_multiplier_pp2_30 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_30_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_30_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_30_1__24_  (.A(u_multiplier_pp2_30 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_30_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_30_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_30_1__25_  (.A(u_multiplier_STAGE3_pp3_29_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_30_1__16_ ),
    .ZN(u_multiplier_pp3_30 [1]));
 NAND2_X2 u_multiplier_STAGE3_E_4_2_pp3_30_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_30_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_30_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_30_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_30_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_30_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_30_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_30_1__17_ ),
    .ZN(u_multiplier_pp3_31 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_30_2__18_  (.A(u_multiplier_STAGE3_pp3_29_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_30_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_30_2__19_  (.A1(u_multiplier_pp2_30 [5]),
    .A2(u_multiplier_pp2_30 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_30_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_30_2__20_  (.A(u_multiplier_pp2_30 [5]),
    .B(u_multiplier_pp2_30 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_30_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_30_2__21_  (.A1(u_multiplier_pp2_30 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_30_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_30_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_30_2__22_  (.A(u_multiplier_pp2_30 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_30_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_30_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_30_2__23_  (.A1(u_multiplier_pp2_30 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_30_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_30_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_30_2__24_  (.A(u_multiplier_pp2_30 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_30_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_30_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_30_2__25_  (.A(u_multiplier_STAGE3_pp3_29_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_30_2__16_ ),
    .ZN(u_multiplier_pp3_30 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_30_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_30_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_30_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_30_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_30_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_30_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_30_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_30_2__17_ ),
    .ZN(u_multiplier_pp3_31 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_31_1__18_  (.A(u_multiplier_STAGE3_pp3_30_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_31_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_31_1__19_  (.A1(u_multiplier_pp2_31 [1]),
    .A2(u_multiplier_pp2_31 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_31_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_31_1__20_  (.A(u_multiplier_pp2_31 [1]),
    .B(u_multiplier_pp2_31 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_31_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_31_1__21_  (.A1(u_multiplier_pp2_31 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_31_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_31_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_31_1__22_  (.A(u_multiplier_pp2_31 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_31_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_31_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_31_1__23_  (.A1(u_multiplier_pp2_31 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_31_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_31_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_31_1__24_  (.A(u_multiplier_pp2_31 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_31_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_31_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_31_1__25_  (.A(u_multiplier_STAGE3_pp3_30_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_31_1__16_ ),
    .ZN(u_multiplier_pp3_31 [1]));
 NAND2_X2 u_multiplier_STAGE3_E_4_2_pp3_31_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_31_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_31_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_31_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_31_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_31_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_31_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_31_1__17_ ),
    .ZN(u_multiplier_pp3_32 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_31_2__18_  (.A(u_multiplier_STAGE3_pp3_30_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_31_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_31_2__19_  (.A1(u_multiplier_pp2_31 [5]),
    .A2(u_multiplier_pp2_31 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_31_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_31_2__20_  (.A(u_multiplier_pp2_31 [5]),
    .B(u_multiplier_pp2_31 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_31_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_31_2__21_  (.A1(u_multiplier_pp2_31 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_31_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_31_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_31_2__22_  (.A(u_multiplier_pp2_31 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_31_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_31_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_31_2__23_  (.A1(u_multiplier_pp2_31 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_31_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_31_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_31_2__24_  (.A(u_multiplier_pp2_31 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_31_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_31_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_31_2__25_  (.A(u_multiplier_STAGE3_pp3_30_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_31_2__16_ ),
    .ZN(u_multiplier_pp3_31 [0]));
 NAND2_X2 u_multiplier_STAGE3_E_4_2_pp3_31_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_31_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_31_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_31_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_31_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_31_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_31_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_31_2__17_ ),
    .ZN(u_multiplier_pp3_32 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_32_1__18_  (.A(u_multiplier_STAGE3_pp3_31_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_32_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_32_1__19_  (.A1(u_multiplier_pp2_32 [1]),
    .A2(u_multiplier_pp2_32 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_32_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_32_1__20_  (.A(u_multiplier_pp2_32 [1]),
    .B(u_multiplier_pp2_32 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_32_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_32_1__21_  (.A1(u_multiplier_pp2_32 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_32_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_32_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_32_1__22_  (.A(u_multiplier_pp2_32 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_32_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_32_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_32_1__23_  (.A1(u_multiplier_pp2_32 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_32_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_32_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_32_1__24_  (.A(u_multiplier_pp2_32 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_32_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_32_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_32_1__25_  (.A(u_multiplier_STAGE3_pp3_31_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_32_1__16_ ),
    .ZN(u_multiplier_pp3_32 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_32_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_32_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_32_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_32_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_32_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_32_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_32_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_32_1__17_ ),
    .ZN(u_multiplier_pp3_33 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_32_2__18_  (.A(u_multiplier_STAGE3_pp3_31_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_32_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_32_2__19_  (.A1(u_multiplier_pp2_32 [5]),
    .A2(u_multiplier_pp2_32 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_32_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_32_2__20_  (.A(u_multiplier_pp2_32 [5]),
    .B(u_multiplier_pp2_32 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_32_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_32_2__21_  (.A1(u_multiplier_pp2_32 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_32_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_32_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_32_2__22_  (.A(u_multiplier_pp2_32 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_32_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_32_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_32_2__23_  (.A1(u_multiplier_pp2_32 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_32_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_32_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_32_2__24_  (.A(u_multiplier_pp2_32 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_32_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_32_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_32_2__25_  (.A(u_multiplier_STAGE3_pp3_31_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_32_2__16_ ),
    .ZN(u_multiplier_pp3_32 [0]));
 NAND2_X2 u_multiplier_STAGE3_E_4_2_pp3_32_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_32_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_32_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_32_e42_2_cout ));
 OAI21_X4 u_multiplier_STAGE3_E_4_2_pp3_32_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_32_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_32_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_32_2__17_ ),
    .ZN(u_multiplier_pp3_33 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_33_1__18_  (.A(u_multiplier_STAGE3_pp3_32_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_33_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_33_1__19_  (.A1(u_multiplier_pp2_33 [1]),
    .A2(u_multiplier_pp2_33 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_33_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_33_1__20_  (.A(u_multiplier_pp2_33 [1]),
    .B(u_multiplier_pp2_33 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_33_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_33_1__21_  (.A1(u_multiplier_pp2_33 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_33_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_33_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_33_1__22_  (.A(u_multiplier_pp2_33 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_33_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_33_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_33_1__23_  (.A1(u_multiplier_pp2_33 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_33_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_33_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_33_1__24_  (.A(u_multiplier_pp2_33 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_33_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_33_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_33_1__25_  (.A(u_multiplier_STAGE3_pp3_32_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_33_1__16_ ),
    .ZN(u_multiplier_pp3_33 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_33_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_33_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_33_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_33_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_33_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_33_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_33_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_33_1__17_ ),
    .ZN(u_multiplier_pp3_34 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_33_2__18_  (.A(u_multiplier_STAGE3_pp3_32_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_33_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_33_2__19_  (.A1(u_multiplier_pp2_33 [5]),
    .A2(u_multiplier_pp2_33 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_33_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_33_2__20_  (.A(u_multiplier_pp2_33 [5]),
    .B(u_multiplier_pp2_33 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_33_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_33_2__21_  (.A1(u_multiplier_pp2_33 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_33_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_33_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_33_2__22_  (.A(u_multiplier_pp2_33 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_33_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_33_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_33_2__23_  (.A1(u_multiplier_pp2_33 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_33_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_33_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_33_2__24_  (.A(u_multiplier_pp2_33 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_33_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_33_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_33_2__25_  (.A(u_multiplier_STAGE3_pp3_32_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_33_2__16_ ),
    .ZN(u_multiplier_pp3_33 [0]));
 NAND2_X2 u_multiplier_STAGE3_E_4_2_pp3_33_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_33_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_33_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_33_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_33_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_33_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_33_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_33_2__17_ ),
    .ZN(u_multiplier_pp3_34 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_34_1__18_  (.A(u_multiplier_STAGE3_pp3_33_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_34_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_34_1__19_  (.A1(u_multiplier_pp2_34 [1]),
    .A2(u_multiplier_pp2_34 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_34_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_34_1__20_  (.A(u_multiplier_pp2_34 [1]),
    .B(u_multiplier_pp2_34 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_34_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_34_1__21_  (.A1(u_multiplier_pp2_34 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_34_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_34_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_34_1__22_  (.A(u_multiplier_pp2_34 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_34_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_34_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_34_1__23_  (.A1(u_multiplier_pp2_34 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_34_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_34_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_34_1__24_  (.A(u_multiplier_pp2_34 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_34_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_34_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_34_1__25_  (.A(u_multiplier_STAGE3_pp3_33_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_34_1__16_ ),
    .ZN(u_multiplier_pp3_34 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_34_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_34_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_34_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_34_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_34_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_34_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_34_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_34_1__17_ ),
    .ZN(u_multiplier_pp3_35 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_34_2__18_  (.A(u_multiplier_STAGE3_pp3_33_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_34_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_34_2__19_  (.A1(u_multiplier_pp2_34 [5]),
    .A2(u_multiplier_pp2_34 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_34_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_34_2__20_  (.A(u_multiplier_pp2_34 [5]),
    .B(u_multiplier_pp2_34 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_34_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_34_2__21_  (.A1(u_multiplier_pp2_34 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_34_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_34_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_34_2__22_  (.A(u_multiplier_pp2_34 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_34_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_34_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_34_2__23_  (.A1(u_multiplier_pp2_34 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_34_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_34_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_34_2__24_  (.A(u_multiplier_pp2_34 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_34_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_34_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_34_2__25_  (.A(u_multiplier_STAGE3_pp3_33_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_34_2__16_ ),
    .ZN(u_multiplier_pp3_34 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_34_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_34_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_34_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_34_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_34_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_34_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_34_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_34_2__17_ ),
    .ZN(u_multiplier_pp3_35 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_35_1__18_  (.A(u_multiplier_STAGE3_pp3_34_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_35_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_35_1__19_  (.A1(u_multiplier_pp2_35 [1]),
    .A2(u_multiplier_pp2_35 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_35_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_35_1__20_  (.A(u_multiplier_pp2_35 [1]),
    .B(u_multiplier_pp2_35 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_35_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_35_1__21_  (.A1(u_multiplier_pp2_35 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_35_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_35_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_35_1__22_  (.A(u_multiplier_pp2_35 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_35_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_35_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_35_1__23_  (.A1(u_multiplier_pp2_35 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_35_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_35_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_35_1__24_  (.A(u_multiplier_pp2_35 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_35_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_35_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_35_1__25_  (.A(u_multiplier_STAGE3_pp3_34_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_35_1__16_ ),
    .ZN(u_multiplier_pp3_35 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_35_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_35_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_35_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_35_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_35_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_35_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_35_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_35_1__17_ ),
    .ZN(u_multiplier_pp3_36 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_35_2__18_  (.A(u_multiplier_STAGE3_pp3_34_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_35_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_35_2__19_  (.A1(u_multiplier_pp2_35 [5]),
    .A2(u_multiplier_pp2_35 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_35_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_35_2__20_  (.A(u_multiplier_pp2_35 [5]),
    .B(u_multiplier_pp2_35 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_35_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_35_2__21_  (.A1(u_multiplier_pp2_35 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_35_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_35_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_35_2__22_  (.A(u_multiplier_pp2_35 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_35_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_35_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_35_2__23_  (.A1(u_multiplier_pp2_35 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_35_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_35_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_35_2__24_  (.A(u_multiplier_pp2_35 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_35_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_35_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_35_2__25_  (.A(u_multiplier_STAGE3_pp3_34_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_35_2__16_ ),
    .ZN(u_multiplier_pp3_35 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_35_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_35_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_35_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_35_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_35_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_35_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_35_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_35_2__17_ ),
    .ZN(u_multiplier_pp3_36 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_36_1__18_  (.A(u_multiplier_STAGE3_pp3_35_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_36_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_36_1__19_  (.A1(u_multiplier_pp2_36 [1]),
    .A2(u_multiplier_pp2_36 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_36_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_36_1__20_  (.A(u_multiplier_pp2_36 [1]),
    .B(u_multiplier_pp2_36 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_36_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_36_1__21_  (.A1(u_multiplier_pp2_36 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_36_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_36_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_36_1__22_  (.A(u_multiplier_pp2_36 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_36_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_36_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_36_1__23_  (.A1(u_multiplier_pp2_36 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_36_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_36_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_36_1__24_  (.A(u_multiplier_pp2_36 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_36_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_36_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_36_1__25_  (.A(u_multiplier_STAGE3_pp3_35_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_36_1__16_ ),
    .ZN(u_multiplier_pp3_36 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_36_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_36_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_36_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_36_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_36_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_36_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_36_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_36_1__17_ ),
    .ZN(u_multiplier_pp3_37 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_36_2__18_  (.A(u_multiplier_STAGE3_pp3_35_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_36_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_36_2__19_  (.A1(u_multiplier_pp2_36 [5]),
    .A2(u_multiplier_pp2_36 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_36_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_36_2__20_  (.A(u_multiplier_pp2_36 [5]),
    .B(u_multiplier_pp2_36 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_36_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_36_2__21_  (.A1(u_multiplier_pp2_36 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_36_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_36_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_36_2__22_  (.A(u_multiplier_pp2_36 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_36_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_36_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_36_2__23_  (.A1(u_multiplier_pp2_36 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_36_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_36_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_36_2__24_  (.A(u_multiplier_pp2_36 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_36_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_36_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_36_2__25_  (.A(u_multiplier_STAGE3_pp3_35_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_36_2__16_ ),
    .ZN(u_multiplier_pp3_36 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_36_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_36_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_36_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_36_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_36_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_36_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_36_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_36_2__17_ ),
    .ZN(u_multiplier_pp3_37 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_37_1__18_  (.A(u_multiplier_STAGE3_pp3_36_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_37_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_37_1__19_  (.A1(u_multiplier_pp2_37 [1]),
    .A2(u_multiplier_pp2_37 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_37_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_37_1__20_  (.A(u_multiplier_pp2_37 [1]),
    .B(u_multiplier_pp2_37 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_37_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_37_1__21_  (.A1(u_multiplier_pp2_37 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_37_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_37_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_37_1__22_  (.A(u_multiplier_pp2_37 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_37_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_37_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_37_1__23_  (.A1(u_multiplier_pp2_37 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_37_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_37_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_37_1__24_  (.A(u_multiplier_pp2_37 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_37_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_37_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_37_1__25_  (.A(u_multiplier_STAGE3_pp3_36_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_37_1__16_ ),
    .ZN(u_multiplier_pp3_37 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_37_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_37_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_37_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_37_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_37_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_37_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_37_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_37_1__17_ ),
    .ZN(u_multiplier_pp3_38 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_37_2__18_  (.A(u_multiplier_STAGE3_pp3_36_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_37_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_37_2__19_  (.A1(u_multiplier_pp2_37 [5]),
    .A2(u_multiplier_pp2_37 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_37_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_37_2__20_  (.A(u_multiplier_pp2_37 [5]),
    .B(u_multiplier_pp2_37 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_37_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_37_2__21_  (.A1(u_multiplier_pp2_37 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_37_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_37_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_37_2__22_  (.A(u_multiplier_pp2_37 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_37_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_37_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_37_2__23_  (.A1(u_multiplier_pp2_37 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_37_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_37_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_37_2__24_  (.A(u_multiplier_pp2_37 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_37_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_37_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_37_2__25_  (.A(u_multiplier_STAGE3_pp3_36_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_37_2__16_ ),
    .ZN(u_multiplier_pp3_37 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_37_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_37_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_37_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_37_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_37_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_37_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_37_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_37_2__17_ ),
    .ZN(u_multiplier_pp3_38 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_38_1__18_  (.A(u_multiplier_STAGE3_pp3_37_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_38_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_38_1__19_  (.A1(u_multiplier_pp2_38 [1]),
    .A2(u_multiplier_pp2_38 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_38_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_38_1__20_  (.A(u_multiplier_pp2_38 [1]),
    .B(u_multiplier_pp2_38 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_38_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_38_1__21_  (.A1(u_multiplier_pp2_38 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_38_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_38_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_38_1__22_  (.A(u_multiplier_pp2_38 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_38_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_38_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_38_1__23_  (.A1(u_multiplier_pp2_38 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_38_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_38_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_38_1__24_  (.A(u_multiplier_pp2_38 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_38_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_38_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_38_1__25_  (.A(u_multiplier_STAGE3_pp3_37_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_38_1__16_ ),
    .ZN(u_multiplier_pp3_38 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_38_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_38_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_38_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_38_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_38_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_38_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_38_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_38_1__17_ ),
    .ZN(u_multiplier_pp3_39 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_38_2__18_  (.A(u_multiplier_STAGE3_pp3_37_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_38_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_38_2__19_  (.A1(u_multiplier_pp2_38 [5]),
    .A2(u_multiplier_pp2_38 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_38_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_38_2__20_  (.A(u_multiplier_pp2_38 [5]),
    .B(u_multiplier_pp2_38 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_38_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_38_2__21_  (.A1(u_multiplier_pp2_38 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_38_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_38_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_38_2__22_  (.A(u_multiplier_pp2_38 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_38_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_38_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_38_2__23_  (.A1(u_multiplier_pp2_38 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_38_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_38_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_38_2__24_  (.A(u_multiplier_pp2_38 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_38_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_38_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_38_2__25_  (.A(u_multiplier_STAGE3_pp3_37_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_38_2__16_ ),
    .ZN(u_multiplier_pp3_38 [0]));
 NAND2_X2 u_multiplier_STAGE3_E_4_2_pp3_38_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_38_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_38_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_38_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_38_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_38_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_38_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_38_2__17_ ),
    .ZN(u_multiplier_pp3_39 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_39_1__18_  (.A(u_multiplier_STAGE3_pp3_38_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_39_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_39_1__19_  (.A1(u_multiplier_pp2_39 [1]),
    .A2(u_multiplier_pp2_39 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_39_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_39_1__20_  (.A(u_multiplier_pp2_39 [1]),
    .B(u_multiplier_pp2_39 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_39_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_39_1__21_  (.A1(u_multiplier_pp2_39 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_39_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_39_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_39_1__22_  (.A(u_multiplier_pp2_39 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_39_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_39_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_39_1__23_  (.A1(u_multiplier_pp2_39 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_39_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_39_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_39_1__24_  (.A(u_multiplier_pp2_39 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_39_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_39_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_39_1__25_  (.A(u_multiplier_STAGE3_pp3_38_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_39_1__16_ ),
    .ZN(u_multiplier_pp3_39 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_39_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_39_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_39_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_39_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_39_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_39_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_39_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_39_1__17_ ),
    .ZN(u_multiplier_pp3_40 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_39_2__18_  (.A(u_multiplier_STAGE3_pp3_38_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_39_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_39_2__19_  (.A1(u_multiplier_pp2_39 [5]),
    .A2(u_multiplier_pp2_39 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_39_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_39_2__20_  (.A(u_multiplier_pp2_39 [5]),
    .B(u_multiplier_pp2_39 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_39_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_39_2__21_  (.A1(u_multiplier_pp2_39 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_39_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_39_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_39_2__22_  (.A(u_multiplier_pp2_39 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_39_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_39_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_39_2__23_  (.A1(u_multiplier_pp2_39 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_39_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_39_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_39_2__24_  (.A(u_multiplier_pp2_39 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_39_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_39_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_39_2__25_  (.A(u_multiplier_STAGE3_pp3_38_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_39_2__16_ ),
    .ZN(u_multiplier_pp3_39 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_39_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_39_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_39_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_39_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_39_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_39_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_39_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_39_2__17_ ),
    .ZN(u_multiplier_pp3_40 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_40_1__18_  (.A(u_multiplier_STAGE3_pp3_39_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_40_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_40_1__19_  (.A1(u_multiplier_pp2_40 [1]),
    .A2(u_multiplier_pp2_40 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_40_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_40_1__20_  (.A(u_multiplier_pp2_40 [1]),
    .B(u_multiplier_pp2_40 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_40_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_40_1__21_  (.A1(u_multiplier_pp2_40 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_40_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_40_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_40_1__22_  (.A(u_multiplier_pp2_40 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_40_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_40_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_40_1__23_  (.A1(u_multiplier_pp2_40 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_40_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_40_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_40_1__24_  (.A(u_multiplier_pp2_40 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_40_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_40_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_40_1__25_  (.A(u_multiplier_STAGE3_pp3_39_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_40_1__16_ ),
    .ZN(u_multiplier_pp3_40 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_40_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_40_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_40_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_40_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_40_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_40_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_40_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_40_1__17_ ),
    .ZN(u_multiplier_pp3_41 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_40_2__18_  (.A(u_multiplier_STAGE3_pp3_39_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_40_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_40_2__19_  (.A1(u_multiplier_pp2_40 [5]),
    .A2(u_multiplier_pp2_40 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_40_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_40_2__20_  (.A(u_multiplier_pp2_40 [5]),
    .B(u_multiplier_pp2_40 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_40_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_40_2__21_  (.A1(u_multiplier_pp2_40 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_40_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_40_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_40_2__22_  (.A(u_multiplier_pp2_40 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_40_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_40_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_40_2__23_  (.A1(u_multiplier_pp2_40 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_40_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_40_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_40_2__24_  (.A(u_multiplier_pp2_40 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_40_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_40_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_40_2__25_  (.A(u_multiplier_STAGE3_pp3_39_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_40_2__16_ ),
    .ZN(u_multiplier_pp3_40 [0]));
 NAND2_X2 u_multiplier_STAGE3_E_4_2_pp3_40_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_40_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_40_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_40_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_40_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_40_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_40_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_40_2__17_ ),
    .ZN(u_multiplier_pp3_41 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_41_1__18_  (.A(u_multiplier_STAGE3_pp3_40_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_41_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_41_1__19_  (.A1(u_multiplier_pp2_41 [1]),
    .A2(u_multiplier_pp2_41 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_41_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_41_1__20_  (.A(u_multiplier_pp2_41 [1]),
    .B(u_multiplier_pp2_41 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_41_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_41_1__21_  (.A1(u_multiplier_pp2_41 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_41_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_41_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_41_1__22_  (.A(u_multiplier_pp2_41 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_41_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_41_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_41_1__23_  (.A1(u_multiplier_pp2_41 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_41_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_41_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_41_1__24_  (.A(u_multiplier_pp2_41 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_41_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_41_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_41_1__25_  (.A(u_multiplier_STAGE3_pp3_40_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_41_1__16_ ),
    .ZN(u_multiplier_pp3_41 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_41_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_41_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_41_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_41_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_41_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_41_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_41_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_41_1__17_ ),
    .ZN(u_multiplier_pp3_42 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_41_2__18_  (.A(u_multiplier_STAGE3_pp3_40_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_41_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_41_2__19_  (.A1(u_multiplier_pp2_41 [5]),
    .A2(u_multiplier_pp2_41 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_41_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_41_2__20_  (.A(u_multiplier_pp2_41 [5]),
    .B(u_multiplier_pp2_41 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_41_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_41_2__21_  (.A1(u_multiplier_pp2_41 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_41_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_41_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_41_2__22_  (.A(u_multiplier_pp2_41 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_41_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_41_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_41_2__23_  (.A1(u_multiplier_pp2_41 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_41_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_41_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_41_2__24_  (.A(u_multiplier_pp2_41 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_41_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_41_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_41_2__25_  (.A(u_multiplier_STAGE3_pp3_40_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_41_2__16_ ),
    .ZN(u_multiplier_pp3_41 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_41_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_41_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_41_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_41_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_41_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_41_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_41_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_41_2__17_ ),
    .ZN(u_multiplier_pp3_42 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_42_1__18_  (.A(u_multiplier_STAGE3_pp3_41_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_42_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_42_1__19_  (.A1(u_multiplier_pp2_42 [1]),
    .A2(u_multiplier_pp2_42 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_42_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_42_1__20_  (.A(u_multiplier_pp2_42 [1]),
    .B(u_multiplier_pp2_42 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_42_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_42_1__21_  (.A1(u_multiplier_pp2_42 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_42_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_42_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_42_1__22_  (.A(u_multiplier_pp2_42 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_42_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_42_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_42_1__23_  (.A1(u_multiplier_pp2_42 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_42_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_42_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_42_1__24_  (.A(u_multiplier_pp2_42 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_42_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_42_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_42_1__25_  (.A(u_multiplier_STAGE3_pp3_41_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_42_1__16_ ),
    .ZN(u_multiplier_pp3_42 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_42_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_42_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_42_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_42_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_42_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_42_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_42_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_42_1__17_ ),
    .ZN(u_multiplier_pp3_43 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_42_2__18_  (.A(u_multiplier_STAGE3_pp3_41_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_42_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_42_2__19_  (.A1(u_multiplier_pp2_42 [5]),
    .A2(u_multiplier_pp2_42 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_42_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_42_2__20_  (.A(u_multiplier_pp2_42 [5]),
    .B(u_multiplier_pp2_42 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_42_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_42_2__21_  (.A1(u_multiplier_pp2_42 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_42_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_42_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_42_2__22_  (.A(u_multiplier_pp2_42 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_42_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_42_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_42_2__23_  (.A1(u_multiplier_pp2_42 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_42_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_42_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_42_2__24_  (.A(u_multiplier_pp2_42 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_42_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_42_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_42_2__25_  (.A(u_multiplier_STAGE3_pp3_41_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_42_2__16_ ),
    .ZN(u_multiplier_pp3_42 [0]));
 NAND2_X2 u_multiplier_STAGE3_E_4_2_pp3_42_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_42_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_42_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_42_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_42_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_42_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_42_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_42_2__17_ ),
    .ZN(u_multiplier_pp3_43 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_43_1__18_  (.A(u_multiplier_STAGE3_pp3_42_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_43_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_43_1__19_  (.A1(u_multiplier_pp2_43 [1]),
    .A2(u_multiplier_pp2_43 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_43_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_43_1__20_  (.A(u_multiplier_pp2_43 [1]),
    .B(u_multiplier_pp2_43 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_43_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_43_1__21_  (.A1(u_multiplier_pp2_43 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_43_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_43_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_43_1__22_  (.A(u_multiplier_pp2_43 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_43_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_43_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_43_1__23_  (.A1(u_multiplier_pp2_43 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_43_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_43_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_43_1__24_  (.A(u_multiplier_pp2_43 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_43_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_43_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_43_1__25_  (.A(u_multiplier_STAGE3_pp3_42_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_43_1__16_ ),
    .ZN(u_multiplier_pp3_43 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_43_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_43_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_43_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_43_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_43_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_43_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_43_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_43_1__17_ ),
    .ZN(u_multiplier_pp3_44 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_43_2__18_  (.A(u_multiplier_STAGE3_pp3_42_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_43_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_43_2__19_  (.A1(u_multiplier_pp2_43 [5]),
    .A2(u_multiplier_pp2_43 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_43_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_43_2__20_  (.A(u_multiplier_pp2_43 [5]),
    .B(u_multiplier_pp2_43 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_43_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_43_2__21_  (.A1(u_multiplier_pp2_43 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_43_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_43_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_43_2__22_  (.A(u_multiplier_pp2_43 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_43_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_43_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_43_2__23_  (.A1(u_multiplier_pp2_43 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_43_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_43_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_43_2__24_  (.A(u_multiplier_pp2_43 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_43_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_43_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_43_2__25_  (.A(u_multiplier_STAGE3_pp3_42_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_43_2__16_ ),
    .ZN(u_multiplier_pp3_43 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_43_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_43_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_43_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_43_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_43_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_43_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_43_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_43_2__17_ ),
    .ZN(u_multiplier_pp3_44 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_44_1__18_  (.A(u_multiplier_STAGE3_pp3_43_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_44_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_44_1__19_  (.A1(u_multiplier_pp2_44 [1]),
    .A2(u_multiplier_pp2_44 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_44_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_44_1__20_  (.A(u_multiplier_pp2_44 [1]),
    .B(u_multiplier_pp2_44 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_44_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_44_1__21_  (.A1(u_multiplier_pp2_44 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_44_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_44_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_44_1__22_  (.A(u_multiplier_pp2_44 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_44_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_44_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_44_1__23_  (.A1(u_multiplier_pp2_44 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_44_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_44_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_44_1__24_  (.A(u_multiplier_pp2_44 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_44_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_44_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_44_1__25_  (.A(u_multiplier_STAGE3_pp3_43_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_44_1__16_ ),
    .ZN(u_multiplier_pp3_44 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_44_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_44_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_44_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_44_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_44_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_44_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_44_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_44_1__17_ ),
    .ZN(u_multiplier_pp3_45 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_44_2__18_  (.A(u_multiplier_STAGE3_pp3_43_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_44_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_44_2__19_  (.A1(u_multiplier_pp2_44 [5]),
    .A2(u_multiplier_pp2_44 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_44_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_44_2__20_  (.A(u_multiplier_pp2_44 [5]),
    .B(u_multiplier_pp2_44 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_44_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_44_2__21_  (.A1(u_multiplier_pp2_44 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_44_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_44_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_44_2__22_  (.A(u_multiplier_pp2_44 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_44_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_44_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_44_2__23_  (.A1(u_multiplier_pp2_44 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_44_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_44_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_44_2__24_  (.A(u_multiplier_pp2_44 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_44_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_44_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_44_2__25_  (.A(u_multiplier_STAGE3_pp3_43_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_44_2__16_ ),
    .ZN(u_multiplier_pp3_44 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_44_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_44_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_44_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_44_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_44_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_44_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_44_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_44_2__17_ ),
    .ZN(u_multiplier_pp3_45 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_45_1__18_  (.A(u_multiplier_STAGE3_pp3_44_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_45_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_45_1__19_  (.A1(u_multiplier_pp2_45 [1]),
    .A2(u_multiplier_pp2_45 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_45_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_45_1__20_  (.A(u_multiplier_pp2_45 [1]),
    .B(u_multiplier_pp2_45 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_45_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_45_1__21_  (.A1(u_multiplier_pp2_45 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_45_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_45_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_45_1__22_  (.A(u_multiplier_pp2_45 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_45_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_45_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_45_1__23_  (.A1(u_multiplier_pp2_45 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_45_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_45_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_45_1__24_  (.A(u_multiplier_pp2_45 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_45_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_45_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_45_1__25_  (.A(u_multiplier_STAGE3_pp3_44_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_45_1__16_ ),
    .ZN(u_multiplier_pp3_45 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_45_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_45_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_45_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_45_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_45_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_45_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_45_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_45_1__17_ ),
    .ZN(u_multiplier_pp3_46 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_45_2__18_  (.A(u_multiplier_STAGE3_pp3_44_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_45_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_45_2__19_  (.A1(u_multiplier_pp2_45 [5]),
    .A2(u_multiplier_pp2_45 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_45_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_45_2__20_  (.A(u_multiplier_pp2_45 [5]),
    .B(u_multiplier_pp2_45 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_45_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_45_2__21_  (.A1(u_multiplier_pp2_45 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_45_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_45_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_45_2__22_  (.A(u_multiplier_pp2_45 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_45_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_45_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_45_2__23_  (.A1(u_multiplier_pp2_45 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_45_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_45_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_45_2__24_  (.A(u_multiplier_pp2_45 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_45_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_45_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_45_2__25_  (.A(u_multiplier_STAGE3_pp3_44_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_45_2__16_ ),
    .ZN(u_multiplier_pp3_45 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_45_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_45_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_45_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_45_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_45_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_45_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_45_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_45_2__17_ ),
    .ZN(u_multiplier_pp3_46 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_46_1__18_  (.A(u_multiplier_STAGE3_pp3_45_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_46_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_46_1__19_  (.A1(u_multiplier_pp2_46 [1]),
    .A2(u_multiplier_pp2_46 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_46_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_46_1__20_  (.A(u_multiplier_pp2_46 [1]),
    .B(u_multiplier_pp2_46 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_46_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_46_1__21_  (.A1(u_multiplier_pp2_46 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_46_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_46_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_46_1__22_  (.A(u_multiplier_pp2_46 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_46_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_46_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_46_1__23_  (.A1(u_multiplier_pp2_46 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_46_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_46_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_46_1__24_  (.A(u_multiplier_pp2_46 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_46_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_46_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_46_1__25_  (.A(u_multiplier_STAGE3_pp3_45_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_46_1__16_ ),
    .ZN(u_multiplier_pp3_46 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_46_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_46_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_46_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_46_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_46_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_46_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_46_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_46_1__17_ ),
    .ZN(u_multiplier_pp3_47 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_46_2__18_  (.A(u_multiplier_STAGE3_pp3_45_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_46_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_46_2__19_  (.A1(u_multiplier_pp2_46 [5]),
    .A2(u_multiplier_pp2_46 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_46_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_46_2__20_  (.A(u_multiplier_pp2_46 [5]),
    .B(u_multiplier_pp2_46 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_46_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_46_2__21_  (.A1(u_multiplier_pp2_46 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_46_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_46_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_46_2__22_  (.A(u_multiplier_pp2_46 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_46_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_46_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_46_2__23_  (.A1(u_multiplier_pp2_46 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_46_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_46_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_46_2__24_  (.A(u_multiplier_pp2_46 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_46_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_46_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_46_2__25_  (.A(u_multiplier_STAGE3_pp3_45_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_46_2__16_ ),
    .ZN(u_multiplier_pp3_46 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_46_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_46_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_46_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_46_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_46_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_46_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_46_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_46_2__17_ ),
    .ZN(u_multiplier_pp3_47 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_47_1__18_  (.A(u_multiplier_STAGE3_pp3_46_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_47_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_47_1__19_  (.A1(u_multiplier_pp2_47 [1]),
    .A2(u_multiplier_pp2_47 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_47_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_47_1__20_  (.A(u_multiplier_pp2_47 [1]),
    .B(u_multiplier_pp2_47 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_47_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_47_1__21_  (.A1(u_multiplier_pp2_47 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_47_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_47_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_47_1__22_  (.A(u_multiplier_pp2_47 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_47_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_47_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_47_1__23_  (.A1(u_multiplier_pp2_47 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_47_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_47_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_47_1__24_  (.A(u_multiplier_pp2_47 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_47_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_47_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_47_1__25_  (.A(u_multiplier_STAGE3_pp3_46_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_47_1__16_ ),
    .ZN(u_multiplier_pp3_47 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_47_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_47_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_47_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_47_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_47_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_47_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_47_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_47_1__17_ ),
    .ZN(u_multiplier_pp3_48 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_47_2__18_  (.A(u_multiplier_STAGE3_pp3_46_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_47_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_47_2__19_  (.A1(u_multiplier_pp2_47 [5]),
    .A2(u_multiplier_pp2_47 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_47_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_47_2__20_  (.A(u_multiplier_pp2_47 [5]),
    .B(u_multiplier_pp2_47 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_47_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_47_2__21_  (.A1(u_multiplier_pp2_47 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_47_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_47_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_47_2__22_  (.A(u_multiplier_pp2_47 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_47_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_47_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_47_2__23_  (.A1(u_multiplier_pp2_47 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_47_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_47_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_47_2__24_  (.A(u_multiplier_pp2_47 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_47_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_47_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_47_2__25_  (.A(u_multiplier_STAGE3_pp3_46_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_47_2__16_ ),
    .ZN(u_multiplier_pp3_47 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_47_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_47_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_47_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_47_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_47_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_47_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_47_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_47_2__17_ ),
    .ZN(u_multiplier_pp3_48 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_48_1__18_  (.A(u_multiplier_STAGE3_pp3_47_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_48_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_48_1__19_  (.A1(u_multiplier_pp2_48 [1]),
    .A2(u_multiplier_pp2_48 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_48_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_48_1__20_  (.A(u_multiplier_pp2_48 [1]),
    .B(u_multiplier_pp2_48 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_48_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_48_1__21_  (.A1(u_multiplier_pp2_48 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_48_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_48_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_48_1__22_  (.A(u_multiplier_pp2_48 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_48_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_48_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_48_1__23_  (.A1(u_multiplier_pp2_48 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_48_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_48_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_48_1__24_  (.A(u_multiplier_pp2_48 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_48_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_48_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_48_1__25_  (.A(u_multiplier_STAGE3_pp3_47_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_48_1__16_ ),
    .ZN(u_multiplier_pp3_48 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_48_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_48_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_48_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_48_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_48_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_48_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_48_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_48_1__17_ ),
    .ZN(u_multiplier_pp3_49 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_48_2__18_  (.A(u_multiplier_STAGE3_pp3_47_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_48_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_48_2__19_  (.A1(u_multiplier_pp2_48 [5]),
    .A2(u_multiplier_pp2_48 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_48_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_48_2__20_  (.A(u_multiplier_pp2_48 [5]),
    .B(u_multiplier_pp2_48 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_48_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_48_2__21_  (.A1(u_multiplier_pp2_48 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_48_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_48_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_48_2__22_  (.A(u_multiplier_pp2_48 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_48_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_48_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_48_2__23_  (.A1(u_multiplier_pp2_48 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_48_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_48_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_48_2__24_  (.A(u_multiplier_pp2_48 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_48_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_48_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_48_2__25_  (.A(u_multiplier_STAGE3_pp3_47_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_48_2__16_ ),
    .ZN(u_multiplier_pp3_48 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_48_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_48_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_48_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_48_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_48_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_48_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_48_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_48_2__17_ ),
    .ZN(u_multiplier_pp3_49 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_49_1__18_  (.A(u_multiplier_STAGE3_pp3_48_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_49_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_49_1__19_  (.A1(u_multiplier_pp2_49 [1]),
    .A2(u_multiplier_pp2_49 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_49_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_49_1__20_  (.A(u_multiplier_pp2_49 [1]),
    .B(u_multiplier_pp2_49 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_49_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_49_1__21_  (.A1(u_multiplier_pp2_49 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_49_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_49_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_49_1__22_  (.A(u_multiplier_pp2_49 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_49_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_49_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_49_1__23_  (.A1(u_multiplier_pp2_49 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_49_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_49_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_49_1__24_  (.A(u_multiplier_pp2_49 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_49_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_49_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_49_1__25_  (.A(u_multiplier_STAGE3_pp3_48_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_49_1__16_ ),
    .ZN(u_multiplier_pp3_49 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_49_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_49_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_49_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_49_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_49_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_49_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_49_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_49_1__17_ ),
    .ZN(u_multiplier_pp3_50 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_49_2__18_  (.A(u_multiplier_STAGE3_pp3_48_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_49_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_49_2__19_  (.A1(u_multiplier_pp2_49 [5]),
    .A2(u_multiplier_pp2_49 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_49_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_49_2__20_  (.A(u_multiplier_pp2_49 [5]),
    .B(u_multiplier_pp2_49 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_49_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_49_2__21_  (.A1(u_multiplier_pp2_49 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_49_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_49_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_49_2__22_  (.A(u_multiplier_pp2_49 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_49_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_49_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_49_2__23_  (.A1(u_multiplier_pp2_49 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_49_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_49_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_49_2__24_  (.A(u_multiplier_pp2_49 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_49_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_49_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_49_2__25_  (.A(u_multiplier_STAGE3_pp3_48_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_49_2__16_ ),
    .ZN(u_multiplier_pp3_49 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_49_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_49_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_49_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_49_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_49_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_49_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_49_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_49_2__17_ ),
    .ZN(u_multiplier_pp3_50 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_50_1__18_  (.A(u_multiplier_STAGE3_pp3_49_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_50_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_50_1__19_  (.A1(u_multiplier_pp2_50 [1]),
    .A2(u_multiplier_pp2_50 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_50_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_50_1__20_  (.A(u_multiplier_pp2_50 [1]),
    .B(u_multiplier_pp2_50 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_50_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_50_1__21_  (.A1(u_multiplier_pp2_50 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_50_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_50_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_50_1__22_  (.A(u_multiplier_pp2_50 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_50_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_50_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_50_1__23_  (.A1(u_multiplier_pp2_50 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_50_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_50_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_50_1__24_  (.A(u_multiplier_pp2_50 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_50_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_50_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_50_1__25_  (.A(u_multiplier_STAGE3_pp3_49_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_50_1__16_ ),
    .ZN(u_multiplier_pp3_50 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_50_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_50_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_50_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_50_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_50_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_50_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_50_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_50_1__17_ ),
    .ZN(u_multiplier_pp3_51 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_50_2__18_  (.A(u_multiplier_STAGE3_pp3_49_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_50_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_50_2__19_  (.A1(u_multiplier_pp2_50 [5]),
    .A2(u_multiplier_pp2_50 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_50_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_50_2__20_  (.A(u_multiplier_pp2_50 [5]),
    .B(u_multiplier_pp2_50 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_50_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_50_2__21_  (.A1(u_multiplier_pp2_50 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_50_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_50_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_50_2__22_  (.A(u_multiplier_pp2_50 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_50_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_50_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_50_2__23_  (.A1(u_multiplier_pp2_50 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_50_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_50_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_50_2__24_  (.A(u_multiplier_pp2_50 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_50_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_50_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_50_2__25_  (.A(u_multiplier_STAGE3_pp3_49_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_50_2__16_ ),
    .ZN(u_multiplier_pp3_50 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_50_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_50_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_50_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_50_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_50_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_50_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_50_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_50_2__17_ ),
    .ZN(u_multiplier_pp3_51 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_51_1__18_  (.A(u_multiplier_STAGE3_pp3_50_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_51_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_51_1__19_  (.A1(u_multiplier_pp2_51 [1]),
    .A2(u_multiplier_pp2_51 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_51_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_51_1__20_  (.A(u_multiplier_pp2_51 [1]),
    .B(u_multiplier_pp2_51 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_51_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_51_1__21_  (.A1(u_multiplier_pp2_51 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_51_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_51_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_51_1__22_  (.A(u_multiplier_pp2_51 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_51_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_51_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_51_1__23_  (.A1(u_multiplier_pp2_51 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_51_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_51_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_51_1__24_  (.A(u_multiplier_pp2_51 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_51_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_51_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_51_1__25_  (.A(u_multiplier_STAGE3_pp3_50_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_51_1__16_ ),
    .ZN(u_multiplier_pp3_51 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_51_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_51_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_51_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_51_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_51_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_51_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_51_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_51_1__17_ ),
    .ZN(u_multiplier_pp3_52 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_51_2__18_  (.A(u_multiplier_STAGE3_pp3_50_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_51_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_51_2__19_  (.A1(u_multiplier_pp2_51 [5]),
    .A2(u_multiplier_pp2_51 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_51_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_51_2__20_  (.A(u_multiplier_pp2_51 [5]),
    .B(u_multiplier_pp2_51 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_51_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_51_2__21_  (.A1(u_multiplier_pp2_51 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_51_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_51_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_51_2__22_  (.A(u_multiplier_pp2_51 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_51_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_51_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_51_2__23_  (.A1(u_multiplier_pp2_51 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_51_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_51_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_51_2__24_  (.A(u_multiplier_pp2_51 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_51_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_51_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_51_2__25_  (.A(u_multiplier_STAGE3_pp3_50_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_51_2__16_ ),
    .ZN(u_multiplier_pp3_51 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_51_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_51_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_51_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_51_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_51_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_51_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_51_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_51_2__17_ ),
    .ZN(u_multiplier_pp3_52 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_52_1__18_  (.A(u_multiplier_STAGE3_pp3_51_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_52_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_52_1__19_  (.A1(u_multiplier_pp2_52 [1]),
    .A2(u_multiplier_pp2_52 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_52_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_52_1__20_  (.A(u_multiplier_pp2_52 [1]),
    .B(u_multiplier_pp2_52 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_52_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_52_1__21_  (.A1(u_multiplier_pp2_52 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_52_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_52_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_52_1__22_  (.A(u_multiplier_pp2_52 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_52_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_52_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_52_1__23_  (.A1(u_multiplier_pp2_52 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_52_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_52_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_52_1__24_  (.A(u_multiplier_pp2_52 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_52_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_52_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_52_1__25_  (.A(u_multiplier_STAGE3_pp3_51_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_52_1__16_ ),
    .ZN(u_multiplier_pp3_52 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_52_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_52_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_52_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_52_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_52_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_52_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_52_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_52_1__17_ ),
    .ZN(u_multiplier_pp3_53 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_52_2__18_  (.A(u_multiplier_STAGE3_pp3_51_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_52_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_52_2__19_  (.A1(u_multiplier_pp2_52 [5]),
    .A2(u_multiplier_pp2_52 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_52_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_52_2__20_  (.A(u_multiplier_pp2_52 [5]),
    .B(u_multiplier_pp2_52 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_52_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_52_2__21_  (.A1(u_multiplier_pp2_52 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_52_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_52_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_52_2__22_  (.A(u_multiplier_pp2_52 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_52_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_52_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_52_2__23_  (.A1(u_multiplier_pp2_52 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_52_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_52_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_52_2__24_  (.A(u_multiplier_pp2_52 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_52_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_52_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_52_2__25_  (.A(u_multiplier_STAGE3_pp3_51_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_52_2__16_ ),
    .ZN(u_multiplier_pp3_52 [0]));
 NAND2_X2 u_multiplier_STAGE3_E_4_2_pp3_52_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_52_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_52_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_52_e42_2_cout ));
 OAI21_X4 u_multiplier_STAGE3_E_4_2_pp3_52_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_52_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_52_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_52_2__17_ ),
    .ZN(u_multiplier_pp3_53 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_53_1__18_  (.A(u_multiplier_STAGE3_pp3_52_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_53_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_53_1__19_  (.A1(u_multiplier_pp2_53 [1]),
    .A2(u_multiplier_pp2_53 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_53_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_53_1__20_  (.A(u_multiplier_pp2_53 [1]),
    .B(u_multiplier_pp2_53 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_53_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_53_1__21_  (.A1(u_multiplier_pp2_53 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_53_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_53_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_53_1__22_  (.A(u_multiplier_pp2_53 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_53_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_53_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_53_1__23_  (.A1(u_multiplier_pp2_53 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_53_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_53_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_53_1__24_  (.A(u_multiplier_pp2_53 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_53_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_53_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_53_1__25_  (.A(u_multiplier_STAGE3_pp3_52_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_53_1__16_ ),
    .ZN(u_multiplier_pp3_53 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_53_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_53_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_53_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_53_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_53_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_53_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_53_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_53_1__17_ ),
    .ZN(u_multiplier_pp3_54 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_53_2__18_  (.A(u_multiplier_STAGE3_pp3_52_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_53_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_53_2__19_  (.A1(u_multiplier_pp2_53 [5]),
    .A2(u_multiplier_pp2_53 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_53_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_53_2__20_  (.A(u_multiplier_pp2_53 [5]),
    .B(u_multiplier_pp2_53 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_53_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_53_2__21_  (.A1(u_multiplier_pp2_53 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_53_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_53_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_53_2__22_  (.A(u_multiplier_pp2_53 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_53_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_53_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_53_2__23_  (.A1(u_multiplier_pp2_53 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_53_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_53_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_53_2__24_  (.A(u_multiplier_pp2_53 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_53_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_53_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_53_2__25_  (.A(u_multiplier_STAGE3_pp3_52_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_53_2__16_ ),
    .ZN(u_multiplier_pp3_53 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_53_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_53_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_53_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_53_e42_2_cout ));
 OAI21_X4 u_multiplier_STAGE3_E_4_2_pp3_53_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_53_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_53_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_53_2__17_ ),
    .ZN(u_multiplier_pp3_54 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_54_1__18_  (.A(u_multiplier_STAGE3_pp3_53_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_54_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_54_1__19_  (.A1(u_multiplier_pp2_54 [1]),
    .A2(u_multiplier_pp2_54 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_54_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_54_1__20_  (.A(u_multiplier_pp2_54 [1]),
    .B(u_multiplier_pp2_54 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_54_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_54_1__21_  (.A1(u_multiplier_pp2_54 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_54_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_54_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_54_1__22_  (.A(u_multiplier_pp2_54 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_54_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_54_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_54_1__23_  (.A1(u_multiplier_pp2_54 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_54_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_54_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_54_1__24_  (.A(u_multiplier_pp2_54 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_54_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_54_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_54_1__25_  (.A(u_multiplier_STAGE3_pp3_53_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_54_1__16_ ),
    .ZN(u_multiplier_pp3_54 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_54_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_54_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_54_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_54_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_54_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_54_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_54_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_54_1__17_ ),
    .ZN(u_multiplier_pp3_55 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_54_2__18_  (.A(u_multiplier_STAGE3_pp3_53_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_54_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_54_2__19_  (.A1(u_multiplier_pp2_54 [5]),
    .A2(u_multiplier_pp2_54 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_54_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_54_2__20_  (.A(u_multiplier_pp2_54 [5]),
    .B(u_multiplier_pp2_54 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_54_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_54_2__21_  (.A1(u_multiplier_pp2_54 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_54_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_54_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_54_2__22_  (.A(u_multiplier_pp2_54 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_54_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_54_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_54_2__23_  (.A1(u_multiplier_pp2_54 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_54_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_54_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_54_2__24_  (.A(u_multiplier_pp2_54 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_54_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_54_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_54_2__25_  (.A(u_multiplier_STAGE3_pp3_53_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_54_2__16_ ),
    .ZN(u_multiplier_pp3_54 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_54_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_54_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_54_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_54_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_54_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_54_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_54_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_54_2__17_ ),
    .ZN(u_multiplier_pp3_55 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_55_1__18_  (.A(u_multiplier_STAGE3_pp3_54_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_55_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_55_1__19_  (.A1(u_multiplier_pp2_55 [1]),
    .A2(u_multiplier_pp2_55 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_55_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_55_1__20_  (.A(u_multiplier_pp2_55 [1]),
    .B(u_multiplier_pp2_55 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_55_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_55_1__21_  (.A1(u_multiplier_pp2_55 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_55_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_55_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_55_1__22_  (.A(u_multiplier_pp2_55 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_55_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_55_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_55_1__23_  (.A1(u_multiplier_pp2_55 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_55_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_55_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_55_1__24_  (.A(u_multiplier_pp2_55 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_55_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_55_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_55_1__25_  (.A(u_multiplier_STAGE3_pp3_54_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_55_1__16_ ),
    .ZN(u_multiplier_pp3_55 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_55_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_55_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_55_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_55_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_55_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_55_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_55_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_55_1__17_ ),
    .ZN(u_multiplier_pp3_56 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_55_2__18_  (.A(u_multiplier_STAGE3_pp3_54_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_55_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_55_2__19_  (.A1(u_multiplier_pp2_55 [5]),
    .A2(u_multiplier_pp2_55 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_55_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_55_2__20_  (.A(u_multiplier_pp2_55 [5]),
    .B(u_multiplier_pp2_55 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_55_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_55_2__21_  (.A1(u_multiplier_pp2_55 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_55_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_55_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_55_2__22_  (.A(u_multiplier_pp2_55 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_55_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_55_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_55_2__23_  (.A1(u_multiplier_pp2_55 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_55_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_55_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_55_2__24_  (.A(u_multiplier_pp2_55 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_55_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_55_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_55_2__25_  (.A(u_multiplier_STAGE3_pp3_54_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_55_2__16_ ),
    .ZN(u_multiplier_pp3_55 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_55_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_55_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_55_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_55_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_55_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_55_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_55_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_55_2__17_ ),
    .ZN(u_multiplier_pp3_56 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_56_1__18_  (.A(u_multiplier_STAGE3_pp3_55_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_56_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_56_1__19_  (.A1(u_multiplier_pp2_56 [1]),
    .A2(u_multiplier_pp2_56 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_56_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_56_1__20_  (.A(u_multiplier_pp2_56 [1]),
    .B(u_multiplier_pp2_56 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_56_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_56_1__21_  (.A1(u_multiplier_pp2_56 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_56_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_56_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_56_1__22_  (.A(u_multiplier_pp2_56 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_56_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_56_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_56_1__23_  (.A1(u_multiplier_pp2_56 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_56_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_56_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_56_1__24_  (.A(u_multiplier_pp2_56 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_56_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_56_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_56_1__25_  (.A(u_multiplier_STAGE3_pp3_55_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_56_1__16_ ),
    .ZN(u_multiplier_pp3_56 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_56_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_56_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_56_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_56_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_56_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_56_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_56_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_56_1__17_ ),
    .ZN(u_multiplier_pp3_57 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_56_2__18_  (.A(u_multiplier_STAGE3_pp3_55_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_56_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_56_2__19_  (.A1(u_multiplier_pp2_56 [5]),
    .A2(u_multiplier_pp2_56 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_56_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_56_2__20_  (.A(u_multiplier_pp2_56 [5]),
    .B(u_multiplier_pp2_56 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_56_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_56_2__21_  (.A1(u_multiplier_pp2_56 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_56_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_56_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_56_2__22_  (.A(u_multiplier_pp2_56 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_56_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_56_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_56_2__23_  (.A1(u_multiplier_pp2_56 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_56_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_56_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_56_2__24_  (.A(u_multiplier_pp2_56 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_56_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_56_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_56_2__25_  (.A(u_multiplier_STAGE3_pp3_55_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_56_2__16_ ),
    .ZN(u_multiplier_pp3_56 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_56_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_56_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_56_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_56_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_56_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_56_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_56_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_56_2__17_ ),
    .ZN(u_multiplier_pp3_57 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_57_1__18_  (.A(u_multiplier_STAGE3_pp3_56_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_57_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_57_1__19_  (.A1(u_multiplier_pp2_57 [1]),
    .A2(u_multiplier_pp2_57 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_57_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_57_1__20_  (.A(u_multiplier_pp2_57 [1]),
    .B(u_multiplier_pp2_57 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_57_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_57_1__21_  (.A1(u_multiplier_pp2_57 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_57_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_57_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_57_1__22_  (.A(u_multiplier_pp2_57 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_57_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_57_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_57_1__23_  (.A1(u_multiplier_pp2_57 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_57_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_57_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_57_1__24_  (.A(u_multiplier_pp2_57 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_57_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_57_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_57_1__25_  (.A(u_multiplier_STAGE3_pp3_56_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_57_1__16_ ),
    .ZN(u_multiplier_pp3_57 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_57_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_57_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_57_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_57_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_57_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_57_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_57_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_57_1__17_ ),
    .ZN(u_multiplier_pp3_58 [1]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_58_1__18_  (.A(u_multiplier_STAGE3_pp3_57_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_58_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_58_1__19_  (.A1(u_multiplier_pp2_58 [1]),
    .A2(u_multiplier_pp2_58 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_58_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_58_1__20_  (.A(u_multiplier_pp2_58 [1]),
    .B(u_multiplier_pp2_58 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_58_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_58_1__21_  (.A1(u_multiplier_pp2_58 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_58_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_58_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_58_1__22_  (.A(u_multiplier_pp2_58 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_58_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_58_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_58_1__23_  (.A1(u_multiplier_pp2_58 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_58_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_58_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_58_1__24_  (.A(u_multiplier_pp2_58 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_58_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_58_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_58_1__25_  (.A(u_multiplier_STAGE3_pp3_57_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_58_1__16_ ),
    .ZN(u_multiplier_pp3_58 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_58_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_58_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_58_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_58_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_58_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_58_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_58_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_58_1__17_ ),
    .ZN(u_multiplier_pp3_59 [1]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_5_1__18_  (.A(net143),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_5_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_5_1__19_  (.A1(u_multiplier_pp2_5 [1]),
    .A2(u_multiplier_pp2_5 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_5_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_5_1__20_  (.A(u_multiplier_pp2_5 [1]),
    .B(u_multiplier_pp2_5 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_5_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_5_1__21_  (.A1(u_multiplier_pp2_5 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_5_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_5_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_5_1__22_  (.A(u_multiplier_pp2_5 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_5_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_5_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_5_1__23_  (.A1(u_multiplier_pp2_5 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_5_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_5_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_5_1__24_  (.A(u_multiplier_pp2_5 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_5_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_5_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_5_1__25_  (.A(net144),
    .B(u_multiplier_STAGE3_E_4_2_pp3_5_1__16_ ),
    .ZN(u_multiplier_pp3_5 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_5_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_5_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_5_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_5_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_5_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_5_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_5_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_5_1__17_ ),
    .ZN(u_multiplier_pp3_6 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_6_1__18_  (.A(u_multiplier_STAGE3_pp3_5_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_6_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_6_1__19_  (.A1(u_multiplier_pp2_6 [1]),
    .A2(u_multiplier_pp2_6 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_6_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_6_1__20_  (.A(u_multiplier_pp2_6 [1]),
    .B(u_multiplier_pp2_6 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_6_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_6_1__21_  (.A1(u_multiplier_pp2_6 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_6_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_6_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_6_1__22_  (.A(u_multiplier_pp2_6 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_6_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_6_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_6_1__23_  (.A1(u_multiplier_pp2_6 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_6_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_6_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_6_1__24_  (.A(u_multiplier_pp2_6 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_6_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_6_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_6_1__25_  (.A(u_multiplier_STAGE3_pp3_5_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_6_1__16_ ),
    .ZN(u_multiplier_pp3_6 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_6_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_6_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_6_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_6_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_6_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_6_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_6_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_6_1__17_ ),
    .ZN(u_multiplier_pp3_7 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_7_1__18_  (.A(u_multiplier_STAGE3_pp3_6_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_7_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_7_1__19_  (.A1(u_multiplier_pp2_7 [1]),
    .A2(u_multiplier_pp2_7 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_7_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_7_1__20_  (.A(u_multiplier_pp2_7 [1]),
    .B(u_multiplier_pp2_7 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_7_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_7_1__21_  (.A1(u_multiplier_pp2_7 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_7_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_7_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_7_1__22_  (.A(u_multiplier_pp2_7 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_7_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_7_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_7_1__23_  (.A1(u_multiplier_pp2_7 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_7_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_7_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_7_1__24_  (.A(u_multiplier_pp2_7 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_7_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_7_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_7_1__25_  (.A(u_multiplier_STAGE3_pp3_6_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_7_1__16_ ),
    .ZN(u_multiplier_pp3_7 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_7_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_7_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_7_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_7_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_7_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_7_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_7_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_7_1__17_ ),
    .ZN(u_multiplier_pp3_8 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_7_2__18_  (.A(net145),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_7_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_7_2__19_  (.A1(u_multiplier_pp2_7 [5]),
    .A2(u_multiplier_pp2_7 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_7_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_7_2__20_  (.A(u_multiplier_pp2_7 [5]),
    .B(u_multiplier_pp2_7 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_7_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_7_2__21_  (.A1(u_multiplier_pp2_7 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_7_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_7_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_7_2__22_  (.A(u_multiplier_pp2_7 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_7_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_7_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_7_2__23_  (.A1(u_multiplier_pp2_7 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_7_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_7_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_7_2__24_  (.A(u_multiplier_pp2_7 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_7_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_7_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_7_2__25_  (.A(net146),
    .B(u_multiplier_STAGE3_E_4_2_pp3_7_2__16_ ),
    .ZN(u_multiplier_pp3_7 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_7_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_7_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_7_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_7_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_7_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_7_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_7_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_7_2__17_ ),
    .ZN(u_multiplier_pp3_8 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_8_1__18_  (.A(u_multiplier_STAGE3_pp3_7_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_8_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_8_1__19_  (.A1(u_multiplier_pp2_8 [1]),
    .A2(u_multiplier_pp2_8 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_8_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_8_1__20_  (.A(u_multiplier_pp2_8 [1]),
    .B(u_multiplier_pp2_8 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_8_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_8_1__21_  (.A1(u_multiplier_pp2_8 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_8_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_8_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_8_1__22_  (.A(u_multiplier_pp2_8 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_8_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_8_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_8_1__23_  (.A1(u_multiplier_pp2_8 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_8_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_8_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_8_1__24_  (.A(u_multiplier_pp2_8 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_8_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_8_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_8_1__25_  (.A(u_multiplier_STAGE3_pp3_7_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_8_1__16_ ),
    .ZN(u_multiplier_pp3_8 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_8_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_8_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_8_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_8_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_8_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_8_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_8_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_8_1__17_ ),
    .ZN(u_multiplier_pp3_9 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_8_2__18_  (.A(u_multiplier_STAGE3_pp3_7_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_8_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_8_2__19_  (.A1(u_multiplier_pp2_8 [5]),
    .A2(u_multiplier_pp2_8 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_8_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_8_2__20_  (.A(u_multiplier_pp2_8 [5]),
    .B(u_multiplier_pp2_8 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_8_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_8_2__21_  (.A1(u_multiplier_pp2_8 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_8_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_8_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_8_2__22_  (.A(u_multiplier_pp2_8 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_8_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_8_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_8_2__23_  (.A1(u_multiplier_pp2_8 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_8_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_8_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_8_2__24_  (.A(u_multiplier_pp2_8 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_8_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_8_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_8_2__25_  (.A(u_multiplier_STAGE3_pp3_7_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_8_2__16_ ),
    .ZN(u_multiplier_pp3_8 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_8_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_8_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_8_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_8_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_8_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_8_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_8_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_8_2__17_ ),
    .ZN(u_multiplier_pp3_9 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_9_1__18_  (.A(u_multiplier_STAGE3_pp3_8_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_9_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_9_1__19_  (.A1(u_multiplier_pp2_9 [1]),
    .A2(u_multiplier_pp2_9 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_9_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_9_1__20_  (.A(u_multiplier_pp2_9 [1]),
    .B(u_multiplier_pp2_9 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_9_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_9_1__21_  (.A1(u_multiplier_pp2_9 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_9_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_9_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_9_1__22_  (.A(u_multiplier_pp2_9 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_9_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_9_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_9_1__23_  (.A1(u_multiplier_pp2_9 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_9_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_9_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_9_1__24_  (.A(u_multiplier_pp2_9 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_9_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_9_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_9_1__25_  (.A(u_multiplier_STAGE3_pp3_8_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_9_1__16_ ),
    .ZN(u_multiplier_pp3_9 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_9_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_9_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_9_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_9_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_9_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_9_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_9_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_9_1__17_ ),
    .ZN(u_multiplier_pp3_10 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_9_2__18_  (.A(u_multiplier_STAGE3_pp3_8_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_9_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_9_2__19_  (.A1(u_multiplier_pp2_9 [5]),
    .A2(u_multiplier_pp2_9 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_9_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_9_2__20_  (.A(u_multiplier_pp2_9 [5]),
    .B(u_multiplier_pp2_9 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_9_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_9_2__21_  (.A1(u_multiplier_pp2_9 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_9_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_9_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_9_2__22_  (.A(u_multiplier_pp2_9 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_9_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_9_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_9_2__23_  (.A1(u_multiplier_pp2_9 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_9_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_9_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_9_2__24_  (.A(u_multiplier_pp2_9 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_9_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_9_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_9_2__25_  (.A(u_multiplier_STAGE3_pp3_8_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_9_2__16_ ),
    .ZN(u_multiplier_pp3_9 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_9_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_9_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_9_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_9_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_9_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_9_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_9_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_9_2__17_ ),
    .ZN(u_multiplier_pp3_10 [2]));
 INV_X1 u_multiplier_STAGE3_Full_adder_pp3_57_1__12_  (.A(u_multiplier_STAGE3_pp3_56_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_Full_adder_pp3_57_1__08_ ));
 NAND3_X2 u_multiplier_STAGE3_Full_adder_pp3_57_1__13_  (.A1(u_multiplier_pp2_57 [5]),
    .A2(u_multiplier_pp2_57 [4]),
    .A3(u_multiplier_STAGE3_pp3_56_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_Full_adder_pp3_57_1__09_ ));
 NOR2_X2 u_multiplier_STAGE3_Full_adder_pp3_57_1__14_  (.A1(u_multiplier_pp2_57 [5]),
    .A2(u_multiplier_pp2_57 [4]),
    .ZN(u_multiplier_STAGE3_Full_adder_pp3_57_1__10_ ));
 AOI21_X1 u_multiplier_STAGE3_Full_adder_pp3_57_1__15_  (.A(u_multiplier_STAGE3_pp3_56_e42_2_cout ),
    .B1(u_multiplier_pp2_57 [4]),
    .B2(u_multiplier_pp2_57 [5]),
    .ZN(u_multiplier_STAGE3_Full_adder_pp3_57_1__11_ ));
 NOR2_X2 u_multiplier_STAGE3_Full_adder_pp3_57_1__16_  (.A1(u_multiplier_STAGE3_Full_adder_pp3_57_1__10_ ),
    .A2(u_multiplier_STAGE3_Full_adder_pp3_57_1__11_ ),
    .ZN(u_multiplier_pp3_58 [2]));
 AOI22_X4 u_multiplier_STAGE3_Full_adder_pp3_57_1__17_  (.A1(u_multiplier_STAGE3_Full_adder_pp3_57_1__08_ ),
    .A2(u_multiplier_STAGE3_Full_adder_pp3_57_1__10_ ),
    .B1(u_multiplier_pp3_58 [2]),
    .B2(u_multiplier_STAGE3_Full_adder_pp3_57_1__09_ ),
    .ZN(u_multiplier_pp3_57 [0]));
 INV_X1 u_multiplier_STAGE3_Full_adder_pp3_59_1__12_  (.A(u_multiplier_STAGE3_pp3_58_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_Full_adder_pp3_59_1__08_ ));
 NAND3_X2 u_multiplier_STAGE3_Full_adder_pp3_59_1__13_  (.A1(u_multiplier_pp2_59 [1]),
    .A2(u_multiplier_pp2_59 [0]),
    .A3(u_multiplier_STAGE3_pp3_58_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_Full_adder_pp3_59_1__09_ ));
 NOR2_X2 u_multiplier_STAGE3_Full_adder_pp3_59_1__14_  (.A1(u_multiplier_pp2_59 [1]),
    .A2(u_multiplier_pp2_59 [0]),
    .ZN(u_multiplier_STAGE3_Full_adder_pp3_59_1__10_ ));
 AOI21_X1 u_multiplier_STAGE3_Full_adder_pp3_59_1__15_  (.A(u_multiplier_STAGE3_pp3_58_e42_1_cout ),
    .B1(u_multiplier_pp2_59 [0]),
    .B2(u_multiplier_pp2_59 [1]),
    .ZN(u_multiplier_STAGE3_Full_adder_pp3_59_1__11_ ));
 NOR2_X2 u_multiplier_STAGE3_Full_adder_pp3_59_1__16_  (.A1(u_multiplier_STAGE3_Full_adder_pp3_59_1__10_ ),
    .A2(u_multiplier_STAGE3_Full_adder_pp3_59_1__11_ ),
    .ZN(u_multiplier_pp3_60 [0]));
 AOI22_X4 u_multiplier_STAGE3_Full_adder_pp3_59_1__17_  (.A1(u_multiplier_STAGE3_Full_adder_pp3_59_1__08_ ),
    .A2(u_multiplier_STAGE3_Full_adder_pp3_59_1__10_ ),
    .B1(u_multiplier_pp3_60 [0]),
    .B2(u_multiplier_STAGE3_Full_adder_pp3_59_1__09_ ),
    .ZN(u_multiplier_pp3_59 [0]));
 AND2_X1 u_multiplier_STAGE3_Half_adder_pp3_4_1__4_  (.A1(u_multiplier_pp2_4 [1]),
    .A2(u_multiplier_pp2_4 [0]),
    .ZN(u_multiplier_pp3_5 [1]));
 XOR2_X2 u_multiplier_STAGE3_Half_adder_pp3_4_1__5_  (.A(u_multiplier_pp2_4 [1]),
    .B(u_multiplier_pp2_4 [0]),
    .Z(u_multiplier_pp3_4 [0]));
 AND2_X1 u_multiplier_STAGE3_Half_adder_pp3_6_1__4_  (.A1(u_multiplier_pp2_6 [5]),
    .A2(u_multiplier_pp2_6 [4]),
    .ZN(u_multiplier_pp3_7 [2]));
 XOR2_X2 u_multiplier_STAGE3_Half_adder_pp3_6_1__5_  (.A(u_multiplier_pp2_6 [5]),
    .B(u_multiplier_pp2_6 [4]),
    .Z(u_multiplier_pp3_6 [0]));
 LOGIC0_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__40__147  (.Z(net147));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_10__18_  (.A(u_multiplier_STAGE4_pp4_9_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_10__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_10__19_  (.A1(u_multiplier_pp3_10 [1]),
    .A2(u_multiplier_pp3_10 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_10__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_10__20_  (.A(u_multiplier_pp3_10 [1]),
    .B(u_multiplier_pp3_10 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_10__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_10__21_  (.A1(u_multiplier_pp3_10 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_10__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_10__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_10__22_  (.A(u_multiplier_pp3_10 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_10__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_10__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_10__23_  (.A1(u_multiplier_pp3_10 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_10__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_10__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_10__24_  (.A(u_multiplier_pp3_10 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_10__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_10__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_10__25_  (.A(u_multiplier_STAGE4_pp4_9_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_10__16_ ),
    .ZN(u_multiplier_A [10]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_10__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_10__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_10__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_10_cout ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_10__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_10__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_10__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_10__17_ ),
    .ZN(u_multiplier_B [11]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_11__18_  (.A(u_multiplier_STAGE4_pp4_10_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_11__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_11__19_  (.A1(u_multiplier_pp3_11 [1]),
    .A2(u_multiplier_pp3_11 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_11__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_11__20_  (.A(u_multiplier_pp3_11 [1]),
    .B(u_multiplier_pp3_11 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_11__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_11__21_  (.A1(u_multiplier_pp3_11 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_11__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_11__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_11__22_  (.A(u_multiplier_pp3_11 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_11__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_11__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_11__23_  (.A1(u_multiplier_pp3_11 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_11__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_11__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_11__24_  (.A(u_multiplier_pp3_11 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_11__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_11__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_11__25_  (.A(u_multiplier_STAGE4_pp4_10_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_11__16_ ),
    .ZN(u_multiplier_A [11]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_11__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_11__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_11__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_11_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_11__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_11__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_11__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_11__17_ ),
    .ZN(u_multiplier_B [12]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_12__18_  (.A(u_multiplier_STAGE4_pp4_11_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_12__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_12__19_  (.A1(u_multiplier_pp3_12 [1]),
    .A2(u_multiplier_pp3_12 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_12__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_12__20_  (.A(u_multiplier_pp3_12 [1]),
    .B(u_multiplier_pp3_12 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_12__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_12__21_  (.A1(u_multiplier_pp3_12 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_12__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_12__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_12__22_  (.A(u_multiplier_pp3_12 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_12__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_12__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_12__23_  (.A1(u_multiplier_pp3_12 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_12__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_12__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_12__24_  (.A(u_multiplier_pp3_12 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_12__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_12__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_12__25_  (.A(u_multiplier_STAGE4_pp4_11_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_12__16_ ),
    .ZN(u_multiplier_A [12]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_12__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_12__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_12__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_12_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_12__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_12__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_12__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_12__17_ ),
    .ZN(u_multiplier_B [13]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_13__18_  (.A(u_multiplier_STAGE4_pp4_12_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_13__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_13__19_  (.A1(u_multiplier_pp3_13 [1]),
    .A2(u_multiplier_pp3_13 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_13__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_13__20_  (.A(u_multiplier_pp3_13 [1]),
    .B(u_multiplier_pp3_13 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_13__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_13__21_  (.A1(u_multiplier_pp3_13 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_13__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_13__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_13__22_  (.A(u_multiplier_pp3_13 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_13__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_13__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_13__23_  (.A1(u_multiplier_pp3_13 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_13__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_13__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_13__24_  (.A(u_multiplier_pp3_13 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_13__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_13__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_13__25_  (.A(u_multiplier_STAGE4_pp4_12_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_13__16_ ),
    .ZN(u_multiplier_A [13]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_13__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_13__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_13__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_13_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_13__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_13__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_13__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_13__17_ ),
    .ZN(u_multiplier_B [14]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_14__18_  (.A(u_multiplier_STAGE4_pp4_13_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_14__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_14__19_  (.A1(u_multiplier_pp3_14 [1]),
    .A2(u_multiplier_pp3_14 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_14__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_14__20_  (.A(u_multiplier_pp3_14 [1]),
    .B(u_multiplier_pp3_14 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_14__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_14__21_  (.A1(u_multiplier_pp3_14 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_14__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_14__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_14__22_  (.A(u_multiplier_pp3_14 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_14__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_14__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_14__23_  (.A1(u_multiplier_pp3_14 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_14__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_14__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_14__24_  (.A(u_multiplier_pp3_14 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_14__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_14__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_14__25_  (.A(u_multiplier_STAGE4_pp4_13_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_14__16_ ),
    .ZN(u_multiplier_A [14]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_14__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_14__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_14__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_14_cout ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_14__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_14__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_14__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_14__17_ ),
    .ZN(u_multiplier_B [15]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_15__18_  (.A(u_multiplier_STAGE4_pp4_14_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_15__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_15__19_  (.A1(u_multiplier_pp3_15 [1]),
    .A2(u_multiplier_pp3_15 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_15__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_15__20_  (.A(u_multiplier_pp3_15 [1]),
    .B(u_multiplier_pp3_15 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_15__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_15__21_  (.A1(u_multiplier_pp3_15 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_15__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_15__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_15__22_  (.A(u_multiplier_pp3_15 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_15__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_15__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_15__23_  (.A1(u_multiplier_pp3_15 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_15__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_15__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_15__24_  (.A(u_multiplier_pp3_15 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_15__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_15__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_15__25_  (.A(u_multiplier_STAGE4_pp4_14_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_15__16_ ),
    .ZN(u_multiplier_A [15]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_15__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_15__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_15__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_15_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_15__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_15__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_15__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_15__17_ ),
    .ZN(u_multiplier_B [16]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_16__18_  (.A(u_multiplier_STAGE4_pp4_15_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_16__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_16__19_  (.A1(u_multiplier_pp3_16 [1]),
    .A2(u_multiplier_pp3_16 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_16__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_16__20_  (.A(u_multiplier_pp3_16 [1]),
    .B(u_multiplier_pp3_16 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_16__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_16__21_  (.A1(u_multiplier_pp3_16 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_16__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_16__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_16__22_  (.A(u_multiplier_pp3_16 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_16__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_16__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_16__23_  (.A1(u_multiplier_pp3_16 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_16__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_16__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_16__24_  (.A(u_multiplier_pp3_16 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_16__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_16__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_16__25_  (.A(u_multiplier_STAGE4_pp4_15_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_16__16_ ),
    .ZN(u_multiplier_A [16]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_16__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_16__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_16__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_16_cout ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_16__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_16__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_16__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_16__17_ ),
    .ZN(u_multiplier_B [17]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_17__18_  (.A(u_multiplier_STAGE4_pp4_16_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_17__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_17__19_  (.A1(u_multiplier_pp3_17 [1]),
    .A2(u_multiplier_pp3_17 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_17__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_17__20_  (.A(u_multiplier_pp3_17 [1]),
    .B(u_multiplier_pp3_17 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_17__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_17__21_  (.A1(u_multiplier_pp3_17 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_17__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_17__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_17__22_  (.A(u_multiplier_pp3_17 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_17__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_17__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_17__23_  (.A1(u_multiplier_pp3_17 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_17__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_17__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_17__24_  (.A(u_multiplier_pp3_17 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_17__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_17__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_17__25_  (.A(u_multiplier_STAGE4_pp4_16_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_17__16_ ),
    .ZN(u_multiplier_A [17]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_17__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_17__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_17__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_17_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_17__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_17__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_17__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_17__17_ ),
    .ZN(u_multiplier_B [18]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_18__18_  (.A(u_multiplier_STAGE4_pp4_17_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_18__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_18__19_  (.A1(u_multiplier_pp3_18 [1]),
    .A2(u_multiplier_pp3_18 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_18__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_18__20_  (.A(u_multiplier_pp3_18 [1]),
    .B(u_multiplier_pp3_18 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_18__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_18__21_  (.A1(u_multiplier_pp3_18 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_18__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_18__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_18__22_  (.A(u_multiplier_pp3_18 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_18__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_18__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_18__23_  (.A1(u_multiplier_pp3_18 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_18__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_18__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_18__24_  (.A(u_multiplier_pp3_18 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_18__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_18__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_18__25_  (.A(u_multiplier_STAGE4_pp4_17_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_18__16_ ),
    .ZN(u_multiplier_A [18]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_18__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_18__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_18__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_18_cout ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_18__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_18__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_18__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_18__17_ ),
    .ZN(u_multiplier_B [19]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_19__18_  (.A(u_multiplier_STAGE4_pp4_18_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_19__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_19__19_  (.A1(u_multiplier_pp3_19 [1]),
    .A2(u_multiplier_pp3_19 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_19__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_19__20_  (.A(u_multiplier_pp3_19 [1]),
    .B(u_multiplier_pp3_19 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_19__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_19__21_  (.A1(u_multiplier_pp3_19 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_19__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_19__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_19__22_  (.A(u_multiplier_pp3_19 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_19__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_19__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_19__23_  (.A1(u_multiplier_pp3_19 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_19__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_19__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_19__24_  (.A(u_multiplier_pp3_19 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_19__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_19__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_19__25_  (.A(u_multiplier_STAGE4_pp4_18_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_19__16_ ),
    .ZN(u_multiplier_A [19]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_19__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_19__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_19__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_19_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_19__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_19__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_19__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_19__17_ ),
    .ZN(u_multiplier_B [20]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_2__18_  (.A(u_multiplier_STAGE4_pp4_1_ha_c ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_2__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_2__19_  (.A1(u_multiplier_pp3_2 [1]),
    .A2(u_multiplier_pp3_2 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_2__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_2__20_  (.A(u_multiplier_pp3_2 [1]),
    .B(u_multiplier_pp3_2 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_2__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_2__21_  (.A1(u_multiplier_pp3_2 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_2__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_2__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_2__22_  (.A(u_multiplier_pp3_2 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_2__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_2__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_2__23_  (.A1(net159),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_2__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_2__24_  (.A(net160),
    .B(u_multiplier_STAGE4_E_4_2_pp4_2__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_2__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_2__25_  (.A(u_multiplier_STAGE4_pp4_1_ha_c ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_2__16_ ),
    .ZN(u_multiplier_A [2]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_2__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_2__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_2__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_2_cout ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_2__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_2__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_2__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_2__17_ ),
    .ZN(u_multiplier_B [3]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_20__18_  (.A(u_multiplier_STAGE4_pp4_19_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_20__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_20__19_  (.A1(u_multiplier_pp3_20 [1]),
    .A2(u_multiplier_pp3_20 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_20__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_20__20_  (.A(u_multiplier_pp3_20 [1]),
    .B(u_multiplier_pp3_20 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_20__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_20__21_  (.A1(u_multiplier_pp3_20 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_20__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_20__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_20__22_  (.A(u_multiplier_pp3_20 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_20__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_20__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_20__23_  (.A1(u_multiplier_pp3_20 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_20__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_20__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_20__24_  (.A(u_multiplier_pp3_20 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_20__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_20__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_20__25_  (.A(u_multiplier_STAGE4_pp4_19_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_20__16_ ),
    .ZN(u_multiplier_A [20]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_20__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_20__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_20__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_20_cout ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_20__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_20__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_20__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_20__17_ ),
    .ZN(u_multiplier_B [21]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_21__18_  (.A(u_multiplier_STAGE4_pp4_20_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_21__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_21__19_  (.A1(u_multiplier_pp3_21 [1]),
    .A2(u_multiplier_pp3_21 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_21__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_21__20_  (.A(u_multiplier_pp3_21 [1]),
    .B(u_multiplier_pp3_21 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_21__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_21__21_  (.A1(u_multiplier_pp3_21 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_21__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_21__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_21__22_  (.A(u_multiplier_pp3_21 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_21__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_21__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_21__23_  (.A1(u_multiplier_pp3_21 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_21__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_21__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_21__24_  (.A(u_multiplier_pp3_21 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_21__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_21__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_21__25_  (.A(u_multiplier_STAGE4_pp4_20_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_21__16_ ),
    .ZN(u_multiplier_A [21]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_21__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_21__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_21__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_21_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_21__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_21__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_21__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_21__17_ ),
    .ZN(u_multiplier_B [22]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_22__18_  (.A(u_multiplier_STAGE4_pp4_21_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_22__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_22__19_  (.A1(u_multiplier_pp3_22 [1]),
    .A2(u_multiplier_pp3_22 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_22__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_22__20_  (.A(u_multiplier_pp3_22 [1]),
    .B(u_multiplier_pp3_22 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_22__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_22__21_  (.A1(u_multiplier_pp3_22 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_22__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_22__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_22__22_  (.A(u_multiplier_pp3_22 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_22__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_22__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_22__23_  (.A1(u_multiplier_pp3_22 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_22__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_22__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_22__24_  (.A(u_multiplier_pp3_22 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_22__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_22__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_22__25_  (.A(u_multiplier_STAGE4_pp4_21_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_22__16_ ),
    .ZN(u_multiplier_A [22]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_22__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_22__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_22__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_22_cout ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_22__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_22__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_22__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_22__17_ ),
    .ZN(u_multiplier_B [23]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_23__18_  (.A(u_multiplier_STAGE4_pp4_22_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_23__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_23__19_  (.A1(u_multiplier_pp3_23 [1]),
    .A2(u_multiplier_pp3_23 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_23__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_23__20_  (.A(u_multiplier_pp3_23 [1]),
    .B(u_multiplier_pp3_23 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_23__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_23__21_  (.A1(u_multiplier_pp3_23 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_23__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_23__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_23__22_  (.A(u_multiplier_pp3_23 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_23__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_23__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_23__23_  (.A1(u_multiplier_pp3_23 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_23__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_23__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_23__24_  (.A(u_multiplier_pp3_23 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_23__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_23__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_23__25_  (.A(u_multiplier_STAGE4_pp4_22_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_23__16_ ),
    .ZN(u_multiplier_A [23]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_23__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_23__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_23__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_23_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_23__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_23__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_23__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_23__17_ ),
    .ZN(u_multiplier_B [24]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_24__18_  (.A(u_multiplier_STAGE4_pp4_23_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_24__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_24__19_  (.A1(u_multiplier_pp3_24 [1]),
    .A2(u_multiplier_pp3_24 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_24__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_24__20_  (.A(u_multiplier_pp3_24 [1]),
    .B(u_multiplier_pp3_24 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_24__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_24__21_  (.A1(u_multiplier_pp3_24 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_24__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_24__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_24__22_  (.A(u_multiplier_pp3_24 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_24__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_24__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_24__23_  (.A1(u_multiplier_pp3_24 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_24__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_24__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_24__24_  (.A(u_multiplier_pp3_24 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_24__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_24__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_24__25_  (.A(u_multiplier_STAGE4_pp4_23_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_24__16_ ),
    .ZN(u_multiplier_A [24]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_24__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_24__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_24__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_24_cout ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_24__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_24__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_24__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_24__17_ ),
    .ZN(u_multiplier_B [25]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_25__18_  (.A(u_multiplier_STAGE4_pp4_24_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_25__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_25__19_  (.A1(u_multiplier_pp3_25 [1]),
    .A2(u_multiplier_pp3_25 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_25__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_25__20_  (.A(u_multiplier_pp3_25 [1]),
    .B(u_multiplier_pp3_25 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_25__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_25__21_  (.A1(u_multiplier_pp3_25 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_25__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_25__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_25__22_  (.A(u_multiplier_pp3_25 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_25__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_25__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_25__23_  (.A1(u_multiplier_pp3_25 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_25__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_25__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_25__24_  (.A(u_multiplier_pp3_25 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_25__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_25__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_25__25_  (.A(u_multiplier_STAGE4_pp4_24_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_25__16_ ),
    .ZN(u_multiplier_A [25]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_25__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_25__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_25__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_25_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_25__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_25__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_25__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_25__17_ ),
    .ZN(u_multiplier_B [26]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_26__18_  (.A(u_multiplier_STAGE4_pp4_25_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_26__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_26__19_  (.A1(u_multiplier_pp3_26 [1]),
    .A2(u_multiplier_pp3_26 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_26__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_26__20_  (.A(u_multiplier_pp3_26 [1]),
    .B(u_multiplier_pp3_26 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_26__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_26__21_  (.A1(u_multiplier_pp3_26 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_26__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_26__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_26__22_  (.A(u_multiplier_pp3_26 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_26__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_26__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_26__23_  (.A1(u_multiplier_pp3_26 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_26__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_26__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_26__24_  (.A(u_multiplier_pp3_26 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_26__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_26__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_26__25_  (.A(u_multiplier_STAGE4_pp4_25_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_26__16_ ),
    .ZN(u_multiplier_A [26]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_26__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_26__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_26__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_26_cout ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_26__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_26__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_26__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_26__17_ ),
    .ZN(u_multiplier_B [27]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_27__18_  (.A(u_multiplier_STAGE4_pp4_26_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_27__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_27__19_  (.A1(u_multiplier_pp3_27 [1]),
    .A2(u_multiplier_pp3_27 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_27__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_27__20_  (.A(u_multiplier_pp3_27 [1]),
    .B(u_multiplier_pp3_27 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_27__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_27__21_  (.A1(u_multiplier_pp3_27 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_27__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_27__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_27__22_  (.A(u_multiplier_pp3_27 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_27__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_27__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_27__23_  (.A1(u_multiplier_pp3_27 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_27__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_27__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_27__24_  (.A(u_multiplier_pp3_27 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_27__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_27__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_27__25_  (.A(u_multiplier_STAGE4_pp4_26_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_27__16_ ),
    .ZN(u_multiplier_A [27]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_27__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_27__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_27__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_27_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_27__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_27__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_27__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_27__17_ ),
    .ZN(u_multiplier_B [28]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_28__18_  (.A(u_multiplier_STAGE4_pp4_27_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_28__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_28__19_  (.A1(u_multiplier_pp3_28 [1]),
    .A2(u_multiplier_pp3_28 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_28__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_28__20_  (.A(u_multiplier_pp3_28 [1]),
    .B(u_multiplier_pp3_28 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_28__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_28__21_  (.A1(u_multiplier_pp3_28 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_28__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_28__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_28__22_  (.A(u_multiplier_pp3_28 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_28__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_28__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_28__23_  (.A1(u_multiplier_pp3_28 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_28__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_28__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_28__24_  (.A(u_multiplier_pp3_28 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_28__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_28__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_28__25_  (.A(u_multiplier_STAGE4_pp4_27_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_28__16_ ),
    .ZN(u_multiplier_A [28]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_28__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_28__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_28__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_28_cout ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_28__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_28__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_28__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_28__17_ ),
    .ZN(u_multiplier_B [29]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_29__18_  (.A(u_multiplier_STAGE4_pp4_28_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_29__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_29__19_  (.A1(u_multiplier_pp3_29 [1]),
    .A2(u_multiplier_pp3_29 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_29__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_29__20_  (.A(u_multiplier_pp3_29 [1]),
    .B(u_multiplier_pp3_29 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_29__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_29__21_  (.A1(u_multiplier_pp3_29 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_29__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_29__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_29__22_  (.A(u_multiplier_pp3_29 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_29__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_29__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_29__23_  (.A1(u_multiplier_pp3_29 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_29__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_29__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_29__24_  (.A(u_multiplier_pp3_29 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_29__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_29__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_29__25_  (.A(u_multiplier_STAGE4_pp4_28_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_29__16_ ),
    .ZN(u_multiplier_A [29]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_29__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_29__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_29__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_29_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_29__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_29__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_29__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_29__17_ ),
    .ZN(u_multiplier_B [30]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_3__18_  (.A(u_multiplier_STAGE4_pp4_2_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_3__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_3__19_  (.A1(u_multiplier_pp3_3 [1]),
    .A2(u_multiplier_pp3_3 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_3__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_3__20_  (.A(u_multiplier_pp3_3 [1]),
    .B(u_multiplier_pp3_3 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_3__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_3__21_  (.A1(u_multiplier_pp3_3 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_3__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_3__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_3__22_  (.A(u_multiplier_pp3_3 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_3__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_3__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_3__23_  (.A1(u_multiplier_pp3_3 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_3__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_3__24_  (.A(u_multiplier_pp3_3 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_3__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_3__25_  (.A(u_multiplier_STAGE4_pp4_2_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_3__16_ ),
    .ZN(u_multiplier_A [3]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_3__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_3__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_3__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_3_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_3__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_3__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_3__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_3__17_ ),
    .ZN(u_multiplier_B [4]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_30__18_  (.A(u_multiplier_STAGE4_pp4_29_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_30__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_30__19_  (.A1(u_multiplier_pp3_30 [1]),
    .A2(u_multiplier_pp3_30 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_30__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_30__20_  (.A(u_multiplier_pp3_30 [1]),
    .B(u_multiplier_pp3_30 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_30__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_30__21_  (.A1(u_multiplier_pp3_30 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_30__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_30__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_30__22_  (.A(u_multiplier_pp3_30 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_30__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_30__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_30__23_  (.A1(u_multiplier_pp3_30 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_30__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_30__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_30__24_  (.A(u_multiplier_pp3_30 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_30__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_30__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_30__25_  (.A(u_multiplier_STAGE4_pp4_29_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_30__16_ ),
    .ZN(u_multiplier_A [30]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_30__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_30__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_30__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_30_cout ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_30__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_30__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_30__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_30__17_ ),
    .ZN(u_multiplier_B [31]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_31__18_  (.A(u_multiplier_STAGE4_pp4_30_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_31__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_31__19_  (.A1(u_multiplier_pp3_31 [1]),
    .A2(u_multiplier_pp3_31 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_31__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_31__20_  (.A(u_multiplier_pp3_31 [1]),
    .B(u_multiplier_pp3_31 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_31__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_31__21_  (.A1(u_multiplier_pp3_31 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_31__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_31__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_31__22_  (.A(u_multiplier_pp3_31 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_31__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_31__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_31__23_  (.A1(u_multiplier_pp3_31 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_31__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_31__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_31__24_  (.A(u_multiplier_pp3_31 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_31__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_31__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_31__25_  (.A(u_multiplier_STAGE4_pp4_30_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_31__16_ ),
    .ZN(u_multiplier_A [31]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_31__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_31__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_31__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_31_cout ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_31__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_31__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_31__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_31__17_ ),
    .ZN(u_multiplier_B [32]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_32__18_  (.A(u_multiplier_STAGE4_pp4_31_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_32__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_32__19_  (.A1(u_multiplier_pp3_32 [1]),
    .A2(u_multiplier_pp3_32 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_32__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_32__20_  (.A(u_multiplier_pp3_32 [1]),
    .B(u_multiplier_pp3_32 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_32__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_32__21_  (.A1(u_multiplier_pp3_32 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_32__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_32__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_32__22_  (.A(u_multiplier_pp3_32 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_32__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_32__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_32__23_  (.A1(u_multiplier_pp3_32 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_32__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_32__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_32__24_  (.A(u_multiplier_pp3_32 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_32__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_32__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_32__25_  (.A(u_multiplier_STAGE4_pp4_31_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_32__16_ ),
    .ZN(u_multiplier_A [32]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_32__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_32__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_32__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_32_cout ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_32__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_32__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_32__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_32__17_ ),
    .ZN(u_multiplier_B [33]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_33__18_  (.A(u_multiplier_STAGE4_pp4_32_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_33__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_33__19_  (.A1(u_multiplier_pp3_33 [1]),
    .A2(u_multiplier_pp3_33 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_33__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_33__20_  (.A(u_multiplier_pp3_33 [1]),
    .B(u_multiplier_pp3_33 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_33__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_33__21_  (.A1(u_multiplier_pp3_33 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_33__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_33__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_33__22_  (.A(u_multiplier_pp3_33 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_33__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_33__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_33__23_  (.A1(u_multiplier_pp3_33 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_33__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_33__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_33__24_  (.A(u_multiplier_pp3_33 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_33__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_33__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_33__25_  (.A(u_multiplier_STAGE4_pp4_32_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_33__16_ ),
    .ZN(u_multiplier_A [33]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_33__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_33__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_33__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_33_cout ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_33__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_33__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_33__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_33__17_ ),
    .ZN(u_multiplier_B [34]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_34__18_  (.A(u_multiplier_STAGE4_pp4_33_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_34__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_34__19_  (.A1(u_multiplier_pp3_34 [1]),
    .A2(u_multiplier_pp3_34 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_34__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_34__20_  (.A(u_multiplier_pp3_34 [1]),
    .B(u_multiplier_pp3_34 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_34__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_34__21_  (.A1(u_multiplier_pp3_34 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_34__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_34__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_34__22_  (.A(u_multiplier_pp3_34 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_34__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_34__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_34__23_  (.A1(u_multiplier_pp3_34 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_34__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_34__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_34__24_  (.A(u_multiplier_pp3_34 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_34__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_34__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_34__25_  (.A(u_multiplier_STAGE4_pp4_33_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_34__16_ ),
    .ZN(u_multiplier_A [34]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_34__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_34__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_34__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_34_cout ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_34__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_34__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_34__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_34__17_ ),
    .ZN(u_multiplier_B [35]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_35__18_  (.A(u_multiplier_STAGE4_pp4_34_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_35__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_35__19_  (.A1(u_multiplier_pp3_35 [1]),
    .A2(u_multiplier_pp3_35 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_35__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_35__20_  (.A(u_multiplier_pp3_35 [1]),
    .B(u_multiplier_pp3_35 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_35__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_35__21_  (.A1(u_multiplier_pp3_35 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_35__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_35__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_35__22_  (.A(u_multiplier_pp3_35 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_35__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_35__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_35__23_  (.A1(u_multiplier_pp3_35 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_35__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_35__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_35__24_  (.A(u_multiplier_pp3_35 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_35__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_35__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_35__25_  (.A(u_multiplier_STAGE4_pp4_34_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_35__16_ ),
    .ZN(u_multiplier_A [35]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_35__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_35__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_35__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_35_cout ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_35__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_35__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_35__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_35__17_ ),
    .ZN(u_multiplier_B [36]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_36__18_  (.A(u_multiplier_STAGE4_pp4_35_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_36__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_36__19_  (.A1(u_multiplier_pp3_36 [1]),
    .A2(u_multiplier_pp3_36 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_36__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_36__20_  (.A(u_multiplier_pp3_36 [1]),
    .B(u_multiplier_pp3_36 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_36__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_36__21_  (.A1(u_multiplier_pp3_36 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_36__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_36__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_36__22_  (.A(u_multiplier_pp3_36 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_36__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_36__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_36__23_  (.A1(u_multiplier_pp3_36 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_36__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_36__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_36__24_  (.A(u_multiplier_pp3_36 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_36__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_36__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_36__25_  (.A(u_multiplier_STAGE4_pp4_35_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_36__16_ ),
    .ZN(u_multiplier_A [36]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_36__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_36__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_36__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_36_cout ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_36__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_36__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_36__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_36__17_ ),
    .ZN(u_multiplier_B [37]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_37__18_  (.A(u_multiplier_STAGE4_pp4_36_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_37__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_37__19_  (.A1(u_multiplier_pp3_37 [1]),
    .A2(u_multiplier_pp3_37 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_37__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_37__20_  (.A(u_multiplier_pp3_37 [1]),
    .B(u_multiplier_pp3_37 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_37__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_37__21_  (.A1(u_multiplier_pp3_37 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_37__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_37__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_37__22_  (.A(u_multiplier_pp3_37 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_37__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_37__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_37__23_  (.A1(u_multiplier_pp3_37 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_37__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_37__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_37__24_  (.A(u_multiplier_pp3_37 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_37__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_37__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_37__25_  (.A(u_multiplier_STAGE4_pp4_36_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_37__16_ ),
    .ZN(u_multiplier_A [37]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_37__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_37__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_37__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_37_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_37__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_37__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_37__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_37__17_ ),
    .ZN(u_multiplier_B [38]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_38__18_  (.A(u_multiplier_STAGE4_pp4_37_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_38__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_38__19_  (.A1(u_multiplier_pp3_38 [1]),
    .A2(u_multiplier_pp3_38 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_38__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_38__20_  (.A(u_multiplier_pp3_38 [1]),
    .B(u_multiplier_pp3_38 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_38__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_38__21_  (.A1(u_multiplier_pp3_38 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_38__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_38__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_38__22_  (.A(u_multiplier_pp3_38 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_38__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_38__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_38__23_  (.A1(u_multiplier_pp3_38 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_38__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_38__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_38__24_  (.A(u_multiplier_pp3_38 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_38__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_38__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_38__25_  (.A(u_multiplier_STAGE4_pp4_37_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_38__16_ ),
    .ZN(u_multiplier_A [38]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_38__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_38__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_38__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_38_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_38__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_38__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_38__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_38__17_ ),
    .ZN(u_multiplier_B [39]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_39__18_  (.A(u_multiplier_STAGE4_pp4_38_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_39__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_39__19_  (.A1(u_multiplier_pp3_39 [1]),
    .A2(u_multiplier_pp3_39 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_39__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_39__20_  (.A(u_multiplier_pp3_39 [1]),
    .B(u_multiplier_pp3_39 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_39__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_39__21_  (.A1(u_multiplier_pp3_39 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_39__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_39__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_39__22_  (.A(u_multiplier_pp3_39 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_39__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_39__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_39__23_  (.A1(u_multiplier_pp3_39 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_39__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_39__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_39__24_  (.A(u_multiplier_pp3_39 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_39__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_39__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_39__25_  (.A(u_multiplier_STAGE4_pp4_38_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_39__16_ ),
    .ZN(u_multiplier_A [39]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_39__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_39__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_39__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_39_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_39__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_39__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_39__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_39__17_ ),
    .ZN(u_multiplier_B [40]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_4__18_  (.A(u_multiplier_STAGE4_pp4_3_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_4__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_4__19_  (.A1(u_multiplier_pp3_4 [1]),
    .A2(u_multiplier_pp3_4 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_4__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_4__20_  (.A(u_multiplier_pp3_4 [1]),
    .B(u_multiplier_pp3_4 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_4__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_4__21_  (.A1(u_multiplier_pp3_4 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_4__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_4__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_4__22_  (.A(u_multiplier_pp3_4 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_4__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_4__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_4__23_  (.A1(u_multiplier_pp3_4 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_4__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_4__24_  (.A(u_multiplier_pp3_4 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_4__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_4__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_4__25_  (.A(u_multiplier_STAGE4_pp4_3_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_4__16_ ),
    .ZN(u_multiplier_A [4]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_4__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_4__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_4__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_4_cout ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_4__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_4__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_4__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_4__17_ ),
    .ZN(u_multiplier_B [5]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_40__18_  (.A(u_multiplier_STAGE4_pp4_39_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_40__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_40__19_  (.A1(u_multiplier_pp3_40 [1]),
    .A2(u_multiplier_pp3_40 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_40__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_40__20_  (.A(u_multiplier_pp3_40 [1]),
    .B(u_multiplier_pp3_40 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_40__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_40__21_  (.A1(u_multiplier_pp3_40 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_40__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_40__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_40__22_  (.A(u_multiplier_pp3_40 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_40__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_40__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_40__23_  (.A1(u_multiplier_pp3_40 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_40__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_40__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_40__24_  (.A(u_multiplier_pp3_40 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_40__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_40__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_40__25_  (.A(u_multiplier_STAGE4_pp4_39_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_40__16_ ),
    .ZN(u_multiplier_A [40]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_40__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_40__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_40__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_40_cout ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_40__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_40__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_40__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_40__17_ ),
    .ZN(u_multiplier_B [41]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_41__18_  (.A(u_multiplier_STAGE4_pp4_40_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_41__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_41__19_  (.A1(u_multiplier_pp3_41 [1]),
    .A2(u_multiplier_pp3_41 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_41__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_41__20_  (.A(u_multiplier_pp3_41 [1]),
    .B(u_multiplier_pp3_41 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_41__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_41__21_  (.A1(u_multiplier_pp3_41 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_41__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_41__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_41__22_  (.A(u_multiplier_pp3_41 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_41__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_41__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_41__23_  (.A1(u_multiplier_pp3_41 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_41__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_41__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_41__24_  (.A(u_multiplier_pp3_41 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_41__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_41__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_41__25_  (.A(u_multiplier_STAGE4_pp4_40_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_41__16_ ),
    .ZN(u_multiplier_A [41]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_41__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_41__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_41__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_41_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_41__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_41__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_41__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_41__17_ ),
    .ZN(u_multiplier_B [42]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_42__18_  (.A(u_multiplier_STAGE4_pp4_41_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_42__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_42__19_  (.A1(u_multiplier_pp3_42 [1]),
    .A2(u_multiplier_pp3_42 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_42__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_42__20_  (.A(u_multiplier_pp3_42 [1]),
    .B(u_multiplier_pp3_42 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_42__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_42__21_  (.A1(u_multiplier_pp3_42 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_42__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_42__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_42__22_  (.A(u_multiplier_pp3_42 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_42__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_42__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_42__23_  (.A1(u_multiplier_pp3_42 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_42__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_42__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_42__24_  (.A(u_multiplier_pp3_42 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_42__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_42__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_42__25_  (.A(u_multiplier_STAGE4_pp4_41_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_42__16_ ),
    .ZN(u_multiplier_A [42]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_42__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_42__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_42__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_42_cout ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_42__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_42__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_42__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_42__17_ ),
    .ZN(u_multiplier_B [43]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_43__18_  (.A(u_multiplier_STAGE4_pp4_42_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_43__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_43__19_  (.A1(u_multiplier_pp3_43 [1]),
    .A2(u_multiplier_pp3_43 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_43__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_43__20_  (.A(u_multiplier_pp3_43 [1]),
    .B(u_multiplier_pp3_43 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_43__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_43__21_  (.A1(u_multiplier_pp3_43 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_43__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_43__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_43__22_  (.A(u_multiplier_pp3_43 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_43__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_43__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_43__23_  (.A1(u_multiplier_pp3_43 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_43__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_43__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_43__24_  (.A(u_multiplier_pp3_43 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_43__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_43__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_43__25_  (.A(u_multiplier_STAGE4_pp4_42_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_43__16_ ),
    .ZN(u_multiplier_A [43]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_43__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_43__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_43__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_43_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_43__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_43__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_43__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_43__17_ ),
    .ZN(u_multiplier_B [44]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_44__18_  (.A(u_multiplier_STAGE4_pp4_43_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_44__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_44__19_  (.A1(u_multiplier_pp3_44 [1]),
    .A2(u_multiplier_pp3_44 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_44__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_44__20_  (.A(u_multiplier_pp3_44 [1]),
    .B(u_multiplier_pp3_44 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_44__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_44__21_  (.A1(u_multiplier_pp3_44 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_44__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_44__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_44__22_  (.A(u_multiplier_pp3_44 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_44__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_44__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_44__23_  (.A1(u_multiplier_pp3_44 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_44__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_44__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_44__24_  (.A(u_multiplier_pp3_44 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_44__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_44__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_44__25_  (.A(u_multiplier_STAGE4_pp4_43_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_44__16_ ),
    .ZN(u_multiplier_A [44]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_44__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_44__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_44__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_44_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_44__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_44__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_44__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_44__17_ ),
    .ZN(u_multiplier_B [45]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_45__18_  (.A(u_multiplier_STAGE4_pp4_44_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_45__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_45__19_  (.A1(u_multiplier_pp3_45 [1]),
    .A2(u_multiplier_pp3_45 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_45__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_45__20_  (.A(u_multiplier_pp3_45 [1]),
    .B(u_multiplier_pp3_45 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_45__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_45__21_  (.A1(u_multiplier_pp3_45 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_45__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_45__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_45__22_  (.A(u_multiplier_pp3_45 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_45__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_45__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_45__23_  (.A1(u_multiplier_pp3_45 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_45__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_45__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_45__24_  (.A(u_multiplier_pp3_45 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_45__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_45__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_45__25_  (.A(u_multiplier_STAGE4_pp4_44_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_45__16_ ),
    .ZN(u_multiplier_A [45]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_45__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_45__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_45__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_45_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_45__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_45__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_45__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_45__17_ ),
    .ZN(u_multiplier_B [46]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_46__18_  (.A(u_multiplier_STAGE4_pp4_45_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_46__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_46__19_  (.A1(u_multiplier_pp3_46 [1]),
    .A2(u_multiplier_pp3_46 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_46__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_46__20_  (.A(u_multiplier_pp3_46 [1]),
    .B(u_multiplier_pp3_46 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_46__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_46__21_  (.A1(u_multiplier_pp3_46 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_46__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_46__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_46__22_  (.A(u_multiplier_pp3_46 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_46__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_46__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_46__23_  (.A1(u_multiplier_pp3_46 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_46__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_46__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_46__24_  (.A(u_multiplier_pp3_46 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_46__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_46__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_46__25_  (.A(u_multiplier_STAGE4_pp4_45_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_46__16_ ),
    .ZN(u_multiplier_A [46]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_46__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_46__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_46__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_46_cout ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_46__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_46__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_46__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_46__17_ ),
    .ZN(u_multiplier_B [47]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_47__18_  (.A(u_multiplier_STAGE4_pp4_46_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_47__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_47__19_  (.A1(u_multiplier_pp3_47 [1]),
    .A2(u_multiplier_pp3_47 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_47__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_47__20_  (.A(u_multiplier_pp3_47 [1]),
    .B(u_multiplier_pp3_47 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_47__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_47__21_  (.A1(u_multiplier_pp3_47 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_47__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_47__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_47__22_  (.A(u_multiplier_pp3_47 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_47__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_47__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_47__23_  (.A1(u_multiplier_pp3_47 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_47__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_47__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_47__24_  (.A(u_multiplier_pp3_47 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_47__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_47__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_47__25_  (.A(u_multiplier_STAGE4_pp4_46_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_47__16_ ),
    .ZN(u_multiplier_A [47]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_47__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_47__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_47__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_47_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_47__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_47__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_47__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_47__17_ ),
    .ZN(u_multiplier_B [48]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_48__18_  (.A(u_multiplier_STAGE4_pp4_47_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_48__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_48__19_  (.A1(u_multiplier_pp3_48 [1]),
    .A2(u_multiplier_pp3_48 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_48__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_48__20_  (.A(u_multiplier_pp3_48 [1]),
    .B(u_multiplier_pp3_48 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_48__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_48__21_  (.A1(u_multiplier_pp3_48 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_48__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_48__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_48__22_  (.A(u_multiplier_pp3_48 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_48__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_48__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_48__23_  (.A1(u_multiplier_pp3_48 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_48__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_48__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_48__24_  (.A(u_multiplier_pp3_48 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_48__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_48__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_48__25_  (.A(u_multiplier_STAGE4_pp4_47_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_48__16_ ),
    .ZN(u_multiplier_A [48]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_48__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_48__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_48__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_48_cout ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_48__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_48__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_48__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_48__17_ ),
    .ZN(u_multiplier_B [49]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_49__18_  (.A(u_multiplier_STAGE4_pp4_48_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_49__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_49__19_  (.A1(u_multiplier_pp3_49 [1]),
    .A2(u_multiplier_pp3_49 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_49__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_49__20_  (.A(u_multiplier_pp3_49 [1]),
    .B(u_multiplier_pp3_49 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_49__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_49__21_  (.A1(u_multiplier_pp3_49 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_49__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_49__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_49__22_  (.A(u_multiplier_pp3_49 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_49__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_49__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_49__23_  (.A1(u_multiplier_pp3_49 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_49__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_49__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_49__24_  (.A(u_multiplier_pp3_49 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_49__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_49__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_49__25_  (.A(u_multiplier_STAGE4_pp4_48_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_49__16_ ),
    .ZN(u_multiplier_A [49]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_49__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_49__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_49__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_49_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_49__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_49__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_49__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_49__17_ ),
    .ZN(u_multiplier_B [50]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_5__18_  (.A(u_multiplier_STAGE4_pp4_4_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_5__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_5__19_  (.A1(u_multiplier_pp3_5 [1]),
    .A2(u_multiplier_pp3_5 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_5__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_5__20_  (.A(u_multiplier_pp3_5 [1]),
    .B(u_multiplier_pp3_5 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_5__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_5__21_  (.A1(u_multiplier_pp3_5 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_5__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_5__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_5__22_  (.A(u_multiplier_pp3_5 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_5__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_5__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_5__23_  (.A1(u_multiplier_pp3_5 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_5__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_5__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_5__24_  (.A(u_multiplier_pp3_5 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_5__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_5__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_5__25_  (.A(u_multiplier_STAGE4_pp4_4_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_5__16_ ),
    .ZN(u_multiplier_A [5]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_5__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_5__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_5__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_5_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_5__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_5__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_5__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_5__17_ ),
    .ZN(u_multiplier_B [6]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_50__18_  (.A(u_multiplier_STAGE4_pp4_49_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_50__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_50__19_  (.A1(u_multiplier_pp3_50 [1]),
    .A2(u_multiplier_pp3_50 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_50__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_50__20_  (.A(u_multiplier_pp3_50 [1]),
    .B(u_multiplier_pp3_50 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_50__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_50__21_  (.A1(u_multiplier_pp3_50 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_50__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_50__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_50__22_  (.A(u_multiplier_pp3_50 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_50__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_50__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_50__23_  (.A1(u_multiplier_pp3_50 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_50__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_50__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_50__24_  (.A(u_multiplier_pp3_50 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_50__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_50__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_50__25_  (.A(u_multiplier_STAGE4_pp4_49_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_50__16_ ),
    .ZN(u_multiplier_A [50]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_50__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_50__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_50__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_50_cout ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_50__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_50__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_50__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_50__17_ ),
    .ZN(u_multiplier_B [51]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_51__18_  (.A(u_multiplier_STAGE4_pp4_50_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_51__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_51__19_  (.A1(u_multiplier_pp3_51 [1]),
    .A2(u_multiplier_pp3_51 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_51__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_51__20_  (.A(u_multiplier_pp3_51 [1]),
    .B(u_multiplier_pp3_51 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_51__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_51__21_  (.A1(u_multiplier_pp3_51 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_51__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_51__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_51__22_  (.A(u_multiplier_pp3_51 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_51__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_51__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_51__23_  (.A1(u_multiplier_pp3_51 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_51__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_51__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_51__24_  (.A(u_multiplier_pp3_51 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_51__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_51__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_51__25_  (.A(u_multiplier_STAGE4_pp4_50_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_51__16_ ),
    .ZN(u_multiplier_A [51]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_51__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_51__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_51__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_51_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_51__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_51__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_51__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_51__17_ ),
    .ZN(u_multiplier_B [52]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_52__18_  (.A(u_multiplier_STAGE4_pp4_51_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_52__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_52__19_  (.A1(u_multiplier_pp3_52 [1]),
    .A2(u_multiplier_pp3_52 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_52__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_52__20_  (.A(u_multiplier_pp3_52 [1]),
    .B(u_multiplier_pp3_52 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_52__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_52__21_  (.A1(u_multiplier_pp3_52 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_52__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_52__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_52__22_  (.A(u_multiplier_pp3_52 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_52__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_52__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_52__23_  (.A1(u_multiplier_pp3_52 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_52__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_52__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_52__24_  (.A(u_multiplier_pp3_52 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_52__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_52__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_52__25_  (.A(u_multiplier_STAGE4_pp4_51_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_52__16_ ),
    .ZN(u_multiplier_A [52]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_52__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_52__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_52__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_52_cout ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_52__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_52__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_52__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_52__17_ ),
    .ZN(u_multiplier_B [53]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_53__18_  (.A(u_multiplier_STAGE4_pp4_52_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_53__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_53__19_  (.A1(u_multiplier_pp3_53 [1]),
    .A2(u_multiplier_pp3_53 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_53__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_53__20_  (.A(u_multiplier_pp3_53 [1]),
    .B(u_multiplier_pp3_53 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_53__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_53__21_  (.A1(u_multiplier_pp3_53 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_53__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_53__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_53__22_  (.A(u_multiplier_pp3_53 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_53__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_53__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_53__23_  (.A1(u_multiplier_pp3_53 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_53__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_53__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_53__24_  (.A(u_multiplier_pp3_53 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_53__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_53__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_53__25_  (.A(u_multiplier_STAGE4_pp4_52_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_53__16_ ),
    .ZN(u_multiplier_A [53]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_53__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_53__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_53__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_53_cout ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_53__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_53__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_53__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_53__17_ ),
    .ZN(u_multiplier_B [54]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_54__18_  (.A(u_multiplier_STAGE4_pp4_53_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_54__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_54__19_  (.A1(u_multiplier_pp3_54 [1]),
    .A2(u_multiplier_pp3_54 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_54__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_54__20_  (.A(u_multiplier_pp3_54 [1]),
    .B(u_multiplier_pp3_54 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_54__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_54__21_  (.A1(u_multiplier_pp3_54 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_54__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_54__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_54__22_  (.A(u_multiplier_pp3_54 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_54__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_54__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_54__23_  (.A1(u_multiplier_pp3_54 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_54__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_54__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_54__24_  (.A(u_multiplier_pp3_54 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_54__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_54__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_54__25_  (.A(u_multiplier_STAGE4_pp4_53_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_54__16_ ),
    .ZN(u_multiplier_A [54]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_54__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_54__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_54__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_54_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_54__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_54__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_54__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_54__17_ ),
    .ZN(u_multiplier_B [55]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_55__18_  (.A(u_multiplier_STAGE4_pp4_54_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_55__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_55__19_  (.A1(u_multiplier_pp3_55 [1]),
    .A2(u_multiplier_pp3_55 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_55__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_55__20_  (.A(u_multiplier_pp3_55 [1]),
    .B(u_multiplier_pp3_55 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_55__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_55__21_  (.A1(u_multiplier_pp3_55 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_55__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_55__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_55__22_  (.A(u_multiplier_pp3_55 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_55__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_55__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_55__23_  (.A1(u_multiplier_pp3_55 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_55__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_55__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_55__24_  (.A(u_multiplier_pp3_55 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_55__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_55__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_55__25_  (.A(u_multiplier_STAGE4_pp4_54_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_55__16_ ),
    .ZN(u_multiplier_A [55]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_55__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_55__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_55__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_55_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_55__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_55__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_55__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_55__17_ ),
    .ZN(u_multiplier_B [56]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_56__18_  (.A(u_multiplier_STAGE4_pp4_55_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_56__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_56__19_  (.A1(u_multiplier_pp3_56 [1]),
    .A2(u_multiplier_pp3_56 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_56__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_56__20_  (.A(u_multiplier_pp3_56 [1]),
    .B(u_multiplier_pp3_56 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_56__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_56__21_  (.A1(u_multiplier_pp3_56 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_56__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_56__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_56__22_  (.A(u_multiplier_pp3_56 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_56__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_56__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_56__23_  (.A1(u_multiplier_pp3_56 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_56__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_56__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_56__24_  (.A(u_multiplier_pp3_56 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_56__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_56__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_56__25_  (.A(u_multiplier_STAGE4_pp4_55_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_56__16_ ),
    .ZN(u_multiplier_A [56]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_56__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_56__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_56__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_56_cout ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_56__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_56__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_56__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_56__17_ ),
    .ZN(u_multiplier_B [57]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_57__18_  (.A(u_multiplier_STAGE4_pp4_56_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_57__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_57__19_  (.A1(u_multiplier_pp3_57 [1]),
    .A2(u_multiplier_pp3_57 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_57__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_57__20_  (.A(u_multiplier_pp3_57 [1]),
    .B(u_multiplier_pp3_57 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_57__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_57__21_  (.A1(u_multiplier_pp3_57 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_57__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_57__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_57__22_  (.A(u_multiplier_pp3_57 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_57__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_57__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_57__23_  (.A1(u_multiplier_pp3_57 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_57__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_57__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_57__24_  (.A(u_multiplier_pp3_57 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_57__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_57__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_57__25_  (.A(u_multiplier_STAGE4_pp4_56_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_57__16_ ),
    .ZN(u_multiplier_A [57]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_57__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_57__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_57__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_57_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_57__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_57__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_57__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_57__17_ ),
    .ZN(u_multiplier_B [58]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_58__18_  (.A(u_multiplier_STAGE4_pp4_57_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_58__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_58__19_  (.A1(u_multiplier_pp3_58 [1]),
    .A2(u_multiplier_pp3_58 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_58__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_58__20_  (.A(u_multiplier_pp3_58 [1]),
    .B(u_multiplier_pp3_58 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_58__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_58__21_  (.A1(u_multiplier_pp3_58 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_58__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_58__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_58__22_  (.A(u_multiplier_pp3_58 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_58__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_58__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_58__23_  (.A1(u_multiplier_pp3_58 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_58__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_58__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_58__24_  (.A(u_multiplier_pp3_58 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_58__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_58__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_58__25_  (.A(u_multiplier_STAGE4_pp4_57_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_58__16_ ),
    .ZN(u_multiplier_A [58]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_58__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_58__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_58__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_58_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_58__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_58__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_58__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_58__17_ ),
    .ZN(u_multiplier_B [59]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_59__18_  (.A(u_multiplier_STAGE4_pp4_58_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_59__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_59__19_  (.A1(u_multiplier_pp3_59 [1]),
    .A2(u_multiplier_pp3_59 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_59__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_59__20_  (.A(u_multiplier_pp3_59 [1]),
    .B(u_multiplier_pp3_59 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_59__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_59__21_  (.A1(u_multiplier_pp3_59 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_59__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_59__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_59__22_  (.A(u_multiplier_pp3_59 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_59__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_59__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_59__23_  (.A1(u_multiplier_pp3_59 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_59__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_59__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_59__24_  (.A(u_multiplier_pp3_59 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_59__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_59__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_59__25_  (.A(u_multiplier_STAGE4_pp4_58_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_59__16_ ),
    .ZN(u_multiplier_A [59]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_59__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_59__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_59__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_59_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_59__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_59__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_59__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_59__17_ ),
    .ZN(u_multiplier_B [60]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_6__18_  (.A(u_multiplier_STAGE4_pp4_5_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_6__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_6__19_  (.A1(u_multiplier_pp3_6 [1]),
    .A2(u_multiplier_pp3_6 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_6__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_6__20_  (.A(u_multiplier_pp3_6 [1]),
    .B(u_multiplier_pp3_6 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_6__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_6__21_  (.A1(u_multiplier_pp3_6 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_6__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_6__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_6__22_  (.A(u_multiplier_pp3_6 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_6__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_6__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_6__23_  (.A1(u_multiplier_pp3_6 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_6__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_6__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_6__24_  (.A(u_multiplier_pp3_6 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_6__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_6__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_6__25_  (.A(u_multiplier_STAGE4_pp4_5_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_6__16_ ),
    .ZN(u_multiplier_A [6]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_6__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_6__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_6__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_6_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_6__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_6__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_6__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_6__17_ ),
    .ZN(u_multiplier_B [7]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_60__18_  (.A(u_multiplier_STAGE4_pp4_59_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_60__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_60__19_  (.A1(u_multiplier_pp3_60 [1]),
    .A2(u_multiplier_pp3_60 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_60__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_60__20_  (.A(u_multiplier_pp3_60 [1]),
    .B(u_multiplier_pp3_60 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_60__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_60__21_  (.A1(u_multiplier_pp3_60 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_60__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_60__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_60__22_  (.A(u_multiplier_pp3_60 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_60__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_60__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_60__23_  (.A1(u_multiplier_pp3_60 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_60__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_60__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_60__24_  (.A(u_multiplier_pp3_60 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_60__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_60__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_60__25_  (.A(u_multiplier_STAGE4_pp4_59_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_60__16_ ),
    .ZN(u_multiplier_A [60]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_60__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_60__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_60__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_60_cout ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_60__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_60__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_60__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_60__17_ ),
    .ZN(u_multiplier_B [61]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_7__18_  (.A(u_multiplier_STAGE4_pp4_6_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_7__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_7__19_  (.A1(u_multiplier_pp3_7 [1]),
    .A2(u_multiplier_pp3_7 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_7__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_7__20_  (.A(u_multiplier_pp3_7 [1]),
    .B(u_multiplier_pp3_7 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_7__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_7__21_  (.A1(u_multiplier_pp3_7 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_7__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_7__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_7__22_  (.A(u_multiplier_pp3_7 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_7__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_7__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_7__23_  (.A1(u_multiplier_pp3_7 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_7__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_7__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_7__24_  (.A(u_multiplier_pp3_7 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_7__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_7__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_7__25_  (.A(u_multiplier_STAGE4_pp4_6_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_7__16_ ),
    .ZN(u_multiplier_A [7]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_7__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_7__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_7__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_7_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_7__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_7__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_7__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_7__17_ ),
    .ZN(u_multiplier_B [8]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_8__18_  (.A(u_multiplier_STAGE4_pp4_7_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_8__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_8__19_  (.A1(u_multiplier_pp3_8 [1]),
    .A2(u_multiplier_pp3_8 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_8__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_8__20_  (.A(u_multiplier_pp3_8 [1]),
    .B(u_multiplier_pp3_8 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_8__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_8__21_  (.A1(u_multiplier_pp3_8 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_8__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_8__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_8__22_  (.A(u_multiplier_pp3_8 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_8__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_8__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_8__23_  (.A1(u_multiplier_pp3_8 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_8__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_8__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_8__24_  (.A(u_multiplier_pp3_8 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_8__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_8__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_8__25_  (.A(u_multiplier_STAGE4_pp4_7_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_8__16_ ),
    .ZN(u_multiplier_A [8]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_8__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_8__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_8__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_8_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_8__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_8__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_8__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_8__17_ ),
    .ZN(u_multiplier_B [9]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_9__18_  (.A(u_multiplier_STAGE4_pp4_8_cout ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_9__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_9__19_  (.A1(u_multiplier_pp3_9 [1]),
    .A2(u_multiplier_pp3_9 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_9__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_9__20_  (.A(u_multiplier_pp3_9 [1]),
    .B(u_multiplier_pp3_9 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_9__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_9__21_  (.A1(u_multiplier_pp3_9 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_9__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_9__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_9__22_  (.A(u_multiplier_pp3_9 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_9__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_9__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_9__23_  (.A1(u_multiplier_pp3_9 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_9__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_9__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_9__24_  (.A(u_multiplier_pp3_9 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_9__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_9__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_9__25_  (.A(u_multiplier_STAGE4_pp4_8_cout ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_9__16_ ),
    .ZN(u_multiplier_A [9]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_9__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_9__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_9__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_9_cout ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_9__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_9__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_9__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_9__17_ ),
    .ZN(u_multiplier_B [10]));
 INV_X1 u_multiplier_STAGE4_Full_adder_pp4_61__12_  (.A(u_multiplier_STAGE4_pp4_60_cout ),
    .ZN(u_multiplier_STAGE4_Full_adder_pp4_61__08_ ));
 NAND3_X2 u_multiplier_STAGE4_Full_adder_pp4_61__13_  (.A1(u_multiplier_pp3_61 [1]),
    .A2(u_multiplier_pp3_61 [0]),
    .A3(u_multiplier_STAGE4_pp4_60_cout ),
    .ZN(u_multiplier_STAGE4_Full_adder_pp4_61__09_ ));
 NOR2_X2 u_multiplier_STAGE4_Full_adder_pp4_61__14_  (.A1(u_multiplier_pp3_61 [1]),
    .A2(u_multiplier_pp3_61 [0]),
    .ZN(u_multiplier_STAGE4_Full_adder_pp4_61__10_ ));
 AOI21_X1 u_multiplier_STAGE4_Full_adder_pp4_61__15_  (.A(u_multiplier_STAGE4_pp4_60_cout ),
    .B1(u_multiplier_pp3_61 [0]),
    .B2(u_multiplier_pp3_61 [1]),
    .ZN(u_multiplier_STAGE4_Full_adder_pp4_61__11_ ));
 NOR2_X2 u_multiplier_STAGE4_Full_adder_pp4_61__16_  (.A1(u_multiplier_STAGE4_Full_adder_pp4_61__10_ ),
    .A2(u_multiplier_STAGE4_Full_adder_pp4_61__11_ ),
    .ZN(u_multiplier_B [62]));
 AOI22_X4 u_multiplier_STAGE4_Full_adder_pp4_61__17_  (.A1(u_multiplier_STAGE4_Full_adder_pp4_61__08_ ),
    .A2(u_multiplier_STAGE4_Full_adder_pp4_61__10_ ),
    .B1(u_multiplier_B [62]),
    .B2(u_multiplier_STAGE4_Full_adder_pp4_61__09_ ),
    .ZN(u_multiplier_A [61]));
 AND2_X1 u_multiplier_STAGE4_Half_adder_pp4_1__4_  (.A1(u_multiplier_pp3_1 [1]),
    .A2(u_multiplier_pp3_1 [0]),
    .ZN(u_multiplier_STAGE4_pp4_1_ha_c ));
 XOR2_X2 u_multiplier_STAGE4_Half_adder_pp4_1__5_  (.A(u_multiplier_pp3_1 [1]),
    .B(u_multiplier_pp3_1 [0]),
    .Z(u_multiplier_A [1]));
 LOGIC0_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__43__161  (.Z(net161));
 CLKBUF_X1 hold163 (.A(net217),
    .Z(net163));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_219_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_220_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_221_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_222_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_223_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_224_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_225_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_226_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_227_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_228_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_229_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_230_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_231_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_232_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_233_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_234_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_235_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_236_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_237_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_2_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_2_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_2_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_2_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_2_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_2_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_2_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_2_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_2_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_2_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_2_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_2_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_2_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_2_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_2_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_2_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_2_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_2_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_2_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_2_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_2_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_2_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_2_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_2_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_2_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_2_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_2_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_2_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_2_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_2_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_2_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_2_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_2_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_2_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_2_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_2_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_2_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_2_Right_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_2_Right_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_2_Right_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_2_Right_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_2_Right_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_2_Right_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_2_Right_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_2_Right_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_2_Right_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_2_Right_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_2_Right_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_2_Right_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_2_Right_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_2_Right_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_2_Right_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_2_Right_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_2_Right_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_2_Right_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_2_Right_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_2_Right_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_2_Right_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_2_Right_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_2_Right_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_2_Right_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_2_Right_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_2_Right_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_2_Right_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_2_Right_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_2_Right_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_2_Right_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_2_Right_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_2_Right_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_2_Right_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_2_Right_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_2_Right_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_2_Right_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_2_Right_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_2_Right_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_2_Right_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_2_Right_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_2_Right_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_2_Right_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_2_Right_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_2_Right_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_2_Right_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_2_Right_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_2_Right_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_2_Right_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_2_Right_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_2_Right_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_2_Right_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_2_Right_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_2_Right_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_2_Right_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_2_Right_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_2_Right_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_2_Right_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_2_Right_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_2_Right_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_2_Right_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_2_Right_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_2_Right_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_2_Right_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_2_Right_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_2_Right_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_2_Right_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_2_Right_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_2_Right_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_2_Right_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_2_Right_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_2_Right_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_2_Right_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_2_Right_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_2_Right_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_2_Right_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_2_Right_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_2_Right_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_2_Right_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_2_Right_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_2_Right_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_2_Right_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_2_Right_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_2_Right_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_2_Right_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_2_Right_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_2_Right_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_2_Right_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_2_Right_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_2_Right_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_2_Right_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_2_Right_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_2_Right_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_2_Right_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_2_Right_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_2_Right_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_2_Right_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_2_Right_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_2_Right_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_2_Right_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_2_Right_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_2_Right_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_2_Right_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_2_Right_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_2_Right_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_2_Right_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_2_Right_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_2_Right_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_2_Right_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_2_Right_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_2_Right_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_2_Right_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_2_Right_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_2_Right_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_2_Right_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_2_Right_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_2_Right_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_2_Right_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_2_Right_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_2_Right_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_2_Right_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_2_Right_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_2_Right_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_2_Right_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_2_Right_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_2_Right_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_2_Right_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_2_Right_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_2_Right_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_2_Right_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_2_Right_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_2_Right_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_265 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_266 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_267 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_268 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_269 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_270 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_271 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_272 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_273 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_274 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_275 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_276 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_277 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_1_Left_278 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_1_Left_279 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_1_Left_280 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_1_Left_281 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_1_Left_282 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_1_Left_283 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_1_Left_284 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_1_Left_285 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_1_Left_286 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_1_Left_287 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_1_Left_288 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_1_Left_289 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_1_Left_290 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_1_Left_291 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_1_Left_292 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_1_Left_293 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_1_Left_294 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_1_Left_295 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_1_Left_296 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_1_Left_297 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_1_Left_298 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_1_Left_299 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_1_Left_300 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_1_Left_301 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_1_Left_302 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_1_Left_303 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_1_Left_304 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_1_Left_305 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_1_Left_306 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_1_Left_307 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_1_Left_308 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_1_Left_309 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_1_Left_310 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_1_Left_311 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_1_Left_312 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_1_Left_313 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_1_Left_314 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_1_Left_315 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_1_Left_316 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_1_Left_317 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_1_Left_318 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_1_Left_319 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_1_Left_320 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_1_Left_321 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_1_Left_322 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_1_Left_323 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_1_Left_324 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_1_Left_325 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_1_Left_326 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_1_Left_327 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_1_Left_328 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_1_Left_329 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_1_Left_330 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_1_Left_331 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_1_Left_332 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_1_Left_333 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_1_Left_334 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_1_Left_335 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_1_Left_336 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_1_Left_337 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_1_Left_338 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_1_Left_339 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_1_Left_340 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_1_Left_341 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_1_Left_342 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_1_Left_343 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_1_Left_344 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_1_Left_345 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_1_Left_346 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_1_Left_347 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_1_Left_348 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_1_Left_349 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_1_Left_350 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_1_Left_351 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_1_Left_352 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_1_Left_353 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_1_Left_354 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_1_Left_355 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_1_Left_356 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_1_Left_357 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_1_Left_358 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_1_Left_359 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_1_Left_360 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_1_Left_361 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_1_Left_362 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_1_Left_363 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_1_Left_364 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_1_Left_365 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_1_Left_366 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_1_Left_367 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_1_Left_368 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_1_Left_369 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_1_Left_370 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_1_Left_371 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_1_Left_372 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_1_Left_373 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_1_Left_374 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_1_Left_375 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_1_Left_376 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_1_Left_377 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_1_Left_378 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_1_Left_379 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_1_Left_380 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_1_Left_381 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_1_Left_382 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_1_Left_383 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_1_Left_384 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_1_Left_385 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_1_Left_386 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_1_Left_387 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_1_Left_388 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_1_Left_389 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_1_Left_390 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_1_Left_391 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_1_Left_392 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_1_Left_393 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_1_Left_394 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_1_Left_395 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_1_Left_396 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_1_Left_397 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_1_Left_398 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_1_Left_399 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_1_Left_400 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_1_Left_401 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_1_Left_402 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_1_Left_403 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_1_Left_404 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_1_Left_405 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_1_Left_406 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_1_Left_407 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_1_Left_408 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_1_Left_409 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_1_Left_410 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_1_Left_411 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_1_Left_412 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_1_Left_413 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_1_Left_414 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_1_Left_415 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_1_Left_416 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_1_Left_417 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_1_Left_418 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_1_Left_419 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_1_Left_420 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_1_Left_421 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_1_Left_422 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_1_Left_423 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_1_Left_424 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_1_Left_425 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_1_Left_426 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_1_Left_427 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_1_Left_428 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_1_Left_429 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_1_Left_430 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_1_Left_431 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_1_Left_432 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_1_Left_433 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_1_Left_434 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_1_Left_435 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_1_Left_436 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_1_Left_437 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_1_Left_438 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_1_Left_439 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_1_Left_440 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_1_Left_441 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_1_Left_442 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_1_Left_443 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_1_Left_444 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Left_445 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Left_446 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Left_447 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Left_448 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Left_449 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Left_450 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Left_451 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Left_452 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Left_453 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Left_454 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Left_455 ();
 TAPCELL_X1 PHY_EDGE_ROW_219_Left_456 ();
 TAPCELL_X1 PHY_EDGE_ROW_220_Left_457 ();
 TAPCELL_X1 PHY_EDGE_ROW_221_Left_458 ();
 TAPCELL_X1 PHY_EDGE_ROW_222_Left_459 ();
 TAPCELL_X1 PHY_EDGE_ROW_223_Left_460 ();
 TAPCELL_X1 PHY_EDGE_ROW_224_Left_461 ();
 TAPCELL_X1 PHY_EDGE_ROW_225_Left_462 ();
 TAPCELL_X1 PHY_EDGE_ROW_226_Left_463 ();
 TAPCELL_X1 PHY_EDGE_ROW_227_Left_464 ();
 TAPCELL_X1 PHY_EDGE_ROW_228_Left_465 ();
 TAPCELL_X1 PHY_EDGE_ROW_229_Left_466 ();
 TAPCELL_X1 PHY_EDGE_ROW_230_Left_467 ();
 TAPCELL_X1 PHY_EDGE_ROW_231_Left_468 ();
 TAPCELL_X1 PHY_EDGE_ROW_232_Left_469 ();
 TAPCELL_X1 PHY_EDGE_ROW_233_Left_470 ();
 TAPCELL_X1 PHY_EDGE_ROW_234_Left_471 ();
 TAPCELL_X1 PHY_EDGE_ROW_235_Left_472 ();
 TAPCELL_X1 PHY_EDGE_ROW_236_Left_473 ();
 TAPCELL_X1 PHY_EDGE_ROW_237_Left_474 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_1_Left_475 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_2_Left_476 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_2_Left_477 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_2_Left_478 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_2_Left_479 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_2_Left_480 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_2_Left_481 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_2_Left_482 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_2_Left_483 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_2_Left_484 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_2_Left_485 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_2_Left_486 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_2_Left_487 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_2_Left_488 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_2_Left_489 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_2_Left_490 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_2_Left_491 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_2_Left_492 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_2_Left_493 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_2_Left_494 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_2_Left_495 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_2_Left_496 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_2_Left_497 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_2_Left_498 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_2_Left_499 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_2_Left_500 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_2_Left_501 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_2_Left_502 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_2_Left_503 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_2_Left_504 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_2_Left_505 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_2_Left_506 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_2_Left_507 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_2_Left_508 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_2_Left_509 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_2_Left_510 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_2_Left_511 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_2_Left_512 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_2_Left_513 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_2_Left_514 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_2_Left_515 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_2_Left_516 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_2_Left_517 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_2_Left_518 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_2_Left_519 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_2_Left_520 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_2_Left_521 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_2_Left_522 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_2_Left_523 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_2_Left_524 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_2_Left_525 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_2_Left_526 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_2_Left_527 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_2_Left_528 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_2_Left_529 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_2_Left_530 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_2_Left_531 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_2_Left_532 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_2_Left_533 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_2_Left_534 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_2_Left_535 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_2_Left_536 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_2_Left_537 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_2_Left_538 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_2_Left_539 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_2_Left_540 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_2_Left_541 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_2_Left_542 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_2_Left_543 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_2_Left_544 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_2_Left_545 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_2_Left_546 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_2_Left_547 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_2_Left_548 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_2_Left_549 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_2_Left_550 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_2_Left_551 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_2_Left_552 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_2_Left_553 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_2_Left_554 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_2_Left_555 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_2_Left_556 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_2_Left_557 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_2_Left_558 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_2_Left_559 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_2_Left_560 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_2_Left_561 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_2_Left_562 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_2_Left_563 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_2_Left_564 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_2_Left_565 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_2_Left_566 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_2_Left_567 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_2_Left_568 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_2_Left_569 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_2_Left_570 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_2_Left_571 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_2_Left_572 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_2_Left_573 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_2_Left_574 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_2_Left_575 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_2_Left_576 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_2_Left_577 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_2_Left_578 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_2_Left_579 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_2_Left_580 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_2_Left_581 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_2_Left_582 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_2_Left_583 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_2_Left_584 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_2_Left_585 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_2_Left_586 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_2_Left_587 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_2_Left_588 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_2_Left_589 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_2_Left_590 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_2_Left_591 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_2_Left_592 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_2_Left_593 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_2_Left_594 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_2_Left_595 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_2_Left_596 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_2_Left_597 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_2_Left_598 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_2_Left_599 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_2_Left_600 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_2_Left_601 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_2_Left_602 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_2_Left_603 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_2_Left_604 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_2_Left_605 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_2_Left_606 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_2_Left_607 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_2_Left_608 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_2_Left_609 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_2_Left_610 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_2_Left_611 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_2_Left_612 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_2_Left_613 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_2_Left_614 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_2_Left_615 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_2_Left_616 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_2_Left_617 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_2_Left_618 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_2_Left_619 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_2_Left_620 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_2_Left_621 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_2_Left_622 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_2_Left_623 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_2_Left_624 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_2_Left_625 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_2_Left_626 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_2_Left_627 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_2_Left_628 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_2_Left_629 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_2_Left_630 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_2_Left_631 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_2_Left_632 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_2_Left_633 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_2_Left_634 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_2_Left_635 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_2_Left_636 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_2_Left_637 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_2_Left_638 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_2_Left_639 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_2_Left_640 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_2_Left_641 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_2_Left_642 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_2_Left_643 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_1_Right_644 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_1_Right_645 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_1_Right_646 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_1_Right_647 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_1_Right_648 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_1_Right_649 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_1_Right_650 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_1_Right_651 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_1_Right_652 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_1_Right_653 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_1_Right_654 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_1_Right_655 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_1_Right_656 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_1_Right_657 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_1_Right_658 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_1_Right_659 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_1_Right_660 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_1_Right_661 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_1_Right_662 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_1_Right_663 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_1_Right_664 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_1_Right_665 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_1_Right_666 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_1_Right_667 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_1_Right_668 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_1_Right_669 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_1_Right_670 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_1_Right_671 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_1_Right_672 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_1_Right_673 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_1_Right_674 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_1_Right_675 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_1_Right_676 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_1_Right_677 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_1_Right_678 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_1_Right_679 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_1_Right_680 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_1_Right_681 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_1_Right_682 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_1_Right_683 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_1_Right_684 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_1_Right_685 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_1_Right_686 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_1_Right_687 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_1_Right_688 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_1_Right_689 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_1_Right_690 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_1_Right_691 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_1_Right_692 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_1_Right_693 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_1_Right_694 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_1_Right_695 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_1_Right_696 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_1_Right_697 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_1_Right_698 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_1_Right_699 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_1_Right_700 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_1_Right_701 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_1_Right_702 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_1_Right_703 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_1_Right_704 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_1_Right_705 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_1_Right_706 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_1_Right_707 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_1_Right_708 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_1_Right_709 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_1_Right_710 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_1_Right_711 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_1_Right_712 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_1_Right_713 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_1_Right_714 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_1_Right_715 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_1_Right_716 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_1_Right_717 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_1_Right_718 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_1_Right_719 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_1_Right_720 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_1_Right_721 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_1_Right_722 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_1_Right_723 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_1_Right_724 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_1_Right_725 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_1_Right_726 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_1_Right_727 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_1_Right_728 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_1_Right_729 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_1_Right_730 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_1_Right_731 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_1_Right_732 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_1_Right_733 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_1_Right_734 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_1_Right_735 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_1_Right_736 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_1_Right_737 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_1_Right_738 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_1_Right_739 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_1_Right_740 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_1_Right_741 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_1_Right_742 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_1_Right_743 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_1_Right_744 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_1_Right_745 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_1_Right_746 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_1_Right_747 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_1_Right_748 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_1_Right_749 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_1_Right_750 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_1_Right_751 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_1_Right_752 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_1_Right_753 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_1_Right_754 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_1_Right_755 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_1_Right_756 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_1_Right_757 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_1_Right_758 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_1_Right_759 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_1_Right_760 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_1_Right_761 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_1_Right_762 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_1_Right_763 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_1_Right_764 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_1_Right_765 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_1_Right_766 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_1_Right_767 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_1_Right_768 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_1_Right_769 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_1_Right_770 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_1_Right_771 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_1_Right_772 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_1_Right_773 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_1_Right_774 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_1_Right_775 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_1_Right_776 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_1_Right_777 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_1_Right_778 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_1_Right_779 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_1_Right_780 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_1_Right_781 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_1_Right_782 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_1_Right_783 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_1_Right_784 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_1_Right_785 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_1_Right_786 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_1_Right_787 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_1_Right_788 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_1_Right_789 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_1_Right_790 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_1_Right_791 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_1_Right_792 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_1_Right_793 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_1_Right_794 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_1_Right_795 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_1_Right_796 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_1_Right_797 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_1_Right_798 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_1_Right_799 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_1_Right_800 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_1_Right_801 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_1_Right_802 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_1_Right_803 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_1_Right_804 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_1_Right_805 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_1_Right_806 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_1_Right_807 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_1_Right_808 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_1_Right_809 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_1_Right_810 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_1_Right_811 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_812 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_813 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_814 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_815 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_816 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_817 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_818 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_819 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_820 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_821 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_822 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_823 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_824 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_825 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_826 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_827 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_828 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_829 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_830 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_831 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_832 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_833 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_834 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_835 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_836 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_837 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_838 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_839 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_840 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_841 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_842 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_843 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_844 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_845 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_846 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_847 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_848 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_849 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_850 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_851 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_852 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_853 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_208_854 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_208_855 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_209_856 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_210_857 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_211_858 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_212_859 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_213_860 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_214_861 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_215_862 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_216_863 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_217_864 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_218_865 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_219_866 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_220_867 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_221_868 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_222_869 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_223_870 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_224_871 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_225_872 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_226_873 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_227_874 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_228_875 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_229_876 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_230_877 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_231_878 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_232_879 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_233_880 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_234_881 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_235_882 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_236_883 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_237_884 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_237_885 ();
 BUF_X16 max_length9 (.A(net10),
    .Z(net9));
 BUF_X16 max_length10 (.A(_0303_),
    .Z(net10));
 BUF_X16 wire11 (.A(net12),
    .Z(net11));
 BUF_X16 wire12 (.A(net47),
    .Z(net12));
 BUF_X4 input13 (.A(data_in[0]),
    .Z(net13));
 BUF_X4 input14 (.A(data_in[10]),
    .Z(net14));
 BUF_X1 input15 (.A(data_in[11]),
    .Z(net15));
 BUF_X2 input16 (.A(data_in[12]),
    .Z(net16));
 BUF_X4 input17 (.A(data_in[13]),
    .Z(net17));
 BUF_X4 input18 (.A(data_in[14]),
    .Z(net18));
 BUF_X1 input19 (.A(data_in[15]),
    .Z(net19));
 BUF_X1 input20 (.A(data_in[16]),
    .Z(net20));
 CLKBUF_X3 input21 (.A(data_in[17]),
    .Z(net21));
 BUF_X1 input22 (.A(data_in[18]),
    .Z(net22));
 BUF_X2 input23 (.A(data_in[19]),
    .Z(net23));
 BUF_X1 input24 (.A(data_in[1]),
    .Z(net24));
 BUF_X1 input25 (.A(data_in[20]),
    .Z(net25));
 BUF_X1 input26 (.A(data_in[21]),
    .Z(net26));
 BUF_X4 input27 (.A(data_in[22]),
    .Z(net27));
 BUF_X4 input28 (.A(data_in[23]),
    .Z(net28));
 BUF_X1 input29 (.A(data_in[24]),
    .Z(net29));
 BUF_X2 input30 (.A(data_in[25]),
    .Z(net30));
 CLKBUF_X3 input31 (.A(data_in[26]),
    .Z(net31));
 CLKBUF_X3 input32 (.A(data_in[27]),
    .Z(net32));
 BUF_X1 input33 (.A(data_in[28]),
    .Z(net33));
 BUF_X1 input34 (.A(data_in[29]),
    .Z(net34));
 BUF_X2 input35 (.A(data_in[2]),
    .Z(net35));
 BUF_X1 input36 (.A(data_in[30]),
    .Z(net36));
 CLKBUF_X3 input37 (.A(data_in[31]),
    .Z(net37));
 BUF_X4 input38 (.A(data_in[3]),
    .Z(net38));
 BUF_X4 input39 (.A(data_in[4]),
    .Z(net39));
 BUF_X4 input40 (.A(data_in[5]),
    .Z(net40));
 BUF_X1 input41 (.A(data_in[6]),
    .Z(net41));
 BUF_X1 input42 (.A(data_in[7]),
    .Z(net42));
 BUF_X4 input43 (.A(data_in[8]),
    .Z(net43));
 BUF_X4 input44 (.A(data_in[9]),
    .Z(net44));
 BUF_X4 input45 (.A(init_enable),
    .Z(net45));
 BUF_X4 input46 (.A(pe_ce),
    .Z(net46));
 BUF_X4 input47 (.A(rst_n),
    .Z(net47));
 BUF_X1 output48 (.A(net48),
    .Z(curr_state[1]));
 BUF_X1 output49 (.A(net49),
    .Z(data_out[0]));
 BUF_X1 output50 (.A(net50),
    .Z(data_out[10]));
 BUF_X1 output51 (.A(net51),
    .Z(data_out[11]));
 BUF_X1 output52 (.A(net52),
    .Z(data_out[12]));
 BUF_X1 output53 (.A(net53),
    .Z(data_out[13]));
 BUF_X1 output54 (.A(net54),
    .Z(data_out[14]));
 BUF_X1 output55 (.A(net55),
    .Z(data_out[15]));
 BUF_X1 output56 (.A(net56),
    .Z(data_out[16]));
 BUF_X1 output57 (.A(net57),
    .Z(data_out[17]));
 BUF_X1 output58 (.A(net58),
    .Z(data_out[18]));
 BUF_X1 output59 (.A(net59),
    .Z(data_out[19]));
 BUF_X1 output60 (.A(net60),
    .Z(data_out[1]));
 BUF_X1 output61 (.A(net61),
    .Z(data_out[20]));
 BUF_X1 output62 (.A(net62),
    .Z(data_out[21]));
 BUF_X1 output63 (.A(net63),
    .Z(data_out[22]));
 BUF_X1 output64 (.A(net64),
    .Z(data_out[23]));
 BUF_X1 output65 (.A(net65),
    .Z(data_out[24]));
 BUF_X1 output66 (.A(net66),
    .Z(data_out[25]));
 BUF_X1 output67 (.A(net67),
    .Z(data_out[26]));
 BUF_X1 output68 (.A(net68),
    .Z(data_out[27]));
 BUF_X1 output69 (.A(net69),
    .Z(data_out[28]));
 BUF_X1 output70 (.A(net70),
    .Z(data_out[29]));
 BUF_X1 output71 (.A(net71),
    .Z(data_out[2]));
 BUF_X1 output72 (.A(net72),
    .Z(data_out[30]));
 BUF_X1 output73 (.A(net73),
    .Z(data_out[31]));
 BUF_X1 output74 (.A(net74),
    .Z(data_out[32]));
 BUF_X1 output75 (.A(net75),
    .Z(data_out[33]));
 BUF_X1 output76 (.A(net76),
    .Z(data_out[34]));
 BUF_X1 output77 (.A(net77),
    .Z(data_out[35]));
 BUF_X1 output78 (.A(net78),
    .Z(data_out[36]));
 BUF_X1 output79 (.A(net79),
    .Z(data_out[37]));
 BUF_X1 output80 (.A(net80),
    .Z(data_out[38]));
 BUF_X1 output81 (.A(net81),
    .Z(data_out[39]));
 BUF_X1 output82 (.A(net82),
    .Z(data_out[3]));
 BUF_X1 output83 (.A(net83),
    .Z(data_out[40]));
 BUF_X1 output84 (.A(net84),
    .Z(data_out[41]));
 BUF_X1 output85 (.A(net85),
    .Z(data_out[42]));
 BUF_X1 output86 (.A(net86),
    .Z(data_out[43]));
 BUF_X1 output87 (.A(net87),
    .Z(data_out[44]));
 BUF_X1 output88 (.A(net88),
    .Z(data_out[45]));
 BUF_X1 output89 (.A(net89),
    .Z(data_out[46]));
 BUF_X1 output90 (.A(net90),
    .Z(data_out[47]));
 BUF_X1 output91 (.A(net91),
    .Z(data_out[48]));
 BUF_X1 output92 (.A(net92),
    .Z(data_out[49]));
 BUF_X1 output93 (.A(net93),
    .Z(data_out[4]));
 BUF_X1 output94 (.A(net94),
    .Z(data_out[50]));
 BUF_X1 output95 (.A(net95),
    .Z(data_out[51]));
 BUF_X1 output96 (.A(net96),
    .Z(data_out[52]));
 BUF_X1 output97 (.A(net97),
    .Z(data_out[53]));
 BUF_X1 output98 (.A(net98),
    .Z(data_out[54]));
 BUF_X1 output99 (.A(net99),
    .Z(data_out[55]));
 BUF_X1 output100 (.A(net100),
    .Z(data_out[56]));
 BUF_X1 output101 (.A(net101),
    .Z(data_out[57]));
 BUF_X1 output102 (.A(net102),
    .Z(data_out[58]));
 BUF_X1 output103 (.A(net103),
    .Z(data_out[59]));
 BUF_X1 output104 (.A(net104),
    .Z(data_out[5]));
 BUF_X1 output105 (.A(net105),
    .Z(data_out[60]));
 BUF_X1 output106 (.A(net106),
    .Z(data_out[61]));
 BUF_X1 output107 (.A(net107),
    .Z(data_out[62]));
 BUF_X1 output108 (.A(net108),
    .Z(data_out[63]));
 BUF_X1 output109 (.A(net109),
    .Z(data_out[6]));
 BUF_X1 output110 (.A(net110),
    .Z(data_out[7]));
 BUF_X1 output111 (.A(net111),
    .Z(data_out[8]));
 BUF_X1 output112 (.A(net112),
    .Z(data_out[9]));
 BUF_X1 output113 (.A(net113),
    .Z(valid_reg_out));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_17_1__18__114  (.Z(net114));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_17_1__25__115  (.Z(net115));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_19_2__18__116  (.Z(net116));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_19_2__25__117  (.Z(net117));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_21_3__18__118  (.Z(net118));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_21_3__25__119  (.Z(net119));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_23_4__18__120  (.Z(net120));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_23_4__25__121  (.Z(net121));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_25_5__18__122  (.Z(net122));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_25_5__25__123  (.Z(net123));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_27_6__18__124  (.Z(net124));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_27_6__25__125  (.Z(net125));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_29_7__18__126  (.Z(net126));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_29_7__25__127  (.Z(net127));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_31_8__18__128  (.Z(net128));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_31_8__25__129  (.Z(net129));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_32_8__23__130  (.Z(net130));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_32_8__24__131  (.Z(net131));
 LOGIC0_X1 u_multiplier_STAGE2_E_4_2_pp2_13_3__18__134  (.Z(net134));
 LOGIC0_X1 u_multiplier_STAGE2_E_4_2_pp2_13_3__25__135  (.Z(net135));
 LOGIC0_X1 u_multiplier_STAGE2_E_4_2_pp2_15_4__18__136  (.Z(net136));
 LOGIC0_X1 u_multiplier_STAGE2_E_4_2_pp2_15_4__25__137  (.Z(net137));
 LOGIC0_X1 u_multiplier_STAGE2_E_4_2_pp2_9_1__18__138  (.Z(net138));
 LOGIC0_X1 u_multiplier_STAGE2_E_4_2_pp2_9_1__25__139  (.Z(net139));
 LOGIC0_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__56__141  (.Z(net141));
 LOGIC0_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__57__142  (.Z(net142));
 LOGIC0_X1 u_multiplier_STAGE3_E_4_2_pp3_5_1__18__143  (.Z(net143));
 LOGIC0_X1 u_multiplier_STAGE3_E_4_2_pp3_5_1__25__144  (.Z(net144));
 LOGIC0_X1 u_multiplier_STAGE3_E_4_2_pp3_7_2__18__145  (.Z(net145));
 LOGIC0_X1 u_multiplier_STAGE3_E_4_2_pp3_7_2__25__146  (.Z(net146));
 LOGIC0_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__41__148  (.Z(net148));
 LOGIC0_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__42__149  (.Z(net149));
 LOGIC0_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__45__150  (.Z(net150));
 LOGIC0_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__46__151  (.Z(net151));
 LOGIC0_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__47__152  (.Z(net152));
 LOGIC0_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__50__153  (.Z(net153));
 LOGIC0_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__51__154  (.Z(net154));
 LOGIC0_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__52__155  (.Z(net155));
 LOGIC0_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__55__156  (.Z(net156));
 LOGIC0_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__56__157  (.Z(net157));
 LOGIC0_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__57__158  (.Z(net158));
 LOGIC0_X1 u_multiplier_STAGE4_E_4_2_pp4_2__23__159  (.Z(net159));
 LOGIC0_X1 u_multiplier_STAGE4_E_4_2_pp4_2__24__160  (.Z(net160));
 LOGIC0_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__44__162  (.Z(net162));
 CLKBUF_X1 hold164 (.A(_0304_),
    .Z(net164));
 CLKBUF_X1 hold165 (.A(net1),
    .Z(net165));
 CLKBUF_X1 hold166 (.A(net184),
    .Z(net166));
 CLKBUF_X1 hold167 (.A(net189),
    .Z(net167));
 CLKBUF_X1 hold168 (.A(net192),
    .Z(net168));
 CLKBUF_X1 hold169 (.A(net3),
    .Z(net169));
 CLKBUF_X1 hold170 (.A(net195),
    .Z(net170));
 CLKBUF_X1 hold171 (.A(net5),
    .Z(net171));
 CLKBUF_X1 hold172 (.A(net182),
    .Z(net172));
 CLKBUF_X1 hold173 (.A(net203),
    .Z(net173));
 CLKBUF_X1 hold174 (.A(net187),
    .Z(net174));
 CLKBUF_X1 hold175 (.A(net198),
    .Z(net175));
 CLKBUF_X1 hold176 (.A(net208),
    .Z(net176));
 CLKBUF_X1 hold177 (.A(net211),
    .Z(net177));
 CLKBUF_X1 hold178 (.A(net213),
    .Z(net178));
 CLKBUF_X1 hold179 (.A(net215),
    .Z(net179));
 CLKBUF_X1 hold180 (.A(net216),
    .Z(net180));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_1_0_0_clk));
 CLKBUF_X3 clkbuf_1_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_1_1_0_clk));
 CLKBUF_X3 clkbuf_2_0_0_clk (.A(clknet_1_0_0_clk),
    .Z(clknet_2_0_0_clk));
 CLKBUF_X3 clkbuf_2_1_0_clk (.A(clknet_1_0_0_clk),
    .Z(clknet_2_1_0_clk));
 CLKBUF_X3 clkbuf_2_2_0_clk (.A(clknet_1_1_0_clk),
    .Z(clknet_2_2_0_clk));
 CLKBUF_X3 clkbuf_2_3_0_clk (.A(clknet_1_1_0_clk),
    .Z(clknet_2_3_0_clk));
 CLKBUF_X3 clkbuf_3_0_0_clk (.A(clknet_2_0_0_clk),
    .Z(clknet_3_0_0_clk));
 CLKBUF_X3 clkbuf_3_1_0_clk (.A(clknet_2_0_0_clk),
    .Z(clknet_3_1_0_clk));
 CLKBUF_X3 clkbuf_3_2_0_clk (.A(clknet_2_1_0_clk),
    .Z(clknet_3_2_0_clk));
 CLKBUF_X3 clkbuf_3_3_0_clk (.A(clknet_2_1_0_clk),
    .Z(clknet_3_3_0_clk));
 CLKBUF_X3 clkbuf_3_4_0_clk (.A(clknet_2_2_0_clk),
    .Z(clknet_3_4_0_clk));
 CLKBUF_X3 clkbuf_3_5_0_clk (.A(clknet_2_2_0_clk),
    .Z(clknet_3_5_0_clk));
 CLKBUF_X3 clkbuf_3_6_0_clk (.A(clknet_2_3_0_clk),
    .Z(clknet_3_6_0_clk));
 CLKBUF_X3 clkbuf_3_7_0_clk (.A(clknet_2_3_0_clk),
    .Z(clknet_3_7_0_clk));
 CLKBUF_X3 clkbuf_4_0__f_clk (.A(clknet_3_0_0_clk),
    .Z(clknet_4_0__leaf_clk));
 CLKBUF_X3 clkbuf_4_1__f_clk (.A(clknet_3_0_0_clk),
    .Z(clknet_4_1__leaf_clk));
 CLKBUF_X3 clkbuf_4_2__f_clk (.A(clknet_3_1_0_clk),
    .Z(clknet_4_2__leaf_clk));
 CLKBUF_X3 clkbuf_4_3__f_clk (.A(clknet_3_1_0_clk),
    .Z(clknet_4_3__leaf_clk));
 CLKBUF_X3 clkbuf_4_4__f_clk (.A(clknet_3_2_0_clk),
    .Z(clknet_4_4__leaf_clk));
 CLKBUF_X3 clkbuf_4_5__f_clk (.A(clknet_3_2_0_clk),
    .Z(clknet_4_5__leaf_clk));
 CLKBUF_X3 clkbuf_4_6__f_clk (.A(clknet_3_3_0_clk),
    .Z(clknet_4_6__leaf_clk));
 CLKBUF_X3 clkbuf_4_7__f_clk (.A(clknet_3_3_0_clk),
    .Z(clknet_4_7__leaf_clk));
 CLKBUF_X3 clkbuf_4_8__f_clk (.A(clknet_3_4_0_clk),
    .Z(clknet_4_8__leaf_clk));
 CLKBUF_X3 clkbuf_4_9__f_clk (.A(clknet_3_4_0_clk),
    .Z(clknet_4_9__leaf_clk));
 CLKBUF_X3 clkbuf_4_10__f_clk (.A(clknet_3_5_0_clk),
    .Z(clknet_4_10__leaf_clk));
 CLKBUF_X3 clkbuf_4_11__f_clk (.A(clknet_3_5_0_clk),
    .Z(clknet_4_11__leaf_clk));
 CLKBUF_X3 clkbuf_4_12__f_clk (.A(clknet_3_6_0_clk),
    .Z(clknet_4_12__leaf_clk));
 CLKBUF_X3 clkbuf_4_13__f_clk (.A(clknet_3_6_0_clk),
    .Z(clknet_4_13__leaf_clk));
 CLKBUF_X3 clkbuf_4_14__f_clk (.A(clknet_3_7_0_clk),
    .Z(clknet_4_14__leaf_clk));
 CLKBUF_X3 clkbuf_4_15__f_clk (.A(clknet_3_7_0_clk),
    .Z(clknet_4_15__leaf_clk));
 INV_X2 clkload0 (.A(clknet_4_1__leaf_clk));
 INV_X2 clkload1 (.A(clknet_4_3__leaf_clk));
 CLKBUF_X1 clkload2 (.A(clknet_4_4__leaf_clk));
 CLKBUF_X1 clkload3 (.A(clknet_4_6__leaf_clk));
 INV_X1 clkload4 (.A(clknet_4_8__leaf_clk));
 INV_X2 clkload5 (.A(clknet_4_11__leaf_clk));
 INV_X2 clkload6 (.A(clknet_4_12__leaf_clk));
 CLKBUF_X1 clkload7 (.A(clknet_4_15__leaf_clk));
 CLKBUF_X1 hold1 (.A(_0651_),
    .Z(net1));
 CLKBUF_X1 hold2 (.A(net165),
    .Z(net2));
 CLKBUF_X1 hold3 (.A(addr_ptr[3]),
    .Z(net3));
 CLKBUF_X1 hold4 (.A(net169),
    .Z(net4));
 CLKBUF_X1 hold5 (.A(addr_ptr[2]),
    .Z(net5));
 CLKBUF_X1 hold6 (.A(net171),
    .Z(net6));
 CLKBUF_X1 hold7 (.A(_0655_),
    .Z(net7));
 CLKBUF_X1 hold8 (.A(_0419_),
    .Z(net8));
 CLKBUF_X1 hold9 (.A(_0168_),
    .Z(net181));
 CLKBUF_X1 hold10 (.A(addr_ptr[4]),
    .Z(net182));
 CLKBUF_X1 hold11 (.A(net172),
    .Z(net183));
 CLKBUF_X1 hold12 (.A(_0656_),
    .Z(net184));
 CLKBUF_X1 hold13 (.A(net166),
    .Z(net185));
 CLKBUF_X1 hold14 (.A(_0265_),
    .Z(net186));
 CLKBUF_X1 hold15 (.A(addr_ptr[5]),
    .Z(net187));
 CLKBUF_X1 hold16 (.A(net174),
    .Z(net188));
 CLKBUF_X1 hold17 (.A(_0661_),
    .Z(net189));
 CLKBUF_X1 hold18 (.A(net167),
    .Z(net190));
 CLKBUF_X1 hold19 (.A(_0270_),
    .Z(net191));
 CLKBUF_X1 hold20 (.A(_0658_),
    .Z(net192));
 CLKBUF_X1 hold21 (.A(net168),
    .Z(net193));
 CLKBUF_X1 hold22 (.A(_0267_),
    .Z(net194));
 CLKBUF_X1 hold23 (.A(_0660_),
    .Z(net195));
 CLKBUF_X1 hold24 (.A(net170),
    .Z(net196));
 CLKBUF_X1 hold25 (.A(_0269_),
    .Z(net197));
 CLKBUF_X1 hold26 (.A(_0657_),
    .Z(net198));
 CLKBUF_X1 hold27 (.A(net175),
    .Z(net199));
 CLKBUF_X1 hold28 (.A(curr_state[0]),
    .Z(net200));
 CLKBUF_X1 hold29 (.A(_0384_),
    .Z(net201));
 CLKBUF_X1 hold30 (.A(_0306_),
    .Z(net202));
 CLKBUF_X1 hold31 (.A(_0659_),
    .Z(net203));
 CLKBUF_X1 hold32 (.A(net173),
    .Z(net204));
 CLKBUF_X1 hold33 (.A(_0268_),
    .Z(net205));
 CLKBUF_X1 hold34 (.A(_0654_),
    .Z(net206));
 CLKBUF_X1 hold35 (.A(_0418_),
    .Z(net207));
 CLKBUF_X1 hold36 (.A(_0650_),
    .Z(net208));
 CLKBUF_X1 hold37 (.A(_0405_),
    .Z(net209));
 CLKBUF_X1 hold38 (.A(_0163_),
    .Z(net210));
 CLKBUF_X1 hold39 (.A(addr_ptr[1]),
    .Z(net211));
 CLKBUF_X1 hold40 (.A(net177),
    .Z(net212));
 CLKBUF_X1 hold41 (.A(_0652_),
    .Z(net213));
 CLKBUF_X1 hold42 (.A(net178),
    .Z(net214));
 CLKBUF_X1 hold43 (.A(addr_ptr[0]),
    .Z(net215));
 CLKBUF_X1 hold44 (.A(_0653_),
    .Z(net216));
 CLKBUF_X1 hold45 (.A(_0518_),
    .Z(net217));
 CLKBUF_X1 hold46 (.A(data_in_reg[15]),
    .Z(net218));
 CLKBUF_X1 hold47 (.A(data_in_reg[6]),
    .Z(net219));
 CLKBUF_X1 hold48 (.A(curr_state[2]),
    .Z(net220));
 CLKBUF_X1 hold49 (.A(data_in_reg[2]),
    .Z(net221));
 CLKBUF_X1 hold50 (.A(data_in_reg[0]),
    .Z(net222));
 CLKBUF_X1 hold51 (.A(data_in_reg[12]),
    .Z(net223));
 CLKBUF_X1 hold52 (.A(data_in_reg[31]),
    .Z(net224));
 CLKBUF_X1 hold53 (.A(data_in_reg[14]),
    .Z(net225));
 CLKBUF_X1 hold54 (.A(data_in_reg[24]),
    .Z(net226));
 CLKBUF_X1 hold55 (.A(data_in_reg[28]),
    .Z(net227));
 CLKBUF_X1 hold56 (.A(data_in_reg[22]),
    .Z(net228));
 CLKBUF_X1 hold57 (.A(data_in_reg[1]),
    .Z(net229));
 CLKBUF_X1 hold58 (.A(data_in_reg[18]),
    .Z(net230));
 CLKBUF_X1 hold59 (.A(data_in_reg[29]),
    .Z(net231));
 CLKBUF_X1 hold60 (.A(data_in_reg[10]),
    .Z(net232));
 CLKBUF_X1 hold61 (.A(init_count[5]),
    .Z(net233));
 CLKBUF_X1 hold62 (.A(init_count[4]),
    .Z(net234));
 FILLCELL_X4 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_8 ();
 FILLCELL_X8 FILLER_0_40 ();
 FILLCELL_X2 FILLER_0_48 ();
 FILLCELL_X16 FILLER_0_53 ();
 FILLCELL_X8 FILLER_0_69 ();
 FILLCELL_X2 FILLER_0_77 ();
 FILLCELL_X1 FILLER_0_79 ();
 FILLCELL_X16 FILLER_0_84 ();
 FILLCELL_X4 FILLER_0_100 ();
 FILLCELL_X2 FILLER_0_104 ();
 FILLCELL_X1 FILLER_0_106 ();
 FILLCELL_X8 FILLER_0_110 ();
 FILLCELL_X1 FILLER_0_118 ();
 FILLCELL_X4 FILLER_0_123 ();
 FILLCELL_X16 FILLER_0_130 ();
 FILLCELL_X4 FILLER_0_146 ();
 FILLCELL_X1 FILLER_0_150 ();
 FILLCELL_X4 FILLER_0_154 ();
 FILLCELL_X2 FILLER_0_158 ();
 FILLCELL_X1 FILLER_0_160 ();
 FILLCELL_X16 FILLER_0_164 ();
 FILLCELL_X8 FILLER_0_180 ();
 FILLCELL_X4 FILLER_0_188 ();
 FILLCELL_X16 FILLER_0_195 ();
 FILLCELL_X8 FILLER_0_211 ();
 FILLCELL_X4 FILLER_0_219 ();
 FILLCELL_X16 FILLER_0_226 ();
 FILLCELL_X2 FILLER_0_242 ();
 FILLCELL_X4 FILLER_0_246 ();
 FILLCELL_X4 FILLER_0_253 ();
 FILLCELL_X1 FILLER_0_257 ();
 FILLCELL_X4 FILLER_0_261 ();
 FILLCELL_X16 FILLER_0_268 ();
 FILLCELL_X8 FILLER_0_284 ();
 FILLCELL_X8 FILLER_0_296 ();
 FILLCELL_X1 FILLER_0_304 ();
 FILLCELL_X8 FILLER_0_309 ();
 FILLCELL_X2 FILLER_0_317 ();
 FILLCELL_X1 FILLER_0_319 ();
 FILLCELL_X8 FILLER_0_323 ();
 FILLCELL_X4 FILLER_0_334 ();
 FILLCELL_X4 FILLER_0_347 ();
 FILLCELL_X1 FILLER_0_351 ();
 FILLCELL_X4 FILLER_0_355 ();
 FILLCELL_X8 FILLER_0_366 ();
 FILLCELL_X2 FILLER_0_374 ();
 FILLCELL_X1 FILLER_0_376 ();
 FILLCELL_X4 FILLER_0_384 ();
 FILLCELL_X2 FILLER_0_388 ();
 FILLCELL_X4 FILLER_0_393 ();
 FILLCELL_X2 FILLER_0_397 ();
 FILLCELL_X4 FILLER_0_402 ();
 FILLCELL_X8 FILLER_0_409 ();
 FILLCELL_X4 FILLER_0_417 ();
 FILLCELL_X2 FILLER_0_421 ();
 FILLCELL_X8 FILLER_0_425 ();
 FILLCELL_X4 FILLER_0_433 ();
 FILLCELL_X1 FILLER_0_437 ();
 FILLCELL_X4 FILLER_0_441 ();
 FILLCELL_X4 FILLER_0_448 ();
 FILLCELL_X1 FILLER_0_452 ();
 FILLCELL_X16 FILLER_0_456 ();
 FILLCELL_X1 FILLER_0_472 ();
 FILLCELL_X4 FILLER_0_479 ();
 FILLCELL_X4 FILLER_0_486 ();
 FILLCELL_X1 FILLER_0_490 ();
 FILLCELL_X16 FILLER_0_495 ();
 FILLCELL_X2 FILLER_0_511 ();
 FILLCELL_X8 FILLER_0_516 ();
 FILLCELL_X16 FILLER_0_528 ();
 FILLCELL_X1 FILLER_0_544 ();
 FILLCELL_X8 FILLER_0_549 ();
 FILLCELL_X1 FILLER_0_557 ();
 FILLCELL_X4 FILLER_0_561 ();
 FILLCELL_X4 FILLER_0_568 ();
 FILLCELL_X1 FILLER_0_572 ();
 FILLCELL_X8 FILLER_0_576 ();
 FILLCELL_X2 FILLER_0_584 ();
 FILLCELL_X1 FILLER_0_586 ();
 FILLCELL_X8 FILLER_0_592 ();
 FILLCELL_X2 FILLER_0_600 ();
 FILLCELL_X4 FILLER_0_605 ();
 FILLCELL_X4 FILLER_0_612 ();
 FILLCELL_X1 FILLER_0_616 ();
 FILLCELL_X4 FILLER_0_620 ();
 FILLCELL_X4 FILLER_0_627 ();
 FILLCELL_X8 FILLER_0_632 ();
 FILLCELL_X2 FILLER_0_640 ();
 FILLCELL_X16 FILLER_0_645 ();
 FILLCELL_X2 FILLER_0_661 ();
 FILLCELL_X1 FILLER_0_663 ();
 FILLCELL_X4 FILLER_0_667 ();
 FILLCELL_X1 FILLER_0_671 ();
 FILLCELL_X8 FILLER_0_676 ();
 FILLCELL_X4 FILLER_0_688 ();
 FILLCELL_X2 FILLER_0_692 ();
 FILLCELL_X1 FILLER_0_694 ();
 FILLCELL_X4 FILLER_0_698 ();
 FILLCELL_X4 FILLER_0_706 ();
 FILLCELL_X8 FILLER_0_717 ();
 FILLCELL_X4 FILLER_0_725 ();
 FILLCELL_X2 FILLER_0_729 ();
 FILLCELL_X1 FILLER_0_731 ();
 FILLCELL_X8 FILLER_0_736 ();
 FILLCELL_X2 FILLER_0_744 ();
 FILLCELL_X4 FILLER_0_749 ();
 FILLCELL_X4 FILLER_0_757 ();
 FILLCELL_X4 FILLER_0_765 ();
 FILLCELL_X2 FILLER_0_769 ();
 FILLCELL_X4 FILLER_0_775 ();
 FILLCELL_X16 FILLER_0_782 ();
 FILLCELL_X2 FILLER_0_798 ();
 FILLCELL_X4 FILLER_0_802 ();
 FILLCELL_X8 FILLER_0_810 ();
 FILLCELL_X4 FILLER_0_823 ();
 FILLCELL_X1 FILLER_0_827 ();
 FILLCELL_X4 FILLER_0_831 ();
 FILLCELL_X1 FILLER_0_835 ();
 FILLCELL_X4 FILLER_0_840 ();
 FILLCELL_X4 FILLER_0_847 ();
 FILLCELL_X1 FILLER_0_851 ();
 FILLCELL_X4 FILLER_0_856 ();
 FILLCELL_X1 FILLER_0_860 ();
 FILLCELL_X4 FILLER_0_868 ();
 FILLCELL_X8 FILLER_0_874 ();
 FILLCELL_X4 FILLER_0_882 ();
 FILLCELL_X2 FILLER_0_886 ();
 FILLCELL_X1 FILLER_0_888 ();
 FILLCELL_X4 FILLER_0_893 ();
 FILLCELL_X2 FILLER_0_897 ();
 FILLCELL_X32 FILLER_0_902 ();
 FILLCELL_X8 FILLER_0_934 ();
 FILLCELL_X4 FILLER_0_942 ();
 FILLCELL_X2 FILLER_0_946 ();
 FILLCELL_X4 FILLER_0_951 ();
 FILLCELL_X8 FILLER_0_959 ();
 FILLCELL_X2 FILLER_0_967 ();
 FILLCELL_X1 FILLER_0_969 ();
 FILLCELL_X4 FILLER_0_974 ();
 FILLCELL_X16 FILLER_0_981 ();
 FILLCELL_X8 FILLER_0_1004 ();
 FILLCELL_X1 FILLER_0_1012 ();
 FILLCELL_X4 FILLER_0_1015 ();
 FILLCELL_X4 FILLER_0_1023 ();
 FILLCELL_X8 FILLER_0_1031 ();
 FILLCELL_X1 FILLER_0_1039 ();
 FILLCELL_X4 FILLER_0_1043 ();
 FILLCELL_X1 FILLER_0_1047 ();
 FILLCELL_X4 FILLER_0_1052 ();
 FILLCELL_X4 FILLER_0_1059 ();
 FILLCELL_X4 FILLER_0_1067 ();
 FILLCELL_X8 FILLER_0_1074 ();
 FILLCELL_X2 FILLER_0_1082 ();
 FILLCELL_X1 FILLER_0_1084 ();
 FILLCELL_X8 FILLER_0_1088 ();
 FILLCELL_X2 FILLER_0_1096 ();
 FILLCELL_X4 FILLER_0_1100 ();
 FILLCELL_X4 FILLER_0_1107 ();
 FILLCELL_X8 FILLER_0_1114 ();
 FILLCELL_X4 FILLER_0_1125 ();
 FILLCELL_X8 FILLER_0_1133 ();
 FILLCELL_X1 FILLER_0_1141 ();
 FILLCELL_X4 FILLER_0_1151 ();
 FILLCELL_X4 FILLER_0_1158 ();
 FILLCELL_X4 FILLER_0_1165 ();
 FILLCELL_X2 FILLER_0_1169 ();
 FILLCELL_X1 FILLER_0_1171 ();
 FILLCELL_X4 FILLER_0_1175 ();
 FILLCELL_X4 FILLER_0_1183 ();
 FILLCELL_X4 FILLER_0_1191 ();
 FILLCELL_X4 FILLER_0_1198 ();
 FILLCELL_X8 FILLER_0_1205 ();
 FILLCELL_X8 FILLER_0_1222 ();
 FILLCELL_X4 FILLER_0_1230 ();
 FILLCELL_X8 FILLER_0_1238 ();
 FILLCELL_X4 FILLER_0_1246 ();
 FILLCELL_X1 FILLER_0_1250 ();
 FILLCELL_X4 FILLER_0_1258 ();
 FILLCELL_X32 FILLER_0_1263 ();
 FILLCELL_X16 FILLER_0_1295 ();
 FILLCELL_X8 FILLER_0_1311 ();
 FILLCELL_X4 FILLER_0_1319 ();
 FILLCELL_X16 FILLER_0_1326 ();
 FILLCELL_X1 FILLER_0_1342 ();
 FILLCELL_X16 FILLER_0_1347 ();
 FILLCELL_X2 FILLER_0_1363 ();
 FILLCELL_X16 FILLER_0_1369 ();
 FILLCELL_X8 FILLER_0_1385 ();
 FILLCELL_X1 FILLER_0_1393 ();
 FILLCELL_X32 FILLER_0_1397 ();
 FILLCELL_X32 FILLER_0_1429 ();
 FILLCELL_X4 FILLER_0_1461 ();
 FILLCELL_X32 FILLER_0_1468 ();
 FILLCELL_X32 FILLER_0_1500 ();
 FILLCELL_X4 FILLER_0_1532 ();
 FILLCELL_X32 FILLER_0_1539 ();
 FILLCELL_X32 FILLER_0_1571 ();
 FILLCELL_X2 FILLER_0_1603 ();
 FILLCELL_X1 FILLER_0_1605 ();
 FILLCELL_X32 FILLER_0_1610 ();
 FILLCELL_X32 FILLER_0_1642 ();
 FILLCELL_X2 FILLER_0_1674 ();
 FILLCELL_X1 FILLER_0_1676 ();
 FILLCELL_X32 FILLER_0_1680 ();
 FILLCELL_X32 FILLER_0_1712 ();
 FILLCELL_X4 FILLER_0_1744 ();
 FILLCELL_X8 FILLER_0_1751 ();
 FILLCELL_X2 FILLER_0_1759 ();
 FILLCELL_X1 FILLER_0_1761 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X16 FILLER_1_33 ();
 FILLCELL_X2 FILLER_1_49 ();
 FILLCELL_X4 FILLER_1_55 ();
 FILLCELL_X4 FILLER_1_78 ();
 FILLCELL_X4 FILLER_1_92 ();
 FILLCELL_X2 FILLER_1_96 ();
 FILLCELL_X1 FILLER_1_98 ();
 FILLCELL_X4 FILLER_1_103 ();
 FILLCELL_X8 FILLER_1_116 ();
 FILLCELL_X1 FILLER_1_124 ();
 FILLCELL_X8 FILLER_1_144 ();
 FILLCELL_X2 FILLER_1_152 ();
 FILLCELL_X4 FILLER_1_163 ();
 FILLCELL_X4 FILLER_1_176 ();
 FILLCELL_X1 FILLER_1_180 ();
 FILLCELL_X4 FILLER_1_185 ();
 FILLCELL_X4 FILLER_1_206 ();
 FILLCELL_X2 FILLER_1_210 ();
 FILLCELL_X4 FILLER_1_216 ();
 FILLCELL_X4 FILLER_1_230 ();
 FILLCELL_X2 FILLER_1_234 ();
 FILLCELL_X4 FILLER_1_243 ();
 FILLCELL_X1 FILLER_1_247 ();
 FILLCELL_X4 FILLER_1_258 ();
 FILLCELL_X8 FILLER_1_271 ();
 FILLCELL_X1 FILLER_1_279 ();
 FILLCELL_X4 FILLER_1_283 ();
 FILLCELL_X4 FILLER_1_291 ();
 FILLCELL_X4 FILLER_1_304 ();
 FILLCELL_X4 FILLER_1_317 ();
 FILLCELL_X2 FILLER_1_321 ();
 FILLCELL_X1 FILLER_1_323 ();
 FILLCELL_X4 FILLER_1_327 ();
 FILLCELL_X8 FILLER_1_341 ();
 FILLCELL_X4 FILLER_1_359 ();
 FILLCELL_X4 FILLER_1_373 ();
 FILLCELL_X2 FILLER_1_377 ();
 FILLCELL_X1 FILLER_1_379 ();
 FILLCELL_X4 FILLER_1_382 ();
 FILLCELL_X8 FILLER_1_396 ();
 FILLCELL_X4 FILLER_1_414 ();
 FILLCELL_X4 FILLER_1_422 ();
 FILLCELL_X1 FILLER_1_426 ();
 FILLCELL_X4 FILLER_1_437 ();
 FILLCELL_X1 FILLER_1_441 ();
 FILLCELL_X8 FILLER_1_451 ();
 FILLCELL_X4 FILLER_1_463 ();
 FILLCELL_X4 FILLER_1_474 ();
 FILLCELL_X2 FILLER_1_478 ();
 FILLCELL_X4 FILLER_1_486 ();
 FILLCELL_X4 FILLER_1_509 ();
 FILLCELL_X4 FILLER_1_522 ();
 FILLCELL_X4 FILLER_1_535 ();
 FILLCELL_X4 FILLER_1_543 ();
 FILLCELL_X4 FILLER_1_556 ();
 FILLCELL_X2 FILLER_1_560 ();
 FILLCELL_X1 FILLER_1_562 ();
 FILLCELL_X4 FILLER_1_567 ();
 FILLCELL_X8 FILLER_1_581 ();
 FILLCELL_X2 FILLER_1_589 ();
 FILLCELL_X1 FILLER_1_591 ();
 FILLCELL_X4 FILLER_1_601 ();
 FILLCELL_X4 FILLER_1_614 ();
 FILLCELL_X4 FILLER_1_628 ();
 FILLCELL_X8 FILLER_1_639 ();
 FILLCELL_X8 FILLER_1_656 ();
 FILLCELL_X2 FILLER_1_664 ();
 FILLCELL_X4 FILLER_1_670 ();
 FILLCELL_X4 FILLER_1_683 ();
 FILLCELL_X4 FILLER_1_696 ();
 FILLCELL_X2 FILLER_1_700 ();
 FILLCELL_X1 FILLER_1_702 ();
 FILLCELL_X4 FILLER_1_713 ();
 FILLCELL_X1 FILLER_1_717 ();
 FILLCELL_X4 FILLER_1_728 ();
 FILLCELL_X4 FILLER_1_751 ();
 FILLCELL_X2 FILLER_1_755 ();
 FILLCELL_X1 FILLER_1_757 ();
 FILLCELL_X8 FILLER_1_767 ();
 FILLCELL_X2 FILLER_1_775 ();
 FILLCELL_X4 FILLER_1_786 ();
 FILLCELL_X2 FILLER_1_790 ();
 FILLCELL_X1 FILLER_1_792 ();
 FILLCELL_X4 FILLER_1_797 ();
 FILLCELL_X4 FILLER_1_805 ();
 FILLCELL_X4 FILLER_1_816 ();
 FILLCELL_X1 FILLER_1_820 ();
 FILLCELL_X4 FILLER_1_824 ();
 FILLCELL_X4 FILLER_1_837 ();
 FILLCELL_X8 FILLER_1_850 ();
 FILLCELL_X4 FILLER_1_868 ();
 FILLCELL_X2 FILLER_1_872 ();
 FILLCELL_X1 FILLER_1_874 ();
 FILLCELL_X8 FILLER_1_885 ();
 FILLCELL_X2 FILLER_1_893 ();
 FILLCELL_X4 FILLER_1_914 ();
 FILLCELL_X8 FILLER_1_921 ();
 FILLCELL_X4 FILLER_1_929 ();
 FILLCELL_X2 FILLER_1_933 ();
 FILLCELL_X4 FILLER_1_939 ();
 FILLCELL_X4 FILLER_1_946 ();
 FILLCELL_X1 FILLER_1_950 ();
 FILLCELL_X4 FILLER_1_955 ();
 FILLCELL_X4 FILLER_1_968 ();
 FILLCELL_X4 FILLER_1_981 ();
 FILLCELL_X4 FILLER_1_989 ();
 FILLCELL_X4 FILLER_1_1003 ();
 FILLCELL_X8 FILLER_1_1017 ();
 FILLCELL_X4 FILLER_1_1030 ();
 FILLCELL_X4 FILLER_1_1038 ();
 FILLCELL_X8 FILLER_1_1046 ();
 FILLCELL_X4 FILLER_1_1063 ();
 FILLCELL_X4 FILLER_1_1076 ();
 FILLCELL_X8 FILLER_1_1084 ();
 FILLCELL_X2 FILLER_1_1092 ();
 FILLCELL_X4 FILLER_1_1098 ();
 FILLCELL_X4 FILLER_1_1112 ();
 FILLCELL_X4 FILLER_1_1126 ();
 FILLCELL_X1 FILLER_1_1130 ();
 FILLCELL_X4 FILLER_1_1140 ();
 FILLCELL_X8 FILLER_1_1147 ();
 FILLCELL_X4 FILLER_1_1165 ();
 FILLCELL_X4 FILLER_1_1179 ();
 FILLCELL_X2 FILLER_1_1183 ();
 FILLCELL_X8 FILLER_1_1194 ();
 FILLCELL_X4 FILLER_1_1205 ();
 FILLCELL_X4 FILLER_1_1218 ();
 FILLCELL_X4 FILLER_1_1226 ();
 FILLCELL_X4 FILLER_1_1249 ();
 FILLCELL_X4 FILLER_1_1257 ();
 FILLCELL_X2 FILLER_1_1261 ();
 FILLCELL_X4 FILLER_1_1264 ();
 FILLCELL_X32 FILLER_1_1287 ();
 FILLCELL_X4 FILLER_1_1328 ();
 FILLCELL_X4 FILLER_1_1335 ();
 FILLCELL_X2 FILLER_1_1339 ();
 FILLCELL_X8 FILLER_1_1360 ();
 FILLCELL_X2 FILLER_1_1368 ();
 FILLCELL_X1 FILLER_1_1370 ();
 FILLCELL_X4 FILLER_1_1380 ();
 FILLCELL_X4 FILLER_1_1387 ();
 FILLCELL_X32 FILLER_1_1394 ();
 FILLCELL_X32 FILLER_1_1426 ();
 FILLCELL_X32 FILLER_1_1458 ();
 FILLCELL_X32 FILLER_1_1490 ();
 FILLCELL_X32 FILLER_1_1522 ();
 FILLCELL_X32 FILLER_1_1554 ();
 FILLCELL_X32 FILLER_1_1586 ();
 FILLCELL_X32 FILLER_1_1618 ();
 FILLCELL_X32 FILLER_1_1650 ();
 FILLCELL_X32 FILLER_1_1682 ();
 FILLCELL_X32 FILLER_1_1714 ();
 FILLCELL_X16 FILLER_1_1746 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X2 FILLER_2_65 ();
 FILLCELL_X4 FILLER_2_71 ();
 FILLCELL_X2 FILLER_2_75 ();
 FILLCELL_X1 FILLER_2_77 ();
 FILLCELL_X4 FILLER_2_81 ();
 FILLCELL_X4 FILLER_2_92 ();
 FILLCELL_X4 FILLER_2_106 ();
 FILLCELL_X4 FILLER_2_114 ();
 FILLCELL_X4 FILLER_2_127 ();
 FILLCELL_X8 FILLER_2_134 ();
 FILLCELL_X4 FILLER_2_142 ();
 FILLCELL_X4 FILLER_2_150 ();
 FILLCELL_X4 FILLER_2_158 ();
 FILLCELL_X8 FILLER_2_166 ();
 FILLCELL_X2 FILLER_2_174 ();
 FILLCELL_X4 FILLER_2_182 ();
 FILLCELL_X8 FILLER_2_192 ();
 FILLCELL_X4 FILLER_2_200 ();
 FILLCELL_X4 FILLER_2_206 ();
 FILLCELL_X4 FILLER_2_214 ();
 FILLCELL_X8 FILLER_2_228 ();
 FILLCELL_X2 FILLER_2_236 ();
 FILLCELL_X4 FILLER_2_248 ();
 FILLCELL_X2 FILLER_2_252 ();
 FILLCELL_X1 FILLER_2_254 ();
 FILLCELL_X8 FILLER_2_265 ();
 FILLCELL_X2 FILLER_2_273 ();
 FILLCELL_X8 FILLER_2_284 ();
 FILLCELL_X2 FILLER_2_292 ();
 FILLCELL_X1 FILLER_2_294 ();
 FILLCELL_X4 FILLER_2_298 ();
 FILLCELL_X4 FILLER_2_305 ();
 FILLCELL_X2 FILLER_2_309 ();
 FILLCELL_X4 FILLER_2_321 ();
 FILLCELL_X4 FILLER_2_334 ();
 FILLCELL_X4 FILLER_2_341 ();
 FILLCELL_X8 FILLER_2_349 ();
 FILLCELL_X4 FILLER_2_357 ();
 FILLCELL_X1 FILLER_2_361 ();
 FILLCELL_X8 FILLER_2_364 ();
 FILLCELL_X4 FILLER_2_375 ();
 FILLCELL_X8 FILLER_2_388 ();
 FILLCELL_X4 FILLER_2_399 ();
 FILLCELL_X4 FILLER_2_406 ();
 FILLCELL_X8 FILLER_2_417 ();
 FILLCELL_X2 FILLER_2_425 ();
 FILLCELL_X4 FILLER_2_434 ();
 FILLCELL_X8 FILLER_2_448 ();
 FILLCELL_X8 FILLER_2_465 ();
 FILLCELL_X2 FILLER_2_473 ();
 FILLCELL_X1 FILLER_2_475 ();
 FILLCELL_X8 FILLER_2_480 ();
 FILLCELL_X2 FILLER_2_488 ();
 FILLCELL_X8 FILLER_2_492 ();
 FILLCELL_X2 FILLER_2_500 ();
 FILLCELL_X1 FILLER_2_502 ();
 FILLCELL_X4 FILLER_2_506 ();
 FILLCELL_X4 FILLER_2_514 ();
 FILLCELL_X4 FILLER_2_522 ();
 FILLCELL_X8 FILLER_2_529 ();
 FILLCELL_X4 FILLER_2_537 ();
 FILLCELL_X2 FILLER_2_541 ();
 FILLCELL_X1 FILLER_2_543 ();
 FILLCELL_X4 FILLER_2_549 ();
 FILLCELL_X2 FILLER_2_553 ();
 FILLCELL_X8 FILLER_2_564 ();
 FILLCELL_X2 FILLER_2_572 ();
 FILLCELL_X1 FILLER_2_574 ();
 FILLCELL_X4 FILLER_2_585 ();
 FILLCELL_X2 FILLER_2_589 ();
 FILLCELL_X1 FILLER_2_591 ();
 FILLCELL_X4 FILLER_2_599 ();
 FILLCELL_X4 FILLER_2_606 ();
 FILLCELL_X8 FILLER_2_612 ();
 FILLCELL_X4 FILLER_2_620 ();
 FILLCELL_X1 FILLER_2_624 ();
 FILLCELL_X4 FILLER_2_627 ();
 FILLCELL_X4 FILLER_2_632 ();
 FILLCELL_X8 FILLER_2_646 ();
 FILLCELL_X2 FILLER_2_654 ();
 FILLCELL_X8 FILLER_2_665 ();
 FILLCELL_X4 FILLER_2_676 ();
 FILLCELL_X4 FILLER_2_683 ();
 FILLCELL_X2 FILLER_2_687 ();
 FILLCELL_X1 FILLER_2_689 ();
 FILLCELL_X8 FILLER_2_693 ();
 FILLCELL_X1 FILLER_2_701 ();
 FILLCELL_X4 FILLER_2_705 ();
 FILLCELL_X4 FILLER_2_712 ();
 FILLCELL_X16 FILLER_2_718 ();
 FILLCELL_X8 FILLER_2_734 ();
 FILLCELL_X4 FILLER_2_742 ();
 FILLCELL_X2 FILLER_2_746 ();
 FILLCELL_X1 FILLER_2_748 ();
 FILLCELL_X4 FILLER_2_752 ();
 FILLCELL_X4 FILLER_2_760 ();
 FILLCELL_X4 FILLER_2_767 ();
 FILLCELL_X2 FILLER_2_771 ();
 FILLCELL_X1 FILLER_2_773 ();
 FILLCELL_X4 FILLER_2_778 ();
 FILLCELL_X4 FILLER_2_792 ();
 FILLCELL_X2 FILLER_2_796 ();
 FILLCELL_X4 FILLER_2_803 ();
 FILLCELL_X4 FILLER_2_824 ();
 FILLCELL_X2 FILLER_2_828 ();
 FILLCELL_X4 FILLER_2_834 ();
 FILLCELL_X16 FILLER_2_842 ();
 FILLCELL_X8 FILLER_2_861 ();
 FILLCELL_X4 FILLER_2_869 ();
 FILLCELL_X2 FILLER_2_873 ();
 FILLCELL_X4 FILLER_2_878 ();
 FILLCELL_X16 FILLER_2_891 ();
 FILLCELL_X1 FILLER_2_907 ();
 FILLCELL_X4 FILLER_2_912 ();
 FILLCELL_X4 FILLER_2_926 ();
 FILLCELL_X4 FILLER_2_934 ();
 FILLCELL_X8 FILLER_2_947 ();
 FILLCELL_X2 FILLER_2_955 ();
 FILLCELL_X4 FILLER_2_960 ();
 FILLCELL_X2 FILLER_2_964 ();
 FILLCELL_X4 FILLER_2_969 ();
 FILLCELL_X1 FILLER_2_973 ();
 FILLCELL_X4 FILLER_2_977 ();
 FILLCELL_X2 FILLER_2_981 ();
 FILLCELL_X4 FILLER_2_987 ();
 FILLCELL_X2 FILLER_2_991 ();
 FILLCELL_X1 FILLER_2_993 ();
 FILLCELL_X4 FILLER_2_997 ();
 FILLCELL_X1 FILLER_2_1001 ();
 FILLCELL_X8 FILLER_2_1004 ();
 FILLCELL_X1 FILLER_2_1012 ();
 FILLCELL_X4 FILLER_2_1018 ();
 FILLCELL_X16 FILLER_2_1031 ();
 FILLCELL_X4 FILLER_2_1047 ();
 FILLCELL_X4 FILLER_2_1055 ();
 FILLCELL_X1 FILLER_2_1059 ();
 FILLCELL_X4 FILLER_2_1063 ();
 FILLCELL_X1 FILLER_2_1067 ();
 FILLCELL_X4 FILLER_2_1072 ();
 FILLCELL_X4 FILLER_2_1085 ();
 FILLCELL_X4 FILLER_2_1098 ();
 FILLCELL_X4 FILLER_2_1105 ();
 FILLCELL_X8 FILLER_2_1116 ();
 FILLCELL_X4 FILLER_2_1124 ();
 FILLCELL_X1 FILLER_2_1128 ();
 FILLCELL_X4 FILLER_2_1133 ();
 FILLCELL_X2 FILLER_2_1137 ();
 FILLCELL_X1 FILLER_2_1139 ();
 FILLCELL_X8 FILLER_2_1144 ();
 FILLCELL_X4 FILLER_2_1152 ();
 FILLCELL_X1 FILLER_2_1156 ();
 FILLCELL_X4 FILLER_2_1164 ();
 FILLCELL_X4 FILLER_2_1171 ();
 FILLCELL_X4 FILLER_2_1177 ();
 FILLCELL_X4 FILLER_2_1185 ();
 FILLCELL_X8 FILLER_2_1198 ();
 FILLCELL_X1 FILLER_2_1206 ();
 FILLCELL_X4 FILLER_2_1211 ();
 FILLCELL_X4 FILLER_2_1219 ();
 FILLCELL_X32 FILLER_2_1226 ();
 FILLCELL_X2 FILLER_2_1258 ();
 FILLCELL_X1 FILLER_2_1260 ();
 FILLCELL_X8 FILLER_2_1270 ();
 FILLCELL_X2 FILLER_2_1278 ();
 FILLCELL_X1 FILLER_2_1280 ();
 FILLCELL_X4 FILLER_2_1300 ();
 FILLCELL_X4 FILLER_2_1308 ();
 FILLCELL_X4 FILLER_2_1315 ();
 FILLCELL_X4 FILLER_2_1328 ();
 FILLCELL_X4 FILLER_2_1336 ();
 FILLCELL_X16 FILLER_2_1344 ();
 FILLCELL_X4 FILLER_2_1367 ();
 FILLCELL_X1 FILLER_2_1371 ();
 FILLCELL_X8 FILLER_2_1381 ();
 FILLCELL_X1 FILLER_2_1389 ();
 FILLCELL_X8 FILLER_2_1393 ();
 FILLCELL_X2 FILLER_2_1401 ();
 FILLCELL_X1 FILLER_2_1403 ();
 FILLCELL_X32 FILLER_2_1407 ();
 FILLCELL_X32 FILLER_2_1439 ();
 FILLCELL_X32 FILLER_2_1471 ();
 FILLCELL_X32 FILLER_2_1503 ();
 FILLCELL_X32 FILLER_2_1535 ();
 FILLCELL_X32 FILLER_2_1567 ();
 FILLCELL_X32 FILLER_2_1599 ();
 FILLCELL_X32 FILLER_2_1631 ();
 FILLCELL_X32 FILLER_2_1663 ();
 FILLCELL_X32 FILLER_2_1695 ();
 FILLCELL_X16 FILLER_2_1727 ();
 FILLCELL_X8 FILLER_2_1743 ();
 FILLCELL_X2 FILLER_2_1751 ();
 FILLCELL_X1 FILLER_2_1753 ();
 FILLCELL_X4 FILLER_2_1758 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X16 FILLER_3_33 ();
 FILLCELL_X4 FILLER_3_49 ();
 FILLCELL_X2 FILLER_3_53 ();
 FILLCELL_X4 FILLER_3_64 ();
 FILLCELL_X16 FILLER_3_77 ();
 FILLCELL_X8 FILLER_3_95 ();
 FILLCELL_X4 FILLER_3_103 ();
 FILLCELL_X4 FILLER_3_110 ();
 FILLCELL_X4 FILLER_3_118 ();
 FILLCELL_X4 FILLER_3_131 ();
 FILLCELL_X16 FILLER_3_138 ();
 FILLCELL_X2 FILLER_3_154 ();
 FILLCELL_X1 FILLER_3_156 ();
 FILLCELL_X4 FILLER_3_160 ();
 FILLCELL_X2 FILLER_3_164 ();
 FILLCELL_X1 FILLER_3_166 ();
 FILLCELL_X4 FILLER_3_171 ();
 FILLCELL_X4 FILLER_3_182 ();
 FILLCELL_X4 FILLER_3_190 ();
 FILLCELL_X1 FILLER_3_194 ();
 FILLCELL_X4 FILLER_3_198 ();
 FILLCELL_X4 FILLER_3_212 ();
 FILLCELL_X4 FILLER_3_220 ();
 FILLCELL_X4 FILLER_3_226 ();
 FILLCELL_X2 FILLER_3_230 ();
 FILLCELL_X4 FILLER_3_236 ();
 FILLCELL_X2 FILLER_3_240 ();
 FILLCELL_X1 FILLER_3_242 ();
 FILLCELL_X4 FILLER_3_250 ();
 FILLCELL_X4 FILLER_3_256 ();
 FILLCELL_X4 FILLER_3_263 ();
 FILLCELL_X2 FILLER_3_267 ();
 FILLCELL_X32 FILLER_3_272 ();
 FILLCELL_X4 FILLER_3_304 ();
 FILLCELL_X1 FILLER_3_308 ();
 FILLCELL_X4 FILLER_3_311 ();
 FILLCELL_X2 FILLER_3_315 ();
 FILLCELL_X1 FILLER_3_317 ();
 FILLCELL_X32 FILLER_3_321 ();
 FILLCELL_X4 FILLER_3_353 ();
 FILLCELL_X1 FILLER_3_357 ();
 FILLCELL_X4 FILLER_3_361 ();
 FILLCELL_X4 FILLER_3_367 ();
 FILLCELL_X4 FILLER_3_381 ();
 FILLCELL_X4 FILLER_3_388 ();
 FILLCELL_X1 FILLER_3_392 ();
 FILLCELL_X4 FILLER_3_402 ();
 FILLCELL_X4 FILLER_3_408 ();
 FILLCELL_X1 FILLER_3_412 ();
 FILLCELL_X4 FILLER_3_419 ();
 FILLCELL_X8 FILLER_3_429 ();
 FILLCELL_X4 FILLER_3_439 ();
 FILLCELL_X16 FILLER_3_445 ();
 FILLCELL_X4 FILLER_3_461 ();
 FILLCELL_X4 FILLER_3_468 ();
 FILLCELL_X4 FILLER_3_482 ();
 FILLCELL_X4 FILLER_3_490 ();
 FILLCELL_X1 FILLER_3_494 ();
 FILLCELL_X4 FILLER_3_498 ();
 FILLCELL_X16 FILLER_3_505 ();
 FILLCELL_X8 FILLER_3_521 ();
 FILLCELL_X2 FILLER_3_529 ();
 FILLCELL_X1 FILLER_3_531 ();
 FILLCELL_X8 FILLER_3_542 ();
 FILLCELL_X1 FILLER_3_550 ();
 FILLCELL_X4 FILLER_3_555 ();
 FILLCELL_X8 FILLER_3_562 ();
 FILLCELL_X2 FILLER_3_570 ();
 FILLCELL_X4 FILLER_3_576 ();
 FILLCELL_X4 FILLER_3_587 ();
 FILLCELL_X2 FILLER_3_591 ();
 FILLCELL_X4 FILLER_3_596 ();
 FILLCELL_X16 FILLER_3_610 ();
 FILLCELL_X8 FILLER_3_626 ();
 FILLCELL_X2 FILLER_3_634 ();
 FILLCELL_X4 FILLER_3_639 ();
 FILLCELL_X4 FILLER_3_647 ();
 FILLCELL_X4 FILLER_3_655 ();
 FILLCELL_X4 FILLER_3_663 ();
 FILLCELL_X8 FILLER_3_670 ();
 FILLCELL_X1 FILLER_3_678 ();
 FILLCELL_X4 FILLER_3_682 ();
 FILLCELL_X8 FILLER_3_690 ();
 FILLCELL_X2 FILLER_3_698 ();
 FILLCELL_X1 FILLER_3_700 ();
 FILLCELL_X4 FILLER_3_704 ();
 FILLCELL_X4 FILLER_3_717 ();
 FILLCELL_X2 FILLER_3_721 ();
 FILLCELL_X4 FILLER_3_727 ();
 FILLCELL_X8 FILLER_3_738 ();
 FILLCELL_X4 FILLER_3_746 ();
 FILLCELL_X2 FILLER_3_750 ();
 FILLCELL_X1 FILLER_3_752 ();
 FILLCELL_X4 FILLER_3_772 ();
 FILLCELL_X1 FILLER_3_776 ();
 FILLCELL_X4 FILLER_3_780 ();
 FILLCELL_X4 FILLER_3_787 ();
 FILLCELL_X16 FILLER_3_798 ();
 FILLCELL_X4 FILLER_3_814 ();
 FILLCELL_X1 FILLER_3_818 ();
 FILLCELL_X4 FILLER_3_823 ();
 FILLCELL_X16 FILLER_3_830 ();
 FILLCELL_X4 FILLER_3_846 ();
 FILLCELL_X2 FILLER_3_850 ();
 FILLCELL_X1 FILLER_3_852 ();
 FILLCELL_X8 FILLER_3_857 ();
 FILLCELL_X1 FILLER_3_865 ();
 FILLCELL_X4 FILLER_3_868 ();
 FILLCELL_X8 FILLER_3_882 ();
 FILLCELL_X4 FILLER_3_900 ();
 FILLCELL_X4 FILLER_3_913 ();
 FILLCELL_X2 FILLER_3_917 ();
 FILLCELL_X8 FILLER_3_926 ();
 FILLCELL_X1 FILLER_3_934 ();
 FILLCELL_X4 FILLER_3_938 ();
 FILLCELL_X4 FILLER_3_946 ();
 FILLCELL_X8 FILLER_3_959 ();
 FILLCELL_X2 FILLER_3_967 ();
 FILLCELL_X4 FILLER_3_972 ();
 FILLCELL_X4 FILLER_3_985 ();
 FILLCELL_X8 FILLER_3_998 ();
 FILLCELL_X4 FILLER_3_1006 ();
 FILLCELL_X2 FILLER_3_1010 ();
 FILLCELL_X1 FILLER_3_1012 ();
 FILLCELL_X4 FILLER_3_1016 ();
 FILLCELL_X8 FILLER_3_1029 ();
 FILLCELL_X4 FILLER_3_1037 ();
 FILLCELL_X1 FILLER_3_1041 ();
 FILLCELL_X16 FILLER_3_1046 ();
 FILLCELL_X8 FILLER_3_1062 ();
 FILLCELL_X4 FILLER_3_1070 ();
 FILLCELL_X8 FILLER_3_1078 ();
 FILLCELL_X1 FILLER_3_1086 ();
 FILLCELL_X16 FILLER_3_1090 ();
 FILLCELL_X8 FILLER_3_1113 ();
 FILLCELL_X2 FILLER_3_1121 ();
 FILLCELL_X16 FILLER_3_1127 ();
 FILLCELL_X8 FILLER_3_1143 ();
 FILLCELL_X4 FILLER_3_1151 ();
 FILLCELL_X4 FILLER_3_1159 ();
 FILLCELL_X1 FILLER_3_1163 ();
 FILLCELL_X8 FILLER_3_1173 ();
 FILLCELL_X4 FILLER_3_1181 ();
 FILLCELL_X2 FILLER_3_1185 ();
 FILLCELL_X8 FILLER_3_1190 ();
 FILLCELL_X4 FILLER_3_1198 ();
 FILLCELL_X2 FILLER_3_1202 ();
 FILLCELL_X4 FILLER_3_1207 ();
 FILLCELL_X1 FILLER_3_1211 ();
 FILLCELL_X4 FILLER_3_1215 ();
 FILLCELL_X4 FILLER_3_1229 ();
 FILLCELL_X2 FILLER_3_1233 ();
 FILLCELL_X1 FILLER_3_1235 ();
 FILLCELL_X4 FILLER_3_1238 ();
 FILLCELL_X2 FILLER_3_1242 ();
 FILLCELL_X4 FILLER_3_1247 ();
 FILLCELL_X8 FILLER_3_1255 ();
 FILLCELL_X4 FILLER_3_1264 ();
 FILLCELL_X4 FILLER_3_1277 ();
 FILLCELL_X4 FILLER_3_1285 ();
 FILLCELL_X16 FILLER_3_1293 ();
 FILLCELL_X8 FILLER_3_1309 ();
 FILLCELL_X4 FILLER_3_1317 ();
 FILLCELL_X2 FILLER_3_1321 ();
 FILLCELL_X1 FILLER_3_1323 ();
 FILLCELL_X4 FILLER_3_1328 ();
 FILLCELL_X8 FILLER_3_1335 ();
 FILLCELL_X2 FILLER_3_1343 ();
 FILLCELL_X1 FILLER_3_1345 ();
 FILLCELL_X4 FILLER_3_1348 ();
 FILLCELL_X4 FILLER_3_1362 ();
 FILLCELL_X4 FILLER_3_1376 ();
 FILLCELL_X4 FILLER_3_1384 ();
 FILLCELL_X8 FILLER_3_1392 ();
 FILLCELL_X2 FILLER_3_1400 ();
 FILLCELL_X4 FILLER_3_1407 ();
 FILLCELL_X1 FILLER_3_1411 ();
 FILLCELL_X32 FILLER_3_1416 ();
 FILLCELL_X32 FILLER_3_1448 ();
 FILLCELL_X32 FILLER_3_1480 ();
 FILLCELL_X32 FILLER_3_1512 ();
 FILLCELL_X32 FILLER_3_1544 ();
 FILLCELL_X32 FILLER_3_1576 ();
 FILLCELL_X32 FILLER_3_1608 ();
 FILLCELL_X32 FILLER_3_1640 ();
 FILLCELL_X32 FILLER_3_1672 ();
 FILLCELL_X32 FILLER_3_1704 ();
 FILLCELL_X16 FILLER_3_1736 ();
 FILLCELL_X8 FILLER_3_1752 ();
 FILLCELL_X2 FILLER_3_1760 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X4 FILLER_4_33 ();
 FILLCELL_X4 FILLER_4_41 ();
 FILLCELL_X2 FILLER_4_45 ();
 FILLCELL_X1 FILLER_4_47 ();
 FILLCELL_X4 FILLER_4_51 ();
 FILLCELL_X4 FILLER_4_58 ();
 FILLCELL_X4 FILLER_4_66 ();
 FILLCELL_X8 FILLER_4_74 ();
 FILLCELL_X4 FILLER_4_82 ();
 FILLCELL_X8 FILLER_4_90 ();
 FILLCELL_X4 FILLER_4_100 ();
 FILLCELL_X8 FILLER_4_114 ();
 FILLCELL_X4 FILLER_4_125 ();
 FILLCELL_X4 FILLER_4_132 ();
 FILLCELL_X4 FILLER_4_145 ();
 FILLCELL_X4 FILLER_4_151 ();
 FILLCELL_X16 FILLER_4_157 ();
 FILLCELL_X8 FILLER_4_173 ();
 FILLCELL_X2 FILLER_4_181 ();
 FILLCELL_X8 FILLER_4_186 ();
 FILLCELL_X2 FILLER_4_194 ();
 FILLCELL_X4 FILLER_4_199 ();
 FILLCELL_X2 FILLER_4_203 ();
 FILLCELL_X4 FILLER_4_208 ();
 FILLCELL_X8 FILLER_4_222 ();
 FILLCELL_X2 FILLER_4_230 ();
 FILLCELL_X1 FILLER_4_232 ();
 FILLCELL_X4 FILLER_4_236 ();
 FILLCELL_X16 FILLER_4_249 ();
 FILLCELL_X4 FILLER_4_265 ();
 FILLCELL_X1 FILLER_4_269 ();
 FILLCELL_X4 FILLER_4_273 ();
 FILLCELL_X8 FILLER_4_287 ();
 FILLCELL_X2 FILLER_4_295 ();
 FILLCELL_X1 FILLER_4_297 ();
 FILLCELL_X4 FILLER_4_305 ();
 FILLCELL_X4 FILLER_4_319 ();
 FILLCELL_X1 FILLER_4_323 ();
 FILLCELL_X4 FILLER_4_327 ();
 FILLCELL_X4 FILLER_4_335 ();
 FILLCELL_X4 FILLER_4_343 ();
 FILLCELL_X1 FILLER_4_347 ();
 FILLCELL_X4 FILLER_4_352 ();
 FILLCELL_X4 FILLER_4_366 ();
 FILLCELL_X16 FILLER_4_377 ();
 FILLCELL_X1 FILLER_4_393 ();
 FILLCELL_X4 FILLER_4_401 ();
 FILLCELL_X2 FILLER_4_405 ();
 FILLCELL_X4 FILLER_4_411 ();
 FILLCELL_X1 FILLER_4_415 ();
 FILLCELL_X4 FILLER_4_420 ();
 FILLCELL_X4 FILLER_4_427 ();
 FILLCELL_X4 FILLER_4_441 ();
 FILLCELL_X2 FILLER_4_445 ();
 FILLCELL_X1 FILLER_4_447 ();
 FILLCELL_X4 FILLER_4_451 ();
 FILLCELL_X4 FILLER_4_465 ();
 FILLCELL_X2 FILLER_4_469 ();
 FILLCELL_X8 FILLER_4_475 ();
 FILLCELL_X4 FILLER_4_485 ();
 FILLCELL_X4 FILLER_4_499 ();
 FILLCELL_X16 FILLER_4_510 ();
 FILLCELL_X2 FILLER_4_526 ();
 FILLCELL_X1 FILLER_4_528 ();
 FILLCELL_X4 FILLER_4_533 ();
 FILLCELL_X8 FILLER_4_540 ();
 FILLCELL_X4 FILLER_4_552 ();
 FILLCELL_X4 FILLER_4_563 ();
 FILLCELL_X8 FILLER_4_569 ();
 FILLCELL_X4 FILLER_4_577 ();
 FILLCELL_X2 FILLER_4_581 ();
 FILLCELL_X8 FILLER_4_593 ();
 FILLCELL_X4 FILLER_4_610 ();
 FILLCELL_X2 FILLER_4_614 ();
 FILLCELL_X1 FILLER_4_616 ();
 FILLCELL_X4 FILLER_4_620 ();
 FILLCELL_X4 FILLER_4_627 ();
 FILLCELL_X4 FILLER_4_632 ();
 FILLCELL_X8 FILLER_4_645 ();
 FILLCELL_X2 FILLER_4_653 ();
 FILLCELL_X4 FILLER_4_662 ();
 FILLCELL_X2 FILLER_4_666 ();
 FILLCELL_X4 FILLER_4_672 ();
 FILLCELL_X4 FILLER_4_685 ();
 FILLCELL_X8 FILLER_4_698 ();
 FILLCELL_X4 FILLER_4_706 ();
 FILLCELL_X8 FILLER_4_719 ();
 FILLCELL_X2 FILLER_4_727 ();
 FILLCELL_X4 FILLER_4_739 ();
 FILLCELL_X32 FILLER_4_745 ();
 FILLCELL_X8 FILLER_4_780 ();
 FILLCELL_X1 FILLER_4_788 ();
 FILLCELL_X4 FILLER_4_798 ();
 FILLCELL_X4 FILLER_4_805 ();
 FILLCELL_X4 FILLER_4_811 ();
 FILLCELL_X8 FILLER_4_819 ();
 FILLCELL_X1 FILLER_4_827 ();
 FILLCELL_X8 FILLER_4_832 ();
 FILLCELL_X4 FILLER_4_840 ();
 FILLCELL_X2 FILLER_4_844 ();
 FILLCELL_X1 FILLER_4_846 ();
 FILLCELL_X4 FILLER_4_850 ();
 FILLCELL_X4 FILLER_4_864 ();
 FILLCELL_X8 FILLER_4_875 ();
 FILLCELL_X2 FILLER_4_883 ();
 FILLCELL_X1 FILLER_4_885 ();
 FILLCELL_X4 FILLER_4_889 ();
 FILLCELL_X4 FILLER_4_896 ();
 FILLCELL_X16 FILLER_4_902 ();
 FILLCELL_X2 FILLER_4_918 ();
 FILLCELL_X1 FILLER_4_920 ();
 FILLCELL_X4 FILLER_4_923 ();
 FILLCELL_X4 FILLER_4_937 ();
 FILLCELL_X2 FILLER_4_941 ();
 FILLCELL_X1 FILLER_4_943 ();
 FILLCELL_X16 FILLER_4_947 ();
 FILLCELL_X4 FILLER_4_963 ();
 FILLCELL_X4 FILLER_4_970 ();
 FILLCELL_X4 FILLER_4_978 ();
 FILLCELL_X16 FILLER_4_986 ();
 FILLCELL_X4 FILLER_4_1002 ();
 FILLCELL_X8 FILLER_4_1010 ();
 FILLCELL_X1 FILLER_4_1018 ();
 FILLCELL_X4 FILLER_4_1022 ();
 FILLCELL_X4 FILLER_4_1029 ();
 FILLCELL_X4 FILLER_4_1036 ();
 FILLCELL_X1 FILLER_4_1040 ();
 FILLCELL_X4 FILLER_4_1051 ();
 FILLCELL_X8 FILLER_4_1058 ();
 FILLCELL_X8 FILLER_4_1069 ();
 FILLCELL_X2 FILLER_4_1077 ();
 FILLCELL_X4 FILLER_4_1083 ();
 FILLCELL_X4 FILLER_4_1090 ();
 FILLCELL_X1 FILLER_4_1094 ();
 FILLCELL_X4 FILLER_4_1098 ();
 FILLCELL_X8 FILLER_4_1112 ();
 FILLCELL_X4 FILLER_4_1130 ();
 FILLCELL_X2 FILLER_4_1134 ();
 FILLCELL_X8 FILLER_4_1143 ();
 FILLCELL_X4 FILLER_4_1154 ();
 FILLCELL_X2 FILLER_4_1158 ();
 FILLCELL_X1 FILLER_4_1160 ();
 FILLCELL_X4 FILLER_4_1164 ();
 FILLCELL_X2 FILLER_4_1168 ();
 FILLCELL_X1 FILLER_4_1170 ();
 FILLCELL_X16 FILLER_4_1180 ();
 FILLCELL_X2 FILLER_4_1196 ();
 FILLCELL_X4 FILLER_4_1201 ();
 FILLCELL_X4 FILLER_4_1209 ();
 FILLCELL_X8 FILLER_4_1216 ();
 FILLCELL_X4 FILLER_4_1231 ();
 FILLCELL_X8 FILLER_4_1245 ();
 FILLCELL_X4 FILLER_4_1253 ();
 FILLCELL_X4 FILLER_4_1261 ();
 FILLCELL_X4 FILLER_4_1268 ();
 FILLCELL_X4 FILLER_4_1275 ();
 FILLCELL_X4 FILLER_4_1282 ();
 FILLCELL_X8 FILLER_4_1293 ();
 FILLCELL_X1 FILLER_4_1301 ();
 FILLCELL_X4 FILLER_4_1306 ();
 FILLCELL_X4 FILLER_4_1329 ();
 FILLCELL_X2 FILLER_4_1333 ();
 FILLCELL_X16 FILLER_4_1339 ();
 FILLCELL_X2 FILLER_4_1355 ();
 FILLCELL_X4 FILLER_4_1361 ();
 FILLCELL_X8 FILLER_4_1368 ();
 FILLCELL_X4 FILLER_4_1376 ();
 FILLCELL_X4 FILLER_4_1384 ();
 FILLCELL_X2 FILLER_4_1388 ();
 FILLCELL_X1 FILLER_4_1390 ();
 FILLCELL_X8 FILLER_4_1400 ();
 FILLCELL_X1 FILLER_4_1408 ();
 FILLCELL_X32 FILLER_4_1418 ();
 FILLCELL_X32 FILLER_4_1450 ();
 FILLCELL_X32 FILLER_4_1482 ();
 FILLCELL_X32 FILLER_4_1514 ();
 FILLCELL_X32 FILLER_4_1546 ();
 FILLCELL_X32 FILLER_4_1578 ();
 FILLCELL_X32 FILLER_4_1610 ();
 FILLCELL_X32 FILLER_4_1642 ();
 FILLCELL_X32 FILLER_4_1674 ();
 FILLCELL_X32 FILLER_4_1706 ();
 FILLCELL_X16 FILLER_4_1738 ();
 FILLCELL_X8 FILLER_4_1754 ();
 FILLCELL_X16 FILLER_5_1 ();
 FILLCELL_X8 FILLER_5_17 ();
 FILLCELL_X4 FILLER_5_25 ();
 FILLCELL_X2 FILLER_5_29 ();
 FILLCELL_X1 FILLER_5_31 ();
 FILLCELL_X4 FILLER_5_36 ();
 FILLCELL_X4 FILLER_5_49 ();
 FILLCELL_X4 FILLER_5_56 ();
 FILLCELL_X2 FILLER_5_60 ();
 FILLCELL_X1 FILLER_5_62 ();
 FILLCELL_X8 FILLER_5_66 ();
 FILLCELL_X4 FILLER_5_77 ();
 FILLCELL_X4 FILLER_5_84 ();
 FILLCELL_X4 FILLER_5_98 ();
 FILLCELL_X16 FILLER_5_109 ();
 FILLCELL_X8 FILLER_5_125 ();
 FILLCELL_X4 FILLER_5_133 ();
 FILLCELL_X4 FILLER_5_140 ();
 FILLCELL_X4 FILLER_5_148 ();
 FILLCELL_X4 FILLER_5_162 ();
 FILLCELL_X4 FILLER_5_172 ();
 FILLCELL_X2 FILLER_5_176 ();
 FILLCELL_X4 FILLER_5_181 ();
 FILLCELL_X8 FILLER_5_194 ();
 FILLCELL_X1 FILLER_5_202 ();
 FILLCELL_X16 FILLER_5_212 ();
 FILLCELL_X4 FILLER_5_228 ();
 FILLCELL_X2 FILLER_5_232 ();
 FILLCELL_X1 FILLER_5_234 ();
 FILLCELL_X16 FILLER_5_238 ();
 FILLCELL_X4 FILLER_5_257 ();
 FILLCELL_X4 FILLER_5_270 ();
 FILLCELL_X2 FILLER_5_274 ();
 FILLCELL_X1 FILLER_5_276 ();
 FILLCELL_X8 FILLER_5_287 ();
 FILLCELL_X2 FILLER_5_295 ();
 FILLCELL_X4 FILLER_5_307 ();
 FILLCELL_X2 FILLER_5_311 ();
 FILLCELL_X4 FILLER_5_315 ();
 FILLCELL_X2 FILLER_5_319 ();
 FILLCELL_X4 FILLER_5_325 ();
 FILLCELL_X4 FILLER_5_338 ();
 FILLCELL_X8 FILLER_5_351 ();
 FILLCELL_X1 FILLER_5_359 ();
 FILLCELL_X4 FILLER_5_363 ();
 FILLCELL_X4 FILLER_5_376 ();
 FILLCELL_X2 FILLER_5_380 ();
 FILLCELL_X4 FILLER_5_391 ();
 FILLCELL_X8 FILLER_5_405 ();
 FILLCELL_X4 FILLER_5_432 ();
 FILLCELL_X1 FILLER_5_436 ();
 FILLCELL_X4 FILLER_5_441 ();
 FILLCELL_X16 FILLER_5_455 ();
 FILLCELL_X2 FILLER_5_471 ();
 FILLCELL_X4 FILLER_5_477 ();
 FILLCELL_X4 FILLER_5_483 ();
 FILLCELL_X2 FILLER_5_487 ();
 FILLCELL_X1 FILLER_5_489 ();
 FILLCELL_X4 FILLER_5_496 ();
 FILLCELL_X4 FILLER_5_506 ();
 FILLCELL_X1 FILLER_5_510 ();
 FILLCELL_X4 FILLER_5_530 ();
 FILLCELL_X4 FILLER_5_543 ();
 FILLCELL_X2 FILLER_5_547 ();
 FILLCELL_X1 FILLER_5_549 ();
 FILLCELL_X4 FILLER_5_560 ();
 FILLCELL_X2 FILLER_5_564 ();
 FILLCELL_X1 FILLER_5_566 ();
 FILLCELL_X4 FILLER_5_577 ();
 FILLCELL_X4 FILLER_5_583 ();
 FILLCELL_X2 FILLER_5_587 ();
 FILLCELL_X4 FILLER_5_591 ();
 FILLCELL_X2 FILLER_5_595 ();
 FILLCELL_X1 FILLER_5_597 ();
 FILLCELL_X4 FILLER_5_601 ();
 FILLCELL_X4 FILLER_5_608 ();
 FILLCELL_X8 FILLER_5_621 ();
 FILLCELL_X4 FILLER_5_632 ();
 FILLCELL_X4 FILLER_5_645 ();
 FILLCELL_X2 FILLER_5_649 ();
 FILLCELL_X1 FILLER_5_651 ();
 FILLCELL_X4 FILLER_5_662 ();
 FILLCELL_X8 FILLER_5_676 ();
 FILLCELL_X16 FILLER_5_687 ();
 FILLCELL_X4 FILLER_5_703 ();
 FILLCELL_X2 FILLER_5_707 ();
 FILLCELL_X1 FILLER_5_709 ();
 FILLCELL_X4 FILLER_5_720 ();
 FILLCELL_X8 FILLER_5_727 ();
 FILLCELL_X2 FILLER_5_735 ();
 FILLCELL_X1 FILLER_5_737 ();
 FILLCELL_X16 FILLER_5_748 ();
 FILLCELL_X2 FILLER_5_764 ();
 FILLCELL_X1 FILLER_5_766 ();
 FILLCELL_X8 FILLER_5_774 ();
 FILLCELL_X1 FILLER_5_782 ();
 FILLCELL_X8 FILLER_5_792 ();
 FILLCELL_X1 FILLER_5_800 ();
 FILLCELL_X8 FILLER_5_811 ();
 FILLCELL_X4 FILLER_5_828 ();
 FILLCELL_X4 FILLER_5_841 ();
 FILLCELL_X2 FILLER_5_845 ();
 FILLCELL_X4 FILLER_5_850 ();
 FILLCELL_X4 FILLER_5_857 ();
 FILLCELL_X8 FILLER_5_870 ();
 FILLCELL_X1 FILLER_5_878 ();
 FILLCELL_X4 FILLER_5_882 ();
 FILLCELL_X16 FILLER_5_890 ();
 FILLCELL_X4 FILLER_5_909 ();
 FILLCELL_X4 FILLER_5_922 ();
 FILLCELL_X16 FILLER_5_929 ();
 FILLCELL_X4 FILLER_5_952 ();
 FILLCELL_X2 FILLER_5_956 ();
 FILLCELL_X1 FILLER_5_958 ();
 FILLCELL_X4 FILLER_5_963 ();
 FILLCELL_X8 FILLER_5_970 ();
 FILLCELL_X4 FILLER_5_981 ();
 FILLCELL_X8 FILLER_5_988 ();
 FILLCELL_X4 FILLER_5_996 ();
 FILLCELL_X4 FILLER_5_1004 ();
 FILLCELL_X4 FILLER_5_1017 ();
 FILLCELL_X4 FILLER_5_1024 ();
 FILLCELL_X2 FILLER_5_1028 ();
 FILLCELL_X1 FILLER_5_1030 ();
 FILLCELL_X4 FILLER_5_1040 ();
 FILLCELL_X4 FILLER_5_1054 ();
 FILLCELL_X1 FILLER_5_1058 ();
 FILLCELL_X4 FILLER_5_1063 ();
 FILLCELL_X4 FILLER_5_1076 ();
 FILLCELL_X8 FILLER_5_1089 ();
 FILLCELL_X2 FILLER_5_1097 ();
 FILLCELL_X1 FILLER_5_1099 ();
 FILLCELL_X8 FILLER_5_1104 ();
 FILLCELL_X2 FILLER_5_1112 ();
 FILLCELL_X4 FILLER_5_1116 ();
 FILLCELL_X1 FILLER_5_1120 ();
 FILLCELL_X4 FILLER_5_1124 ();
 FILLCELL_X4 FILLER_5_1138 ();
 FILLCELL_X4 FILLER_5_1152 ();
 FILLCELL_X4 FILLER_5_1166 ();
 FILLCELL_X16 FILLER_5_1173 ();
 FILLCELL_X4 FILLER_5_1193 ();
 FILLCELL_X1 FILLER_5_1197 ();
 FILLCELL_X4 FILLER_5_1208 ();
 FILLCELL_X8 FILLER_5_1221 ();
 FILLCELL_X4 FILLER_5_1232 ();
 FILLCELL_X16 FILLER_5_1246 ();
 FILLCELL_X1 FILLER_5_1262 ();
 FILLCELL_X4 FILLER_5_1264 ();
 FILLCELL_X4 FILLER_5_1271 ();
 FILLCELL_X1 FILLER_5_1275 ();
 FILLCELL_X4 FILLER_5_1280 ();
 FILLCELL_X4 FILLER_5_1294 ();
 FILLCELL_X4 FILLER_5_1300 ();
 FILLCELL_X4 FILLER_5_1308 ();
 FILLCELL_X4 FILLER_5_1316 ();
 FILLCELL_X1 FILLER_5_1320 ();
 FILLCELL_X8 FILLER_5_1324 ();
 FILLCELL_X4 FILLER_5_1351 ();
 FILLCELL_X2 FILLER_5_1355 ();
 FILLCELL_X4 FILLER_5_1361 ();
 FILLCELL_X8 FILLER_5_1370 ();
 FILLCELL_X4 FILLER_5_1378 ();
 FILLCELL_X2 FILLER_5_1382 ();
 FILLCELL_X4 FILLER_5_1387 ();
 FILLCELL_X8 FILLER_5_1394 ();
 FILLCELL_X4 FILLER_5_1404 ();
 FILLCELL_X4 FILLER_5_1411 ();
 FILLCELL_X32 FILLER_5_1425 ();
 FILLCELL_X32 FILLER_5_1457 ();
 FILLCELL_X32 FILLER_5_1489 ();
 FILLCELL_X32 FILLER_5_1521 ();
 FILLCELL_X32 FILLER_5_1553 ();
 FILLCELL_X32 FILLER_5_1585 ();
 FILLCELL_X32 FILLER_5_1617 ();
 FILLCELL_X32 FILLER_5_1649 ();
 FILLCELL_X32 FILLER_5_1681 ();
 FILLCELL_X32 FILLER_5_1713 ();
 FILLCELL_X16 FILLER_5_1745 ();
 FILLCELL_X1 FILLER_5_1761 ();
 FILLCELL_X4 FILLER_6_1 ();
 FILLCELL_X8 FILLER_6_8 ();
 FILLCELL_X2 FILLER_6_16 ();
 FILLCELL_X4 FILLER_6_21 ();
 FILLCELL_X4 FILLER_6_29 ();
 FILLCELL_X4 FILLER_6_42 ();
 FILLCELL_X4 FILLER_6_50 ();
 FILLCELL_X4 FILLER_6_57 ();
 FILLCELL_X4 FILLER_6_70 ();
 FILLCELL_X4 FILLER_6_78 ();
 FILLCELL_X1 FILLER_6_82 ();
 FILLCELL_X4 FILLER_6_87 ();
 FILLCELL_X2 FILLER_6_91 ();
 FILLCELL_X1 FILLER_6_93 ();
 FILLCELL_X4 FILLER_6_103 ();
 FILLCELL_X4 FILLER_6_110 ();
 FILLCELL_X1 FILLER_6_114 ();
 FILLCELL_X4 FILLER_6_121 ();
 FILLCELL_X4 FILLER_6_131 ();
 FILLCELL_X2 FILLER_6_135 ();
 FILLCELL_X4 FILLER_6_147 ();
 FILLCELL_X16 FILLER_6_158 ();
 FILLCELL_X4 FILLER_6_174 ();
 FILLCELL_X1 FILLER_6_178 ();
 FILLCELL_X4 FILLER_6_189 ();
 FILLCELL_X2 FILLER_6_193 ();
 FILLCELL_X1 FILLER_6_195 ();
 FILLCELL_X4 FILLER_6_198 ();
 FILLCELL_X8 FILLER_6_212 ();
 FILLCELL_X2 FILLER_6_220 ();
 FILLCELL_X4 FILLER_6_225 ();
 FILLCELL_X4 FILLER_6_232 ();
 FILLCELL_X4 FILLER_6_240 ();
 FILLCELL_X4 FILLER_6_248 ();
 FILLCELL_X1 FILLER_6_252 ();
 FILLCELL_X4 FILLER_6_257 ();
 FILLCELL_X2 FILLER_6_261 ();
 FILLCELL_X1 FILLER_6_263 ();
 FILLCELL_X8 FILLER_6_268 ();
 FILLCELL_X4 FILLER_6_283 ();
 FILLCELL_X2 FILLER_6_287 ();
 FILLCELL_X4 FILLER_6_293 ();
 FILLCELL_X1 FILLER_6_297 ();
 FILLCELL_X4 FILLER_6_301 ();
 FILLCELL_X2 FILLER_6_305 ();
 FILLCELL_X4 FILLER_6_311 ();
 FILLCELL_X2 FILLER_6_315 ();
 FILLCELL_X8 FILLER_6_327 ();
 FILLCELL_X4 FILLER_6_338 ();
 FILLCELL_X16 FILLER_6_345 ();
 FILLCELL_X4 FILLER_6_361 ();
 FILLCELL_X1 FILLER_6_365 ();
 FILLCELL_X4 FILLER_6_369 ();
 FILLCELL_X2 FILLER_6_373 ();
 FILLCELL_X1 FILLER_6_375 ();
 FILLCELL_X8 FILLER_6_379 ();
 FILLCELL_X4 FILLER_6_387 ();
 FILLCELL_X4 FILLER_6_394 ();
 FILLCELL_X16 FILLER_6_408 ();
 FILLCELL_X8 FILLER_6_424 ();
 FILLCELL_X2 FILLER_6_432 ();
 FILLCELL_X4 FILLER_6_444 ();
 FILLCELL_X8 FILLER_6_451 ();
 FILLCELL_X4 FILLER_6_459 ();
 FILLCELL_X4 FILLER_6_468 ();
 FILLCELL_X4 FILLER_6_479 ();
 FILLCELL_X4 FILLER_6_487 ();
 FILLCELL_X2 FILLER_6_491 ();
 FILLCELL_X8 FILLER_6_496 ();
 FILLCELL_X2 FILLER_6_504 ();
 FILLCELL_X1 FILLER_6_506 ();
 FILLCELL_X8 FILLER_6_511 ();
 FILLCELL_X4 FILLER_6_522 ();
 FILLCELL_X4 FILLER_6_535 ();
 FILLCELL_X2 FILLER_6_539 ();
 FILLCELL_X1 FILLER_6_541 ();
 FILLCELL_X4 FILLER_6_545 ();
 FILLCELL_X4 FILLER_6_554 ();
 FILLCELL_X8 FILLER_6_561 ();
 FILLCELL_X4 FILLER_6_576 ();
 FILLCELL_X4 FILLER_6_590 ();
 FILLCELL_X1 FILLER_6_594 ();
 FILLCELL_X4 FILLER_6_602 ();
 FILLCELL_X8 FILLER_6_616 ();
 FILLCELL_X4 FILLER_6_627 ();
 FILLCELL_X4 FILLER_6_632 ();
 FILLCELL_X4 FILLER_6_646 ();
 FILLCELL_X8 FILLER_6_654 ();
 FILLCELL_X4 FILLER_6_664 ();
 FILLCELL_X4 FILLER_6_678 ();
 FILLCELL_X8 FILLER_6_685 ();
 FILLCELL_X1 FILLER_6_693 ();
 FILLCELL_X8 FILLER_6_697 ();
 FILLCELL_X4 FILLER_6_708 ();
 FILLCELL_X4 FILLER_6_722 ();
 FILLCELL_X4 FILLER_6_728 ();
 FILLCELL_X1 FILLER_6_732 ();
 FILLCELL_X4 FILLER_6_736 ();
 FILLCELL_X4 FILLER_6_749 ();
 FILLCELL_X4 FILLER_6_756 ();
 FILLCELL_X4 FILLER_6_770 ();
 FILLCELL_X8 FILLER_6_784 ();
 FILLCELL_X2 FILLER_6_792 ();
 FILLCELL_X4 FILLER_6_799 ();
 FILLCELL_X1 FILLER_6_803 ();
 FILLCELL_X4 FILLER_6_813 ();
 FILLCELL_X2 FILLER_6_817 ();
 FILLCELL_X4 FILLER_6_822 ();
 FILLCELL_X8 FILLER_6_829 ();
 FILLCELL_X4 FILLER_6_837 ();
 FILLCELL_X2 FILLER_6_841 ();
 FILLCELL_X1 FILLER_6_843 ();
 FILLCELL_X4 FILLER_6_847 ();
 FILLCELL_X4 FILLER_6_860 ();
 FILLCELL_X2 FILLER_6_864 ();
 FILLCELL_X4 FILLER_6_870 ();
 FILLCELL_X4 FILLER_6_884 ();
 FILLCELL_X4 FILLER_6_898 ();
 FILLCELL_X2 FILLER_6_902 ();
 FILLCELL_X4 FILLER_6_911 ();
 FILLCELL_X4 FILLER_6_920 ();
 FILLCELL_X4 FILLER_6_926 ();
 FILLCELL_X2 FILLER_6_930 ();
 FILLCELL_X1 FILLER_6_932 ();
 FILLCELL_X4 FILLER_6_936 ();
 FILLCELL_X4 FILLER_6_950 ();
 FILLCELL_X1 FILLER_6_954 ();
 FILLCELL_X4 FILLER_6_965 ();
 FILLCELL_X8 FILLER_6_973 ();
 FILLCELL_X2 FILLER_6_981 ();
 FILLCELL_X4 FILLER_6_992 ();
 FILLCELL_X4 FILLER_6_1005 ();
 FILLCELL_X4 FILLER_6_1013 ();
 FILLCELL_X16 FILLER_6_1026 ();
 FILLCELL_X4 FILLER_6_1042 ();
 FILLCELL_X4 FILLER_6_1050 ();
 FILLCELL_X2 FILLER_6_1054 ();
 FILLCELL_X4 FILLER_6_1058 ();
 FILLCELL_X2 FILLER_6_1062 ();
 FILLCELL_X4 FILLER_6_1068 ();
 FILLCELL_X8 FILLER_6_1075 ();
 FILLCELL_X4 FILLER_6_1083 ();
 FILLCELL_X2 FILLER_6_1087 ();
 FILLCELL_X1 FILLER_6_1089 ();
 FILLCELL_X4 FILLER_6_1093 ();
 FILLCELL_X4 FILLER_6_1106 ();
 FILLCELL_X4 FILLER_6_1113 ();
 FILLCELL_X16 FILLER_6_1119 ();
 FILLCELL_X4 FILLER_6_1137 ();
 FILLCELL_X2 FILLER_6_1141 ();
 FILLCELL_X4 FILLER_6_1146 ();
 FILLCELL_X1 FILLER_6_1150 ();
 FILLCELL_X4 FILLER_6_1158 ();
 FILLCELL_X4 FILLER_6_1172 ();
 FILLCELL_X16 FILLER_6_1195 ();
 FILLCELL_X4 FILLER_6_1214 ();
 FILLCELL_X2 FILLER_6_1218 ();
 FILLCELL_X1 FILLER_6_1220 ();
 FILLCELL_X16 FILLER_6_1230 ();
 FILLCELL_X4 FILLER_6_1249 ();
 FILLCELL_X4 FILLER_6_1257 ();
 FILLCELL_X4 FILLER_6_1270 ();
 FILLCELL_X4 FILLER_6_1283 ();
 FILLCELL_X2 FILLER_6_1287 ();
 FILLCELL_X1 FILLER_6_1289 ();
 FILLCELL_X8 FILLER_6_1300 ();
 FILLCELL_X2 FILLER_6_1308 ();
 FILLCELL_X8 FILLER_6_1319 ();
 FILLCELL_X2 FILLER_6_1327 ();
 FILLCELL_X4 FILLER_6_1348 ();
 FILLCELL_X1 FILLER_6_1352 ();
 FILLCELL_X4 FILLER_6_1357 ();
 FILLCELL_X4 FILLER_6_1368 ();
 FILLCELL_X4 FILLER_6_1377 ();
 FILLCELL_X4 FILLER_6_1385 ();
 FILLCELL_X8 FILLER_6_1398 ();
 FILLCELL_X4 FILLER_6_1416 ();
 FILLCELL_X4 FILLER_6_1427 ();
 FILLCELL_X4 FILLER_6_1435 ();
 FILLCELL_X32 FILLER_6_1441 ();
 FILLCELL_X32 FILLER_6_1473 ();
 FILLCELL_X32 FILLER_6_1505 ();
 FILLCELL_X32 FILLER_6_1537 ();
 FILLCELL_X32 FILLER_6_1569 ();
 FILLCELL_X32 FILLER_6_1601 ();
 FILLCELL_X32 FILLER_6_1633 ();
 FILLCELL_X32 FILLER_6_1665 ();
 FILLCELL_X32 FILLER_6_1697 ();
 FILLCELL_X32 FILLER_6_1729 ();
 FILLCELL_X1 FILLER_6_1761 ();
 FILLCELL_X16 FILLER_7_1 ();
 FILLCELL_X8 FILLER_7_17 ();
 FILLCELL_X4 FILLER_7_25 ();
 FILLCELL_X1 FILLER_7_29 ();
 FILLCELL_X4 FILLER_7_33 ();
 FILLCELL_X16 FILLER_7_56 ();
 FILLCELL_X8 FILLER_7_81 ();
 FILLCELL_X2 FILLER_7_89 ();
 FILLCELL_X1 FILLER_7_91 ();
 FILLCELL_X16 FILLER_7_96 ();
 FILLCELL_X1 FILLER_7_112 ();
 FILLCELL_X4 FILLER_7_116 ();
 FILLCELL_X4 FILLER_7_127 ();
 FILLCELL_X16 FILLER_7_134 ();
 FILLCELL_X4 FILLER_7_150 ();
 FILLCELL_X2 FILLER_7_154 ();
 FILLCELL_X1 FILLER_7_156 ();
 FILLCELL_X4 FILLER_7_176 ();
 FILLCELL_X4 FILLER_7_182 ();
 FILLCELL_X2 FILLER_7_186 ();
 FILLCELL_X4 FILLER_7_192 ();
 FILLCELL_X8 FILLER_7_199 ();
 FILLCELL_X1 FILLER_7_207 ();
 FILLCELL_X4 FILLER_7_210 ();
 FILLCELL_X4 FILLER_7_217 ();
 FILLCELL_X4 FILLER_7_230 ();
 FILLCELL_X1 FILLER_7_234 ();
 FILLCELL_X4 FILLER_7_238 ();
 FILLCELL_X4 FILLER_7_251 ();
 FILLCELL_X4 FILLER_7_264 ();
 FILLCELL_X1 FILLER_7_268 ();
 FILLCELL_X4 FILLER_7_278 ();
 FILLCELL_X1 FILLER_7_282 ();
 FILLCELL_X4 FILLER_7_286 ();
 FILLCELL_X4 FILLER_7_292 ();
 FILLCELL_X4 FILLER_7_299 ();
 FILLCELL_X4 FILLER_7_313 ();
 FILLCELL_X2 FILLER_7_317 ();
 FILLCELL_X1 FILLER_7_319 ();
 FILLCELL_X8 FILLER_7_323 ();
 FILLCELL_X4 FILLER_7_331 ();
 FILLCELL_X1 FILLER_7_335 ();
 FILLCELL_X4 FILLER_7_339 ();
 FILLCELL_X8 FILLER_7_347 ();
 FILLCELL_X1 FILLER_7_355 ();
 FILLCELL_X4 FILLER_7_359 ();
 FILLCELL_X8 FILLER_7_367 ();
 FILLCELL_X2 FILLER_7_375 ();
 FILLCELL_X1 FILLER_7_377 ();
 FILLCELL_X8 FILLER_7_382 ();
 FILLCELL_X4 FILLER_7_390 ();
 FILLCELL_X1 FILLER_7_394 ();
 FILLCELL_X4 FILLER_7_398 ();
 FILLCELL_X16 FILLER_7_405 ();
 FILLCELL_X8 FILLER_7_421 ();
 FILLCELL_X8 FILLER_7_431 ();
 FILLCELL_X2 FILLER_7_439 ();
 FILLCELL_X4 FILLER_7_444 ();
 FILLCELL_X8 FILLER_7_457 ();
 FILLCELL_X1 FILLER_7_465 ();
 FILLCELL_X4 FILLER_7_483 ();
 FILLCELL_X4 FILLER_7_491 ();
 FILLCELL_X2 FILLER_7_495 ();
 FILLCELL_X1 FILLER_7_497 ();
 FILLCELL_X8 FILLER_7_508 ();
 FILLCELL_X4 FILLER_7_519 ();
 FILLCELL_X4 FILLER_7_527 ();
 FILLCELL_X4 FILLER_7_535 ();
 FILLCELL_X2 FILLER_7_539 ();
 FILLCELL_X4 FILLER_7_544 ();
 FILLCELL_X4 FILLER_7_557 ();
 FILLCELL_X16 FILLER_7_570 ();
 FILLCELL_X8 FILLER_7_586 ();
 FILLCELL_X4 FILLER_7_597 ();
 FILLCELL_X4 FILLER_7_611 ();
 FILLCELL_X2 FILLER_7_615 ();
 FILLCELL_X1 FILLER_7_617 ();
 FILLCELL_X8 FILLER_7_620 ();
 FILLCELL_X1 FILLER_7_628 ();
 FILLCELL_X8 FILLER_7_632 ();
 FILLCELL_X4 FILLER_7_640 ();
 FILLCELL_X2 FILLER_7_644 ();
 FILLCELL_X1 FILLER_7_646 ();
 FILLCELL_X8 FILLER_7_650 ();
 FILLCELL_X1 FILLER_7_658 ();
 FILLCELL_X16 FILLER_7_661 ();
 FILLCELL_X4 FILLER_7_677 ();
 FILLCELL_X2 FILLER_7_681 ();
 FILLCELL_X1 FILLER_7_683 ();
 FILLCELL_X4 FILLER_7_694 ();
 FILLCELL_X4 FILLER_7_707 ();
 FILLCELL_X4 FILLER_7_718 ();
 FILLCELL_X8 FILLER_7_724 ();
 FILLCELL_X4 FILLER_7_732 ();
 FILLCELL_X2 FILLER_7_736 ();
 FILLCELL_X1 FILLER_7_738 ();
 FILLCELL_X4 FILLER_7_742 ();
 FILLCELL_X2 FILLER_7_746 ();
 FILLCELL_X1 FILLER_7_748 ();
 FILLCELL_X4 FILLER_7_751 ();
 FILLCELL_X8 FILLER_7_764 ();
 FILLCELL_X1 FILLER_7_772 ();
 FILLCELL_X4 FILLER_7_776 ();
 FILLCELL_X4 FILLER_7_783 ();
 FILLCELL_X8 FILLER_7_794 ();
 FILLCELL_X1 FILLER_7_802 ();
 FILLCELL_X8 FILLER_7_806 ();
 FILLCELL_X1 FILLER_7_814 ();
 FILLCELL_X4 FILLER_7_818 ();
 FILLCELL_X1 FILLER_7_822 ();
 FILLCELL_X4 FILLER_7_826 ();
 FILLCELL_X8 FILLER_7_834 ();
 FILLCELL_X1 FILLER_7_842 ();
 FILLCELL_X4 FILLER_7_846 ();
 FILLCELL_X16 FILLER_7_859 ();
 FILLCELL_X8 FILLER_7_875 ();
 FILLCELL_X4 FILLER_7_883 ();
 FILLCELL_X2 FILLER_7_887 ();
 FILLCELL_X1 FILLER_7_889 ();
 FILLCELL_X4 FILLER_7_893 ();
 FILLCELL_X4 FILLER_7_899 ();
 FILLCELL_X2 FILLER_7_903 ();
 FILLCELL_X4 FILLER_7_914 ();
 FILLCELL_X4 FILLER_7_928 ();
 FILLCELL_X8 FILLER_7_941 ();
 FILLCELL_X1 FILLER_7_949 ();
 FILLCELL_X4 FILLER_7_955 ();
 FILLCELL_X4 FILLER_7_968 ();
 FILLCELL_X8 FILLER_7_974 ();
 FILLCELL_X2 FILLER_7_982 ();
 FILLCELL_X4 FILLER_7_987 ();
 FILLCELL_X4 FILLER_7_995 ();
 FILLCELL_X4 FILLER_7_1003 ();
 FILLCELL_X4 FILLER_7_1010 ();
 FILLCELL_X8 FILLER_7_1017 ();
 FILLCELL_X4 FILLER_7_1025 ();
 FILLCELL_X4 FILLER_7_1032 ();
 FILLCELL_X2 FILLER_7_1036 ();
 FILLCELL_X4 FILLER_7_1041 ();
 FILLCELL_X32 FILLER_7_1055 ();
 FILLCELL_X2 FILLER_7_1087 ();
 FILLCELL_X4 FILLER_7_1098 ();
 FILLCELL_X4 FILLER_7_1105 ();
 FILLCELL_X1 FILLER_7_1109 ();
 FILLCELL_X4 FILLER_7_1117 ();
 FILLCELL_X4 FILLER_7_1131 ();
 FILLCELL_X8 FILLER_7_1138 ();
 FILLCELL_X2 FILLER_7_1146 ();
 FILLCELL_X4 FILLER_7_1157 ();
 FILLCELL_X2 FILLER_7_1161 ();
 FILLCELL_X4 FILLER_7_1165 ();
 FILLCELL_X2 FILLER_7_1169 ();
 FILLCELL_X8 FILLER_7_1175 ();
 FILLCELL_X4 FILLER_7_1183 ();
 FILLCELL_X2 FILLER_7_1187 ();
 FILLCELL_X1 FILLER_7_1189 ();
 FILLCELL_X4 FILLER_7_1192 ();
 FILLCELL_X2 FILLER_7_1196 ();
 FILLCELL_X1 FILLER_7_1198 ();
 FILLCELL_X4 FILLER_7_1201 ();
 FILLCELL_X4 FILLER_7_1212 ();
 FILLCELL_X1 FILLER_7_1216 ();
 FILLCELL_X4 FILLER_7_1220 ();
 FILLCELL_X4 FILLER_7_1227 ();
 FILLCELL_X2 FILLER_7_1231 ();
 FILLCELL_X1 FILLER_7_1233 ();
 FILLCELL_X4 FILLER_7_1236 ();
 FILLCELL_X16 FILLER_7_1247 ();
 FILLCELL_X4 FILLER_7_1264 ();
 FILLCELL_X8 FILLER_7_1272 ();
 FILLCELL_X4 FILLER_7_1280 ();
 FILLCELL_X4 FILLER_7_1287 ();
 FILLCELL_X8 FILLER_7_1294 ();
 FILLCELL_X2 FILLER_7_1302 ();
 FILLCELL_X1 FILLER_7_1304 ();
 FILLCELL_X4 FILLER_7_1308 ();
 FILLCELL_X8 FILLER_7_1315 ();
 FILLCELL_X2 FILLER_7_1323 ();
 FILLCELL_X16 FILLER_7_1329 ();
 FILLCELL_X8 FILLER_7_1345 ();
 FILLCELL_X2 FILLER_7_1353 ();
 FILLCELL_X1 FILLER_7_1355 ();
 FILLCELL_X4 FILLER_7_1358 ();
 FILLCELL_X4 FILLER_7_1379 ();
 FILLCELL_X2 FILLER_7_1383 ();
 FILLCELL_X4 FILLER_7_1394 ();
 FILLCELL_X4 FILLER_7_1401 ();
 FILLCELL_X16 FILLER_7_1408 ();
 FILLCELL_X8 FILLER_7_1424 ();
 FILLCELL_X4 FILLER_7_1435 ();
 FILLCELL_X1 FILLER_7_1439 ();
 FILLCELL_X16 FILLER_7_1447 ();
 FILLCELL_X2 FILLER_7_1463 ();
 FILLCELL_X1 FILLER_7_1465 ();
 FILLCELL_X32 FILLER_7_1485 ();
 FILLCELL_X32 FILLER_7_1517 ();
 FILLCELL_X32 FILLER_7_1549 ();
 FILLCELL_X32 FILLER_7_1581 ();
 FILLCELL_X32 FILLER_7_1613 ();
 FILLCELL_X32 FILLER_7_1645 ();
 FILLCELL_X32 FILLER_7_1677 ();
 FILLCELL_X32 FILLER_7_1709 ();
 FILLCELL_X16 FILLER_7_1741 ();
 FILLCELL_X4 FILLER_7_1757 ();
 FILLCELL_X1 FILLER_7_1761 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X16 FILLER_8_33 ();
 FILLCELL_X8 FILLER_8_49 ();
 FILLCELL_X4 FILLER_8_57 ();
 FILLCELL_X1 FILLER_8_61 ();
 FILLCELL_X4 FILLER_8_65 ();
 FILLCELL_X4 FILLER_8_73 ();
 FILLCELL_X4 FILLER_8_80 ();
 FILLCELL_X4 FILLER_8_87 ();
 FILLCELL_X4 FILLER_8_94 ();
 FILLCELL_X4 FILLER_8_107 ();
 FILLCELL_X8 FILLER_8_120 ();
 FILLCELL_X4 FILLER_8_128 ();
 FILLCELL_X1 FILLER_8_132 ();
 FILLCELL_X4 FILLER_8_135 ();
 FILLCELL_X4 FILLER_8_142 ();
 FILLCELL_X8 FILLER_8_156 ();
 FILLCELL_X4 FILLER_8_164 ();
 FILLCELL_X4 FILLER_8_171 ();
 FILLCELL_X8 FILLER_8_185 ();
 FILLCELL_X1 FILLER_8_193 ();
 FILLCELL_X8 FILLER_8_204 ();
 FILLCELL_X8 FILLER_8_222 ();
 FILLCELL_X2 FILLER_8_230 ();
 FILLCELL_X8 FILLER_8_241 ();
 FILLCELL_X8 FILLER_8_252 ();
 FILLCELL_X4 FILLER_8_260 ();
 FILLCELL_X2 FILLER_8_264 ();
 FILLCELL_X1 FILLER_8_266 ();
 FILLCELL_X4 FILLER_8_270 ();
 FILLCELL_X1 FILLER_8_274 ();
 FILLCELL_X4 FILLER_8_279 ();
 FILLCELL_X4 FILLER_8_293 ();
 FILLCELL_X8 FILLER_8_299 ();
 FILLCELL_X4 FILLER_8_307 ();
 FILLCELL_X2 FILLER_8_311 ();
 FILLCELL_X8 FILLER_8_316 ();
 FILLCELL_X1 FILLER_8_324 ();
 FILLCELL_X4 FILLER_8_334 ();
 FILLCELL_X1 FILLER_8_338 ();
 FILLCELL_X4 FILLER_8_343 ();
 FILLCELL_X8 FILLER_8_356 ();
 FILLCELL_X4 FILLER_8_373 ();
 FILLCELL_X2 FILLER_8_377 ();
 FILLCELL_X1 FILLER_8_379 ();
 FILLCELL_X8 FILLER_8_390 ();
 FILLCELL_X2 FILLER_8_398 ();
 FILLCELL_X8 FILLER_8_409 ();
 FILLCELL_X2 FILLER_8_417 ();
 FILLCELL_X8 FILLER_8_426 ();
 FILLCELL_X4 FILLER_8_444 ();
 FILLCELL_X2 FILLER_8_448 ();
 FILLCELL_X1 FILLER_8_450 ();
 FILLCELL_X8 FILLER_8_460 ();
 FILLCELL_X4 FILLER_8_468 ();
 FILLCELL_X1 FILLER_8_472 ();
 FILLCELL_X8 FILLER_8_478 ();
 FILLCELL_X2 FILLER_8_486 ();
 FILLCELL_X1 FILLER_8_488 ();
 FILLCELL_X32 FILLER_8_508 ();
 FILLCELL_X4 FILLER_8_540 ();
 FILLCELL_X2 FILLER_8_544 ();
 FILLCELL_X1 FILLER_8_546 ();
 FILLCELL_X4 FILLER_8_550 ();
 FILLCELL_X2 FILLER_8_554 ();
 FILLCELL_X1 FILLER_8_556 ();
 FILLCELL_X4 FILLER_8_564 ();
 FILLCELL_X1 FILLER_8_568 ();
 FILLCELL_X4 FILLER_8_572 ();
 FILLCELL_X4 FILLER_8_585 ();
 FILLCELL_X4 FILLER_8_592 ();
 FILLCELL_X2 FILLER_8_596 ();
 FILLCELL_X1 FILLER_8_598 ();
 FILLCELL_X4 FILLER_8_602 ();
 FILLCELL_X2 FILLER_8_606 ();
 FILLCELL_X1 FILLER_8_608 ();
 FILLCELL_X4 FILLER_8_613 ();
 FILLCELL_X4 FILLER_8_619 ();
 FILLCELL_X4 FILLER_8_627 ();
 FILLCELL_X4 FILLER_8_632 ();
 FILLCELL_X8 FILLER_8_645 ();
 FILLCELL_X8 FILLER_8_656 ();
 FILLCELL_X4 FILLER_8_667 ();
 FILLCELL_X4 FILLER_8_681 ();
 FILLCELL_X4 FILLER_8_692 ();
 FILLCELL_X8 FILLER_8_699 ();
 FILLCELL_X4 FILLER_8_710 ();
 FILLCELL_X8 FILLER_8_718 ();
 FILLCELL_X4 FILLER_8_736 ();
 FILLCELL_X1 FILLER_8_740 ();
 FILLCELL_X4 FILLER_8_745 ();
 FILLCELL_X8 FILLER_8_758 ();
 FILLCELL_X1 FILLER_8_766 ();
 FILLCELL_X4 FILLER_8_771 ();
 FILLCELL_X4 FILLER_8_785 ();
 FILLCELL_X1 FILLER_8_789 ();
 FILLCELL_X4 FILLER_8_792 ();
 FILLCELL_X4 FILLER_8_806 ();
 FILLCELL_X4 FILLER_8_819 ();
 FILLCELL_X2 FILLER_8_823 ();
 FILLCELL_X1 FILLER_8_825 ();
 FILLCELL_X4 FILLER_8_830 ();
 FILLCELL_X4 FILLER_8_843 ();
 FILLCELL_X2 FILLER_8_847 ();
 FILLCELL_X4 FILLER_8_853 ();
 FILLCELL_X2 FILLER_8_857 ();
 FILLCELL_X4 FILLER_8_862 ();
 FILLCELL_X2 FILLER_8_866 ();
 FILLCELL_X1 FILLER_8_868 ();
 FILLCELL_X4 FILLER_8_878 ();
 FILLCELL_X8 FILLER_8_889 ();
 FILLCELL_X4 FILLER_8_900 ();
 FILLCELL_X8 FILLER_8_914 ();
 FILLCELL_X4 FILLER_8_922 ();
 FILLCELL_X1 FILLER_8_926 ();
 FILLCELL_X4 FILLER_8_930 ();
 FILLCELL_X4 FILLER_8_943 ();
 FILLCELL_X4 FILLER_8_950 ();
 FILLCELL_X4 FILLER_8_957 ();
 FILLCELL_X16 FILLER_8_964 ();
 FILLCELL_X4 FILLER_8_980 ();
 FILLCELL_X1 FILLER_8_984 ();
 FILLCELL_X8 FILLER_8_989 ();
 FILLCELL_X4 FILLER_8_1006 ();
 FILLCELL_X4 FILLER_8_1015 ();
 FILLCELL_X1 FILLER_8_1019 ();
 FILLCELL_X4 FILLER_8_1024 ();
 FILLCELL_X8 FILLER_8_1038 ();
 FILLCELL_X4 FILLER_8_1053 ();
 FILLCELL_X8 FILLER_8_1067 ();
 FILLCELL_X1 FILLER_8_1075 ();
 FILLCELL_X4 FILLER_8_1078 ();
 FILLCELL_X8 FILLER_8_1092 ();
 FILLCELL_X4 FILLER_8_1104 ();
 FILLCELL_X8 FILLER_8_1118 ();
 FILLCELL_X4 FILLER_8_1129 ();
 FILLCELL_X8 FILLER_8_1142 ();
 FILLCELL_X2 FILLER_8_1150 ();
 FILLCELL_X1 FILLER_8_1152 ();
 FILLCELL_X4 FILLER_8_1156 ();
 FILLCELL_X4 FILLER_8_1170 ();
 FILLCELL_X2 FILLER_8_1174 ();
 FILLCELL_X4 FILLER_8_1183 ();
 FILLCELL_X8 FILLER_8_1196 ();
 FILLCELL_X1 FILLER_8_1204 ();
 FILLCELL_X4 FILLER_8_1215 ();
 FILLCELL_X2 FILLER_8_1219 ();
 FILLCELL_X1 FILLER_8_1221 ();
 FILLCELL_X4 FILLER_8_1232 ();
 FILLCELL_X4 FILLER_8_1238 ();
 FILLCELL_X4 FILLER_8_1252 ();
 FILLCELL_X2 FILLER_8_1256 ();
 FILLCELL_X4 FILLER_8_1261 ();
 FILLCELL_X1 FILLER_8_1265 ();
 FILLCELL_X8 FILLER_8_1270 ();
 FILLCELL_X4 FILLER_8_1278 ();
 FILLCELL_X1 FILLER_8_1282 ();
 FILLCELL_X4 FILLER_8_1286 ();
 FILLCELL_X4 FILLER_8_1299 ();
 FILLCELL_X2 FILLER_8_1303 ();
 FILLCELL_X1 FILLER_8_1305 ();
 FILLCELL_X4 FILLER_8_1310 ();
 FILLCELL_X8 FILLER_8_1323 ();
 FILLCELL_X4 FILLER_8_1331 ();
 FILLCELL_X4 FILLER_8_1342 ();
 FILLCELL_X4 FILLER_8_1349 ();
 FILLCELL_X1 FILLER_8_1353 ();
 FILLCELL_X4 FILLER_8_1363 ();
 FILLCELL_X8 FILLER_8_1370 ();
 FILLCELL_X2 FILLER_8_1378 ();
 FILLCELL_X1 FILLER_8_1380 ();
 FILLCELL_X4 FILLER_8_1391 ();
 FILLCELL_X8 FILLER_8_1398 ();
 FILLCELL_X4 FILLER_8_1406 ();
 FILLCELL_X8 FILLER_8_1414 ();
 FILLCELL_X4 FILLER_8_1422 ();
 FILLCELL_X2 FILLER_8_1426 ();
 FILLCELL_X1 FILLER_8_1428 ();
 FILLCELL_X4 FILLER_8_1439 ();
 FILLCELL_X8 FILLER_8_1453 ();
 FILLCELL_X4 FILLER_8_1461 ();
 FILLCELL_X1 FILLER_8_1465 ();
 FILLCELL_X4 FILLER_8_1470 ();
 FILLCELL_X2 FILLER_8_1474 ();
 FILLCELL_X32 FILLER_8_1480 ();
 FILLCELL_X32 FILLER_8_1512 ();
 FILLCELL_X32 FILLER_8_1544 ();
 FILLCELL_X32 FILLER_8_1576 ();
 FILLCELL_X32 FILLER_8_1608 ();
 FILLCELL_X32 FILLER_8_1640 ();
 FILLCELL_X32 FILLER_8_1672 ();
 FILLCELL_X32 FILLER_8_1704 ();
 FILLCELL_X16 FILLER_8_1736 ();
 FILLCELL_X8 FILLER_8_1752 ();
 FILLCELL_X2 FILLER_8_1760 ();
 FILLCELL_X16 FILLER_9_1 ();
 FILLCELL_X8 FILLER_9_17 ();
 FILLCELL_X4 FILLER_9_25 ();
 FILLCELL_X2 FILLER_9_29 ();
 FILLCELL_X1 FILLER_9_31 ();
 FILLCELL_X4 FILLER_9_34 ();
 FILLCELL_X2 FILLER_9_38 ();
 FILLCELL_X4 FILLER_9_49 ();
 FILLCELL_X8 FILLER_9_56 ();
 FILLCELL_X8 FILLER_9_74 ();
 FILLCELL_X8 FILLER_9_85 ();
 FILLCELL_X4 FILLER_9_93 ();
 FILLCELL_X2 FILLER_9_97 ();
 FILLCELL_X4 FILLER_9_102 ();
 FILLCELL_X8 FILLER_9_109 ();
 FILLCELL_X4 FILLER_9_117 ();
 FILLCELL_X4 FILLER_9_128 ();
 FILLCELL_X16 FILLER_9_142 ();
 FILLCELL_X1 FILLER_9_158 ();
 FILLCELL_X8 FILLER_9_163 ();
 FILLCELL_X4 FILLER_9_171 ();
 FILLCELL_X8 FILLER_9_182 ();
 FILLCELL_X2 FILLER_9_190 ();
 FILLCELL_X1 FILLER_9_192 ();
 FILLCELL_X4 FILLER_9_197 ();
 FILLCELL_X1 FILLER_9_201 ();
 FILLCELL_X16 FILLER_9_206 ();
 FILLCELL_X2 FILLER_9_222 ();
 FILLCELL_X4 FILLER_9_227 ();
 FILLCELL_X2 FILLER_9_231 ();
 FILLCELL_X1 FILLER_9_233 ();
 FILLCELL_X16 FILLER_9_236 ();
 FILLCELL_X4 FILLER_9_252 ();
 FILLCELL_X1 FILLER_9_256 ();
 FILLCELL_X4 FILLER_9_260 ();
 FILLCELL_X4 FILLER_9_267 ();
 FILLCELL_X4 FILLER_9_280 ();
 FILLCELL_X1 FILLER_9_284 ();
 FILLCELL_X8 FILLER_9_292 ();
 FILLCELL_X1 FILLER_9_300 ();
 FILLCELL_X4 FILLER_9_311 ();
 FILLCELL_X2 FILLER_9_315 ();
 FILLCELL_X1 FILLER_9_317 ();
 FILLCELL_X4 FILLER_9_327 ();
 FILLCELL_X8 FILLER_9_334 ();
 FILLCELL_X4 FILLER_9_342 ();
 FILLCELL_X4 FILLER_9_349 ();
 FILLCELL_X2 FILLER_9_353 ();
 FILLCELL_X4 FILLER_9_359 ();
 FILLCELL_X2 FILLER_9_363 ();
 FILLCELL_X1 FILLER_9_365 ();
 FILLCELL_X8 FILLER_9_370 ();
 FILLCELL_X1 FILLER_9_378 ();
 FILLCELL_X4 FILLER_9_382 ();
 FILLCELL_X4 FILLER_9_393 ();
 FILLCELL_X8 FILLER_9_406 ();
 FILLCELL_X4 FILLER_9_424 ();
 FILLCELL_X8 FILLER_9_438 ();
 FILLCELL_X2 FILLER_9_446 ();
 FILLCELL_X4 FILLER_9_451 ();
 FILLCELL_X16 FILLER_9_458 ();
 FILLCELL_X4 FILLER_9_474 ();
 FILLCELL_X4 FILLER_9_482 ();
 FILLCELL_X4 FILLER_9_490 ();
 FILLCELL_X4 FILLER_9_497 ();
 FILLCELL_X4 FILLER_9_504 ();
 FILLCELL_X2 FILLER_9_508 ();
 FILLCELL_X4 FILLER_9_513 ();
 FILLCELL_X4 FILLER_9_521 ();
 FILLCELL_X1 FILLER_9_525 ();
 FILLCELL_X4 FILLER_9_530 ();
 FILLCELL_X2 FILLER_9_534 ();
 FILLCELL_X1 FILLER_9_536 ();
 FILLCELL_X4 FILLER_9_541 ();
 FILLCELL_X4 FILLER_9_555 ();
 FILLCELL_X1 FILLER_9_559 ();
 FILLCELL_X4 FILLER_9_562 ();
 FILLCELL_X8 FILLER_9_576 ();
 FILLCELL_X4 FILLER_9_593 ();
 FILLCELL_X8 FILLER_9_607 ();
 FILLCELL_X1 FILLER_9_615 ();
 FILLCELL_X4 FILLER_9_626 ();
 FILLCELL_X4 FILLER_9_634 ();
 FILLCELL_X4 FILLER_9_647 ();
 FILLCELL_X8 FILLER_9_661 ();
 FILLCELL_X2 FILLER_9_669 ();
 FILLCELL_X8 FILLER_9_675 ();
 FILLCELL_X4 FILLER_9_685 ();
 FILLCELL_X2 FILLER_9_689 ();
 FILLCELL_X1 FILLER_9_691 ();
 FILLCELL_X4 FILLER_9_695 ();
 FILLCELL_X4 FILLER_9_702 ();
 FILLCELL_X4 FILLER_9_709 ();
 FILLCELL_X8 FILLER_9_717 ();
 FILLCELL_X2 FILLER_9_725 ();
 FILLCELL_X1 FILLER_9_727 ();
 FILLCELL_X4 FILLER_9_733 ();
 FILLCELL_X4 FILLER_9_746 ();
 FILLCELL_X4 FILLER_9_753 ();
 FILLCELL_X4 FILLER_9_761 ();
 FILLCELL_X2 FILLER_9_765 ();
 FILLCELL_X4 FILLER_9_771 ();
 FILLCELL_X8 FILLER_9_780 ();
 FILLCELL_X2 FILLER_9_788 ();
 FILLCELL_X4 FILLER_9_793 ();
 FILLCELL_X2 FILLER_9_797 ();
 FILLCELL_X1 FILLER_9_799 ();
 FILLCELL_X8 FILLER_9_803 ();
 FILLCELL_X4 FILLER_9_813 ();
 FILLCELL_X8 FILLER_9_821 ();
 FILLCELL_X4 FILLER_9_829 ();
 FILLCELL_X16 FILLER_9_836 ();
 FILLCELL_X1 FILLER_9_852 ();
 FILLCELL_X4 FILLER_9_863 ();
 FILLCELL_X4 FILLER_9_877 ();
 FILLCELL_X2 FILLER_9_881 ();
 FILLCELL_X4 FILLER_9_893 ();
 FILLCELL_X4 FILLER_9_899 ();
 FILLCELL_X2 FILLER_9_903 ();
 FILLCELL_X1 FILLER_9_905 ();
 FILLCELL_X4 FILLER_9_913 ();
 FILLCELL_X8 FILLER_9_919 ();
 FILLCELL_X4 FILLER_9_927 ();
 FILLCELL_X4 FILLER_9_935 ();
 FILLCELL_X4 FILLER_9_942 ();
 FILLCELL_X2 FILLER_9_946 ();
 FILLCELL_X1 FILLER_9_948 ();
 FILLCELL_X4 FILLER_9_953 ();
 FILLCELL_X4 FILLER_9_966 ();
 FILLCELL_X2 FILLER_9_970 ();
 FILLCELL_X4 FILLER_9_982 ();
 FILLCELL_X4 FILLER_9_995 ();
 FILLCELL_X2 FILLER_9_999 ();
 FILLCELL_X1 FILLER_9_1001 ();
 FILLCELL_X8 FILLER_9_1005 ();
 FILLCELL_X4 FILLER_9_1013 ();
 FILLCELL_X2 FILLER_9_1017 ();
 FILLCELL_X1 FILLER_9_1019 ();
 FILLCELL_X8 FILLER_9_1023 ();
 FILLCELL_X1 FILLER_9_1031 ();
 FILLCELL_X4 FILLER_9_1039 ();
 FILLCELL_X8 FILLER_9_1046 ();
 FILLCELL_X16 FILLER_9_1056 ();
 FILLCELL_X4 FILLER_9_1072 ();
 FILLCELL_X1 FILLER_9_1076 ();
 FILLCELL_X4 FILLER_9_1087 ();
 FILLCELL_X4 FILLER_9_1098 ();
 FILLCELL_X4 FILLER_9_1105 ();
 FILLCELL_X4 FILLER_9_1112 ();
 FILLCELL_X2 FILLER_9_1116 ();
 FILLCELL_X8 FILLER_9_1122 ();
 FILLCELL_X1 FILLER_9_1130 ();
 FILLCELL_X8 FILLER_9_1134 ();
 FILLCELL_X4 FILLER_9_1142 ();
 FILLCELL_X1 FILLER_9_1146 ();
 FILLCELL_X8 FILLER_9_1150 ();
 FILLCELL_X1 FILLER_9_1158 ();
 FILLCELL_X4 FILLER_9_1162 ();
 FILLCELL_X2 FILLER_9_1166 ();
 FILLCELL_X1 FILLER_9_1168 ();
 FILLCELL_X4 FILLER_9_1172 ();
 FILLCELL_X8 FILLER_9_1185 ();
 FILLCELL_X4 FILLER_9_1193 ();
 FILLCELL_X1 FILLER_9_1197 ();
 FILLCELL_X8 FILLER_9_1208 ();
 FILLCELL_X2 FILLER_9_1216 ();
 FILLCELL_X4 FILLER_9_1225 ();
 FILLCELL_X4 FILLER_9_1232 ();
 FILLCELL_X4 FILLER_9_1239 ();
 FILLCELL_X4 FILLER_9_1246 ();
 FILLCELL_X1 FILLER_9_1250 ();
 FILLCELL_X8 FILLER_9_1255 ();
 FILLCELL_X4 FILLER_9_1264 ();
 FILLCELL_X4 FILLER_9_1278 ();
 FILLCELL_X4 FILLER_9_1292 ();
 FILLCELL_X4 FILLER_9_1305 ();
 FILLCELL_X2 FILLER_9_1309 ();
 FILLCELL_X1 FILLER_9_1311 ();
 FILLCELL_X4 FILLER_9_1316 ();
 FILLCELL_X8 FILLER_9_1323 ();
 FILLCELL_X1 FILLER_9_1331 ();
 FILLCELL_X4 FILLER_9_1342 ();
 FILLCELL_X4 FILLER_9_1356 ();
 FILLCELL_X1 FILLER_9_1360 ();
 FILLCELL_X4 FILLER_9_1364 ();
 FILLCELL_X1 FILLER_9_1368 ();
 FILLCELL_X4 FILLER_9_1371 ();
 FILLCELL_X4 FILLER_9_1379 ();
 FILLCELL_X8 FILLER_9_1387 ();
 FILLCELL_X4 FILLER_9_1395 ();
 FILLCELL_X1 FILLER_9_1399 ();
 FILLCELL_X4 FILLER_9_1410 ();
 FILLCELL_X4 FILLER_9_1418 ();
 FILLCELL_X4 FILLER_9_1425 ();
 FILLCELL_X8 FILLER_9_1432 ();
 FILLCELL_X4 FILLER_9_1443 ();
 FILLCELL_X8 FILLER_9_1450 ();
 FILLCELL_X2 FILLER_9_1458 ();
 FILLCELL_X4 FILLER_9_1466 ();
 FILLCELL_X4 FILLER_9_1476 ();
 FILLCELL_X32 FILLER_9_1484 ();
 FILLCELL_X32 FILLER_9_1516 ();
 FILLCELL_X32 FILLER_9_1548 ();
 FILLCELL_X32 FILLER_9_1580 ();
 FILLCELL_X32 FILLER_9_1612 ();
 FILLCELL_X32 FILLER_9_1644 ();
 FILLCELL_X32 FILLER_9_1676 ();
 FILLCELL_X32 FILLER_9_1708 ();
 FILLCELL_X16 FILLER_9_1740 ();
 FILLCELL_X4 FILLER_9_1756 ();
 FILLCELL_X2 FILLER_9_1760 ();
 FILLCELL_X16 FILLER_10_1 ();
 FILLCELL_X4 FILLER_10_17 ();
 FILLCELL_X2 FILLER_10_21 ();
 FILLCELL_X1 FILLER_10_23 ();
 FILLCELL_X4 FILLER_10_27 ();
 FILLCELL_X1 FILLER_10_31 ();
 FILLCELL_X4 FILLER_10_42 ();
 FILLCELL_X2 FILLER_10_46 ();
 FILLCELL_X4 FILLER_10_57 ();
 FILLCELL_X4 FILLER_10_71 ();
 FILLCELL_X4 FILLER_10_82 ();
 FILLCELL_X1 FILLER_10_86 ();
 FILLCELL_X8 FILLER_10_96 ();
 FILLCELL_X4 FILLER_10_114 ();
 FILLCELL_X8 FILLER_10_124 ();
 FILLCELL_X2 FILLER_10_132 ();
 FILLCELL_X1 FILLER_10_134 ();
 FILLCELL_X4 FILLER_10_145 ();
 FILLCELL_X2 FILLER_10_149 ();
 FILLCELL_X4 FILLER_10_160 ();
 FILLCELL_X4 FILLER_10_168 ();
 FILLCELL_X4 FILLER_10_175 ();
 FILLCELL_X2 FILLER_10_179 ();
 FILLCELL_X1 FILLER_10_181 ();
 FILLCELL_X8 FILLER_10_191 ();
 FILLCELL_X8 FILLER_10_209 ();
 FILLCELL_X4 FILLER_10_221 ();
 FILLCELL_X4 FILLER_10_232 ();
 FILLCELL_X2 FILLER_10_236 ();
 FILLCELL_X4 FILLER_10_241 ();
 FILLCELL_X4 FILLER_10_249 ();
 FILLCELL_X32 FILLER_10_257 ();
 FILLCELL_X8 FILLER_10_289 ();
 FILLCELL_X4 FILLER_10_300 ();
 FILLCELL_X8 FILLER_10_311 ();
 FILLCELL_X2 FILLER_10_319 ();
 FILLCELL_X1 FILLER_10_321 ();
 FILLCELL_X16 FILLER_10_325 ();
 FILLCELL_X4 FILLER_10_344 ();
 FILLCELL_X4 FILLER_10_352 ();
 FILLCELL_X4 FILLER_10_365 ();
 FILLCELL_X16 FILLER_10_378 ();
 FILLCELL_X2 FILLER_10_394 ();
 FILLCELL_X1 FILLER_10_396 ();
 FILLCELL_X8 FILLER_10_400 ();
 FILLCELL_X2 FILLER_10_408 ();
 FILLCELL_X4 FILLER_10_414 ();
 FILLCELL_X4 FILLER_10_421 ();
 FILLCELL_X4 FILLER_10_427 ();
 FILLCELL_X2 FILLER_10_431 ();
 FILLCELL_X1 FILLER_10_433 ();
 FILLCELL_X8 FILLER_10_444 ();
 FILLCELL_X4 FILLER_10_452 ();
 FILLCELL_X4 FILLER_10_460 ();
 FILLCELL_X8 FILLER_10_473 ();
 FILLCELL_X2 FILLER_10_481 ();
 FILLCELL_X1 FILLER_10_483 ();
 FILLCELL_X4 FILLER_10_488 ();
 FILLCELL_X1 FILLER_10_492 ();
 FILLCELL_X8 FILLER_10_497 ();
 FILLCELL_X2 FILLER_10_505 ();
 FILLCELL_X1 FILLER_10_507 ();
 FILLCELL_X4 FILLER_10_512 ();
 FILLCELL_X4 FILLER_10_525 ();
 FILLCELL_X16 FILLER_10_538 ();
 FILLCELL_X8 FILLER_10_554 ();
 FILLCELL_X2 FILLER_10_562 ();
 FILLCELL_X8 FILLER_10_571 ();
 FILLCELL_X8 FILLER_10_582 ();
 FILLCELL_X4 FILLER_10_590 ();
 FILLCELL_X16 FILLER_10_598 ();
 FILLCELL_X2 FILLER_10_614 ();
 FILLCELL_X1 FILLER_10_616 ();
 FILLCELL_X4 FILLER_10_620 ();
 FILLCELL_X4 FILLER_10_627 ();
 FILLCELL_X4 FILLER_10_632 ();
 FILLCELL_X4 FILLER_10_640 ();
 FILLCELL_X2 FILLER_10_644 ();
 FILLCELL_X1 FILLER_10_646 ();
 FILLCELL_X4 FILLER_10_651 ();
 FILLCELL_X16 FILLER_10_674 ();
 FILLCELL_X2 FILLER_10_690 ();
 FILLCELL_X4 FILLER_10_696 ();
 FILLCELL_X4 FILLER_10_709 ();
 FILLCELL_X4 FILLER_10_722 ();
 FILLCELL_X4 FILLER_10_729 ();
 FILLCELL_X4 FILLER_10_737 ();
 FILLCELL_X4 FILLER_10_745 ();
 FILLCELL_X1 FILLER_10_749 ();
 FILLCELL_X4 FILLER_10_755 ();
 FILLCELL_X4 FILLER_10_768 ();
 FILLCELL_X8 FILLER_10_781 ();
 FILLCELL_X4 FILLER_10_799 ();
 FILLCELL_X4 FILLER_10_810 ();
 FILLCELL_X2 FILLER_10_814 ();
 FILLCELL_X1 FILLER_10_816 ();
 FILLCELL_X4 FILLER_10_827 ();
 FILLCELL_X8 FILLER_10_834 ();
 FILLCELL_X4 FILLER_10_844 ();
 FILLCELL_X1 FILLER_10_848 ();
 FILLCELL_X8 FILLER_10_859 ();
 FILLCELL_X2 FILLER_10_867 ();
 FILLCELL_X8 FILLER_10_872 ();
 FILLCELL_X4 FILLER_10_880 ();
 FILLCELL_X2 FILLER_10_884 ();
 FILLCELL_X8 FILLER_10_890 ();
 FILLCELL_X4 FILLER_10_898 ();
 FILLCELL_X2 FILLER_10_902 ();
 FILLCELL_X1 FILLER_10_904 ();
 FILLCELL_X4 FILLER_10_915 ();
 FILLCELL_X8 FILLER_10_929 ();
 FILLCELL_X8 FILLER_10_947 ();
 FILLCELL_X4 FILLER_10_965 ();
 FILLCELL_X1 FILLER_10_969 ();
 FILLCELL_X8 FILLER_10_979 ();
 FILLCELL_X4 FILLER_10_987 ();
 FILLCELL_X2 FILLER_10_991 ();
 FILLCELL_X1 FILLER_10_993 ();
 FILLCELL_X4 FILLER_10_997 ();
 FILLCELL_X4 FILLER_10_1011 ();
 FILLCELL_X2 FILLER_10_1015 ();
 FILLCELL_X1 FILLER_10_1017 ();
 FILLCELL_X4 FILLER_10_1021 ();
 FILLCELL_X4 FILLER_10_1034 ();
 FILLCELL_X2 FILLER_10_1038 ();
 FILLCELL_X4 FILLER_10_1050 ();
 FILLCELL_X4 FILLER_10_1073 ();
 FILLCELL_X4 FILLER_10_1086 ();
 FILLCELL_X4 FILLER_10_1094 ();
 FILLCELL_X8 FILLER_10_1102 ();
 FILLCELL_X2 FILLER_10_1110 ();
 FILLCELL_X8 FILLER_10_1116 ();
 FILLCELL_X1 FILLER_10_1124 ();
 FILLCELL_X4 FILLER_10_1134 ();
 FILLCELL_X4 FILLER_10_1141 ();
 FILLCELL_X4 FILLER_10_1148 ();
 FILLCELL_X1 FILLER_10_1152 ();
 FILLCELL_X4 FILLER_10_1157 ();
 FILLCELL_X2 FILLER_10_1161 ();
 FILLCELL_X1 FILLER_10_1163 ();
 FILLCELL_X4 FILLER_10_1174 ();
 FILLCELL_X2 FILLER_10_1178 ();
 FILLCELL_X4 FILLER_10_1185 ();
 FILLCELL_X4 FILLER_10_1192 ();
 FILLCELL_X16 FILLER_10_1199 ();
 FILLCELL_X8 FILLER_10_1225 ();
 FILLCELL_X1 FILLER_10_1233 ();
 FILLCELL_X4 FILLER_10_1243 ();
 FILLCELL_X8 FILLER_10_1250 ();
 FILLCELL_X1 FILLER_10_1258 ();
 FILLCELL_X8 FILLER_10_1266 ();
 FILLCELL_X2 FILLER_10_1274 ();
 FILLCELL_X1 FILLER_10_1276 ();
 FILLCELL_X8 FILLER_10_1280 ();
 FILLCELL_X4 FILLER_10_1291 ();
 FILLCELL_X2 FILLER_10_1295 ();
 FILLCELL_X1 FILLER_10_1297 ();
 FILLCELL_X4 FILLER_10_1315 ();
 FILLCELL_X4 FILLER_10_1329 ();
 FILLCELL_X2 FILLER_10_1333 ();
 FILLCELL_X4 FILLER_10_1337 ();
 FILLCELL_X4 FILLER_10_1345 ();
 FILLCELL_X2 FILLER_10_1349 ();
 FILLCELL_X1 FILLER_10_1351 ();
 FILLCELL_X8 FILLER_10_1355 ();
 FILLCELL_X4 FILLER_10_1363 ();
 FILLCELL_X2 FILLER_10_1367 ();
 FILLCELL_X1 FILLER_10_1369 ();
 FILLCELL_X8 FILLER_10_1380 ();
 FILLCELL_X4 FILLER_10_1388 ();
 FILLCELL_X2 FILLER_10_1392 ();
 FILLCELL_X4 FILLER_10_1396 ();
 FILLCELL_X2 FILLER_10_1400 ();
 FILLCELL_X8 FILLER_10_1406 ();
 FILLCELL_X4 FILLER_10_1423 ();
 FILLCELL_X4 FILLER_10_1436 ();
 FILLCELL_X8 FILLER_10_1449 ();
 FILLCELL_X2 FILLER_10_1457 ();
 FILLCELL_X4 FILLER_10_1465 ();
 FILLCELL_X4 FILLER_10_1476 ();
 FILLCELL_X32 FILLER_10_1484 ();
 FILLCELL_X32 FILLER_10_1516 ();
 FILLCELL_X32 FILLER_10_1548 ();
 FILLCELL_X32 FILLER_10_1580 ();
 FILLCELL_X32 FILLER_10_1612 ();
 FILLCELL_X32 FILLER_10_1644 ();
 FILLCELL_X32 FILLER_10_1676 ();
 FILLCELL_X32 FILLER_10_1708 ();
 FILLCELL_X16 FILLER_10_1740 ();
 FILLCELL_X4 FILLER_10_1756 ();
 FILLCELL_X2 FILLER_10_1760 ();
 FILLCELL_X8 FILLER_11_1 ();
 FILLCELL_X4 FILLER_11_9 ();
 FILLCELL_X4 FILLER_11_17 ();
 FILLCELL_X4 FILLER_11_31 ();
 FILLCELL_X8 FILLER_11_42 ();
 FILLCELL_X2 FILLER_11_50 ();
 FILLCELL_X4 FILLER_11_55 ();
 FILLCELL_X4 FILLER_11_62 ();
 FILLCELL_X8 FILLER_11_68 ();
 FILLCELL_X2 FILLER_11_76 ();
 FILLCELL_X1 FILLER_11_78 ();
 FILLCELL_X4 FILLER_11_81 ();
 FILLCELL_X8 FILLER_11_95 ();
 FILLCELL_X4 FILLER_11_107 ();
 FILLCELL_X4 FILLER_11_117 ();
 FILLCELL_X4 FILLER_11_128 ();
 FILLCELL_X4 FILLER_11_136 ();
 FILLCELL_X8 FILLER_11_143 ();
 FILLCELL_X2 FILLER_11_151 ();
 FILLCELL_X4 FILLER_11_156 ();
 FILLCELL_X4 FILLER_11_163 ();
 FILLCELL_X4 FILLER_11_176 ();
 FILLCELL_X8 FILLER_11_184 ();
 FILLCELL_X4 FILLER_11_192 ();
 FILLCELL_X2 FILLER_11_196 ();
 FILLCELL_X1 FILLER_11_198 ();
 FILLCELL_X4 FILLER_11_202 ();
 FILLCELL_X4 FILLER_11_210 ();
 FILLCELL_X4 FILLER_11_219 ();
 FILLCELL_X4 FILLER_11_240 ();
 FILLCELL_X4 FILLER_11_253 ();
 FILLCELL_X4 FILLER_11_266 ();
 FILLCELL_X4 FILLER_11_274 ();
 FILLCELL_X4 FILLER_11_285 ();
 FILLCELL_X4 FILLER_11_291 ();
 FILLCELL_X4 FILLER_11_305 ();
 FILLCELL_X1 FILLER_11_309 ();
 FILLCELL_X4 FILLER_11_320 ();
 FILLCELL_X2 FILLER_11_324 ();
 FILLCELL_X1 FILLER_11_326 ();
 FILLCELL_X4 FILLER_11_331 ();
 FILLCELL_X16 FILLER_11_339 ();
 FILLCELL_X4 FILLER_11_358 ();
 FILLCELL_X16 FILLER_11_365 ();
 FILLCELL_X2 FILLER_11_381 ();
 FILLCELL_X16 FILLER_11_387 ();
 FILLCELL_X4 FILLER_11_403 ();
 FILLCELL_X4 FILLER_11_414 ();
 FILLCELL_X4 FILLER_11_420 ();
 FILLCELL_X2 FILLER_11_424 ();
 FILLCELL_X1 FILLER_11_426 ();
 FILLCELL_X4 FILLER_11_430 ();
 FILLCELL_X4 FILLER_11_437 ();
 FILLCELL_X2 FILLER_11_441 ();
 FILLCELL_X4 FILLER_11_446 ();
 FILLCELL_X4 FILLER_11_454 ();
 FILLCELL_X4 FILLER_11_467 ();
 FILLCELL_X8 FILLER_11_475 ();
 FILLCELL_X4 FILLER_11_492 ();
 FILLCELL_X8 FILLER_11_505 ();
 FILLCELL_X4 FILLER_11_513 ();
 FILLCELL_X4 FILLER_11_520 ();
 FILLCELL_X16 FILLER_11_527 ();
 FILLCELL_X4 FILLER_11_543 ();
 FILLCELL_X2 FILLER_11_547 ();
 FILLCELL_X4 FILLER_11_552 ();
 FILLCELL_X8 FILLER_11_566 ();
 FILLCELL_X1 FILLER_11_574 ();
 FILLCELL_X16 FILLER_11_585 ();
 FILLCELL_X4 FILLER_11_601 ();
 FILLCELL_X8 FILLER_11_624 ();
 FILLCELL_X4 FILLER_11_632 ();
 FILLCELL_X4 FILLER_11_639 ();
 FILLCELL_X8 FILLER_11_649 ();
 FILLCELL_X2 FILLER_11_657 ();
 FILLCELL_X4 FILLER_11_663 ();
 FILLCELL_X16 FILLER_11_671 ();
 FILLCELL_X2 FILLER_11_687 ();
 FILLCELL_X4 FILLER_11_692 ();
 FILLCELL_X1 FILLER_11_696 ();
 FILLCELL_X4 FILLER_11_701 ();
 FILLCELL_X16 FILLER_11_707 ();
 FILLCELL_X4 FILLER_11_723 ();
 FILLCELL_X1 FILLER_11_727 ();
 FILLCELL_X16 FILLER_11_731 ();
 FILLCELL_X2 FILLER_11_747 ();
 FILLCELL_X1 FILLER_11_749 ();
 FILLCELL_X4 FILLER_11_753 ();
 FILLCELL_X4 FILLER_11_761 ();
 FILLCELL_X8 FILLER_11_768 ();
 FILLCELL_X4 FILLER_11_776 ();
 FILLCELL_X2 FILLER_11_780 ();
 FILLCELL_X1 FILLER_11_782 ();
 FILLCELL_X16 FILLER_11_787 ();
 FILLCELL_X4 FILLER_11_803 ();
 FILLCELL_X4 FILLER_11_817 ();
 FILLCELL_X8 FILLER_11_825 ();
 FILLCELL_X1 FILLER_11_833 ();
 FILLCELL_X4 FILLER_11_844 ();
 FILLCELL_X8 FILLER_11_851 ();
 FILLCELL_X4 FILLER_11_859 ();
 FILLCELL_X2 FILLER_11_863 ();
 FILLCELL_X1 FILLER_11_865 ();
 FILLCELL_X8 FILLER_11_869 ();
 FILLCELL_X4 FILLER_11_877 ();
 FILLCELL_X1 FILLER_11_881 ();
 FILLCELL_X4 FILLER_11_892 ();
 FILLCELL_X4 FILLER_11_906 ();
 FILLCELL_X8 FILLER_11_912 ();
 FILLCELL_X4 FILLER_11_920 ();
 FILLCELL_X2 FILLER_11_924 ();
 FILLCELL_X1 FILLER_11_926 ();
 FILLCELL_X4 FILLER_11_930 ();
 FILLCELL_X2 FILLER_11_934 ();
 FILLCELL_X1 FILLER_11_936 ();
 FILLCELL_X4 FILLER_11_950 ();
 FILLCELL_X1 FILLER_11_954 ();
 FILLCELL_X4 FILLER_11_958 ();
 FILLCELL_X4 FILLER_11_969 ();
 FILLCELL_X8 FILLER_11_975 ();
 FILLCELL_X2 FILLER_11_983 ();
 FILLCELL_X1 FILLER_11_985 ();
 FILLCELL_X4 FILLER_11_989 ();
 FILLCELL_X1 FILLER_11_993 ();
 FILLCELL_X16 FILLER_11_1003 ();
 FILLCELL_X4 FILLER_11_1019 ();
 FILLCELL_X2 FILLER_11_1023 ();
 FILLCELL_X1 FILLER_11_1025 ();
 FILLCELL_X4 FILLER_11_1035 ();
 FILLCELL_X16 FILLER_11_1041 ();
 FILLCELL_X4 FILLER_11_1057 ();
 FILLCELL_X2 FILLER_11_1061 ();
 FILLCELL_X4 FILLER_11_1066 ();
 FILLCELL_X4 FILLER_11_1073 ();
 FILLCELL_X8 FILLER_11_1080 ();
 FILLCELL_X4 FILLER_11_1091 ();
 FILLCELL_X16 FILLER_11_1105 ();
 FILLCELL_X1 FILLER_11_1121 ();
 FILLCELL_X4 FILLER_11_1126 ();
 FILLCELL_X4 FILLER_11_1133 ();
 FILLCELL_X2 FILLER_11_1137 ();
 FILLCELL_X1 FILLER_11_1139 ();
 FILLCELL_X4 FILLER_11_1144 ();
 FILLCELL_X4 FILLER_11_1157 ();
 FILLCELL_X4 FILLER_11_1170 ();
 FILLCELL_X8 FILLER_11_1178 ();
 FILLCELL_X1 FILLER_11_1186 ();
 FILLCELL_X8 FILLER_11_1194 ();
 FILLCELL_X4 FILLER_11_1202 ();
 FILLCELL_X4 FILLER_11_1215 ();
 FILLCELL_X2 FILLER_11_1219 ();
 FILLCELL_X8 FILLER_11_1224 ();
 FILLCELL_X1 FILLER_11_1232 ();
 FILLCELL_X4 FILLER_11_1242 ();
 FILLCELL_X8 FILLER_11_1249 ();
 FILLCELL_X4 FILLER_11_1259 ();
 FILLCELL_X4 FILLER_11_1264 ();
 FILLCELL_X16 FILLER_11_1278 ();
 FILLCELL_X1 FILLER_11_1294 ();
 FILLCELL_X4 FILLER_11_1297 ();
 FILLCELL_X4 FILLER_11_1306 ();
 FILLCELL_X4 FILLER_11_1315 ();
 FILLCELL_X1 FILLER_11_1319 ();
 FILLCELL_X16 FILLER_11_1327 ();
 FILLCELL_X1 FILLER_11_1343 ();
 FILLCELL_X16 FILLER_11_1349 ();
 FILLCELL_X8 FILLER_11_1365 ();
 FILLCELL_X2 FILLER_11_1373 ();
 FILLCELL_X8 FILLER_11_1378 ();
 FILLCELL_X16 FILLER_11_1396 ();
 FILLCELL_X2 FILLER_11_1412 ();
 FILLCELL_X1 FILLER_11_1414 ();
 FILLCELL_X4 FILLER_11_1424 ();
 FILLCELL_X4 FILLER_11_1431 ();
 FILLCELL_X8 FILLER_11_1438 ();
 FILLCELL_X4 FILLER_11_1446 ();
 FILLCELL_X1 FILLER_11_1450 ();
 FILLCELL_X4 FILLER_11_1453 ();
 FILLCELL_X4 FILLER_11_1467 ();
 FILLCELL_X4 FILLER_11_1478 ();
 FILLCELL_X2 FILLER_11_1482 ();
 FILLCELL_X32 FILLER_11_1501 ();
 FILLCELL_X32 FILLER_11_1533 ();
 FILLCELL_X32 FILLER_11_1565 ();
 FILLCELL_X32 FILLER_11_1597 ();
 FILLCELL_X32 FILLER_11_1629 ();
 FILLCELL_X32 FILLER_11_1661 ();
 FILLCELL_X32 FILLER_11_1693 ();
 FILLCELL_X16 FILLER_11_1725 ();
 FILLCELL_X8 FILLER_11_1741 ();
 FILLCELL_X4 FILLER_11_1749 ();
 FILLCELL_X2 FILLER_11_1753 ();
 FILLCELL_X4 FILLER_11_1758 ();
 FILLCELL_X8 FILLER_12_1 ();
 FILLCELL_X16 FILLER_12_12 ();
 FILLCELL_X8 FILLER_12_28 ();
 FILLCELL_X2 FILLER_12_36 ();
 FILLCELL_X4 FILLER_12_48 ();
 FILLCELL_X8 FILLER_12_54 ();
 FILLCELL_X2 FILLER_12_62 ();
 FILLCELL_X1 FILLER_12_64 ();
 FILLCELL_X16 FILLER_12_67 ();
 FILLCELL_X2 FILLER_12_83 ();
 FILLCELL_X8 FILLER_12_92 ();
 FILLCELL_X1 FILLER_12_100 ();
 FILLCELL_X4 FILLER_12_105 ();
 FILLCELL_X4 FILLER_12_111 ();
 FILLCELL_X32 FILLER_12_119 ();
 FILLCELL_X4 FILLER_12_161 ();
 FILLCELL_X4 FILLER_12_167 ();
 FILLCELL_X4 FILLER_12_174 ();
 FILLCELL_X4 FILLER_12_181 ();
 FILLCELL_X2 FILLER_12_185 ();
 FILLCELL_X1 FILLER_12_187 ();
 FILLCELL_X4 FILLER_12_192 ();
 FILLCELL_X16 FILLER_12_205 ();
 FILLCELL_X2 FILLER_12_221 ();
 FILLCELL_X1 FILLER_12_223 ();
 FILLCELL_X4 FILLER_12_229 ();
 FILLCELL_X8 FILLER_12_237 ();
 FILLCELL_X1 FILLER_12_245 ();
 FILLCELL_X4 FILLER_12_250 ();
 FILLCELL_X2 FILLER_12_254 ();
 FILLCELL_X1 FILLER_12_256 ();
 FILLCELL_X4 FILLER_12_260 ();
 FILLCELL_X2 FILLER_12_264 ();
 FILLCELL_X1 FILLER_12_266 ();
 FILLCELL_X4 FILLER_12_270 ();
 FILLCELL_X4 FILLER_12_284 ();
 FILLCELL_X2 FILLER_12_288 ();
 FILLCELL_X1 FILLER_12_290 ();
 FILLCELL_X4 FILLER_12_295 ();
 FILLCELL_X8 FILLER_12_309 ();
 FILLCELL_X4 FILLER_12_321 ();
 FILLCELL_X4 FILLER_12_334 ();
 FILLCELL_X8 FILLER_12_347 ();
 FILLCELL_X4 FILLER_12_355 ();
 FILLCELL_X2 FILLER_12_359 ();
 FILLCELL_X4 FILLER_12_363 ();
 FILLCELL_X1 FILLER_12_367 ();
 FILLCELL_X4 FILLER_12_371 ();
 FILLCELL_X4 FILLER_12_378 ();
 FILLCELL_X4 FILLER_12_392 ();
 FILLCELL_X4 FILLER_12_400 ();
 FILLCELL_X8 FILLER_12_414 ();
 FILLCELL_X1 FILLER_12_422 ();
 FILLCELL_X4 FILLER_12_432 ();
 FILLCELL_X2 FILLER_12_436 ();
 FILLCELL_X1 FILLER_12_438 ();
 FILLCELL_X8 FILLER_12_444 ();
 FILLCELL_X4 FILLER_12_452 ();
 FILLCELL_X4 FILLER_12_459 ();
 FILLCELL_X4 FILLER_12_466 ();
 FILLCELL_X4 FILLER_12_473 ();
 FILLCELL_X4 FILLER_12_481 ();
 FILLCELL_X4 FILLER_12_489 ();
 FILLCELL_X4 FILLER_12_496 ();
 FILLCELL_X2 FILLER_12_500 ();
 FILLCELL_X4 FILLER_12_506 ();
 FILLCELL_X8 FILLER_12_529 ();
 FILLCELL_X4 FILLER_12_537 ();
 FILLCELL_X4 FILLER_12_547 ();
 FILLCELL_X1 FILLER_12_551 ();
 FILLCELL_X8 FILLER_12_556 ();
 FILLCELL_X4 FILLER_12_564 ();
 FILLCELL_X2 FILLER_12_568 ();
 FILLCELL_X1 FILLER_12_570 ();
 FILLCELL_X16 FILLER_12_573 ();
 FILLCELL_X4 FILLER_12_589 ();
 FILLCELL_X2 FILLER_12_593 ();
 FILLCELL_X4 FILLER_12_601 ();
 FILLCELL_X1 FILLER_12_605 ();
 FILLCELL_X16 FILLER_12_610 ();
 FILLCELL_X4 FILLER_12_626 ();
 FILLCELL_X1 FILLER_12_630 ();
 FILLCELL_X4 FILLER_12_632 ();
 FILLCELL_X4 FILLER_12_643 ();
 FILLCELL_X8 FILLER_12_653 ();
 FILLCELL_X2 FILLER_12_661 ();
 FILLCELL_X1 FILLER_12_663 ();
 FILLCELL_X4 FILLER_12_671 ();
 FILLCELL_X4 FILLER_12_684 ();
 FILLCELL_X8 FILLER_12_698 ();
 FILLCELL_X4 FILLER_12_709 ();
 FILLCELL_X8 FILLER_12_720 ();
 FILLCELL_X4 FILLER_12_731 ();
 FILLCELL_X8 FILLER_12_744 ();
 FILLCELL_X1 FILLER_12_752 ();
 FILLCELL_X4 FILLER_12_760 ();
 FILLCELL_X16 FILLER_12_774 ();
 FILLCELL_X8 FILLER_12_790 ();
 FILLCELL_X4 FILLER_12_798 ();
 FILLCELL_X2 FILLER_12_802 ();
 FILLCELL_X4 FILLER_12_813 ();
 FILLCELL_X4 FILLER_12_820 ();
 FILLCELL_X2 FILLER_12_824 ();
 FILLCELL_X1 FILLER_12_826 ();
 FILLCELL_X4 FILLER_12_829 ();
 FILLCELL_X2 FILLER_12_833 ();
 FILLCELL_X8 FILLER_12_839 ();
 FILLCELL_X4 FILLER_12_847 ();
 FILLCELL_X1 FILLER_12_851 ();
 FILLCELL_X4 FILLER_12_855 ();
 FILLCELL_X2 FILLER_12_859 ();
 FILLCELL_X4 FILLER_12_864 ();
 FILLCELL_X4 FILLER_12_881 ();
 FILLCELL_X2 FILLER_12_885 ();
 FILLCELL_X4 FILLER_12_890 ();
 FILLCELL_X4 FILLER_12_898 ();
 FILLCELL_X4 FILLER_12_906 ();
 FILLCELL_X2 FILLER_12_910 ();
 FILLCELL_X1 FILLER_12_912 ();
 FILLCELL_X4 FILLER_12_923 ();
 FILLCELL_X4 FILLER_12_936 ();
 FILLCELL_X32 FILLER_12_942 ();
 FILLCELL_X4 FILLER_12_978 ();
 FILLCELL_X4 FILLER_12_985 ();
 FILLCELL_X2 FILLER_12_989 ();
 FILLCELL_X1 FILLER_12_991 ();
 FILLCELL_X8 FILLER_12_996 ();
 FILLCELL_X2 FILLER_12_1004 ();
 FILLCELL_X1 FILLER_12_1006 ();
 FILLCELL_X4 FILLER_12_1011 ();
 FILLCELL_X4 FILLER_12_1017 ();
 FILLCELL_X4 FILLER_12_1023 ();
 FILLCELL_X4 FILLER_12_1034 ();
 FILLCELL_X4 FILLER_12_1048 ();
 FILLCELL_X8 FILLER_12_1056 ();
 FILLCELL_X2 FILLER_12_1064 ();
 FILLCELL_X1 FILLER_12_1066 ();
 FILLCELL_X16 FILLER_12_1076 ();
 FILLCELL_X4 FILLER_12_1092 ();
 FILLCELL_X1 FILLER_12_1096 ();
 FILLCELL_X4 FILLER_12_1099 ();
 FILLCELL_X4 FILLER_12_1113 ();
 FILLCELL_X1 FILLER_12_1117 ();
 FILLCELL_X4 FILLER_12_1128 ();
 FILLCELL_X4 FILLER_12_1141 ();
 FILLCELL_X4 FILLER_12_1149 ();
 FILLCELL_X4 FILLER_12_1156 ();
 FILLCELL_X2 FILLER_12_1160 ();
 FILLCELL_X1 FILLER_12_1162 ();
 FILLCELL_X8 FILLER_12_1170 ();
 FILLCELL_X2 FILLER_12_1178 ();
 FILLCELL_X4 FILLER_12_1190 ();
 FILLCELL_X1 FILLER_12_1194 ();
 FILLCELL_X4 FILLER_12_1205 ();
 FILLCELL_X8 FILLER_12_1218 ();
 FILLCELL_X1 FILLER_12_1226 ();
 FILLCELL_X4 FILLER_12_1236 ();
 FILLCELL_X1 FILLER_12_1240 ();
 FILLCELL_X4 FILLER_12_1244 ();
 FILLCELL_X1 FILLER_12_1248 ();
 FILLCELL_X8 FILLER_12_1258 ();
 FILLCELL_X4 FILLER_12_1275 ();
 FILLCELL_X4 FILLER_12_1286 ();
 FILLCELL_X2 FILLER_12_1290 ();
 FILLCELL_X4 FILLER_12_1296 ();
 FILLCELL_X4 FILLER_12_1307 ();
 FILLCELL_X4 FILLER_12_1315 ();
 FILLCELL_X1 FILLER_12_1319 ();
 FILLCELL_X8 FILLER_12_1329 ();
 FILLCELL_X4 FILLER_12_1340 ();
 FILLCELL_X4 FILLER_12_1353 ();
 FILLCELL_X8 FILLER_12_1361 ();
 FILLCELL_X4 FILLER_12_1378 ();
 FILLCELL_X8 FILLER_12_1385 ();
 FILLCELL_X1 FILLER_12_1393 ();
 FILLCELL_X4 FILLER_12_1401 ();
 FILLCELL_X8 FILLER_12_1407 ();
 FILLCELL_X2 FILLER_12_1415 ();
 FILLCELL_X1 FILLER_12_1417 ();
 FILLCELL_X8 FILLER_12_1421 ();
 FILLCELL_X1 FILLER_12_1429 ();
 FILLCELL_X4 FILLER_12_1433 ();
 FILLCELL_X8 FILLER_12_1447 ();
 FILLCELL_X4 FILLER_12_1455 ();
 FILLCELL_X2 FILLER_12_1459 ();
 FILLCELL_X8 FILLER_12_1464 ();
 FILLCELL_X4 FILLER_12_1475 ();
 FILLCELL_X32 FILLER_12_1485 ();
 FILLCELL_X32 FILLER_12_1517 ();
 FILLCELL_X32 FILLER_12_1549 ();
 FILLCELL_X32 FILLER_12_1581 ();
 FILLCELL_X32 FILLER_12_1613 ();
 FILLCELL_X32 FILLER_12_1645 ();
 FILLCELL_X32 FILLER_12_1677 ();
 FILLCELL_X32 FILLER_12_1709 ();
 FILLCELL_X16 FILLER_12_1741 ();
 FILLCELL_X4 FILLER_12_1757 ();
 FILLCELL_X1 FILLER_12_1761 ();
 FILLCELL_X4 FILLER_13_1 ();
 FILLCELL_X4 FILLER_13_8 ();
 FILLCELL_X16 FILLER_13_21 ();
 FILLCELL_X2 FILLER_13_37 ();
 FILLCELL_X4 FILLER_13_46 ();
 FILLCELL_X1 FILLER_13_50 ();
 FILLCELL_X4 FILLER_13_60 ();
 FILLCELL_X4 FILLER_13_74 ();
 FILLCELL_X4 FILLER_13_88 ();
 FILLCELL_X8 FILLER_13_102 ();
 FILLCELL_X4 FILLER_13_110 ();
 FILLCELL_X2 FILLER_13_114 ();
 FILLCELL_X4 FILLER_13_120 ();
 FILLCELL_X8 FILLER_13_128 ();
 FILLCELL_X4 FILLER_13_136 ();
 FILLCELL_X1 FILLER_13_140 ();
 FILLCELL_X4 FILLER_13_145 ();
 FILLCELL_X2 FILLER_13_149 ();
 FILLCELL_X1 FILLER_13_151 ();
 FILLCELL_X4 FILLER_13_159 ();
 FILLCELL_X2 FILLER_13_163 ();
 FILLCELL_X1 FILLER_13_165 ();
 FILLCELL_X4 FILLER_13_169 ();
 FILLCELL_X8 FILLER_13_182 ();
 FILLCELL_X4 FILLER_13_193 ();
 FILLCELL_X4 FILLER_13_206 ();
 FILLCELL_X16 FILLER_13_213 ();
 FILLCELL_X4 FILLER_13_229 ();
 FILLCELL_X1 FILLER_13_233 ();
 FILLCELL_X4 FILLER_13_236 ();
 FILLCELL_X2 FILLER_13_240 ();
 FILLCELL_X4 FILLER_13_245 ();
 FILLCELL_X4 FILLER_13_253 ();
 FILLCELL_X4 FILLER_13_261 ();
 FILLCELL_X1 FILLER_13_265 ();
 FILLCELL_X4 FILLER_13_270 ();
 FILLCELL_X16 FILLER_13_277 ();
 FILLCELL_X2 FILLER_13_293 ();
 FILLCELL_X1 FILLER_13_295 ();
 FILLCELL_X8 FILLER_13_299 ();
 FILLCELL_X2 FILLER_13_307 ();
 FILLCELL_X1 FILLER_13_309 ();
 FILLCELL_X4 FILLER_13_312 ();
 FILLCELL_X8 FILLER_13_318 ();
 FILLCELL_X4 FILLER_13_326 ();
 FILLCELL_X1 FILLER_13_330 ();
 FILLCELL_X4 FILLER_13_334 ();
 FILLCELL_X8 FILLER_13_341 ();
 FILLCELL_X4 FILLER_13_359 ();
 FILLCELL_X4 FILLER_13_367 ();
 FILLCELL_X4 FILLER_13_381 ();
 FILLCELL_X2 FILLER_13_385 ();
 FILLCELL_X1 FILLER_13_387 ();
 FILLCELL_X4 FILLER_13_391 ();
 FILLCELL_X2 FILLER_13_395 ();
 FILLCELL_X4 FILLER_13_401 ();
 FILLCELL_X8 FILLER_13_408 ();
 FILLCELL_X4 FILLER_13_416 ();
 FILLCELL_X2 FILLER_13_420 ();
 FILLCELL_X1 FILLER_13_422 ();
 FILLCELL_X4 FILLER_13_427 ();
 FILLCELL_X4 FILLER_13_440 ();
 FILLCELL_X4 FILLER_13_448 ();
 FILLCELL_X2 FILLER_13_452 ();
 FILLCELL_X1 FILLER_13_454 ();
 FILLCELL_X8 FILLER_13_459 ();
 FILLCELL_X2 FILLER_13_467 ();
 FILLCELL_X8 FILLER_13_474 ();
 FILLCELL_X1 FILLER_13_482 ();
 FILLCELL_X4 FILLER_13_488 ();
 FILLCELL_X4 FILLER_13_495 ();
 FILLCELL_X8 FILLER_13_508 ();
 FILLCELL_X4 FILLER_13_516 ();
 FILLCELL_X2 FILLER_13_520 ();
 FILLCELL_X4 FILLER_13_524 ();
 FILLCELL_X1 FILLER_13_528 ();
 FILLCELL_X4 FILLER_13_533 ();
 FILLCELL_X4 FILLER_13_544 ();
 FILLCELL_X1 FILLER_13_548 ();
 FILLCELL_X4 FILLER_13_555 ();
 FILLCELL_X4 FILLER_13_563 ();
 FILLCELL_X4 FILLER_13_584 ();
 FILLCELL_X4 FILLER_13_594 ();
 FILLCELL_X4 FILLER_13_611 ();
 FILLCELL_X16 FILLER_13_619 ();
 FILLCELL_X1 FILLER_13_635 ();
 FILLCELL_X8 FILLER_13_639 ();
 FILLCELL_X4 FILLER_13_647 ();
 FILLCELL_X8 FILLER_13_657 ();
 FILLCELL_X2 FILLER_13_665 ();
 FILLCELL_X8 FILLER_13_673 ();
 FILLCELL_X1 FILLER_13_681 ();
 FILLCELL_X4 FILLER_13_686 ();
 FILLCELL_X8 FILLER_13_700 ();
 FILLCELL_X1 FILLER_13_708 ();
 FILLCELL_X4 FILLER_13_719 ();
 FILLCELL_X8 FILLER_13_733 ();
 FILLCELL_X4 FILLER_13_741 ();
 FILLCELL_X2 FILLER_13_745 ();
 FILLCELL_X1 FILLER_13_747 ();
 FILLCELL_X8 FILLER_13_758 ();
 FILLCELL_X2 FILLER_13_766 ();
 FILLCELL_X8 FILLER_13_787 ();
 FILLCELL_X4 FILLER_13_795 ();
 FILLCELL_X4 FILLER_13_802 ();
 FILLCELL_X2 FILLER_13_806 ();
 FILLCELL_X1 FILLER_13_808 ();
 FILLCELL_X8 FILLER_13_812 ();
 FILLCELL_X2 FILLER_13_820 ();
 FILLCELL_X1 FILLER_13_822 ();
 FILLCELL_X8 FILLER_13_833 ();
 FILLCELL_X4 FILLER_13_845 ();
 FILLCELL_X4 FILLER_13_859 ();
 FILLCELL_X16 FILLER_13_869 ();
 FILLCELL_X4 FILLER_13_885 ();
 FILLCELL_X1 FILLER_13_889 ();
 FILLCELL_X4 FILLER_13_894 ();
 FILLCELL_X8 FILLER_13_911 ();
 FILLCELL_X4 FILLER_13_919 ();
 FILLCELL_X2 FILLER_13_923 ();
 FILLCELL_X8 FILLER_13_928 ();
 FILLCELL_X2 FILLER_13_936 ();
 FILLCELL_X1 FILLER_13_938 ();
 FILLCELL_X16 FILLER_13_942 ();
 FILLCELL_X4 FILLER_13_965 ();
 FILLCELL_X4 FILLER_13_973 ();
 FILLCELL_X4 FILLER_13_986 ();
 FILLCELL_X8 FILLER_13_1000 ();
 FILLCELL_X4 FILLER_13_1012 ();
 FILLCELL_X4 FILLER_13_1026 ();
 FILLCELL_X4 FILLER_13_1040 ();
 FILLCELL_X8 FILLER_13_1054 ();
 FILLCELL_X4 FILLER_13_1062 ();
 FILLCELL_X1 FILLER_13_1066 ();
 FILLCELL_X16 FILLER_13_1070 ();
 FILLCELL_X1 FILLER_13_1086 ();
 FILLCELL_X4 FILLER_13_1091 ();
 FILLCELL_X4 FILLER_13_1102 ();
 FILLCELL_X4 FILLER_13_1113 ();
 FILLCELL_X8 FILLER_13_1119 ();
 FILLCELL_X2 FILLER_13_1127 ();
 FILLCELL_X1 FILLER_13_1129 ();
 FILLCELL_X4 FILLER_13_1132 ();
 FILLCELL_X1 FILLER_13_1136 ();
 FILLCELL_X16 FILLER_13_1144 ();
 FILLCELL_X2 FILLER_13_1160 ();
 FILLCELL_X1 FILLER_13_1162 ();
 FILLCELL_X4 FILLER_13_1173 ();
 FILLCELL_X8 FILLER_13_1179 ();
 FILLCELL_X4 FILLER_13_1187 ();
 FILLCELL_X2 FILLER_13_1191 ();
 FILLCELL_X4 FILLER_13_1195 ();
 FILLCELL_X2 FILLER_13_1199 ();
 FILLCELL_X1 FILLER_13_1201 ();
 FILLCELL_X4 FILLER_13_1205 ();
 FILLCELL_X8 FILLER_13_1212 ();
 FILLCELL_X8 FILLER_13_1230 ();
 FILLCELL_X4 FILLER_13_1241 ();
 FILLCELL_X8 FILLER_13_1255 ();
 FILLCELL_X4 FILLER_13_1264 ();
 FILLCELL_X8 FILLER_13_1271 ();
 FILLCELL_X4 FILLER_13_1289 ();
 FILLCELL_X4 FILLER_13_1295 ();
 FILLCELL_X2 FILLER_13_1299 ();
 FILLCELL_X8 FILLER_13_1305 ();
 FILLCELL_X2 FILLER_13_1313 ();
 FILLCELL_X4 FILLER_13_1318 ();
 FILLCELL_X4 FILLER_13_1332 ();
 FILLCELL_X4 FILLER_13_1341 ();
 FILLCELL_X4 FILLER_13_1354 ();
 FILLCELL_X1 FILLER_13_1358 ();
 FILLCELL_X4 FILLER_13_1368 ();
 FILLCELL_X4 FILLER_13_1375 ();
 FILLCELL_X1 FILLER_13_1379 ();
 FILLCELL_X4 FILLER_13_1390 ();
 FILLCELL_X4 FILLER_13_1404 ();
 FILLCELL_X4 FILLER_13_1411 ();
 FILLCELL_X8 FILLER_13_1418 ();
 FILLCELL_X8 FILLER_13_1430 ();
 FILLCELL_X8 FILLER_13_1448 ();
 FILLCELL_X2 FILLER_13_1456 ();
 FILLCELL_X8 FILLER_13_1467 ();
 FILLCELL_X2 FILLER_13_1475 ();
 FILLCELL_X4 FILLER_13_1483 ();
 FILLCELL_X32 FILLER_13_1490 ();
 FILLCELL_X32 FILLER_13_1522 ();
 FILLCELL_X32 FILLER_13_1554 ();
 FILLCELL_X32 FILLER_13_1586 ();
 FILLCELL_X32 FILLER_13_1618 ();
 FILLCELL_X32 FILLER_13_1650 ();
 FILLCELL_X32 FILLER_13_1682 ();
 FILLCELL_X32 FILLER_13_1714 ();
 FILLCELL_X16 FILLER_13_1746 ();
 FILLCELL_X8 FILLER_14_1 ();
 FILLCELL_X4 FILLER_14_13 ();
 FILLCELL_X4 FILLER_14_21 ();
 FILLCELL_X4 FILLER_14_29 ();
 FILLCELL_X4 FILLER_14_43 ();
 FILLCELL_X4 FILLER_14_56 ();
 FILLCELL_X4 FILLER_14_63 ();
 FILLCELL_X2 FILLER_14_67 ();
 FILLCELL_X8 FILLER_14_76 ();
 FILLCELL_X1 FILLER_14_84 ();
 FILLCELL_X4 FILLER_14_88 ();
 FILLCELL_X4 FILLER_14_95 ();
 FILLCELL_X4 FILLER_14_103 ();
 FILLCELL_X4 FILLER_14_111 ();
 FILLCELL_X4 FILLER_14_124 ();
 FILLCELL_X4 FILLER_14_137 ();
 FILLCELL_X1 FILLER_14_141 ();
 FILLCELL_X8 FILLER_14_152 ();
 FILLCELL_X1 FILLER_14_160 ();
 FILLCELL_X16 FILLER_14_171 ();
 FILLCELL_X4 FILLER_14_190 ();
 FILLCELL_X2 FILLER_14_194 ();
 FILLCELL_X1 FILLER_14_196 ();
 FILLCELL_X4 FILLER_14_201 ();
 FILLCELL_X8 FILLER_14_209 ();
 FILLCELL_X4 FILLER_14_217 ();
 FILLCELL_X1 FILLER_14_221 ();
 FILLCELL_X4 FILLER_14_229 ();
 FILLCELL_X8 FILLER_14_243 ();
 FILLCELL_X2 FILLER_14_251 ();
 FILLCELL_X4 FILLER_14_262 ();
 FILLCELL_X8 FILLER_14_275 ();
 FILLCELL_X4 FILLER_14_283 ();
 FILLCELL_X2 FILLER_14_287 ();
 FILLCELL_X1 FILLER_14_289 ();
 FILLCELL_X4 FILLER_14_294 ();
 FILLCELL_X2 FILLER_14_298 ();
 FILLCELL_X1 FILLER_14_300 ();
 FILLCELL_X4 FILLER_14_304 ();
 FILLCELL_X1 FILLER_14_308 ();
 FILLCELL_X4 FILLER_14_314 ();
 FILLCELL_X2 FILLER_14_318 ();
 FILLCELL_X8 FILLER_14_329 ();
 FILLCELL_X4 FILLER_14_337 ();
 FILLCELL_X2 FILLER_14_341 ();
 FILLCELL_X1 FILLER_14_343 ();
 FILLCELL_X4 FILLER_14_347 ();
 FILLCELL_X1 FILLER_14_351 ();
 FILLCELL_X8 FILLER_14_355 ();
 FILLCELL_X1 FILLER_14_363 ();
 FILLCELL_X4 FILLER_14_366 ();
 FILLCELL_X2 FILLER_14_370 ();
 FILLCELL_X8 FILLER_14_376 ();
 FILLCELL_X1 FILLER_14_384 ();
 FILLCELL_X8 FILLER_14_395 ();
 FILLCELL_X16 FILLER_14_413 ();
 FILLCELL_X4 FILLER_14_429 ();
 FILLCELL_X4 FILLER_14_437 ();
 FILLCELL_X2 FILLER_14_441 ();
 FILLCELL_X1 FILLER_14_443 ();
 FILLCELL_X8 FILLER_14_453 ();
 FILLCELL_X4 FILLER_14_470 ();
 FILLCELL_X2 FILLER_14_474 ();
 FILLCELL_X16 FILLER_14_485 ();
 FILLCELL_X4 FILLER_14_501 ();
 FILLCELL_X4 FILLER_14_515 ();
 FILLCELL_X4 FILLER_14_526 ();
 FILLCELL_X4 FILLER_14_536 ();
 FILLCELL_X16 FILLER_14_544 ();
 FILLCELL_X8 FILLER_14_560 ();
 FILLCELL_X8 FILLER_14_572 ();
 FILLCELL_X4 FILLER_14_590 ();
 FILLCELL_X4 FILLER_14_596 ();
 FILLCELL_X4 FILLER_14_604 ();
 FILLCELL_X4 FILLER_14_627 ();
 FILLCELL_X8 FILLER_14_632 ();
 FILLCELL_X2 FILLER_14_640 ();
 FILLCELL_X1 FILLER_14_642 ();
 FILLCELL_X4 FILLER_14_647 ();
 FILLCELL_X4 FILLER_14_654 ();
 FILLCELL_X2 FILLER_14_658 ();
 FILLCELL_X1 FILLER_14_660 ();
 FILLCELL_X4 FILLER_14_664 ();
 FILLCELL_X4 FILLER_14_671 ();
 FILLCELL_X8 FILLER_14_681 ();
 FILLCELL_X2 FILLER_14_689 ();
 FILLCELL_X1 FILLER_14_691 ();
 FILLCELL_X8 FILLER_14_695 ();
 FILLCELL_X2 FILLER_14_703 ();
 FILLCELL_X1 FILLER_14_705 ();
 FILLCELL_X4 FILLER_14_708 ();
 FILLCELL_X4 FILLER_14_716 ();
 FILLCELL_X4 FILLER_14_722 ();
 FILLCELL_X1 FILLER_14_726 ();
 FILLCELL_X4 FILLER_14_730 ();
 FILLCELL_X8 FILLER_14_743 ();
 FILLCELL_X4 FILLER_14_751 ();
 FILLCELL_X4 FILLER_14_757 ();
 FILLCELL_X2 FILLER_14_761 ();
 FILLCELL_X8 FILLER_14_766 ();
 FILLCELL_X4 FILLER_14_774 ();
 FILLCELL_X2 FILLER_14_778 ();
 FILLCELL_X1 FILLER_14_780 ();
 FILLCELL_X8 FILLER_14_800 ();
 FILLCELL_X2 FILLER_14_808 ();
 FILLCELL_X4 FILLER_14_813 ();
 FILLCELL_X4 FILLER_14_820 ();
 FILLCELL_X4 FILLER_14_827 ();
 FILLCELL_X4 FILLER_14_841 ();
 FILLCELL_X4 FILLER_14_847 ();
 FILLCELL_X2 FILLER_14_851 ();
 FILLCELL_X16 FILLER_14_859 ();
 FILLCELL_X8 FILLER_14_888 ();
 FILLCELL_X2 FILLER_14_896 ();
 FILLCELL_X1 FILLER_14_898 ();
 FILLCELL_X16 FILLER_14_905 ();
 FILLCELL_X4 FILLER_14_921 ();
 FILLCELL_X2 FILLER_14_925 ();
 FILLCELL_X4 FILLER_14_930 ();
 FILLCELL_X4 FILLER_14_937 ();
 FILLCELL_X4 FILLER_14_950 ();
 FILLCELL_X4 FILLER_14_964 ();
 FILLCELL_X4 FILLER_14_978 ();
 FILLCELL_X4 FILLER_14_985 ();
 FILLCELL_X2 FILLER_14_989 ();
 FILLCELL_X1 FILLER_14_991 ();
 FILLCELL_X8 FILLER_14_995 ();
 FILLCELL_X8 FILLER_14_1013 ();
 FILLCELL_X4 FILLER_14_1021 ();
 FILLCELL_X2 FILLER_14_1025 ();
 FILLCELL_X4 FILLER_14_1030 ();
 FILLCELL_X2 FILLER_14_1034 ();
 FILLCELL_X8 FILLER_14_1038 ();
 FILLCELL_X2 FILLER_14_1046 ();
 FILLCELL_X4 FILLER_14_1051 ();
 FILLCELL_X8 FILLER_14_1064 ();
 FILLCELL_X4 FILLER_14_1082 ();
 FILLCELL_X2 FILLER_14_1086 ();
 FILLCELL_X1 FILLER_14_1088 ();
 FILLCELL_X4 FILLER_14_1099 ();
 FILLCELL_X8 FILLER_14_1107 ();
 FILLCELL_X4 FILLER_14_1119 ();
 FILLCELL_X4 FILLER_14_1126 ();
 FILLCELL_X8 FILLER_14_1140 ();
 FILLCELL_X4 FILLER_14_1158 ();
 FILLCELL_X16 FILLER_14_1165 ();
 FILLCELL_X8 FILLER_14_1181 ();
 FILLCELL_X1 FILLER_14_1189 ();
 FILLCELL_X8 FILLER_14_1193 ();
 FILLCELL_X2 FILLER_14_1201 ();
 FILLCELL_X1 FILLER_14_1203 ();
 FILLCELL_X4 FILLER_14_1207 ();
 FILLCELL_X1 FILLER_14_1211 ();
 FILLCELL_X32 FILLER_14_1215 ();
 FILLCELL_X8 FILLER_14_1247 ();
 FILLCELL_X4 FILLER_14_1255 ();
 FILLCELL_X2 FILLER_14_1259 ();
 FILLCELL_X1 FILLER_14_1261 ();
 FILLCELL_X4 FILLER_14_1265 ();
 FILLCELL_X4 FILLER_14_1272 ();
 FILLCELL_X2 FILLER_14_1276 ();
 FILLCELL_X4 FILLER_14_1281 ();
 FILLCELL_X16 FILLER_14_1295 ();
 FILLCELL_X8 FILLER_14_1311 ();
 FILLCELL_X4 FILLER_14_1322 ();
 FILLCELL_X8 FILLER_14_1328 ();
 FILLCELL_X2 FILLER_14_1336 ();
 FILLCELL_X1 FILLER_14_1338 ();
 FILLCELL_X4 FILLER_14_1342 ();
 FILLCELL_X4 FILLER_14_1350 ();
 FILLCELL_X32 FILLER_14_1358 ();
 FILLCELL_X4 FILLER_14_1390 ();
 FILLCELL_X1 FILLER_14_1394 ();
 FILLCELL_X4 FILLER_14_1399 ();
 FILLCELL_X1 FILLER_14_1403 ();
 FILLCELL_X4 FILLER_14_1413 ();
 FILLCELL_X4 FILLER_14_1421 ();
 FILLCELL_X8 FILLER_14_1428 ();
 FILLCELL_X4 FILLER_14_1439 ();
 FILLCELL_X1 FILLER_14_1443 ();
 FILLCELL_X4 FILLER_14_1451 ();
 FILLCELL_X4 FILLER_14_1457 ();
 FILLCELL_X1 FILLER_14_1461 ();
 FILLCELL_X8 FILLER_14_1465 ();
 FILLCELL_X2 FILLER_14_1473 ();
 FILLCELL_X1 FILLER_14_1475 ();
 FILLCELL_X32 FILLER_14_1483 ();
 FILLCELL_X32 FILLER_14_1515 ();
 FILLCELL_X32 FILLER_14_1547 ();
 FILLCELL_X32 FILLER_14_1579 ();
 FILLCELL_X32 FILLER_14_1611 ();
 FILLCELL_X32 FILLER_14_1643 ();
 FILLCELL_X32 FILLER_14_1675 ();
 FILLCELL_X32 FILLER_14_1707 ();
 FILLCELL_X16 FILLER_14_1739 ();
 FILLCELL_X4 FILLER_14_1755 ();
 FILLCELL_X2 FILLER_14_1759 ();
 FILLCELL_X1 FILLER_14_1761 ();
 FILLCELL_X8 FILLER_15_1 ();
 FILLCELL_X1 FILLER_15_9 ();
 FILLCELL_X4 FILLER_15_19 ();
 FILLCELL_X8 FILLER_15_27 ();
 FILLCELL_X1 FILLER_15_35 ();
 FILLCELL_X4 FILLER_15_39 ();
 FILLCELL_X2 FILLER_15_43 ();
 FILLCELL_X8 FILLER_15_48 ();
 FILLCELL_X8 FILLER_15_59 ();
 FILLCELL_X2 FILLER_15_67 ();
 FILLCELL_X8 FILLER_15_72 ();
 FILLCELL_X4 FILLER_15_89 ();
 FILLCELL_X4 FILLER_15_112 ();
 FILLCELL_X1 FILLER_15_116 ();
 FILLCELL_X4 FILLER_15_120 ();
 FILLCELL_X16 FILLER_15_127 ();
 FILLCELL_X4 FILLER_15_143 ();
 FILLCELL_X4 FILLER_15_154 ();
 FILLCELL_X4 FILLER_15_161 ();
 FILLCELL_X8 FILLER_15_167 ();
 FILLCELL_X2 FILLER_15_175 ();
 FILLCELL_X4 FILLER_15_187 ();
 FILLCELL_X4 FILLER_15_193 ();
 FILLCELL_X2 FILLER_15_197 ();
 FILLCELL_X1 FILLER_15_199 ();
 FILLCELL_X4 FILLER_15_203 ();
 FILLCELL_X4 FILLER_15_211 ();
 FILLCELL_X4 FILLER_15_224 ();
 FILLCELL_X4 FILLER_15_238 ();
 FILLCELL_X4 FILLER_15_245 ();
 FILLCELL_X2 FILLER_15_249 ();
 FILLCELL_X1 FILLER_15_251 ();
 FILLCELL_X4 FILLER_15_255 ();
 FILLCELL_X8 FILLER_15_262 ();
 FILLCELL_X4 FILLER_15_270 ();
 FILLCELL_X1 FILLER_15_274 ();
 FILLCELL_X4 FILLER_15_279 ();
 FILLCELL_X4 FILLER_15_292 ();
 FILLCELL_X4 FILLER_15_305 ();
 FILLCELL_X4 FILLER_15_318 ();
 FILLCELL_X4 FILLER_15_339 ();
 FILLCELL_X8 FILLER_15_352 ();
 FILLCELL_X1 FILLER_15_360 ();
 FILLCELL_X8 FILLER_15_371 ();
 FILLCELL_X1 FILLER_15_379 ();
 FILLCELL_X4 FILLER_15_382 ();
 FILLCELL_X1 FILLER_15_386 ();
 FILLCELL_X8 FILLER_15_394 ();
 FILLCELL_X4 FILLER_15_415 ();
 FILLCELL_X2 FILLER_15_419 ();
 FILLCELL_X1 FILLER_15_421 ();
 FILLCELL_X4 FILLER_15_425 ();
 FILLCELL_X4 FILLER_15_434 ();
 FILLCELL_X2 FILLER_15_438 ();
 FILLCELL_X1 FILLER_15_440 ();
 FILLCELL_X4 FILLER_15_444 ();
 FILLCELL_X16 FILLER_15_458 ();
 FILLCELL_X8 FILLER_15_474 ();
 FILLCELL_X8 FILLER_15_485 ();
 FILLCELL_X1 FILLER_15_493 ();
 FILLCELL_X4 FILLER_15_501 ();
 FILLCELL_X1 FILLER_15_505 ();
 FILLCELL_X16 FILLER_15_509 ();
 FILLCELL_X2 FILLER_15_525 ();
 FILLCELL_X4 FILLER_15_530 ();
 FILLCELL_X4 FILLER_15_537 ();
 FILLCELL_X4 FILLER_15_544 ();
 FILLCELL_X1 FILLER_15_548 ();
 FILLCELL_X8 FILLER_15_558 ();
 FILLCELL_X1 FILLER_15_566 ();
 FILLCELL_X4 FILLER_15_577 ();
 FILLCELL_X4 FILLER_15_584 ();
 FILLCELL_X4 FILLER_15_590 ();
 FILLCELL_X2 FILLER_15_594 ();
 FILLCELL_X4 FILLER_15_600 ();
 FILLCELL_X16 FILLER_15_607 ();
 FILLCELL_X4 FILLER_15_623 ();
 FILLCELL_X2 FILLER_15_627 ();
 FILLCELL_X1 FILLER_15_629 ();
 FILLCELL_X8 FILLER_15_632 ();
 FILLCELL_X1 FILLER_15_640 ();
 FILLCELL_X4 FILLER_15_647 ();
 FILLCELL_X4 FILLER_15_653 ();
 FILLCELL_X4 FILLER_15_660 ();
 FILLCELL_X8 FILLER_15_673 ();
 FILLCELL_X4 FILLER_15_681 ();
 FILLCELL_X2 FILLER_15_685 ();
 FILLCELL_X1 FILLER_15_687 ();
 FILLCELL_X4 FILLER_15_695 ();
 FILLCELL_X4 FILLER_15_702 ();
 FILLCELL_X2 FILLER_15_706 ();
 FILLCELL_X4 FILLER_15_714 ();
 FILLCELL_X8 FILLER_15_724 ();
 FILLCELL_X16 FILLER_15_735 ();
 FILLCELL_X4 FILLER_15_751 ();
 FILLCELL_X4 FILLER_15_759 ();
 FILLCELL_X8 FILLER_15_767 ();
 FILLCELL_X1 FILLER_15_775 ();
 FILLCELL_X4 FILLER_15_778 ();
 FILLCELL_X4 FILLER_15_791 ();
 FILLCELL_X16 FILLER_15_799 ();
 FILLCELL_X4 FILLER_15_815 ();
 FILLCELL_X2 FILLER_15_819 ();
 FILLCELL_X1 FILLER_15_821 ();
 FILLCELL_X8 FILLER_15_831 ();
 FILLCELL_X4 FILLER_15_839 ();
 FILLCELL_X4 FILLER_15_853 ();
 FILLCELL_X1 FILLER_15_857 ();
 FILLCELL_X8 FILLER_15_860 ();
 FILLCELL_X4 FILLER_15_872 ();
 FILLCELL_X4 FILLER_15_886 ();
 FILLCELL_X16 FILLER_15_893 ();
 FILLCELL_X1 FILLER_15_909 ();
 FILLCELL_X8 FILLER_15_916 ();
 FILLCELL_X4 FILLER_15_931 ();
 FILLCELL_X4 FILLER_15_941 ();
 FILLCELL_X4 FILLER_15_951 ();
 FILLCELL_X4 FILLER_15_959 ();
 FILLCELL_X4 FILLER_15_966 ();
 FILLCELL_X4 FILLER_15_974 ();
 FILLCELL_X4 FILLER_15_981 ();
 FILLCELL_X4 FILLER_15_988 ();
 FILLCELL_X4 FILLER_15_995 ();
 FILLCELL_X4 FILLER_15_1002 ();
 FILLCELL_X1 FILLER_15_1006 ();
 FILLCELL_X4 FILLER_15_1014 ();
 FILLCELL_X2 FILLER_15_1018 ();
 FILLCELL_X1 FILLER_15_1020 ();
 FILLCELL_X4 FILLER_15_1023 ();
 FILLCELL_X4 FILLER_15_1033 ();
 FILLCELL_X2 FILLER_15_1037 ();
 FILLCELL_X1 FILLER_15_1039 ();
 FILLCELL_X8 FILLER_15_1046 ();
 FILLCELL_X8 FILLER_15_1057 ();
 FILLCELL_X4 FILLER_15_1068 ();
 FILLCELL_X4 FILLER_15_1081 ();
 FILLCELL_X8 FILLER_15_1088 ();
 FILLCELL_X2 FILLER_15_1096 ();
 FILLCELL_X1 FILLER_15_1098 ();
 FILLCELL_X4 FILLER_15_1109 ();
 FILLCELL_X16 FILLER_15_1117 ();
 FILLCELL_X2 FILLER_15_1133 ();
 FILLCELL_X1 FILLER_15_1135 ();
 FILLCELL_X8 FILLER_15_1138 ();
 FILLCELL_X4 FILLER_15_1148 ();
 FILLCELL_X1 FILLER_15_1152 ();
 FILLCELL_X4 FILLER_15_1156 ();
 FILLCELL_X2 FILLER_15_1160 ();
 FILLCELL_X1 FILLER_15_1162 ();
 FILLCELL_X4 FILLER_15_1172 ();
 FILLCELL_X2 FILLER_15_1176 ();
 FILLCELL_X1 FILLER_15_1178 ();
 FILLCELL_X4 FILLER_15_1183 ();
 FILLCELL_X8 FILLER_15_1190 ();
 FILLCELL_X8 FILLER_15_1207 ();
 FILLCELL_X2 FILLER_15_1215 ();
 FILLCELL_X4 FILLER_15_1221 ();
 FILLCELL_X4 FILLER_15_1229 ();
 FILLCELL_X4 FILLER_15_1236 ();
 FILLCELL_X4 FILLER_15_1242 ();
 FILLCELL_X8 FILLER_15_1253 ();
 FILLCELL_X2 FILLER_15_1261 ();
 FILLCELL_X4 FILLER_15_1264 ();
 FILLCELL_X4 FILLER_15_1277 ();
 FILLCELL_X8 FILLER_15_1288 ();
 FILLCELL_X4 FILLER_15_1296 ();
 FILLCELL_X1 FILLER_15_1300 ();
 FILLCELL_X4 FILLER_15_1305 ();
 FILLCELL_X8 FILLER_15_1316 ();
 FILLCELL_X1 FILLER_15_1324 ();
 FILLCELL_X4 FILLER_15_1328 ();
 FILLCELL_X2 FILLER_15_1332 ();
 FILLCELL_X1 FILLER_15_1334 ();
 FILLCELL_X4 FILLER_15_1339 ();
 FILLCELL_X4 FILLER_15_1347 ();
 FILLCELL_X8 FILLER_15_1354 ();
 FILLCELL_X4 FILLER_15_1362 ();
 FILLCELL_X1 FILLER_15_1366 ();
 FILLCELL_X4 FILLER_15_1376 ();
 FILLCELL_X4 FILLER_15_1384 ();
 FILLCELL_X4 FILLER_15_1391 ();
 FILLCELL_X2 FILLER_15_1395 ();
 FILLCELL_X1 FILLER_15_1397 ();
 FILLCELL_X4 FILLER_15_1402 ();
 FILLCELL_X8 FILLER_15_1415 ();
 FILLCELL_X2 FILLER_15_1423 ();
 FILLCELL_X4 FILLER_15_1429 ();
 FILLCELL_X4 FILLER_15_1442 ();
 FILLCELL_X8 FILLER_15_1448 ();
 FILLCELL_X4 FILLER_15_1456 ();
 FILLCELL_X32 FILLER_15_1469 ();
 FILLCELL_X32 FILLER_15_1501 ();
 FILLCELL_X32 FILLER_15_1533 ();
 FILLCELL_X32 FILLER_15_1565 ();
 FILLCELL_X32 FILLER_15_1597 ();
 FILLCELL_X32 FILLER_15_1629 ();
 FILLCELL_X32 FILLER_15_1661 ();
 FILLCELL_X32 FILLER_15_1693 ();
 FILLCELL_X32 FILLER_15_1725 ();
 FILLCELL_X4 FILLER_15_1757 ();
 FILLCELL_X1 FILLER_15_1761 ();
 FILLCELL_X8 FILLER_16_1 ();
 FILLCELL_X2 FILLER_16_9 ();
 FILLCELL_X4 FILLER_16_14 ();
 FILLCELL_X8 FILLER_16_21 ();
 FILLCELL_X4 FILLER_16_29 ();
 FILLCELL_X1 FILLER_16_33 ();
 FILLCELL_X4 FILLER_16_43 ();
 FILLCELL_X1 FILLER_16_47 ();
 FILLCELL_X8 FILLER_16_52 ();
 FILLCELL_X4 FILLER_16_60 ();
 FILLCELL_X2 FILLER_16_64 ();
 FILLCELL_X4 FILLER_16_76 ();
 FILLCELL_X4 FILLER_16_83 ();
 FILLCELL_X16 FILLER_16_89 ();
 FILLCELL_X8 FILLER_16_105 ();
 FILLCELL_X1 FILLER_16_113 ();
 FILLCELL_X4 FILLER_16_117 ();
 FILLCELL_X4 FILLER_16_123 ();
 FILLCELL_X2 FILLER_16_127 ();
 FILLCELL_X8 FILLER_16_132 ();
 FILLCELL_X4 FILLER_16_149 ();
 FILLCELL_X8 FILLER_16_163 ();
 FILLCELL_X4 FILLER_16_178 ();
 FILLCELL_X4 FILLER_16_192 ();
 FILLCELL_X4 FILLER_16_200 ();
 FILLCELL_X2 FILLER_16_204 ();
 FILLCELL_X4 FILLER_16_210 ();
 FILLCELL_X8 FILLER_16_217 ();
 FILLCELL_X4 FILLER_16_225 ();
 FILLCELL_X16 FILLER_16_233 ();
 FILLCELL_X8 FILLER_16_249 ();
 FILLCELL_X4 FILLER_16_257 ();
 FILLCELL_X4 FILLER_16_264 ();
 FILLCELL_X1 FILLER_16_268 ();
 FILLCELL_X8 FILLER_16_272 ();
 FILLCELL_X2 FILLER_16_280 ();
 FILLCELL_X4 FILLER_16_285 ();
 FILLCELL_X8 FILLER_16_293 ();
 FILLCELL_X2 FILLER_16_301 ();
 FILLCELL_X4 FILLER_16_308 ();
 FILLCELL_X4 FILLER_16_319 ();
 FILLCELL_X8 FILLER_16_330 ();
 FILLCELL_X2 FILLER_16_338 ();
 FILLCELL_X4 FILLER_16_349 ();
 FILLCELL_X4 FILLER_16_356 ();
 FILLCELL_X4 FILLER_16_369 ();
 FILLCELL_X8 FILLER_16_376 ();
 FILLCELL_X4 FILLER_16_394 ();
 FILLCELL_X4 FILLER_16_400 ();
 FILLCELL_X4 FILLER_16_407 ();
 FILLCELL_X4 FILLER_16_420 ();
 FILLCELL_X4 FILLER_16_433 ();
 FILLCELL_X4 FILLER_16_444 ();
 FILLCELL_X2 FILLER_16_448 ();
 FILLCELL_X4 FILLER_16_454 ();
 FILLCELL_X8 FILLER_16_461 ();
 FILLCELL_X2 FILLER_16_469 ();
 FILLCELL_X1 FILLER_16_471 ();
 FILLCELL_X4 FILLER_16_476 ();
 FILLCELL_X4 FILLER_16_490 ();
 FILLCELL_X4 FILLER_16_496 ();
 FILLCELL_X4 FILLER_16_510 ();
 FILLCELL_X8 FILLER_16_517 ();
 FILLCELL_X4 FILLER_16_525 ();
 FILLCELL_X1 FILLER_16_529 ();
 FILLCELL_X4 FILLER_16_540 ();
 FILLCELL_X8 FILLER_16_553 ();
 FILLCELL_X1 FILLER_16_561 ();
 FILLCELL_X8 FILLER_16_566 ();
 FILLCELL_X2 FILLER_16_574 ();
 FILLCELL_X4 FILLER_16_583 ();
 FILLCELL_X8 FILLER_16_589 ();
 FILLCELL_X2 FILLER_16_597 ();
 FILLCELL_X4 FILLER_16_602 ();
 FILLCELL_X4 FILLER_16_615 ();
 FILLCELL_X8 FILLER_16_622 ();
 FILLCELL_X1 FILLER_16_630 ();
 FILLCELL_X4 FILLER_16_632 ();
 FILLCELL_X8 FILLER_16_645 ();
 FILLCELL_X1 FILLER_16_653 ();
 FILLCELL_X4 FILLER_16_658 ();
 FILLCELL_X4 FILLER_16_672 ();
 FILLCELL_X4 FILLER_16_678 ();
 FILLCELL_X2 FILLER_16_682 ();
 FILLCELL_X4 FILLER_16_690 ();
 FILLCELL_X4 FILLER_16_700 ();
 FILLCELL_X8 FILLER_16_711 ();
 FILLCELL_X1 FILLER_16_719 ();
 FILLCELL_X4 FILLER_16_727 ();
 FILLCELL_X1 FILLER_16_731 ();
 FILLCELL_X4 FILLER_16_742 ();
 FILLCELL_X1 FILLER_16_746 ();
 FILLCELL_X4 FILLER_16_750 ();
 FILLCELL_X4 FILLER_16_758 ();
 FILLCELL_X2 FILLER_16_762 ();
 FILLCELL_X1 FILLER_16_764 ();
 FILLCELL_X4 FILLER_16_768 ();
 FILLCELL_X2 FILLER_16_772 ();
 FILLCELL_X1 FILLER_16_774 ();
 FILLCELL_X8 FILLER_16_779 ();
 FILLCELL_X2 FILLER_16_787 ();
 FILLCELL_X4 FILLER_16_792 ();
 FILLCELL_X8 FILLER_16_805 ();
 FILLCELL_X1 FILLER_16_813 ();
 FILLCELL_X16 FILLER_16_833 ();
 FILLCELL_X2 FILLER_16_849 ();
 FILLCELL_X8 FILLER_16_855 ();
 FILLCELL_X2 FILLER_16_863 ();
 FILLCELL_X4 FILLER_16_868 ();
 FILLCELL_X2 FILLER_16_872 ();
 FILLCELL_X1 FILLER_16_874 ();
 FILLCELL_X4 FILLER_16_879 ();
 FILLCELL_X4 FILLER_16_892 ();
 FILLCELL_X1 FILLER_16_896 ();
 FILLCELL_X4 FILLER_16_901 ();
 FILLCELL_X32 FILLER_16_909 ();
 FILLCELL_X8 FILLER_16_941 ();
 FILLCELL_X1 FILLER_16_949 ();
 FILLCELL_X4 FILLER_16_954 ();
 FILLCELL_X1 FILLER_16_958 ();
 FILLCELL_X4 FILLER_16_961 ();
 FILLCELL_X4 FILLER_16_969 ();
 FILLCELL_X4 FILLER_16_982 ();
 FILLCELL_X2 FILLER_16_986 ();
 FILLCELL_X1 FILLER_16_988 ();
 FILLCELL_X4 FILLER_16_998 ();
 FILLCELL_X4 FILLER_16_1006 ();
 FILLCELL_X16 FILLER_16_1014 ();
 FILLCELL_X4 FILLER_16_1030 ();
 FILLCELL_X4 FILLER_16_1040 ();
 FILLCELL_X4 FILLER_16_1051 ();
 FILLCELL_X8 FILLER_16_1059 ();
 FILLCELL_X2 FILLER_16_1067 ();
 FILLCELL_X8 FILLER_16_1073 ();
 FILLCELL_X4 FILLER_16_1081 ();
 FILLCELL_X2 FILLER_16_1085 ();
 FILLCELL_X8 FILLER_16_1090 ();
 FILLCELL_X2 FILLER_16_1098 ();
 FILLCELL_X8 FILLER_16_1103 ();
 FILLCELL_X4 FILLER_16_1111 ();
 FILLCELL_X4 FILLER_16_1119 ();
 FILLCELL_X8 FILLER_16_1126 ();
 FILLCELL_X4 FILLER_16_1134 ();
 FILLCELL_X4 FILLER_16_1148 ();
 FILLCELL_X8 FILLER_16_1162 ();
 FILLCELL_X2 FILLER_16_1170 ();
 FILLCELL_X4 FILLER_16_1176 ();
 FILLCELL_X4 FILLER_16_1189 ();
 FILLCELL_X4 FILLER_16_1196 ();
 FILLCELL_X8 FILLER_16_1203 ();
 FILLCELL_X4 FILLER_16_1217 ();
 FILLCELL_X8 FILLER_16_1227 ();
 FILLCELL_X1 FILLER_16_1235 ();
 FILLCELL_X4 FILLER_16_1246 ();
 FILLCELL_X4 FILLER_16_1260 ();
 FILLCELL_X4 FILLER_16_1266 ();
 FILLCELL_X1 FILLER_16_1270 ();
 FILLCELL_X4 FILLER_16_1273 ();
 FILLCELL_X4 FILLER_16_1287 ();
 FILLCELL_X4 FILLER_16_1294 ();
 FILLCELL_X2 FILLER_16_1298 ();
 FILLCELL_X1 FILLER_16_1300 ();
 FILLCELL_X4 FILLER_16_1303 ();
 FILLCELL_X4 FILLER_16_1317 ();
 FILLCELL_X8 FILLER_16_1331 ();
 FILLCELL_X2 FILLER_16_1339 ();
 FILLCELL_X4 FILLER_16_1350 ();
 FILLCELL_X4 FILLER_16_1358 ();
 FILLCELL_X4 FILLER_16_1365 ();
 FILLCELL_X4 FILLER_16_1378 ();
 FILLCELL_X4 FILLER_16_1385 ();
 FILLCELL_X8 FILLER_16_1392 ();
 FILLCELL_X4 FILLER_16_1400 ();
 FILLCELL_X8 FILLER_16_1408 ();
 FILLCELL_X1 FILLER_16_1416 ();
 FILLCELL_X4 FILLER_16_1420 ();
 FILLCELL_X1 FILLER_16_1424 ();
 FILLCELL_X4 FILLER_16_1434 ();
 FILLCELL_X8 FILLER_16_1441 ();
 FILLCELL_X1 FILLER_16_1449 ();
 FILLCELL_X4 FILLER_16_1460 ();
 FILLCELL_X4 FILLER_16_1467 ();
 FILLCELL_X32 FILLER_16_1474 ();
 FILLCELL_X32 FILLER_16_1506 ();
 FILLCELL_X32 FILLER_16_1538 ();
 FILLCELL_X32 FILLER_16_1570 ();
 FILLCELL_X32 FILLER_16_1602 ();
 FILLCELL_X32 FILLER_16_1634 ();
 FILLCELL_X32 FILLER_16_1666 ();
 FILLCELL_X32 FILLER_16_1698 ();
 FILLCELL_X32 FILLER_16_1730 ();
 FILLCELL_X4 FILLER_17_1 ();
 FILLCELL_X16 FILLER_17_9 ();
 FILLCELL_X1 FILLER_17_25 ();
 FILLCELL_X4 FILLER_17_29 ();
 FILLCELL_X4 FILLER_17_37 ();
 FILLCELL_X4 FILLER_17_50 ();
 FILLCELL_X8 FILLER_17_58 ();
 FILLCELL_X1 FILLER_17_66 ();
 FILLCELL_X8 FILLER_17_76 ();
 FILLCELL_X8 FILLER_17_94 ();
 FILLCELL_X2 FILLER_17_102 ();
 FILLCELL_X4 FILLER_17_108 ();
 FILLCELL_X8 FILLER_17_117 ();
 FILLCELL_X8 FILLER_17_128 ();
 FILLCELL_X2 FILLER_17_136 ();
 FILLCELL_X8 FILLER_17_141 ();
 FILLCELL_X4 FILLER_17_149 ();
 FILLCELL_X2 FILLER_17_153 ();
 FILLCELL_X8 FILLER_17_158 ();
 FILLCELL_X4 FILLER_17_170 ();
 FILLCELL_X4 FILLER_17_177 ();
 FILLCELL_X2 FILLER_17_181 ();
 FILLCELL_X8 FILLER_17_186 ();
 FILLCELL_X4 FILLER_17_194 ();
 FILLCELL_X2 FILLER_17_198 ();
 FILLCELL_X4 FILLER_17_204 ();
 FILLCELL_X8 FILLER_17_217 ();
 FILLCELL_X4 FILLER_17_229 ();
 FILLCELL_X4 FILLER_17_240 ();
 FILLCELL_X4 FILLER_17_247 ();
 FILLCELL_X1 FILLER_17_251 ();
 FILLCELL_X4 FILLER_17_261 ();
 FILLCELL_X4 FILLER_17_269 ();
 FILLCELL_X2 FILLER_17_273 ();
 FILLCELL_X1 FILLER_17_275 ();
 FILLCELL_X4 FILLER_17_279 ();
 FILLCELL_X4 FILLER_17_293 ();
 FILLCELL_X8 FILLER_17_301 ();
 FILLCELL_X1 FILLER_17_309 ();
 FILLCELL_X4 FILLER_17_313 ();
 FILLCELL_X4 FILLER_17_336 ();
 FILLCELL_X4 FILLER_17_343 ();
 FILLCELL_X8 FILLER_17_357 ();
 FILLCELL_X2 FILLER_17_365 ();
 FILLCELL_X4 FILLER_17_369 ();
 FILLCELL_X16 FILLER_17_383 ();
 FILLCELL_X8 FILLER_17_399 ();
 FILLCELL_X2 FILLER_17_407 ();
 FILLCELL_X1 FILLER_17_409 ();
 FILLCELL_X4 FILLER_17_412 ();
 FILLCELL_X4 FILLER_17_420 ();
 FILLCELL_X1 FILLER_17_424 ();
 FILLCELL_X4 FILLER_17_429 ();
 FILLCELL_X8 FILLER_17_436 ();
 FILLCELL_X2 FILLER_17_444 ();
 FILLCELL_X4 FILLER_17_450 ();
 FILLCELL_X4 FILLER_17_458 ();
 FILLCELL_X4 FILLER_17_466 ();
 FILLCELL_X4 FILLER_17_474 ();
 FILLCELL_X8 FILLER_17_487 ();
 FILLCELL_X2 FILLER_17_495 ();
 FILLCELL_X1 FILLER_17_497 ();
 FILLCELL_X4 FILLER_17_501 ();
 FILLCELL_X4 FILLER_17_512 ();
 FILLCELL_X16 FILLER_17_525 ();
 FILLCELL_X4 FILLER_17_541 ();
 FILLCELL_X2 FILLER_17_545 ();
 FILLCELL_X1 FILLER_17_547 ();
 FILLCELL_X8 FILLER_17_552 ();
 FILLCELL_X4 FILLER_17_560 ();
 FILLCELL_X4 FILLER_17_567 ();
 FILLCELL_X4 FILLER_17_581 ();
 FILLCELL_X8 FILLER_17_595 ();
 FILLCELL_X2 FILLER_17_603 ();
 FILLCELL_X8 FILLER_17_624 ();
 FILLCELL_X4 FILLER_17_639 ();
 FILLCELL_X4 FILLER_17_653 ();
 FILLCELL_X2 FILLER_17_657 ();
 FILLCELL_X1 FILLER_17_659 ();
 FILLCELL_X4 FILLER_17_670 ();
 FILLCELL_X1 FILLER_17_674 ();
 FILLCELL_X4 FILLER_17_694 ();
 FILLCELL_X4 FILLER_17_702 ();
 FILLCELL_X4 FILLER_17_710 ();
 FILLCELL_X8 FILLER_17_720 ();
 FILLCELL_X4 FILLER_17_731 ();
 FILLCELL_X4 FILLER_17_739 ();
 FILLCELL_X2 FILLER_17_743 ();
 FILLCELL_X1 FILLER_17_745 ();
 FILLCELL_X4 FILLER_17_755 ();
 FILLCELL_X4 FILLER_17_768 ();
 FILLCELL_X4 FILLER_17_775 ();
 FILLCELL_X4 FILLER_17_782 ();
 FILLCELL_X8 FILLER_17_789 ();
 FILLCELL_X4 FILLER_17_797 ();
 FILLCELL_X8 FILLER_17_810 ();
 FILLCELL_X8 FILLER_17_828 ();
 FILLCELL_X4 FILLER_17_839 ();
 FILLCELL_X2 FILLER_17_843 ();
 FILLCELL_X1 FILLER_17_845 ();
 FILLCELL_X4 FILLER_17_863 ();
 FILLCELL_X2 FILLER_17_867 ();
 FILLCELL_X1 FILLER_17_869 ();
 FILLCELL_X4 FILLER_17_874 ();
 FILLCELL_X4 FILLER_17_881 ();
 FILLCELL_X2 FILLER_17_885 ();
 FILLCELL_X4 FILLER_17_906 ();
 FILLCELL_X4 FILLER_17_929 ();
 FILLCELL_X32 FILLER_17_937 ();
 FILLCELL_X2 FILLER_17_969 ();
 FILLCELL_X8 FILLER_17_990 ();
 FILLCELL_X4 FILLER_17_998 ();
 FILLCELL_X16 FILLER_17_1021 ();
 FILLCELL_X8 FILLER_17_1037 ();
 FILLCELL_X16 FILLER_17_1049 ();
 FILLCELL_X4 FILLER_17_1069 ();
 FILLCELL_X4 FILLER_17_1082 ();
 FILLCELL_X4 FILLER_17_1089 ();
 FILLCELL_X16 FILLER_17_1096 ();
 FILLCELL_X4 FILLER_17_1116 ();
 FILLCELL_X4 FILLER_17_1129 ();
 FILLCELL_X4 FILLER_17_1136 ();
 FILLCELL_X16 FILLER_17_1143 ();
 FILLCELL_X2 FILLER_17_1159 ();
 FILLCELL_X4 FILLER_17_1164 ();
 FILLCELL_X2 FILLER_17_1168 ();
 FILLCELL_X4 FILLER_17_1174 ();
 FILLCELL_X8 FILLER_17_1187 ();
 FILLCELL_X4 FILLER_17_1198 ();
 FILLCELL_X4 FILLER_17_1209 ();
 FILLCELL_X4 FILLER_17_1219 ();
 FILLCELL_X4 FILLER_17_1229 ();
 FILLCELL_X4 FILLER_17_1235 ();
 FILLCELL_X1 FILLER_17_1239 ();
 FILLCELL_X4 FILLER_17_1243 ();
 FILLCELL_X4 FILLER_17_1256 ();
 FILLCELL_X2 FILLER_17_1260 ();
 FILLCELL_X1 FILLER_17_1262 ();
 FILLCELL_X16 FILLER_17_1264 ();
 FILLCELL_X1 FILLER_17_1280 ();
 FILLCELL_X4 FILLER_17_1290 ();
 FILLCELL_X8 FILLER_17_1303 ();
 FILLCELL_X1 FILLER_17_1311 ();
 FILLCELL_X4 FILLER_17_1315 ();
 FILLCELL_X16 FILLER_17_1322 ();
 FILLCELL_X2 FILLER_17_1338 ();
 FILLCELL_X4 FILLER_17_1343 ();
 FILLCELL_X8 FILLER_17_1356 ();
 FILLCELL_X4 FILLER_17_1368 ();
 FILLCELL_X8 FILLER_17_1376 ();
 FILLCELL_X1 FILLER_17_1384 ();
 FILLCELL_X4 FILLER_17_1389 ();
 FILLCELL_X4 FILLER_17_1398 ();
 FILLCELL_X8 FILLER_17_1406 ();
 FILLCELL_X2 FILLER_17_1414 ();
 FILLCELL_X4 FILLER_17_1420 ();
 FILLCELL_X4 FILLER_17_1428 ();
 FILLCELL_X8 FILLER_17_1435 ();
 FILLCELL_X1 FILLER_17_1443 ();
 FILLCELL_X4 FILLER_17_1451 ();
 FILLCELL_X4 FILLER_17_1465 ();
 FILLCELL_X4 FILLER_17_1471 ();
 FILLCELL_X32 FILLER_17_1485 ();
 FILLCELL_X32 FILLER_17_1517 ();
 FILLCELL_X32 FILLER_17_1549 ();
 FILLCELL_X32 FILLER_17_1581 ();
 FILLCELL_X32 FILLER_17_1613 ();
 FILLCELL_X32 FILLER_17_1645 ();
 FILLCELL_X32 FILLER_17_1677 ();
 FILLCELL_X32 FILLER_17_1709 ();
 FILLCELL_X16 FILLER_17_1741 ();
 FILLCELL_X4 FILLER_17_1757 ();
 FILLCELL_X1 FILLER_17_1761 ();
 FILLCELL_X8 FILLER_18_1 ();
 FILLCELL_X4 FILLER_18_28 ();
 FILLCELL_X1 FILLER_18_32 ();
 FILLCELL_X4 FILLER_18_36 ();
 FILLCELL_X2 FILLER_18_40 ();
 FILLCELL_X16 FILLER_18_45 ();
 FILLCELL_X1 FILLER_18_61 ();
 FILLCELL_X8 FILLER_18_72 ();
 FILLCELL_X1 FILLER_18_80 ();
 FILLCELL_X4 FILLER_18_84 ();
 FILLCELL_X4 FILLER_18_91 ();
 FILLCELL_X2 FILLER_18_95 ();
 FILLCELL_X4 FILLER_18_101 ();
 FILLCELL_X4 FILLER_18_110 ();
 FILLCELL_X4 FILLER_18_123 ();
 FILLCELL_X2 FILLER_18_127 ();
 FILLCELL_X1 FILLER_18_129 ();
 FILLCELL_X4 FILLER_18_139 ();
 FILLCELL_X8 FILLER_18_149 ();
 FILLCELL_X4 FILLER_18_161 ();
 FILLCELL_X4 FILLER_18_174 ();
 FILLCELL_X16 FILLER_18_187 ();
 FILLCELL_X4 FILLER_18_203 ();
 FILLCELL_X16 FILLER_18_210 ();
 FILLCELL_X4 FILLER_18_226 ();
 FILLCELL_X2 FILLER_18_230 ();
 FILLCELL_X8 FILLER_18_242 ();
 FILLCELL_X4 FILLER_18_259 ();
 FILLCELL_X4 FILLER_18_272 ();
 FILLCELL_X8 FILLER_18_283 ();
 FILLCELL_X4 FILLER_18_291 ();
 FILLCELL_X2 FILLER_18_295 ();
 FILLCELL_X1 FILLER_18_297 ();
 FILLCELL_X4 FILLER_18_301 ();
 FILLCELL_X8 FILLER_18_309 ();
 FILLCELL_X1 FILLER_18_317 ();
 FILLCELL_X4 FILLER_18_324 ();
 FILLCELL_X4 FILLER_18_332 ();
 FILLCELL_X16 FILLER_18_339 ();
 FILLCELL_X8 FILLER_18_355 ();
 FILLCELL_X2 FILLER_18_363 ();
 FILLCELL_X8 FILLER_18_368 ();
 FILLCELL_X1 FILLER_18_376 ();
 FILLCELL_X8 FILLER_18_381 ();
 FILLCELL_X1 FILLER_18_389 ();
 FILLCELL_X8 FILLER_18_394 ();
 FILLCELL_X2 FILLER_18_402 ();
 FILLCELL_X4 FILLER_18_408 ();
 FILLCELL_X8 FILLER_18_419 ();
 FILLCELL_X4 FILLER_18_427 ();
 FILLCELL_X2 FILLER_18_431 ();
 FILLCELL_X1 FILLER_18_433 ();
 FILLCELL_X4 FILLER_18_437 ();
 FILLCELL_X4 FILLER_18_445 ();
 FILLCELL_X4 FILLER_18_458 ();
 FILLCELL_X8 FILLER_18_471 ();
 FILLCELL_X1 FILLER_18_479 ();
 FILLCELL_X4 FILLER_18_483 ();
 FILLCELL_X2 FILLER_18_487 ();
 FILLCELL_X1 FILLER_18_489 ();
 FILLCELL_X4 FILLER_18_493 ();
 FILLCELL_X4 FILLER_18_500 ();
 FILLCELL_X8 FILLER_18_513 ();
 FILLCELL_X8 FILLER_18_530 ();
 FILLCELL_X4 FILLER_18_538 ();
 FILLCELL_X2 FILLER_18_542 ();
 FILLCELL_X4 FILLER_18_547 ();
 FILLCELL_X4 FILLER_18_560 ();
 FILLCELL_X4 FILLER_18_574 ();
 FILLCELL_X2 FILLER_18_578 ();
 FILLCELL_X4 FILLER_18_590 ();
 FILLCELL_X1 FILLER_18_594 ();
 FILLCELL_X8 FILLER_18_598 ();
 FILLCELL_X4 FILLER_18_606 ();
 FILLCELL_X1 FILLER_18_610 ();
 FILLCELL_X4 FILLER_18_614 ();
 FILLCELL_X4 FILLER_18_627 ();
 FILLCELL_X4 FILLER_18_632 ();
 FILLCELL_X8 FILLER_18_646 ();
 FILLCELL_X1 FILLER_18_654 ();
 FILLCELL_X16 FILLER_18_658 ();
 FILLCELL_X8 FILLER_18_674 ();
 FILLCELL_X2 FILLER_18_682 ();
 FILLCELL_X16 FILLER_18_688 ();
 FILLCELL_X8 FILLER_18_704 ();
 FILLCELL_X4 FILLER_18_712 ();
 FILLCELL_X1 FILLER_18_716 ();
 FILLCELL_X4 FILLER_18_720 ();
 FILLCELL_X1 FILLER_18_724 ();
 FILLCELL_X4 FILLER_18_727 ();
 FILLCELL_X4 FILLER_18_735 ();
 FILLCELL_X16 FILLER_18_749 ();
 FILLCELL_X4 FILLER_18_768 ();
 FILLCELL_X2 FILLER_18_772 ();
 FILLCELL_X1 FILLER_18_774 ();
 FILLCELL_X8 FILLER_18_785 ();
 FILLCELL_X1 FILLER_18_793 ();
 FILLCELL_X4 FILLER_18_798 ();
 FILLCELL_X4 FILLER_18_806 ();
 FILLCELL_X4 FILLER_18_814 ();
 FILLCELL_X4 FILLER_18_820 ();
 FILLCELL_X4 FILLER_18_831 ();
 FILLCELL_X8 FILLER_18_845 ();
 FILLCELL_X4 FILLER_18_853 ();
 FILLCELL_X1 FILLER_18_857 ();
 FILLCELL_X4 FILLER_18_861 ();
 FILLCELL_X4 FILLER_18_869 ();
 FILLCELL_X4 FILLER_18_882 ();
 FILLCELL_X2 FILLER_18_886 ();
 FILLCELL_X4 FILLER_18_892 ();
 FILLCELL_X16 FILLER_18_900 ();
 FILLCELL_X8 FILLER_18_916 ();
 FILLCELL_X4 FILLER_18_924 ();
 FILLCELL_X2 FILLER_18_928 ();
 FILLCELL_X16 FILLER_18_949 ();
 FILLCELL_X1 FILLER_18_965 ();
 FILLCELL_X32 FILLER_18_970 ();
 FILLCELL_X8 FILLER_18_1002 ();
 FILLCELL_X4 FILLER_18_1012 ();
 FILLCELL_X4 FILLER_18_1035 ();
 FILLCELL_X2 FILLER_18_1039 ();
 FILLCELL_X4 FILLER_18_1044 ();
 FILLCELL_X1 FILLER_18_1048 ();
 FILLCELL_X4 FILLER_18_1053 ();
 FILLCELL_X16 FILLER_18_1060 ();
 FILLCELL_X4 FILLER_18_1080 ();
 FILLCELL_X4 FILLER_18_1093 ();
 FILLCELL_X4 FILLER_18_1100 ();
 FILLCELL_X8 FILLER_18_1106 ();
 FILLCELL_X4 FILLER_18_1114 ();
 FILLCELL_X1 FILLER_18_1118 ();
 FILLCELL_X4 FILLER_18_1123 ();
 FILLCELL_X16 FILLER_18_1136 ();
 FILLCELL_X4 FILLER_18_1152 ();
 FILLCELL_X4 FILLER_18_1159 ();
 FILLCELL_X1 FILLER_18_1163 ();
 FILLCELL_X8 FILLER_18_1167 ();
 FILLCELL_X2 FILLER_18_1175 ();
 FILLCELL_X32 FILLER_18_1180 ();
 FILLCELL_X4 FILLER_18_1212 ();
 FILLCELL_X4 FILLER_18_1220 ();
 FILLCELL_X16 FILLER_18_1230 ();
 FILLCELL_X1 FILLER_18_1246 ();
 FILLCELL_X4 FILLER_18_1250 ();
 FILLCELL_X4 FILLER_18_1257 ();
 FILLCELL_X4 FILLER_18_1264 ();
 FILLCELL_X8 FILLER_18_1271 ();
 FILLCELL_X4 FILLER_18_1279 ();
 FILLCELL_X2 FILLER_18_1283 ();
 FILLCELL_X4 FILLER_18_1288 ();
 FILLCELL_X8 FILLER_18_1295 ();
 FILLCELL_X4 FILLER_18_1303 ();
 FILLCELL_X4 FILLER_18_1311 ();
 FILLCELL_X4 FILLER_18_1324 ();
 FILLCELL_X4 FILLER_18_1333 ();
 FILLCELL_X8 FILLER_18_1340 ();
 FILLCELL_X1 FILLER_18_1348 ();
 FILLCELL_X16 FILLER_18_1353 ();
 FILLCELL_X8 FILLER_18_1369 ();
 FILLCELL_X2 FILLER_18_1377 ();
 FILLCELL_X1 FILLER_18_1379 ();
 FILLCELL_X4 FILLER_18_1384 ();
 FILLCELL_X4 FILLER_18_1395 ();
 FILLCELL_X4 FILLER_18_1416 ();
 FILLCELL_X2 FILLER_18_1420 ();
 FILLCELL_X1 FILLER_18_1422 ();
 FILLCELL_X4 FILLER_18_1427 ();
 FILLCELL_X1 FILLER_18_1431 ();
 FILLCELL_X4 FILLER_18_1435 ();
 FILLCELL_X4 FILLER_18_1449 ();
 FILLCELL_X4 FILLER_18_1456 ();
 FILLCELL_X4 FILLER_18_1462 ();
 FILLCELL_X1 FILLER_18_1466 ();
 FILLCELL_X4 FILLER_18_1470 ();
 FILLCELL_X4 FILLER_18_1484 ();
 FILLCELL_X32 FILLER_18_1492 ();
 FILLCELL_X32 FILLER_18_1524 ();
 FILLCELL_X32 FILLER_18_1556 ();
 FILLCELL_X32 FILLER_18_1588 ();
 FILLCELL_X32 FILLER_18_1620 ();
 FILLCELL_X32 FILLER_18_1652 ();
 FILLCELL_X32 FILLER_18_1684 ();
 FILLCELL_X32 FILLER_18_1716 ();
 FILLCELL_X8 FILLER_18_1748 ();
 FILLCELL_X4 FILLER_18_1756 ();
 FILLCELL_X2 FILLER_18_1760 ();
 FILLCELL_X4 FILLER_19_1 ();
 FILLCELL_X8 FILLER_19_24 ();
 FILLCELL_X4 FILLER_19_41 ();
 FILLCELL_X8 FILLER_19_47 ();
 FILLCELL_X4 FILLER_19_55 ();
 FILLCELL_X2 FILLER_19_59 ();
 FILLCELL_X4 FILLER_19_63 ();
 FILLCELL_X8 FILLER_19_74 ();
 FILLCELL_X2 FILLER_19_82 ();
 FILLCELL_X4 FILLER_19_91 ();
 FILLCELL_X4 FILLER_19_99 ();
 FILLCELL_X4 FILLER_19_105 ();
 FILLCELL_X1 FILLER_19_109 ();
 FILLCELL_X4 FILLER_19_114 ();
 FILLCELL_X8 FILLER_19_122 ();
 FILLCELL_X4 FILLER_19_130 ();
 FILLCELL_X2 FILLER_19_134 ();
 FILLCELL_X1 FILLER_19_136 ();
 FILLCELL_X4 FILLER_19_144 ();
 FILLCELL_X4 FILLER_19_154 ();
 FILLCELL_X8 FILLER_19_161 ();
 FILLCELL_X4 FILLER_19_172 ();
 FILLCELL_X2 FILLER_19_176 ();
 FILLCELL_X4 FILLER_19_182 ();
 FILLCELL_X4 FILLER_19_189 ();
 FILLCELL_X8 FILLER_19_210 ();
 FILLCELL_X1 FILLER_19_218 ();
 FILLCELL_X4 FILLER_19_221 ();
 FILLCELL_X4 FILLER_19_235 ();
 FILLCELL_X4 FILLER_19_241 ();
 FILLCELL_X2 FILLER_19_245 ();
 FILLCELL_X4 FILLER_19_257 ();
 FILLCELL_X4 FILLER_19_264 ();
 FILLCELL_X4 FILLER_19_271 ();
 FILLCELL_X4 FILLER_19_277 ();
 FILLCELL_X4 FILLER_19_285 ();
 FILLCELL_X4 FILLER_19_298 ();
 FILLCELL_X4 FILLER_19_311 ();
 FILLCELL_X4 FILLER_19_318 ();
 FILLCELL_X2 FILLER_19_322 ();
 FILLCELL_X4 FILLER_19_330 ();
 FILLCELL_X4 FILLER_19_347 ();
 FILLCELL_X1 FILLER_19_351 ();
 FILLCELL_X4 FILLER_19_356 ();
 FILLCELL_X8 FILLER_19_363 ();
 FILLCELL_X4 FILLER_19_375 ();
 FILLCELL_X4 FILLER_19_388 ();
 FILLCELL_X4 FILLER_19_401 ();
 FILLCELL_X2 FILLER_19_405 ();
 FILLCELL_X4 FILLER_19_417 ();
 FILLCELL_X8 FILLER_19_431 ();
 FILLCELL_X4 FILLER_19_439 ();
 FILLCELL_X2 FILLER_19_443 ();
 FILLCELL_X4 FILLER_19_454 ();
 FILLCELL_X8 FILLER_19_461 ();
 FILLCELL_X1 FILLER_19_469 ();
 FILLCELL_X4 FILLER_19_474 ();
 FILLCELL_X4 FILLER_19_488 ();
 FILLCELL_X2 FILLER_19_492 ();
 FILLCELL_X1 FILLER_19_494 ();
 FILLCELL_X4 FILLER_19_505 ();
 FILLCELL_X4 FILLER_19_511 ();
 FILLCELL_X8 FILLER_19_518 ();
 FILLCELL_X2 FILLER_19_526 ();
 FILLCELL_X1 FILLER_19_528 ();
 FILLCELL_X4 FILLER_19_531 ();
 FILLCELL_X1 FILLER_19_535 ();
 FILLCELL_X4 FILLER_19_538 ();
 FILLCELL_X4 FILLER_19_546 ();
 FILLCELL_X8 FILLER_19_554 ();
 FILLCELL_X4 FILLER_19_565 ();
 FILLCELL_X4 FILLER_19_573 ();
 FILLCELL_X8 FILLER_19_579 ();
 FILLCELL_X4 FILLER_19_587 ();
 FILLCELL_X2 FILLER_19_591 ();
 FILLCELL_X4 FILLER_19_596 ();
 FILLCELL_X8 FILLER_19_609 ();
 FILLCELL_X8 FILLER_19_621 ();
 FILLCELL_X4 FILLER_19_633 ();
 FILLCELL_X2 FILLER_19_637 ();
 FILLCELL_X1 FILLER_19_639 ();
 FILLCELL_X4 FILLER_19_643 ();
 FILLCELL_X4 FILLER_19_651 ();
 FILLCELL_X16 FILLER_19_659 ();
 FILLCELL_X4 FILLER_19_675 ();
 FILLCELL_X2 FILLER_19_679 ();
 FILLCELL_X1 FILLER_19_681 ();
 FILLCELL_X4 FILLER_19_685 ();
 FILLCELL_X4 FILLER_19_692 ();
 FILLCELL_X4 FILLER_19_699 ();
 FILLCELL_X4 FILLER_19_707 ();
 FILLCELL_X4 FILLER_19_715 ();
 FILLCELL_X4 FILLER_19_722 ();
 FILLCELL_X16 FILLER_19_736 ();
 FILLCELL_X1 FILLER_19_752 ();
 FILLCELL_X4 FILLER_19_755 ();
 FILLCELL_X8 FILLER_19_763 ();
 FILLCELL_X4 FILLER_19_775 ();
 FILLCELL_X4 FILLER_19_783 ();
 FILLCELL_X4 FILLER_19_794 ();
 FILLCELL_X8 FILLER_19_800 ();
 FILLCELL_X4 FILLER_19_808 ();
 FILLCELL_X2 FILLER_19_812 ();
 FILLCELL_X4 FILLER_19_817 ();
 FILLCELL_X8 FILLER_19_825 ();
 FILLCELL_X4 FILLER_19_833 ();
 FILLCELL_X2 FILLER_19_837 ();
 FILLCELL_X16 FILLER_19_843 ();
 FILLCELL_X8 FILLER_19_859 ();
 FILLCELL_X4 FILLER_19_867 ();
 FILLCELL_X8 FILLER_19_875 ();
 FILLCELL_X1 FILLER_19_883 ();
 FILLCELL_X8 FILLER_19_893 ();
 FILLCELL_X1 FILLER_19_901 ();
 FILLCELL_X8 FILLER_19_906 ();
 FILLCELL_X4 FILLER_19_914 ();
 FILLCELL_X2 FILLER_19_918 ();
 FILLCELL_X4 FILLER_19_923 ();
 FILLCELL_X4 FILLER_19_931 ();
 FILLCELL_X16 FILLER_19_939 ();
 FILLCELL_X2 FILLER_19_955 ();
 FILLCELL_X4 FILLER_19_961 ();
 FILLCELL_X2 FILLER_19_965 ();
 FILLCELL_X1 FILLER_19_967 ();
 FILLCELL_X16 FILLER_19_977 ();
 FILLCELL_X4 FILLER_19_993 ();
 FILLCELL_X4 FILLER_19_1001 ();
 FILLCELL_X4 FILLER_19_1009 ();
 FILLCELL_X2 FILLER_19_1013 ();
 FILLCELL_X1 FILLER_19_1015 ();
 FILLCELL_X4 FILLER_19_1021 ();
 FILLCELL_X4 FILLER_19_1029 ();
 FILLCELL_X8 FILLER_19_1037 ();
 FILLCELL_X1 FILLER_19_1045 ();
 FILLCELL_X4 FILLER_19_1055 ();
 FILLCELL_X4 FILLER_19_1063 ();
 FILLCELL_X4 FILLER_19_1073 ();
 FILLCELL_X4 FILLER_19_1080 ();
 FILLCELL_X2 FILLER_19_1084 ();
 FILLCELL_X1 FILLER_19_1086 ();
 FILLCELL_X4 FILLER_19_1091 ();
 FILLCELL_X4 FILLER_19_1105 ();
 FILLCELL_X8 FILLER_19_1116 ();
 FILLCELL_X4 FILLER_19_1128 ();
 FILLCELL_X2 FILLER_19_1132 ();
 FILLCELL_X1 FILLER_19_1134 ();
 FILLCELL_X8 FILLER_19_1145 ();
 FILLCELL_X4 FILLER_19_1162 ();
 FILLCELL_X2 FILLER_19_1166 ();
 FILLCELL_X4 FILLER_19_1172 ();
 FILLCELL_X8 FILLER_19_1186 ();
 FILLCELL_X4 FILLER_19_1194 ();
 FILLCELL_X8 FILLER_19_1202 ();
 FILLCELL_X4 FILLER_19_1210 ();
 FILLCELL_X1 FILLER_19_1214 ();
 FILLCELL_X8 FILLER_19_1222 ();
 FILLCELL_X4 FILLER_19_1230 ();
 FILLCELL_X1 FILLER_19_1234 ();
 FILLCELL_X4 FILLER_19_1245 ();
 FILLCELL_X1 FILLER_19_1249 ();
 FILLCELL_X4 FILLER_19_1259 ();
 FILLCELL_X4 FILLER_19_1264 ();
 FILLCELL_X2 FILLER_19_1268 ();
 FILLCELL_X1 FILLER_19_1270 ();
 FILLCELL_X8 FILLER_19_1281 ();
 FILLCELL_X2 FILLER_19_1289 ();
 FILLCELL_X1 FILLER_19_1291 ();
 FILLCELL_X4 FILLER_19_1296 ();
 FILLCELL_X1 FILLER_19_1300 ();
 FILLCELL_X8 FILLER_19_1304 ();
 FILLCELL_X2 FILLER_19_1312 ();
 FILLCELL_X4 FILLER_19_1318 ();
 FILLCELL_X4 FILLER_19_1331 ();
 FILLCELL_X1 FILLER_19_1335 ();
 FILLCELL_X4 FILLER_19_1343 ();
 FILLCELL_X4 FILLER_19_1357 ();
 FILLCELL_X4 FILLER_19_1364 ();
 FILLCELL_X16 FILLER_19_1372 ();
 FILLCELL_X8 FILLER_19_1388 ();
 FILLCELL_X4 FILLER_19_1401 ();
 FILLCELL_X16 FILLER_19_1407 ();
 FILLCELL_X1 FILLER_19_1423 ();
 FILLCELL_X4 FILLER_19_1428 ();
 FILLCELL_X4 FILLER_19_1436 ();
 FILLCELL_X1 FILLER_19_1440 ();
 FILLCELL_X8 FILLER_19_1445 ();
 FILLCELL_X2 FILLER_19_1453 ();
 FILLCELL_X32 FILLER_19_1462 ();
 FILLCELL_X32 FILLER_19_1494 ();
 FILLCELL_X32 FILLER_19_1526 ();
 FILLCELL_X32 FILLER_19_1558 ();
 FILLCELL_X32 FILLER_19_1590 ();
 FILLCELL_X32 FILLER_19_1622 ();
 FILLCELL_X32 FILLER_19_1654 ();
 FILLCELL_X32 FILLER_19_1686 ();
 FILLCELL_X32 FILLER_19_1718 ();
 FILLCELL_X8 FILLER_19_1750 ();
 FILLCELL_X4 FILLER_19_1758 ();
 FILLCELL_X4 FILLER_20_1 ();
 FILLCELL_X2 FILLER_20_5 ();
 FILLCELL_X1 FILLER_20_7 ();
 FILLCELL_X16 FILLER_20_12 ();
 FILLCELL_X1 FILLER_20_28 ();
 FILLCELL_X4 FILLER_20_32 ();
 FILLCELL_X1 FILLER_20_36 ();
 FILLCELL_X4 FILLER_20_47 ();
 FILLCELL_X8 FILLER_20_54 ();
 FILLCELL_X2 FILLER_20_62 ();
 FILLCELL_X4 FILLER_20_74 ();
 FILLCELL_X2 FILLER_20_78 ();
 FILLCELL_X4 FILLER_20_90 ();
 FILLCELL_X4 FILLER_20_104 ();
 FILLCELL_X8 FILLER_20_111 ();
 FILLCELL_X4 FILLER_20_119 ();
 FILLCELL_X8 FILLER_20_133 ();
 FILLCELL_X4 FILLER_20_141 ();
 FILLCELL_X1 FILLER_20_145 ();
 FILLCELL_X32 FILLER_20_165 ();
 FILLCELL_X8 FILLER_20_201 ();
 FILLCELL_X1 FILLER_20_209 ();
 FILLCELL_X16 FILLER_20_214 ();
 FILLCELL_X1 FILLER_20_230 ();
 FILLCELL_X8 FILLER_20_237 ();
 FILLCELL_X1 FILLER_20_245 ();
 FILLCELL_X8 FILLER_20_253 ();
 FILLCELL_X4 FILLER_20_261 ();
 FILLCELL_X2 FILLER_20_265 ();
 FILLCELL_X4 FILLER_20_274 ();
 FILLCELL_X1 FILLER_20_278 ();
 FILLCELL_X16 FILLER_20_282 ();
 FILLCELL_X4 FILLER_20_298 ();
 FILLCELL_X2 FILLER_20_302 ();
 FILLCELL_X1 FILLER_20_304 ();
 FILLCELL_X16 FILLER_20_309 ();
 FILLCELL_X8 FILLER_20_325 ();
 FILLCELL_X1 FILLER_20_333 ();
 FILLCELL_X8 FILLER_20_337 ();
 FILLCELL_X2 FILLER_20_345 ();
 FILLCELL_X4 FILLER_20_351 ();
 FILLCELL_X4 FILLER_20_364 ();
 FILLCELL_X8 FILLER_20_372 ();
 FILLCELL_X4 FILLER_20_383 ();
 FILLCELL_X8 FILLER_20_390 ();
 FILLCELL_X4 FILLER_20_398 ();
 FILLCELL_X1 FILLER_20_402 ();
 FILLCELL_X4 FILLER_20_406 ();
 FILLCELL_X4 FILLER_20_412 ();
 FILLCELL_X4 FILLER_20_419 ();
 FILLCELL_X4 FILLER_20_426 ();
 FILLCELL_X4 FILLER_20_439 ();
 FILLCELL_X32 FILLER_20_446 ();
 FILLCELL_X8 FILLER_20_478 ();
 FILLCELL_X4 FILLER_20_486 ();
 FILLCELL_X1 FILLER_20_490 ();
 FILLCELL_X4 FILLER_20_498 ();
 FILLCELL_X16 FILLER_20_505 ();
 FILLCELL_X1 FILLER_20_521 ();
 FILLCELL_X4 FILLER_20_526 ();
 FILLCELL_X8 FILLER_20_540 ();
 FILLCELL_X4 FILLER_20_557 ();
 FILLCELL_X8 FILLER_20_564 ();
 FILLCELL_X1 FILLER_20_572 ();
 FILLCELL_X4 FILLER_20_577 ();
 FILLCELL_X4 FILLER_20_584 ();
 FILLCELL_X1 FILLER_20_588 ();
 FILLCELL_X4 FILLER_20_593 ();
 FILLCELL_X4 FILLER_20_600 ();
 FILLCELL_X4 FILLER_20_614 ();
 FILLCELL_X8 FILLER_20_620 ();
 FILLCELL_X2 FILLER_20_628 ();
 FILLCELL_X1 FILLER_20_630 ();
 FILLCELL_X4 FILLER_20_632 ();
 FILLCELL_X2 FILLER_20_636 ();
 FILLCELL_X4 FILLER_20_642 ();
 FILLCELL_X4 FILLER_20_655 ();
 FILLCELL_X8 FILLER_20_668 ();
 FILLCELL_X1 FILLER_20_676 ();
 FILLCELL_X4 FILLER_20_681 ();
 FILLCELL_X8 FILLER_20_694 ();
 FILLCELL_X4 FILLER_20_711 ();
 FILLCELL_X4 FILLER_20_719 ();
 FILLCELL_X4 FILLER_20_725 ();
 FILLCELL_X4 FILLER_20_732 ();
 FILLCELL_X4 FILLER_20_743 ();
 FILLCELL_X4 FILLER_20_751 ();
 FILLCELL_X4 FILLER_20_764 ();
 FILLCELL_X4 FILLER_20_777 ();
 FILLCELL_X2 FILLER_20_781 ();
 FILLCELL_X1 FILLER_20_783 ();
 FILLCELL_X4 FILLER_20_788 ();
 FILLCELL_X4 FILLER_20_802 ();
 FILLCELL_X2 FILLER_20_806 ();
 FILLCELL_X1 FILLER_20_808 ();
 FILLCELL_X4 FILLER_20_818 ();
 FILLCELL_X4 FILLER_20_825 ();
 FILLCELL_X8 FILLER_20_833 ();
 FILLCELL_X4 FILLER_20_841 ();
 FILLCELL_X4 FILLER_20_854 ();
 FILLCELL_X8 FILLER_20_861 ();
 FILLCELL_X16 FILLER_20_879 ();
 FILLCELL_X4 FILLER_20_904 ();
 FILLCELL_X4 FILLER_20_911 ();
 FILLCELL_X4 FILLER_20_924 ();
 FILLCELL_X4 FILLER_20_937 ();
 FILLCELL_X4 FILLER_20_944 ();
 FILLCELL_X1 FILLER_20_948 ();
 FILLCELL_X4 FILLER_20_953 ();
 FILLCELL_X8 FILLER_20_966 ();
 FILLCELL_X4 FILLER_20_979 ();
 FILLCELL_X8 FILLER_20_987 ();
 FILLCELL_X2 FILLER_20_995 ();
 FILLCELL_X1 FILLER_20_997 ();
 FILLCELL_X4 FILLER_20_1007 ();
 FILLCELL_X4 FILLER_20_1014 ();
 FILLCELL_X4 FILLER_20_1022 ();
 FILLCELL_X4 FILLER_20_1029 ();
 FILLCELL_X8 FILLER_20_1042 ();
 FILLCELL_X2 FILLER_20_1050 ();
 FILLCELL_X4 FILLER_20_1058 ();
 FILLCELL_X4 FILLER_20_1069 ();
 FILLCELL_X16 FILLER_20_1083 ();
 FILLCELL_X2 FILLER_20_1099 ();
 FILLCELL_X8 FILLER_20_1111 ();
 FILLCELL_X4 FILLER_20_1119 ();
 FILLCELL_X2 FILLER_20_1123 ();
 FILLCELL_X4 FILLER_20_1129 ();
 FILLCELL_X8 FILLER_20_1136 ();
 FILLCELL_X4 FILLER_20_1151 ();
 FILLCELL_X8 FILLER_20_1164 ();
 FILLCELL_X1 FILLER_20_1172 ();
 FILLCELL_X8 FILLER_20_1180 ();
 FILLCELL_X2 FILLER_20_1188 ();
 FILLCELL_X4 FILLER_20_1209 ();
 FILLCELL_X4 FILLER_20_1219 ();
 FILLCELL_X8 FILLER_20_1227 ();
 FILLCELL_X2 FILLER_20_1235 ();
 FILLCELL_X4 FILLER_20_1240 ();
 FILLCELL_X4 FILLER_20_1248 ();
 FILLCELL_X2 FILLER_20_1252 ();
 FILLCELL_X1 FILLER_20_1254 ();
 FILLCELL_X4 FILLER_20_1265 ();
 FILLCELL_X2 FILLER_20_1269 ();
 FILLCELL_X1 FILLER_20_1271 ();
 FILLCELL_X4 FILLER_20_1276 ();
 FILLCELL_X4 FILLER_20_1282 ();
 FILLCELL_X4 FILLER_20_1290 ();
 FILLCELL_X4 FILLER_20_1303 ();
 FILLCELL_X4 FILLER_20_1311 ();
 FILLCELL_X4 FILLER_20_1318 ();
 FILLCELL_X2 FILLER_20_1322 ();
 FILLCELL_X8 FILLER_20_1333 ();
 FILLCELL_X4 FILLER_20_1351 ();
 FILLCELL_X8 FILLER_20_1357 ();
 FILLCELL_X1 FILLER_20_1365 ();
 FILLCELL_X8 FILLER_20_1385 ();
 FILLCELL_X4 FILLER_20_1393 ();
 FILLCELL_X4 FILLER_20_1400 ();
 FILLCELL_X2 FILLER_20_1404 ();
 FILLCELL_X4 FILLER_20_1415 ();
 FILLCELL_X8 FILLER_20_1423 ();
 FILLCELL_X2 FILLER_20_1431 ();
 FILLCELL_X4 FILLER_20_1442 ();
 FILLCELL_X2 FILLER_20_1446 ();
 FILLCELL_X4 FILLER_20_1458 ();
 FILLCELL_X4 FILLER_20_1471 ();
 FILLCELL_X1 FILLER_20_1475 ();
 FILLCELL_X32 FILLER_20_1482 ();
 FILLCELL_X32 FILLER_20_1514 ();
 FILLCELL_X32 FILLER_20_1546 ();
 FILLCELL_X32 FILLER_20_1578 ();
 FILLCELL_X32 FILLER_20_1610 ();
 FILLCELL_X32 FILLER_20_1642 ();
 FILLCELL_X32 FILLER_20_1674 ();
 FILLCELL_X32 FILLER_20_1706 ();
 FILLCELL_X16 FILLER_20_1738 ();
 FILLCELL_X8 FILLER_20_1754 ();
 FILLCELL_X4 FILLER_21_1 ();
 FILLCELL_X4 FILLER_21_15 ();
 FILLCELL_X8 FILLER_21_28 ();
 FILLCELL_X4 FILLER_21_43 ();
 FILLCELL_X4 FILLER_21_57 ();
 FILLCELL_X8 FILLER_21_65 ();
 FILLCELL_X2 FILLER_21_73 ();
 FILLCELL_X1 FILLER_21_75 ();
 FILLCELL_X8 FILLER_21_79 ();
 FILLCELL_X4 FILLER_21_87 ();
 FILLCELL_X2 FILLER_21_91 ();
 FILLCELL_X1 FILLER_21_93 ();
 FILLCELL_X8 FILLER_21_101 ();
 FILLCELL_X4 FILLER_21_109 ();
 FILLCELL_X2 FILLER_21_113 ();
 FILLCELL_X1 FILLER_21_115 ();
 FILLCELL_X4 FILLER_21_123 ();
 FILLCELL_X4 FILLER_21_129 ();
 FILLCELL_X2 FILLER_21_133 ();
 FILLCELL_X1 FILLER_21_135 ();
 FILLCELL_X4 FILLER_21_139 ();
 FILLCELL_X4 FILLER_21_147 ();
 FILLCELL_X4 FILLER_21_156 ();
 FILLCELL_X2 FILLER_21_160 ();
 FILLCELL_X4 FILLER_21_166 ();
 FILLCELL_X4 FILLER_21_187 ();
 FILLCELL_X4 FILLER_21_197 ();
 FILLCELL_X4 FILLER_21_207 ();
 FILLCELL_X4 FILLER_21_224 ();
 FILLCELL_X4 FILLER_21_231 ();
 FILLCELL_X1 FILLER_21_235 ();
 FILLCELL_X8 FILLER_21_239 ();
 FILLCELL_X4 FILLER_21_247 ();
 FILLCELL_X2 FILLER_21_251 ();
 FILLCELL_X1 FILLER_21_253 ();
 FILLCELL_X4 FILLER_21_258 ();
 FILLCELL_X2 FILLER_21_262 ();
 FILLCELL_X4 FILLER_21_274 ();
 FILLCELL_X4 FILLER_21_288 ();
 FILLCELL_X4 FILLER_21_296 ();
 FILLCELL_X32 FILLER_21_303 ();
 FILLCELL_X16 FILLER_21_335 ();
 FILLCELL_X1 FILLER_21_351 ();
 FILLCELL_X4 FILLER_21_355 ();
 FILLCELL_X4 FILLER_21_362 ();
 FILLCELL_X4 FILLER_21_375 ();
 FILLCELL_X4 FILLER_21_382 ();
 FILLCELL_X2 FILLER_21_386 ();
 FILLCELL_X1 FILLER_21_388 ();
 FILLCELL_X4 FILLER_21_392 ();
 FILLCELL_X4 FILLER_21_398 ();
 FILLCELL_X2 FILLER_21_402 ();
 FILLCELL_X4 FILLER_21_414 ();
 FILLCELL_X1 FILLER_21_418 ();
 FILLCELL_X16 FILLER_21_422 ();
 FILLCELL_X2 FILLER_21_438 ();
 FILLCELL_X1 FILLER_21_440 ();
 FILLCELL_X8 FILLER_21_444 ();
 FILLCELL_X4 FILLER_21_456 ();
 FILLCELL_X16 FILLER_21_467 ();
 FILLCELL_X4 FILLER_21_486 ();
 FILLCELL_X8 FILLER_21_499 ();
 FILLCELL_X4 FILLER_21_516 ();
 FILLCELL_X1 FILLER_21_520 ();
 FILLCELL_X4 FILLER_21_531 ();
 FILLCELL_X8 FILLER_21_538 ();
 FILLCELL_X2 FILLER_21_546 ();
 FILLCELL_X8 FILLER_21_551 ();
 FILLCELL_X4 FILLER_21_559 ();
 FILLCELL_X2 FILLER_21_563 ();
 FILLCELL_X4 FILLER_21_584 ();
 FILLCELL_X2 FILLER_21_588 ();
 FILLCELL_X1 FILLER_21_590 ();
 FILLCELL_X8 FILLER_21_600 ();
 FILLCELL_X4 FILLER_21_618 ();
 FILLCELL_X1 FILLER_21_622 ();
 FILLCELL_X8 FILLER_21_626 ();
 FILLCELL_X1 FILLER_21_634 ();
 FILLCELL_X4 FILLER_21_638 ();
 FILLCELL_X4 FILLER_21_645 ();
 FILLCELL_X4 FILLER_21_652 ();
 FILLCELL_X8 FILLER_21_659 ();
 FILLCELL_X2 FILLER_21_667 ();
 FILLCELL_X4 FILLER_21_673 ();
 FILLCELL_X16 FILLER_21_686 ();
 FILLCELL_X4 FILLER_21_702 ();
 FILLCELL_X4 FILLER_21_709 ();
 FILLCELL_X4 FILLER_21_722 ();
 FILLCELL_X4 FILLER_21_736 ();
 FILLCELL_X2 FILLER_21_740 ();
 FILLCELL_X1 FILLER_21_742 ();
 FILLCELL_X8 FILLER_21_753 ();
 FILLCELL_X1 FILLER_21_761 ();
 FILLCELL_X4 FILLER_21_765 ();
 FILLCELL_X16 FILLER_21_772 ();
 FILLCELL_X4 FILLER_21_788 ();
 FILLCELL_X2 FILLER_21_792 ();
 FILLCELL_X8 FILLER_21_797 ();
 FILLCELL_X4 FILLER_21_805 ();
 FILLCELL_X1 FILLER_21_809 ();
 FILLCELL_X4 FILLER_21_814 ();
 FILLCELL_X8 FILLER_21_827 ();
 FILLCELL_X2 FILLER_21_835 ();
 FILLCELL_X4 FILLER_21_841 ();
 FILLCELL_X4 FILLER_21_854 ();
 FILLCELL_X4 FILLER_21_862 ();
 FILLCELL_X4 FILLER_21_868 ();
 FILLCELL_X4 FILLER_21_875 ();
 FILLCELL_X8 FILLER_21_882 ();
 FILLCELL_X4 FILLER_21_890 ();
 FILLCELL_X2 FILLER_21_894 ();
 FILLCELL_X1 FILLER_21_896 ();
 FILLCELL_X4 FILLER_21_900 ();
 FILLCELL_X8 FILLER_21_907 ();
 FILLCELL_X1 FILLER_21_915 ();
 FILLCELL_X4 FILLER_21_920 ();
 FILLCELL_X4 FILLER_21_926 ();
 FILLCELL_X4 FILLER_21_935 ();
 FILLCELL_X2 FILLER_21_939 ();
 FILLCELL_X1 FILLER_21_941 ();
 FILLCELL_X4 FILLER_21_945 ();
 FILLCELL_X4 FILLER_21_959 ();
 FILLCELL_X2 FILLER_21_963 ();
 FILLCELL_X4 FILLER_21_968 ();
 FILLCELL_X4 FILLER_21_975 ();
 FILLCELL_X1 FILLER_21_979 ();
 FILLCELL_X8 FILLER_21_984 ();
 FILLCELL_X4 FILLER_21_992 ();
 FILLCELL_X1 FILLER_21_996 ();
 FILLCELL_X4 FILLER_21_1006 ();
 FILLCELL_X8 FILLER_21_1014 ();
 FILLCELL_X2 FILLER_21_1022 ();
 FILLCELL_X8 FILLER_21_1034 ();
 FILLCELL_X2 FILLER_21_1042 ();
 FILLCELL_X1 FILLER_21_1044 ();
 FILLCELL_X4 FILLER_21_1051 ();
 FILLCELL_X8 FILLER_21_1058 ();
 FILLCELL_X4 FILLER_21_1066 ();
 FILLCELL_X2 FILLER_21_1070 ();
 FILLCELL_X8 FILLER_21_1075 ();
 FILLCELL_X4 FILLER_21_1083 ();
 FILLCELL_X2 FILLER_21_1087 ();
 FILLCELL_X4 FILLER_21_1099 ();
 FILLCELL_X8 FILLER_21_1105 ();
 FILLCELL_X4 FILLER_21_1113 ();
 FILLCELL_X4 FILLER_21_1127 ();
 FILLCELL_X4 FILLER_21_1138 ();
 FILLCELL_X4 FILLER_21_1145 ();
 FILLCELL_X8 FILLER_21_1151 ();
 FILLCELL_X4 FILLER_21_1159 ();
 FILLCELL_X2 FILLER_21_1163 ();
 FILLCELL_X4 FILLER_21_1168 ();
 FILLCELL_X2 FILLER_21_1172 ();
 FILLCELL_X1 FILLER_21_1174 ();
 FILLCELL_X4 FILLER_21_1185 ();
 FILLCELL_X16 FILLER_21_1191 ();
 FILLCELL_X2 FILLER_21_1207 ();
 FILLCELL_X8 FILLER_21_1216 ();
 FILLCELL_X4 FILLER_21_1224 ();
 FILLCELL_X2 FILLER_21_1228 ();
 FILLCELL_X1 FILLER_21_1230 ();
 FILLCELL_X4 FILLER_21_1233 ();
 FILLCELL_X4 FILLER_21_1247 ();
 FILLCELL_X4 FILLER_21_1258 ();
 FILLCELL_X1 FILLER_21_1262 ();
 FILLCELL_X8 FILLER_21_1264 ();
 FILLCELL_X4 FILLER_21_1282 ();
 FILLCELL_X4 FILLER_21_1289 ();
 FILLCELL_X2 FILLER_21_1293 ();
 FILLCELL_X1 FILLER_21_1295 ();
 FILLCELL_X4 FILLER_21_1299 ();
 FILLCELL_X2 FILLER_21_1303 ();
 FILLCELL_X16 FILLER_21_1314 ();
 FILLCELL_X4 FILLER_21_1330 ();
 FILLCELL_X1 FILLER_21_1334 ();
 FILLCELL_X8 FILLER_21_1339 ();
 FILLCELL_X4 FILLER_21_1347 ();
 FILLCELL_X2 FILLER_21_1351 ();
 FILLCELL_X1 FILLER_21_1353 ();
 FILLCELL_X4 FILLER_21_1358 ();
 FILLCELL_X4 FILLER_21_1366 ();
 FILLCELL_X8 FILLER_21_1373 ();
 FILLCELL_X4 FILLER_21_1381 ();
 FILLCELL_X2 FILLER_21_1385 ();
 FILLCELL_X4 FILLER_21_1391 ();
 FILLCELL_X4 FILLER_21_1404 ();
 FILLCELL_X4 FILLER_21_1412 ();
 FILLCELL_X4 FILLER_21_1419 ();
 FILLCELL_X1 FILLER_21_1423 ();
 FILLCELL_X4 FILLER_21_1433 ();
 FILLCELL_X16 FILLER_21_1440 ();
 FILLCELL_X4 FILLER_21_1456 ();
 FILLCELL_X1 FILLER_21_1460 ();
 FILLCELL_X4 FILLER_21_1465 ();
 FILLCELL_X32 FILLER_21_1488 ();
 FILLCELL_X32 FILLER_21_1520 ();
 FILLCELL_X32 FILLER_21_1552 ();
 FILLCELL_X32 FILLER_21_1584 ();
 FILLCELL_X32 FILLER_21_1616 ();
 FILLCELL_X32 FILLER_21_1648 ();
 FILLCELL_X32 FILLER_21_1680 ();
 FILLCELL_X32 FILLER_21_1712 ();
 FILLCELL_X8 FILLER_21_1744 ();
 FILLCELL_X2 FILLER_21_1752 ();
 FILLCELL_X1 FILLER_21_1754 ();
 FILLCELL_X4 FILLER_21_1758 ();
 FILLCELL_X8 FILLER_22_1 ();
 FILLCELL_X4 FILLER_22_9 ();
 FILLCELL_X2 FILLER_22_13 ();
 FILLCELL_X4 FILLER_22_25 ();
 FILLCELL_X4 FILLER_22_32 ();
 FILLCELL_X1 FILLER_22_36 ();
 FILLCELL_X8 FILLER_22_46 ();
 FILLCELL_X4 FILLER_22_54 ();
 FILLCELL_X2 FILLER_22_58 ();
 FILLCELL_X1 FILLER_22_60 ();
 FILLCELL_X16 FILLER_22_64 ();
 FILLCELL_X1 FILLER_22_80 ();
 FILLCELL_X4 FILLER_22_84 ();
 FILLCELL_X8 FILLER_22_98 ();
 FILLCELL_X2 FILLER_22_106 ();
 FILLCELL_X1 FILLER_22_108 ();
 FILLCELL_X4 FILLER_22_113 ();
 FILLCELL_X16 FILLER_22_127 ();
 FILLCELL_X1 FILLER_22_143 ();
 FILLCELL_X8 FILLER_22_150 ();
 FILLCELL_X2 FILLER_22_158 ();
 FILLCELL_X1 FILLER_22_160 ();
 FILLCELL_X4 FILLER_22_167 ();
 FILLCELL_X8 FILLER_22_178 ();
 FILLCELL_X4 FILLER_22_186 ();
 FILLCELL_X4 FILLER_22_192 ();
 FILLCELL_X8 FILLER_22_200 ();
 FILLCELL_X2 FILLER_22_208 ();
 FILLCELL_X8 FILLER_22_214 ();
 FILLCELL_X2 FILLER_22_222 ();
 FILLCELL_X1 FILLER_22_224 ();
 FILLCELL_X8 FILLER_22_234 ();
 FILLCELL_X1 FILLER_22_242 ();
 FILLCELL_X4 FILLER_22_253 ();
 FILLCELL_X1 FILLER_22_257 ();
 FILLCELL_X4 FILLER_22_260 ();
 FILLCELL_X1 FILLER_22_264 ();
 FILLCELL_X16 FILLER_22_268 ();
 FILLCELL_X1 FILLER_22_284 ();
 FILLCELL_X4 FILLER_22_289 ();
 FILLCELL_X8 FILLER_22_297 ();
 FILLCELL_X4 FILLER_22_308 ();
 FILLCELL_X4 FILLER_22_316 ();
 FILLCELL_X4 FILLER_22_329 ();
 FILLCELL_X4 FILLER_22_337 ();
 FILLCELL_X2 FILLER_22_341 ();
 FILLCELL_X1 FILLER_22_343 ();
 FILLCELL_X4 FILLER_22_351 ();
 FILLCELL_X8 FILLER_22_357 ();
 FILLCELL_X2 FILLER_22_365 ();
 FILLCELL_X1 FILLER_22_367 ();
 FILLCELL_X8 FILLER_22_370 ();
 FILLCELL_X1 FILLER_22_378 ();
 FILLCELL_X4 FILLER_22_383 ();
 FILLCELL_X8 FILLER_22_397 ();
 FILLCELL_X2 FILLER_22_405 ();
 FILLCELL_X1 FILLER_22_407 ();
 FILLCELL_X8 FILLER_22_417 ();
 FILLCELL_X4 FILLER_22_434 ();
 FILLCELL_X1 FILLER_22_438 ();
 FILLCELL_X4 FILLER_22_449 ();
 FILLCELL_X4 FILLER_22_463 ();
 FILLCELL_X4 FILLER_22_477 ();
 FILLCELL_X8 FILLER_22_490 ();
 FILLCELL_X1 FILLER_22_498 ();
 FILLCELL_X8 FILLER_22_508 ();
 FILLCELL_X4 FILLER_22_516 ();
 FILLCELL_X2 FILLER_22_520 ();
 FILLCELL_X1 FILLER_22_522 ();
 FILLCELL_X4 FILLER_22_530 ();
 FILLCELL_X2 FILLER_22_534 ();
 FILLCELL_X4 FILLER_22_540 ();
 FILLCELL_X4 FILLER_22_548 ();
 FILLCELL_X16 FILLER_22_556 ();
 FILLCELL_X8 FILLER_22_572 ();
 FILLCELL_X4 FILLER_22_583 ();
 FILLCELL_X4 FILLER_22_590 ();
 FILLCELL_X2 FILLER_22_594 ();
 FILLCELL_X1 FILLER_22_596 ();
 FILLCELL_X4 FILLER_22_601 ();
 FILLCELL_X4 FILLER_22_612 ();
 FILLCELL_X4 FILLER_22_619 ();
 FILLCELL_X4 FILLER_22_627 ();
 FILLCELL_X4 FILLER_22_632 ();
 FILLCELL_X4 FILLER_22_645 ();
 FILLCELL_X4 FILLER_22_653 ();
 FILLCELL_X8 FILLER_22_660 ();
 FILLCELL_X4 FILLER_22_668 ();
 FILLCELL_X4 FILLER_22_676 ();
 FILLCELL_X8 FILLER_22_690 ();
 FILLCELL_X4 FILLER_22_698 ();
 FILLCELL_X2 FILLER_22_702 ();
 FILLCELL_X1 FILLER_22_704 ();
 FILLCELL_X8 FILLER_22_714 ();
 FILLCELL_X4 FILLER_22_722 ();
 FILLCELL_X4 FILLER_22_729 ();
 FILLCELL_X2 FILLER_22_733 ();
 FILLCELL_X4 FILLER_22_741 ();
 FILLCELL_X32 FILLER_22_748 ();
 FILLCELL_X2 FILLER_22_780 ();
 FILLCELL_X1 FILLER_22_782 ();
 FILLCELL_X4 FILLER_22_787 ();
 FILLCELL_X16 FILLER_22_795 ();
 FILLCELL_X8 FILLER_22_811 ();
 FILLCELL_X1 FILLER_22_819 ();
 FILLCELL_X16 FILLER_22_823 ();
 FILLCELL_X2 FILLER_22_839 ();
 FILLCELL_X1 FILLER_22_841 ();
 FILLCELL_X4 FILLER_22_847 ();
 FILLCELL_X4 FILLER_22_855 ();
 FILLCELL_X4 FILLER_22_862 ();
 FILLCELL_X1 FILLER_22_866 ();
 FILLCELL_X4 FILLER_22_874 ();
 FILLCELL_X2 FILLER_22_878 ();
 FILLCELL_X1 FILLER_22_880 ();
 FILLCELL_X8 FILLER_22_884 ();
 FILLCELL_X4 FILLER_22_892 ();
 FILLCELL_X16 FILLER_22_899 ();
 FILLCELL_X8 FILLER_22_915 ();
 FILLCELL_X4 FILLER_22_923 ();
 FILLCELL_X1 FILLER_22_927 ();
 FILLCELL_X8 FILLER_22_938 ();
 FILLCELL_X1 FILLER_22_946 ();
 FILLCELL_X16 FILLER_22_954 ();
 FILLCELL_X1 FILLER_22_970 ();
 FILLCELL_X4 FILLER_22_974 ();
 FILLCELL_X4 FILLER_22_987 ();
 FILLCELL_X4 FILLER_22_995 ();
 FILLCELL_X2 FILLER_22_999 ();
 FILLCELL_X4 FILLER_22_1004 ();
 FILLCELL_X8 FILLER_22_1011 ();
 FILLCELL_X2 FILLER_22_1019 ();
 FILLCELL_X4 FILLER_22_1023 ();
 FILLCELL_X4 FILLER_22_1034 ();
 FILLCELL_X2 FILLER_22_1038 ();
 FILLCELL_X4 FILLER_22_1046 ();
 FILLCELL_X4 FILLER_22_1057 ();
 FILLCELL_X8 FILLER_22_1065 ();
 FILLCELL_X4 FILLER_22_1076 ();
 FILLCELL_X4 FILLER_22_1083 ();
 FILLCELL_X4 FILLER_22_1090 ();
 FILLCELL_X4 FILLER_22_1097 ();
 FILLCELL_X2 FILLER_22_1101 ();
 FILLCELL_X1 FILLER_22_1103 ();
 FILLCELL_X4 FILLER_22_1108 ();
 FILLCELL_X4 FILLER_22_1119 ();
 FILLCELL_X2 FILLER_22_1123 ();
 FILLCELL_X4 FILLER_22_1129 ();
 FILLCELL_X4 FILLER_22_1136 ();
 FILLCELL_X2 FILLER_22_1140 ();
 FILLCELL_X4 FILLER_22_1152 ();
 FILLCELL_X4 FILLER_22_1165 ();
 FILLCELL_X2 FILLER_22_1169 ();
 FILLCELL_X1 FILLER_22_1171 ();
 FILLCELL_X4 FILLER_22_1181 ();
 FILLCELL_X8 FILLER_22_1188 ();
 FILLCELL_X1 FILLER_22_1196 ();
 FILLCELL_X4 FILLER_22_1207 ();
 FILLCELL_X4 FILLER_22_1220 ();
 FILLCELL_X8 FILLER_22_1227 ();
 FILLCELL_X1 FILLER_22_1235 ();
 FILLCELL_X4 FILLER_22_1246 ();
 FILLCELL_X2 FILLER_22_1250 ();
 FILLCELL_X4 FILLER_22_1259 ();
 FILLCELL_X4 FILLER_22_1273 ();
 FILLCELL_X4 FILLER_22_1280 ();
 FILLCELL_X4 FILLER_22_1287 ();
 FILLCELL_X4 FILLER_22_1294 ();
 FILLCELL_X8 FILLER_22_1301 ();
 FILLCELL_X1 FILLER_22_1309 ();
 FILLCELL_X4 FILLER_22_1314 ();
 FILLCELL_X4 FILLER_22_1321 ();
 FILLCELL_X4 FILLER_22_1328 ();
 FILLCELL_X1 FILLER_22_1332 ();
 FILLCELL_X8 FILLER_22_1352 ();
 FILLCELL_X4 FILLER_22_1369 ();
 FILLCELL_X16 FILLER_22_1376 ();
 FILLCELL_X8 FILLER_22_1392 ();
 FILLCELL_X1 FILLER_22_1400 ();
 FILLCELL_X8 FILLER_22_1404 ();
 FILLCELL_X4 FILLER_22_1412 ();
 FILLCELL_X2 FILLER_22_1416 ();
 FILLCELL_X1 FILLER_22_1418 ();
 FILLCELL_X4 FILLER_22_1422 ();
 FILLCELL_X2 FILLER_22_1426 ();
 FILLCELL_X1 FILLER_22_1428 ();
 FILLCELL_X16 FILLER_22_1432 ();
 FILLCELL_X8 FILLER_22_1448 ();
 FILLCELL_X2 FILLER_22_1456 ();
 FILLCELL_X1 FILLER_22_1458 ();
 FILLCELL_X8 FILLER_22_1462 ();
 FILLCELL_X4 FILLER_22_1476 ();
 FILLCELL_X4 FILLER_22_1487 ();
 FILLCELL_X32 FILLER_22_1495 ();
 FILLCELL_X32 FILLER_22_1527 ();
 FILLCELL_X32 FILLER_22_1559 ();
 FILLCELL_X32 FILLER_22_1591 ();
 FILLCELL_X32 FILLER_22_1623 ();
 FILLCELL_X32 FILLER_22_1655 ();
 FILLCELL_X32 FILLER_22_1687 ();
 FILLCELL_X32 FILLER_22_1719 ();
 FILLCELL_X8 FILLER_22_1751 ();
 FILLCELL_X2 FILLER_22_1759 ();
 FILLCELL_X1 FILLER_22_1761 ();
 FILLCELL_X8 FILLER_23_1 ();
 FILLCELL_X4 FILLER_23_11 ();
 FILLCELL_X2 FILLER_23_15 ();
 FILLCELL_X1 FILLER_23_17 ();
 FILLCELL_X4 FILLER_23_21 ();
 FILLCELL_X16 FILLER_23_27 ();
 FILLCELL_X2 FILLER_23_43 ();
 FILLCELL_X1 FILLER_23_45 ();
 FILLCELL_X4 FILLER_23_56 ();
 FILLCELL_X1 FILLER_23_60 ();
 FILLCELL_X4 FILLER_23_70 ();
 FILLCELL_X8 FILLER_23_78 ();
 FILLCELL_X8 FILLER_23_89 ();
 FILLCELL_X8 FILLER_23_106 ();
 FILLCELL_X4 FILLER_23_114 ();
 FILLCELL_X4 FILLER_23_121 ();
 FILLCELL_X2 FILLER_23_125 ();
 FILLCELL_X8 FILLER_23_131 ();
 FILLCELL_X1 FILLER_23_139 ();
 FILLCELL_X4 FILLER_23_146 ();
 FILLCELL_X8 FILLER_23_157 ();
 FILLCELL_X1 FILLER_23_165 ();
 FILLCELL_X8 FILLER_23_172 ();
 FILLCELL_X1 FILLER_23_180 ();
 FILLCELL_X4 FILLER_23_191 ();
 FILLCELL_X8 FILLER_23_205 ();
 FILLCELL_X1 FILLER_23_213 ();
 FILLCELL_X4 FILLER_23_223 ();
 FILLCELL_X16 FILLER_23_230 ();
 FILLCELL_X2 FILLER_23_246 ();
 FILLCELL_X1 FILLER_23_248 ();
 FILLCELL_X4 FILLER_23_251 ();
 FILLCELL_X4 FILLER_23_265 ();
 FILLCELL_X2 FILLER_23_269 ();
 FILLCELL_X8 FILLER_23_281 ();
 FILLCELL_X2 FILLER_23_289 ();
 FILLCELL_X4 FILLER_23_300 ();
 FILLCELL_X4 FILLER_23_309 ();
 FILLCELL_X4 FILLER_23_322 ();
 FILLCELL_X4 FILLER_23_330 ();
 FILLCELL_X8 FILLER_23_344 ();
 FILLCELL_X4 FILLER_23_362 ();
 FILLCELL_X2 FILLER_23_366 ();
 FILLCELL_X4 FILLER_23_370 ();
 FILLCELL_X8 FILLER_23_384 ();
 FILLCELL_X4 FILLER_23_392 ();
 FILLCELL_X2 FILLER_23_396 ();
 FILLCELL_X1 FILLER_23_398 ();
 FILLCELL_X4 FILLER_23_406 ();
 FILLCELL_X1 FILLER_23_410 ();
 FILLCELL_X4 FILLER_23_414 ();
 FILLCELL_X2 FILLER_23_418 ();
 FILLCELL_X4 FILLER_23_424 ();
 FILLCELL_X4 FILLER_23_438 ();
 FILLCELL_X8 FILLER_23_449 ();
 FILLCELL_X1 FILLER_23_457 ();
 FILLCELL_X4 FILLER_23_461 ();
 FILLCELL_X1 FILLER_23_465 ();
 FILLCELL_X4 FILLER_23_468 ();
 FILLCELL_X4 FILLER_23_475 ();
 FILLCELL_X4 FILLER_23_482 ();
 FILLCELL_X4 FILLER_23_489 ();
 FILLCELL_X4 FILLER_23_497 ();
 FILLCELL_X8 FILLER_23_504 ();
 FILLCELL_X2 FILLER_23_512 ();
 FILLCELL_X8 FILLER_23_521 ();
 FILLCELL_X1 FILLER_23_529 ();
 FILLCELL_X4 FILLER_23_533 ();
 FILLCELL_X4 FILLER_23_546 ();
 FILLCELL_X16 FILLER_23_559 ();
 FILLCELL_X4 FILLER_23_579 ();
 FILLCELL_X4 FILLER_23_592 ();
 FILLCELL_X2 FILLER_23_596 ();
 FILLCELL_X4 FILLER_23_600 ();
 FILLCELL_X2 FILLER_23_604 ();
 FILLCELL_X1 FILLER_23_606 ();
 FILLCELL_X4 FILLER_23_610 ();
 FILLCELL_X4 FILLER_23_619 ();
 FILLCELL_X2 FILLER_23_623 ();
 FILLCELL_X1 FILLER_23_625 ();
 FILLCELL_X8 FILLER_23_629 ();
 FILLCELL_X8 FILLER_23_641 ();
 FILLCELL_X2 FILLER_23_649 ();
 FILLCELL_X4 FILLER_23_655 ();
 FILLCELL_X2 FILLER_23_659 ();
 FILLCELL_X1 FILLER_23_661 ();
 FILLCELL_X16 FILLER_23_665 ();
 FILLCELL_X1 FILLER_23_681 ();
 FILLCELL_X8 FILLER_23_685 ();
 FILLCELL_X2 FILLER_23_693 ();
 FILLCELL_X1 FILLER_23_695 ();
 FILLCELL_X4 FILLER_23_699 ();
 FILLCELL_X4 FILLER_23_713 ();
 FILLCELL_X8 FILLER_23_721 ();
 FILLCELL_X2 FILLER_23_729 ();
 FILLCELL_X4 FILLER_23_738 ();
 FILLCELL_X4 FILLER_23_748 ();
 FILLCELL_X4 FILLER_23_758 ();
 FILLCELL_X4 FILLER_23_769 ();
 FILLCELL_X8 FILLER_23_779 ();
 FILLCELL_X2 FILLER_23_787 ();
 FILLCELL_X8 FILLER_23_798 ();
 FILLCELL_X2 FILLER_23_806 ();
 FILLCELL_X1 FILLER_23_808 ();
 FILLCELL_X4 FILLER_23_813 ();
 FILLCELL_X4 FILLER_23_821 ();
 FILLCELL_X4 FILLER_23_829 ();
 FILLCELL_X8 FILLER_23_836 ();
 FILLCELL_X4 FILLER_23_844 ();
 FILLCELL_X2 FILLER_23_848 ();
 FILLCELL_X1 FILLER_23_850 ();
 FILLCELL_X8 FILLER_23_861 ();
 FILLCELL_X4 FILLER_23_878 ();
 FILLCELL_X2 FILLER_23_882 ();
 FILLCELL_X4 FILLER_23_891 ();
 FILLCELL_X4 FILLER_23_905 ();
 FILLCELL_X4 FILLER_23_913 ();
 FILLCELL_X4 FILLER_23_919 ();
 FILLCELL_X4 FILLER_23_933 ();
 FILLCELL_X8 FILLER_23_940 ();
 FILLCELL_X8 FILLER_23_950 ();
 FILLCELL_X4 FILLER_23_958 ();
 FILLCELL_X4 FILLER_23_966 ();
 FILLCELL_X4 FILLER_23_979 ();
 FILLCELL_X16 FILLER_23_986 ();
 FILLCELL_X4 FILLER_23_1002 ();
 FILLCELL_X1 FILLER_23_1006 ();
 FILLCELL_X8 FILLER_23_1017 ();
 FILLCELL_X8 FILLER_23_1035 ();
 FILLCELL_X4 FILLER_23_1043 ();
 FILLCELL_X4 FILLER_23_1051 ();
 FILLCELL_X2 FILLER_23_1055 ();
 FILLCELL_X4 FILLER_23_1064 ();
 FILLCELL_X4 FILLER_23_1077 ();
 FILLCELL_X4 FILLER_23_1090 ();
 FILLCELL_X2 FILLER_23_1094 ();
 FILLCELL_X4 FILLER_23_1100 ();
 FILLCELL_X4 FILLER_23_1113 ();
 FILLCELL_X4 FILLER_23_1127 ();
 FILLCELL_X16 FILLER_23_1134 ();
 FILLCELL_X2 FILLER_23_1150 ();
 FILLCELL_X4 FILLER_23_1162 ();
 FILLCELL_X8 FILLER_23_1169 ();
 FILLCELL_X8 FILLER_23_1180 ();
 FILLCELL_X4 FILLER_23_1188 ();
 FILLCELL_X2 FILLER_23_1192 ();
 FILLCELL_X8 FILLER_23_1204 ();
 FILLCELL_X2 FILLER_23_1212 ();
 FILLCELL_X4 FILLER_23_1217 ();
 FILLCELL_X2 FILLER_23_1221 ();
 FILLCELL_X4 FILLER_23_1226 ();
 FILLCELL_X2 FILLER_23_1230 ();
 FILLCELL_X4 FILLER_23_1235 ();
 FILLCELL_X1 FILLER_23_1239 ();
 FILLCELL_X4 FILLER_23_1243 ();
 FILLCELL_X1 FILLER_23_1247 ();
 FILLCELL_X4 FILLER_23_1257 ();
 FILLCELL_X2 FILLER_23_1261 ();
 FILLCELL_X4 FILLER_23_1264 ();
 FILLCELL_X8 FILLER_23_1271 ();
 FILLCELL_X4 FILLER_23_1288 ();
 FILLCELL_X2 FILLER_23_1292 ();
 FILLCELL_X1 FILLER_23_1294 ();
 FILLCELL_X4 FILLER_23_1305 ();
 FILLCELL_X4 FILLER_23_1319 ();
 FILLCELL_X8 FILLER_23_1333 ();
 FILLCELL_X1 FILLER_23_1341 ();
 FILLCELL_X8 FILLER_23_1346 ();
 FILLCELL_X4 FILLER_23_1354 ();
 FILLCELL_X1 FILLER_23_1358 ();
 FILLCELL_X16 FILLER_23_1362 ();
 FILLCELL_X8 FILLER_23_1378 ();
 FILLCELL_X2 FILLER_23_1386 ();
 FILLCELL_X1 FILLER_23_1388 ();
 FILLCELL_X8 FILLER_23_1392 ();
 FILLCELL_X1 FILLER_23_1400 ();
 FILLCELL_X4 FILLER_23_1404 ();
 FILLCELL_X4 FILLER_23_1418 ();
 FILLCELL_X1 FILLER_23_1422 ();
 FILLCELL_X4 FILLER_23_1427 ();
 FILLCELL_X4 FILLER_23_1436 ();
 FILLCELL_X4 FILLER_23_1444 ();
 FILLCELL_X2 FILLER_23_1448 ();
 FILLCELL_X4 FILLER_23_1459 ();
 FILLCELL_X4 FILLER_23_1466 ();
 FILLCELL_X8 FILLER_23_1473 ();
 FILLCELL_X32 FILLER_23_1485 ();
 FILLCELL_X32 FILLER_23_1517 ();
 FILLCELL_X32 FILLER_23_1549 ();
 FILLCELL_X32 FILLER_23_1581 ();
 FILLCELL_X32 FILLER_23_1613 ();
 FILLCELL_X32 FILLER_23_1645 ();
 FILLCELL_X32 FILLER_23_1677 ();
 FILLCELL_X32 FILLER_23_1709 ();
 FILLCELL_X16 FILLER_23_1741 ();
 FILLCELL_X4 FILLER_23_1757 ();
 FILLCELL_X1 FILLER_23_1761 ();
 FILLCELL_X4 FILLER_24_1 ();
 FILLCELL_X16 FILLER_24_8 ();
 FILLCELL_X1 FILLER_24_24 ();
 FILLCELL_X4 FILLER_24_34 ();
 FILLCELL_X8 FILLER_24_41 ();
 FILLCELL_X8 FILLER_24_56 ();
 FILLCELL_X2 FILLER_24_64 ();
 FILLCELL_X8 FILLER_24_75 ();
 FILLCELL_X1 FILLER_24_83 ();
 FILLCELL_X4 FILLER_24_93 ();
 FILLCELL_X2 FILLER_24_97 ();
 FILLCELL_X1 FILLER_24_99 ();
 FILLCELL_X4 FILLER_24_103 ();
 FILLCELL_X4 FILLER_24_110 ();
 FILLCELL_X2 FILLER_24_114 ();
 FILLCELL_X8 FILLER_24_125 ();
 FILLCELL_X4 FILLER_24_143 ();
 FILLCELL_X1 FILLER_24_147 ();
 FILLCELL_X4 FILLER_24_152 ();
 FILLCELL_X2 FILLER_24_156 ();
 FILLCELL_X1 FILLER_24_158 ();
 FILLCELL_X8 FILLER_24_163 ();
 FILLCELL_X4 FILLER_24_174 ();
 FILLCELL_X16 FILLER_24_181 ();
 FILLCELL_X4 FILLER_24_197 ();
 FILLCELL_X1 FILLER_24_201 ();
 FILLCELL_X4 FILLER_24_205 ();
 FILLCELL_X4 FILLER_24_216 ();
 FILLCELL_X2 FILLER_24_220 ();
 FILLCELL_X4 FILLER_24_225 ();
 FILLCELL_X2 FILLER_24_229 ();
 FILLCELL_X4 FILLER_24_235 ();
 FILLCELL_X4 FILLER_24_243 ();
 FILLCELL_X1 FILLER_24_247 ();
 FILLCELL_X4 FILLER_24_251 ();
 FILLCELL_X4 FILLER_24_258 ();
 FILLCELL_X16 FILLER_24_265 ();
 FILLCELL_X8 FILLER_24_281 ();
 FILLCELL_X4 FILLER_24_289 ();
 FILLCELL_X8 FILLER_24_296 ();
 FILLCELL_X1 FILLER_24_304 ();
 FILLCELL_X4 FILLER_24_307 ();
 FILLCELL_X8 FILLER_24_315 ();
 FILLCELL_X1 FILLER_24_323 ();
 FILLCELL_X8 FILLER_24_328 ();
 FILLCELL_X4 FILLER_24_339 ();
 FILLCELL_X2 FILLER_24_343 ();
 FILLCELL_X1 FILLER_24_345 ();
 FILLCELL_X4 FILLER_24_350 ();
 FILLCELL_X4 FILLER_24_364 ();
 FILLCELL_X4 FILLER_24_375 ();
 FILLCELL_X2 FILLER_24_379 ();
 FILLCELL_X4 FILLER_24_384 ();
 FILLCELL_X1 FILLER_24_388 ();
 FILLCELL_X4 FILLER_24_393 ();
 FILLCELL_X4 FILLER_24_401 ();
 FILLCELL_X4 FILLER_24_408 ();
 FILLCELL_X8 FILLER_24_416 ();
 FILLCELL_X4 FILLER_24_424 ();
 FILLCELL_X1 FILLER_24_428 ();
 FILLCELL_X4 FILLER_24_432 ();
 FILLCELL_X2 FILLER_24_436 ();
 FILLCELL_X4 FILLER_24_440 ();
 FILLCELL_X4 FILLER_24_446 ();
 FILLCELL_X8 FILLER_24_460 ();
 FILLCELL_X16 FILLER_24_470 ();
 FILLCELL_X1 FILLER_24_486 ();
 FILLCELL_X4 FILLER_24_490 ();
 FILLCELL_X4 FILLER_24_497 ();
 FILLCELL_X2 FILLER_24_501 ();
 FILLCELL_X1 FILLER_24_503 ();
 FILLCELL_X4 FILLER_24_507 ();
 FILLCELL_X4 FILLER_24_521 ();
 FILLCELL_X4 FILLER_24_535 ();
 FILLCELL_X2 FILLER_24_539 ();
 FILLCELL_X1 FILLER_24_541 ();
 FILLCELL_X4 FILLER_24_545 ();
 FILLCELL_X8 FILLER_24_552 ();
 FILLCELL_X2 FILLER_24_560 ();
 FILLCELL_X1 FILLER_24_562 ();
 FILLCELL_X4 FILLER_24_567 ();
 FILLCELL_X4 FILLER_24_581 ();
 FILLCELL_X1 FILLER_24_585 ();
 FILLCELL_X4 FILLER_24_593 ();
 FILLCELL_X1 FILLER_24_597 ();
 FILLCELL_X8 FILLER_24_608 ();
 FILLCELL_X2 FILLER_24_616 ();
 FILLCELL_X4 FILLER_24_627 ();
 FILLCELL_X8 FILLER_24_632 ();
 FILLCELL_X1 FILLER_24_640 ();
 FILLCELL_X4 FILLER_24_650 ();
 FILLCELL_X4 FILLER_24_663 ();
 FILLCELL_X4 FILLER_24_671 ();
 FILLCELL_X1 FILLER_24_675 ();
 FILLCELL_X4 FILLER_24_683 ();
 FILLCELL_X4 FILLER_24_691 ();
 FILLCELL_X2 FILLER_24_695 ();
 FILLCELL_X1 FILLER_24_697 ();
 FILLCELL_X4 FILLER_24_700 ();
 FILLCELL_X4 FILLER_24_707 ();
 FILLCELL_X16 FILLER_24_721 ();
 FILLCELL_X1 FILLER_24_737 ();
 FILLCELL_X4 FILLER_24_742 ();
 FILLCELL_X8 FILLER_24_748 ();
 FILLCELL_X4 FILLER_24_756 ();
 FILLCELL_X1 FILLER_24_760 ();
 FILLCELL_X4 FILLER_24_765 ();
 FILLCELL_X8 FILLER_24_773 ();
 FILLCELL_X4 FILLER_24_781 ();
 FILLCELL_X1 FILLER_24_785 ();
 FILLCELL_X8 FILLER_24_790 ();
 FILLCELL_X4 FILLER_24_798 ();
 FILLCELL_X2 FILLER_24_802 ();
 FILLCELL_X4 FILLER_24_807 ();
 FILLCELL_X4 FILLER_24_820 ();
 FILLCELL_X4 FILLER_24_833 ();
 FILLCELL_X1 FILLER_24_837 ();
 FILLCELL_X4 FILLER_24_840 ();
 FILLCELL_X1 FILLER_24_844 ();
 FILLCELL_X8 FILLER_24_854 ();
 FILLCELL_X1 FILLER_24_862 ();
 FILLCELL_X4 FILLER_24_866 ();
 FILLCELL_X4 FILLER_24_880 ();
 FILLCELL_X4 FILLER_24_893 ();
 FILLCELL_X8 FILLER_24_900 ();
 FILLCELL_X8 FILLER_24_918 ();
 FILLCELL_X1 FILLER_24_926 ();
 FILLCELL_X4 FILLER_24_936 ();
 FILLCELL_X1 FILLER_24_940 ();
 FILLCELL_X4 FILLER_24_944 ();
 FILLCELL_X4 FILLER_24_958 ();
 FILLCELL_X8 FILLER_24_969 ();
 FILLCELL_X2 FILLER_24_977 ();
 FILLCELL_X4 FILLER_24_981 ();
 FILLCELL_X4 FILLER_24_990 ();
 FILLCELL_X2 FILLER_24_994 ();
 FILLCELL_X1 FILLER_24_996 ();
 FILLCELL_X4 FILLER_24_999 ();
 FILLCELL_X4 FILLER_24_1006 ();
 FILLCELL_X16 FILLER_24_1020 ();
 FILLCELL_X8 FILLER_24_1036 ();
 FILLCELL_X2 FILLER_24_1044 ();
 FILLCELL_X4 FILLER_24_1052 ();
 FILLCELL_X8 FILLER_24_1066 ();
 FILLCELL_X4 FILLER_24_1074 ();
 FILLCELL_X2 FILLER_24_1078 ();
 FILLCELL_X4 FILLER_24_1090 ();
 FILLCELL_X16 FILLER_24_1096 ();
 FILLCELL_X1 FILLER_24_1112 ();
 FILLCELL_X4 FILLER_24_1116 ();
 FILLCELL_X2 FILLER_24_1120 ();
 FILLCELL_X1 FILLER_24_1122 ();
 FILLCELL_X4 FILLER_24_1126 ();
 FILLCELL_X4 FILLER_24_1133 ();
 FILLCELL_X2 FILLER_24_1137 ();
 FILLCELL_X1 FILLER_24_1139 ();
 FILLCELL_X8 FILLER_24_1143 ();
 FILLCELL_X4 FILLER_24_1151 ();
 FILLCELL_X2 FILLER_24_1155 ();
 FILLCELL_X1 FILLER_24_1157 ();
 FILLCELL_X8 FILLER_24_1160 ();
 FILLCELL_X4 FILLER_24_1168 ();
 FILLCELL_X1 FILLER_24_1172 ();
 FILLCELL_X4 FILLER_24_1182 ();
 FILLCELL_X4 FILLER_24_1189 ();
 FILLCELL_X1 FILLER_24_1193 ();
 FILLCELL_X4 FILLER_24_1197 ();
 FILLCELL_X2 FILLER_24_1201 ();
 FILLCELL_X4 FILLER_24_1205 ();
 FILLCELL_X1 FILLER_24_1209 ();
 FILLCELL_X4 FILLER_24_1217 ();
 FILLCELL_X4 FILLER_24_1231 ();
 FILLCELL_X8 FILLER_24_1244 ();
 FILLCELL_X1 FILLER_24_1252 ();
 FILLCELL_X4 FILLER_24_1263 ();
 FILLCELL_X4 FILLER_24_1269 ();
 FILLCELL_X1 FILLER_24_1273 ();
 FILLCELL_X4 FILLER_24_1277 ();
 FILLCELL_X8 FILLER_24_1290 ();
 FILLCELL_X4 FILLER_24_1298 ();
 FILLCELL_X4 FILLER_24_1304 ();
 FILLCELL_X2 FILLER_24_1308 ();
 FILLCELL_X4 FILLER_24_1314 ();
 FILLCELL_X16 FILLER_24_1325 ();
 FILLCELL_X4 FILLER_24_1341 ();
 FILLCELL_X1 FILLER_24_1345 ();
 FILLCELL_X8 FILLER_24_1349 ();
 FILLCELL_X2 FILLER_24_1357 ();
 FILLCELL_X1 FILLER_24_1359 ();
 FILLCELL_X4 FILLER_24_1369 ();
 FILLCELL_X1 FILLER_24_1373 ();
 FILLCELL_X4 FILLER_24_1378 ();
 FILLCELL_X1 FILLER_24_1382 ();
 FILLCELL_X4 FILLER_24_1387 ();
 FILLCELL_X1 FILLER_24_1391 ();
 FILLCELL_X4 FILLER_24_1396 ();
 FILLCELL_X4 FILLER_24_1410 ();
 FILLCELL_X2 FILLER_24_1414 ();
 FILLCELL_X4 FILLER_24_1420 ();
 FILLCELL_X4 FILLER_24_1431 ();
 FILLCELL_X8 FILLER_24_1452 ();
 FILLCELL_X4 FILLER_24_1463 ();
 FILLCELL_X1 FILLER_24_1467 ();
 FILLCELL_X8 FILLER_24_1474 ();
 FILLCELL_X2 FILLER_24_1482 ();
 FILLCELL_X1 FILLER_24_1484 ();
 FILLCELL_X32 FILLER_24_1504 ();
 FILLCELL_X32 FILLER_24_1536 ();
 FILLCELL_X32 FILLER_24_1568 ();
 FILLCELL_X32 FILLER_24_1600 ();
 FILLCELL_X32 FILLER_24_1632 ();
 FILLCELL_X32 FILLER_24_1664 ();
 FILLCELL_X32 FILLER_24_1696 ();
 FILLCELL_X32 FILLER_24_1728 ();
 FILLCELL_X2 FILLER_24_1760 ();
 FILLCELL_X4 FILLER_25_1 ();
 FILLCELL_X2 FILLER_25_5 ();
 FILLCELL_X4 FILLER_25_14 ();
 FILLCELL_X4 FILLER_25_25 ();
 FILLCELL_X4 FILLER_25_32 ();
 FILLCELL_X4 FILLER_25_39 ();
 FILLCELL_X8 FILLER_25_45 ();
 FILLCELL_X2 FILLER_25_53 ();
 FILLCELL_X1 FILLER_25_55 ();
 FILLCELL_X4 FILLER_25_59 ();
 FILLCELL_X4 FILLER_25_66 ();
 FILLCELL_X4 FILLER_25_74 ();
 FILLCELL_X4 FILLER_25_82 ();
 FILLCELL_X1 FILLER_25_86 ();
 FILLCELL_X4 FILLER_25_90 ();
 FILLCELL_X4 FILLER_25_97 ();
 FILLCELL_X4 FILLER_25_110 ();
 FILLCELL_X4 FILLER_25_117 ();
 FILLCELL_X4 FILLER_25_130 ();
 FILLCELL_X2 FILLER_25_134 ();
 FILLCELL_X4 FILLER_25_140 ();
 FILLCELL_X1 FILLER_25_144 ();
 FILLCELL_X4 FILLER_25_147 ();
 FILLCELL_X16 FILLER_25_153 ();
 FILLCELL_X4 FILLER_25_169 ();
 FILLCELL_X4 FILLER_25_176 ();
 FILLCELL_X4 FILLER_25_183 ();
 FILLCELL_X4 FILLER_25_197 ();
 FILLCELL_X4 FILLER_25_203 ();
 FILLCELL_X2 FILLER_25_207 ();
 FILLCELL_X1 FILLER_25_209 ();
 FILLCELL_X4 FILLER_25_220 ();
 FILLCELL_X2 FILLER_25_224 ();
 FILLCELL_X4 FILLER_25_229 ();
 FILLCELL_X4 FILLER_25_242 ();
 FILLCELL_X1 FILLER_25_246 ();
 FILLCELL_X4 FILLER_25_256 ();
 FILLCELL_X8 FILLER_25_269 ();
 FILLCELL_X2 FILLER_25_277 ();
 FILLCELL_X1 FILLER_25_279 ();
 FILLCELL_X4 FILLER_25_284 ();
 FILLCELL_X8 FILLER_25_297 ();
 FILLCELL_X2 FILLER_25_305 ();
 FILLCELL_X1 FILLER_25_307 ();
 FILLCELL_X4 FILLER_25_310 ();
 FILLCELL_X4 FILLER_25_317 ();
 FILLCELL_X4 FILLER_25_325 ();
 FILLCELL_X4 FILLER_25_332 ();
 FILLCELL_X4 FILLER_25_345 ();
 FILLCELL_X8 FILLER_25_352 ();
 FILLCELL_X4 FILLER_25_360 ();
 FILLCELL_X4 FILLER_25_367 ();
 FILLCELL_X4 FILLER_25_380 ();
 FILLCELL_X8 FILLER_25_393 ();
 FILLCELL_X4 FILLER_25_410 ();
 FILLCELL_X4 FILLER_25_423 ();
 FILLCELL_X2 FILLER_25_427 ();
 FILLCELL_X1 FILLER_25_429 ();
 FILLCELL_X4 FILLER_25_433 ();
 FILLCELL_X4 FILLER_25_447 ();
 FILLCELL_X4 FILLER_25_455 ();
 FILLCELL_X2 FILLER_25_459 ();
 FILLCELL_X1 FILLER_25_461 ();
 FILLCELL_X4 FILLER_25_465 ();
 FILLCELL_X2 FILLER_25_469 ();
 FILLCELL_X1 FILLER_25_471 ();
 FILLCELL_X8 FILLER_25_482 ();
 FILLCELL_X4 FILLER_25_494 ();
 FILLCELL_X4 FILLER_25_507 ();
 FILLCELL_X2 FILLER_25_511 ();
 FILLCELL_X1 FILLER_25_513 ();
 FILLCELL_X4 FILLER_25_518 ();
 FILLCELL_X16 FILLER_25_524 ();
 FILLCELL_X2 FILLER_25_540 ();
 FILLCELL_X1 FILLER_25_542 ();
 FILLCELL_X4 FILLER_25_547 ();
 FILLCELL_X8 FILLER_25_556 ();
 FILLCELL_X1 FILLER_25_564 ();
 FILLCELL_X4 FILLER_25_569 ();
 FILLCELL_X8 FILLER_25_592 ();
 FILLCELL_X1 FILLER_25_600 ();
 FILLCELL_X4 FILLER_25_605 ();
 FILLCELL_X1 FILLER_25_609 ();
 FILLCELL_X4 FILLER_25_614 ();
 FILLCELL_X8 FILLER_25_623 ();
 FILLCELL_X1 FILLER_25_631 ();
 FILLCELL_X4 FILLER_25_636 ();
 FILLCELL_X16 FILLER_25_644 ();
 FILLCELL_X4 FILLER_25_660 ();
 FILLCELL_X4 FILLER_25_674 ();
 FILLCELL_X4 FILLER_25_680 ();
 FILLCELL_X2 FILLER_25_684 ();
 FILLCELL_X1 FILLER_25_686 ();
 FILLCELL_X4 FILLER_25_697 ();
 FILLCELL_X4 FILLER_25_703 ();
 FILLCELL_X8 FILLER_25_710 ();
 FILLCELL_X4 FILLER_25_718 ();
 FILLCELL_X1 FILLER_25_722 ();
 FILLCELL_X4 FILLER_25_726 ();
 FILLCELL_X8 FILLER_25_736 ();
 FILLCELL_X8 FILLER_25_750 ();
 FILLCELL_X4 FILLER_25_758 ();
 FILLCELL_X2 FILLER_25_762 ();
 FILLCELL_X4 FILLER_25_768 ();
 FILLCELL_X8 FILLER_25_782 ();
 FILLCELL_X2 FILLER_25_790 ();
 FILLCELL_X1 FILLER_25_792 ();
 FILLCELL_X4 FILLER_25_795 ();
 FILLCELL_X4 FILLER_25_809 ();
 FILLCELL_X2 FILLER_25_813 ();
 FILLCELL_X4 FILLER_25_818 ();
 FILLCELL_X4 FILLER_25_825 ();
 FILLCELL_X4 FILLER_25_832 ();
 FILLCELL_X8 FILLER_25_839 ();
 FILLCELL_X1 FILLER_25_847 ();
 FILLCELL_X4 FILLER_25_857 ();
 FILLCELL_X8 FILLER_25_864 ();
 FILLCELL_X2 FILLER_25_872 ();
 FILLCELL_X1 FILLER_25_874 ();
 FILLCELL_X4 FILLER_25_877 ();
 FILLCELL_X16 FILLER_25_883 ();
 FILLCELL_X2 FILLER_25_899 ();
 FILLCELL_X1 FILLER_25_901 ();
 FILLCELL_X4 FILLER_25_905 ();
 FILLCELL_X4 FILLER_25_918 ();
 FILLCELL_X4 FILLER_25_929 ();
 FILLCELL_X8 FILLER_25_938 ();
 FILLCELL_X4 FILLER_25_956 ();
 FILLCELL_X4 FILLER_25_963 ();
 FILLCELL_X4 FILLER_25_977 ();
 FILLCELL_X2 FILLER_25_981 ();
 FILLCELL_X4 FILLER_25_987 ();
 FILLCELL_X4 FILLER_25_1001 ();
 FILLCELL_X4 FILLER_25_1008 ();
 FILLCELL_X4 FILLER_25_1019 ();
 FILLCELL_X8 FILLER_25_1026 ();
 FILLCELL_X4 FILLER_25_1043 ();
 FILLCELL_X4 FILLER_25_1054 ();
 FILLCELL_X1 FILLER_25_1058 ();
 FILLCELL_X4 FILLER_25_1062 ();
 FILLCELL_X16 FILLER_25_1068 ();
 FILLCELL_X2 FILLER_25_1084 ();
 FILLCELL_X4 FILLER_25_1093 ();
 FILLCELL_X4 FILLER_25_1107 ();
 FILLCELL_X4 FILLER_25_1113 ();
 FILLCELL_X4 FILLER_25_1121 ();
 FILLCELL_X1 FILLER_25_1125 ();
 FILLCELL_X4 FILLER_25_1135 ();
 FILLCELL_X4 FILLER_25_1149 ();
 FILLCELL_X4 FILLER_25_1163 ();
 FILLCELL_X4 FILLER_25_1174 ();
 FILLCELL_X4 FILLER_25_1182 ();
 FILLCELL_X4 FILLER_25_1189 ();
 FILLCELL_X8 FILLER_25_1202 ();
 FILLCELL_X2 FILLER_25_1210 ();
 FILLCELL_X4 FILLER_25_1219 ();
 FILLCELL_X8 FILLER_25_1226 ();
 FILLCELL_X2 FILLER_25_1234 ();
 FILLCELL_X4 FILLER_25_1243 ();
 FILLCELL_X1 FILLER_25_1247 ();
 FILLCELL_X8 FILLER_25_1250 ();
 FILLCELL_X4 FILLER_25_1258 ();
 FILLCELL_X1 FILLER_25_1262 ();
 FILLCELL_X4 FILLER_25_1264 ();
 FILLCELL_X2 FILLER_25_1268 ();
 FILLCELL_X4 FILLER_25_1273 ();
 FILLCELL_X2 FILLER_25_1277 ();
 FILLCELL_X4 FILLER_25_1286 ();
 FILLCELL_X16 FILLER_25_1293 ();
 FILLCELL_X4 FILLER_25_1309 ();
 FILLCELL_X2 FILLER_25_1313 ();
 FILLCELL_X1 FILLER_25_1315 ();
 FILLCELL_X8 FILLER_25_1326 ();
 FILLCELL_X4 FILLER_25_1338 ();
 FILLCELL_X4 FILLER_25_1346 ();
 FILLCELL_X4 FILLER_25_1354 ();
 FILLCELL_X8 FILLER_25_1361 ();
 FILLCELL_X4 FILLER_25_1373 ();
 FILLCELL_X4 FILLER_25_1386 ();
 FILLCELL_X8 FILLER_25_1399 ();
 FILLCELL_X4 FILLER_25_1414 ();
 FILLCELL_X8 FILLER_25_1420 ();
 FILLCELL_X4 FILLER_25_1428 ();
 FILLCELL_X2 FILLER_25_1432 ();
 FILLCELL_X4 FILLER_25_1439 ();
 FILLCELL_X4 FILLER_25_1445 ();
 FILLCELL_X2 FILLER_25_1449 ();
 FILLCELL_X4 FILLER_25_1455 ();
 FILLCELL_X8 FILLER_25_1465 ();
 FILLCELL_X2 FILLER_25_1473 ();
 FILLCELL_X4 FILLER_25_1481 ();
 FILLCELL_X4 FILLER_25_1489 ();
 FILLCELL_X32 FILLER_25_1497 ();
 FILLCELL_X32 FILLER_25_1529 ();
 FILLCELL_X32 FILLER_25_1561 ();
 FILLCELL_X32 FILLER_25_1593 ();
 FILLCELL_X32 FILLER_25_1625 ();
 FILLCELL_X32 FILLER_25_1657 ();
 FILLCELL_X32 FILLER_25_1689 ();
 FILLCELL_X32 FILLER_25_1721 ();
 FILLCELL_X8 FILLER_25_1753 ();
 FILLCELL_X1 FILLER_25_1761 ();
 FILLCELL_X4 FILLER_26_1 ();
 FILLCELL_X4 FILLER_26_8 ();
 FILLCELL_X4 FILLER_26_22 ();
 FILLCELL_X4 FILLER_26_30 ();
 FILLCELL_X2 FILLER_26_34 ();
 FILLCELL_X1 FILLER_26_36 ();
 FILLCELL_X4 FILLER_26_41 ();
 FILLCELL_X2 FILLER_26_45 ();
 FILLCELL_X4 FILLER_26_57 ();
 FILLCELL_X16 FILLER_26_64 ();
 FILLCELL_X1 FILLER_26_80 ();
 FILLCELL_X4 FILLER_26_90 ();
 FILLCELL_X8 FILLER_26_97 ();
 FILLCELL_X4 FILLER_26_105 ();
 FILLCELL_X4 FILLER_26_111 ();
 FILLCELL_X4 FILLER_26_118 ();
 FILLCELL_X1 FILLER_26_122 ();
 FILLCELL_X4 FILLER_26_126 ();
 FILLCELL_X4 FILLER_26_134 ();
 FILLCELL_X4 FILLER_26_142 ();
 FILLCELL_X1 FILLER_26_146 ();
 FILLCELL_X4 FILLER_26_153 ();
 FILLCELL_X4 FILLER_26_164 ();
 FILLCELL_X4 FILLER_26_171 ();
 FILLCELL_X8 FILLER_26_184 ();
 FILLCELL_X4 FILLER_26_195 ();
 FILLCELL_X2 FILLER_26_199 ();
 FILLCELL_X1 FILLER_26_201 ();
 FILLCELL_X4 FILLER_26_209 ();
 FILLCELL_X16 FILLER_26_217 ();
 FILLCELL_X4 FILLER_26_233 ();
 FILLCELL_X4 FILLER_26_240 ();
 FILLCELL_X4 FILLER_26_247 ();
 FILLCELL_X2 FILLER_26_251 ();
 FILLCELL_X1 FILLER_26_253 ();
 FILLCELL_X4 FILLER_26_256 ();
 FILLCELL_X8 FILLER_26_270 ();
 FILLCELL_X2 FILLER_26_278 ();
 FILLCELL_X4 FILLER_26_290 ();
 FILLCELL_X4 FILLER_26_298 ();
 FILLCELL_X1 FILLER_26_302 ();
 FILLCELL_X4 FILLER_26_307 ();
 FILLCELL_X8 FILLER_26_318 ();
 FILLCELL_X1 FILLER_26_326 ();
 FILLCELL_X4 FILLER_26_336 ();
 FILLCELL_X4 FILLER_26_344 ();
 FILLCELL_X2 FILLER_26_348 ();
 FILLCELL_X4 FILLER_26_354 ();
 FILLCELL_X8 FILLER_26_367 ();
 FILLCELL_X4 FILLER_26_375 ();
 FILLCELL_X2 FILLER_26_379 ();
 FILLCELL_X16 FILLER_26_384 ();
 FILLCELL_X8 FILLER_26_400 ();
 FILLCELL_X2 FILLER_26_408 ();
 FILLCELL_X4 FILLER_26_413 ();
 FILLCELL_X8 FILLER_26_420 ();
 FILLCELL_X4 FILLER_26_428 ();
 FILLCELL_X2 FILLER_26_432 ();
 FILLCELL_X1 FILLER_26_434 ();
 FILLCELL_X8 FILLER_26_438 ();
 FILLCELL_X2 FILLER_26_446 ();
 FILLCELL_X4 FILLER_26_457 ();
 FILLCELL_X8 FILLER_26_471 ();
 FILLCELL_X2 FILLER_26_479 ();
 FILLCELL_X4 FILLER_26_485 ();
 FILLCELL_X4 FILLER_26_498 ();
 FILLCELL_X8 FILLER_26_505 ();
 FILLCELL_X4 FILLER_26_513 ();
 FILLCELL_X2 FILLER_26_517 ();
 FILLCELL_X4 FILLER_26_522 ();
 FILLCELL_X2 FILLER_26_526 ();
 FILLCELL_X4 FILLER_26_532 ();
 FILLCELL_X4 FILLER_26_540 ();
 FILLCELL_X4 FILLER_26_553 ();
 FILLCELL_X8 FILLER_26_560 ();
 FILLCELL_X4 FILLER_26_568 ();
 FILLCELL_X1 FILLER_26_572 ();
 FILLCELL_X16 FILLER_26_576 ();
 FILLCELL_X4 FILLER_26_592 ();
 FILLCELL_X1 FILLER_26_596 ();
 FILLCELL_X4 FILLER_26_606 ();
 FILLCELL_X4 FILLER_26_619 ();
 FILLCELL_X4 FILLER_26_627 ();
 FILLCELL_X8 FILLER_26_632 ();
 FILLCELL_X4 FILLER_26_640 ();
 FILLCELL_X2 FILLER_26_644 ();
 FILLCELL_X4 FILLER_26_653 ();
 FILLCELL_X4 FILLER_26_660 ();
 FILLCELL_X2 FILLER_26_664 ();
 FILLCELL_X1 FILLER_26_666 ();
 FILLCELL_X4 FILLER_26_670 ();
 FILLCELL_X2 FILLER_26_674 ();
 FILLCELL_X4 FILLER_26_686 ();
 FILLCELL_X2 FILLER_26_690 ();
 FILLCELL_X1 FILLER_26_692 ();
 FILLCELL_X8 FILLER_26_702 ();
 FILLCELL_X2 FILLER_26_710 ();
 FILLCELL_X16 FILLER_26_721 ();
 FILLCELL_X1 FILLER_26_737 ();
 FILLCELL_X4 FILLER_26_740 ();
 FILLCELL_X4 FILLER_26_747 ();
 FILLCELL_X4 FILLER_26_754 ();
 FILLCELL_X4 FILLER_26_767 ();
 FILLCELL_X2 FILLER_26_771 ();
 FILLCELL_X1 FILLER_26_773 ();
 FILLCELL_X4 FILLER_26_777 ();
 FILLCELL_X4 FILLER_26_783 ();
 FILLCELL_X1 FILLER_26_787 ();
 FILLCELL_X4 FILLER_26_792 ();
 FILLCELL_X4 FILLER_26_800 ();
 FILLCELL_X4 FILLER_26_813 ();
 FILLCELL_X2 FILLER_26_817 ();
 FILLCELL_X1 FILLER_26_819 ();
 FILLCELL_X4 FILLER_26_824 ();
 FILLCELL_X8 FILLER_26_838 ();
 FILLCELL_X4 FILLER_26_846 ();
 FILLCELL_X2 FILLER_26_850 ();
 FILLCELL_X8 FILLER_26_855 ();
 FILLCELL_X4 FILLER_26_863 ();
 FILLCELL_X2 FILLER_26_867 ();
 FILLCELL_X4 FILLER_26_872 ();
 FILLCELL_X4 FILLER_26_886 ();
 FILLCELL_X1 FILLER_26_890 ();
 FILLCELL_X4 FILLER_26_900 ();
 FILLCELL_X4 FILLER_26_907 ();
 FILLCELL_X8 FILLER_26_914 ();
 FILLCELL_X2 FILLER_26_922 ();
 FILLCELL_X1 FILLER_26_924 ();
 FILLCELL_X16 FILLER_26_928 ();
 FILLCELL_X2 FILLER_26_944 ();
 FILLCELL_X4 FILLER_26_955 ();
 FILLCELL_X8 FILLER_26_962 ();
 FILLCELL_X4 FILLER_26_970 ();
 FILLCELL_X8 FILLER_26_984 ();
 FILLCELL_X8 FILLER_26_999 ();
 FILLCELL_X2 FILLER_26_1007 ();
 FILLCELL_X1 FILLER_26_1009 ();
 FILLCELL_X4 FILLER_26_1020 ();
 FILLCELL_X4 FILLER_26_1033 ();
 FILLCELL_X4 FILLER_26_1047 ();
 FILLCELL_X4 FILLER_26_1054 ();
 FILLCELL_X4 FILLER_26_1060 ();
 FILLCELL_X4 FILLER_26_1071 ();
 FILLCELL_X1 FILLER_26_1075 ();
 FILLCELL_X4 FILLER_26_1079 ();
 FILLCELL_X2 FILLER_26_1083 ();
 FILLCELL_X4 FILLER_26_1095 ();
 FILLCELL_X8 FILLER_26_1102 ();
 FILLCELL_X4 FILLER_26_1114 ();
 FILLCELL_X16 FILLER_26_1127 ();
 FILLCELL_X2 FILLER_26_1143 ();
 FILLCELL_X4 FILLER_26_1155 ();
 FILLCELL_X4 FILLER_26_1161 ();
 FILLCELL_X2 FILLER_26_1165 ();
 FILLCELL_X1 FILLER_26_1167 ();
 FILLCELL_X4 FILLER_26_1172 ();
 FILLCELL_X4 FILLER_26_1185 ();
 FILLCELL_X4 FILLER_26_1192 ();
 FILLCELL_X1 FILLER_26_1196 ();
 FILLCELL_X4 FILLER_26_1207 ();
 FILLCELL_X8 FILLER_26_1221 ();
 FILLCELL_X1 FILLER_26_1229 ();
 FILLCELL_X4 FILLER_26_1240 ();
 FILLCELL_X4 FILLER_26_1254 ();
 FILLCELL_X1 FILLER_26_1258 ();
 FILLCELL_X4 FILLER_26_1261 ();
 FILLCELL_X2 FILLER_26_1265 ();
 FILLCELL_X8 FILLER_26_1277 ();
 FILLCELL_X4 FILLER_26_1285 ();
 FILLCELL_X1 FILLER_26_1289 ();
 FILLCELL_X4 FILLER_26_1299 ();
 FILLCELL_X16 FILLER_26_1306 ();
 FILLCELL_X4 FILLER_26_1322 ();
 FILLCELL_X2 FILLER_26_1326 ();
 FILLCELL_X8 FILLER_26_1330 ();
 FILLCELL_X4 FILLER_26_1338 ();
 FILLCELL_X1 FILLER_26_1342 ();
 FILLCELL_X4 FILLER_26_1352 ();
 FILLCELL_X8 FILLER_26_1365 ();
 FILLCELL_X4 FILLER_26_1373 ();
 FILLCELL_X2 FILLER_26_1377 ();
 FILLCELL_X4 FILLER_26_1382 ();
 FILLCELL_X4 FILLER_26_1389 ();
 FILLCELL_X1 FILLER_26_1393 ();
 FILLCELL_X32 FILLER_26_1396 ();
 FILLCELL_X8 FILLER_26_1428 ();
 FILLCELL_X2 FILLER_26_1436 ();
 FILLCELL_X1 FILLER_26_1438 ();
 FILLCELL_X8 FILLER_26_1448 ();
 FILLCELL_X8 FILLER_26_1458 ();
 FILLCELL_X2 FILLER_26_1466 ();
 FILLCELL_X32 FILLER_26_1474 ();
 FILLCELL_X32 FILLER_26_1506 ();
 FILLCELL_X32 FILLER_26_1538 ();
 FILLCELL_X32 FILLER_26_1570 ();
 FILLCELL_X32 FILLER_26_1602 ();
 FILLCELL_X32 FILLER_26_1634 ();
 FILLCELL_X32 FILLER_26_1666 ();
 FILLCELL_X32 FILLER_26_1698 ();
 FILLCELL_X32 FILLER_26_1730 ();
 FILLCELL_X4 FILLER_27_1 ();
 FILLCELL_X2 FILLER_27_5 ();
 FILLCELL_X1 FILLER_27_7 ();
 FILLCELL_X4 FILLER_27_18 ();
 FILLCELL_X16 FILLER_27_25 ();
 FILLCELL_X4 FILLER_27_41 ();
 FILLCELL_X2 FILLER_27_45 ();
 FILLCELL_X1 FILLER_27_47 ();
 FILLCELL_X8 FILLER_27_58 ();
 FILLCELL_X2 FILLER_27_66 ();
 FILLCELL_X8 FILLER_27_78 ();
 FILLCELL_X1 FILLER_27_86 ();
 FILLCELL_X4 FILLER_27_90 ();
 FILLCELL_X8 FILLER_27_96 ();
 FILLCELL_X2 FILLER_27_104 ();
 FILLCELL_X8 FILLER_27_116 ();
 FILLCELL_X4 FILLER_27_127 ();
 FILLCELL_X8 FILLER_27_141 ();
 FILLCELL_X4 FILLER_27_149 ();
 FILLCELL_X2 FILLER_27_153 ();
 FILLCELL_X8 FILLER_27_165 ();
 FILLCELL_X2 FILLER_27_173 ();
 FILLCELL_X1 FILLER_27_175 ();
 FILLCELL_X4 FILLER_27_186 ();
 FILLCELL_X8 FILLER_27_200 ();
 FILLCELL_X4 FILLER_27_208 ();
 FILLCELL_X4 FILLER_27_219 ();
 FILLCELL_X2 FILLER_27_223 ();
 FILLCELL_X4 FILLER_27_229 ();
 FILLCELL_X4 FILLER_27_242 ();
 FILLCELL_X4 FILLER_27_250 ();
 FILLCELL_X1 FILLER_27_254 ();
 FILLCELL_X4 FILLER_27_258 ();
 FILLCELL_X4 FILLER_27_265 ();
 FILLCELL_X4 FILLER_27_276 ();
 FILLCELL_X4 FILLER_27_283 ();
 FILLCELL_X1 FILLER_27_287 ();
 FILLCELL_X8 FILLER_27_290 ();
 FILLCELL_X2 FILLER_27_298 ();
 FILLCELL_X4 FILLER_27_310 ();
 FILLCELL_X4 FILLER_27_324 ();
 FILLCELL_X4 FILLER_27_331 ();
 FILLCELL_X4 FILLER_27_338 ();
 FILLCELL_X2 FILLER_27_342 ();
 FILLCELL_X4 FILLER_27_348 ();
 FILLCELL_X4 FILLER_27_361 ();
 FILLCELL_X8 FILLER_27_374 ();
 FILLCELL_X2 FILLER_27_382 ();
 FILLCELL_X1 FILLER_27_384 ();
 FILLCELL_X8 FILLER_27_395 ();
 FILLCELL_X4 FILLER_27_405 ();
 FILLCELL_X4 FILLER_27_419 ();
 FILLCELL_X4 FILLER_27_433 ();
 FILLCELL_X4 FILLER_27_446 ();
 FILLCELL_X16 FILLER_27_453 ();
 FILLCELL_X4 FILLER_27_469 ();
 FILLCELL_X8 FILLER_27_477 ();
 FILLCELL_X2 FILLER_27_485 ();
 FILLCELL_X16 FILLER_27_491 ();
 FILLCELL_X2 FILLER_27_507 ();
 FILLCELL_X4 FILLER_27_513 ();
 FILLCELL_X8 FILLER_27_527 ();
 FILLCELL_X4 FILLER_27_535 ();
 FILLCELL_X4 FILLER_27_548 ();
 FILLCELL_X8 FILLER_27_555 ();
 FILLCELL_X4 FILLER_27_563 ();
 FILLCELL_X4 FILLER_27_571 ();
 FILLCELL_X4 FILLER_27_579 ();
 FILLCELL_X1 FILLER_27_583 ();
 FILLCELL_X4 FILLER_27_587 ();
 FILLCELL_X4 FILLER_27_594 ();
 FILLCELL_X4 FILLER_27_601 ();
 FILLCELL_X2 FILLER_27_605 ();
 FILLCELL_X1 FILLER_27_607 ();
 FILLCELL_X4 FILLER_27_611 ();
 FILLCELL_X8 FILLER_27_618 ();
 FILLCELL_X8 FILLER_27_629 ();
 FILLCELL_X4 FILLER_27_641 ();
 FILLCELL_X4 FILLER_27_655 ();
 FILLCELL_X2 FILLER_27_659 ();
 FILLCELL_X4 FILLER_27_664 ();
 FILLCELL_X4 FILLER_27_671 ();
 FILLCELL_X8 FILLER_27_678 ();
 FILLCELL_X2 FILLER_27_686 ();
 FILLCELL_X4 FILLER_27_691 ();
 FILLCELL_X4 FILLER_27_698 ();
 FILLCELL_X8 FILLER_27_704 ();
 FILLCELL_X4 FILLER_27_712 ();
 FILLCELL_X1 FILLER_27_716 ();
 FILLCELL_X8 FILLER_27_724 ();
 FILLCELL_X4 FILLER_27_732 ();
 FILLCELL_X2 FILLER_27_736 ();
 FILLCELL_X1 FILLER_27_738 ();
 FILLCELL_X4 FILLER_27_742 ();
 FILLCELL_X16 FILLER_27_755 ();
 FILLCELL_X4 FILLER_27_771 ();
 FILLCELL_X4 FILLER_27_785 ();
 FILLCELL_X4 FILLER_27_799 ();
 FILLCELL_X4 FILLER_27_805 ();
 FILLCELL_X4 FILLER_27_812 ();
 FILLCELL_X4 FILLER_27_819 ();
 FILLCELL_X2 FILLER_27_823 ();
 FILLCELL_X1 FILLER_27_825 ();
 FILLCELL_X4 FILLER_27_833 ();
 FILLCELL_X4 FILLER_27_839 ();
 FILLCELL_X1 FILLER_27_843 ();
 FILLCELL_X4 FILLER_27_846 ();
 FILLCELL_X4 FILLER_27_860 ();
 FILLCELL_X8 FILLER_27_871 ();
 FILLCELL_X4 FILLER_27_889 ();
 FILLCELL_X2 FILLER_27_893 ();
 FILLCELL_X4 FILLER_27_904 ();
 FILLCELL_X2 FILLER_27_908 ();
 FILLCELL_X16 FILLER_27_914 ();
 FILLCELL_X4 FILLER_27_930 ();
 FILLCELL_X1 FILLER_27_934 ();
 FILLCELL_X8 FILLER_27_944 ();
 FILLCELL_X2 FILLER_27_952 ();
 FILLCELL_X4 FILLER_27_961 ();
 FILLCELL_X4 FILLER_27_968 ();
 FILLCELL_X8 FILLER_27_975 ();
 FILLCELL_X2 FILLER_27_983 ();
 FILLCELL_X4 FILLER_27_989 ();
 FILLCELL_X8 FILLER_27_995 ();
 FILLCELL_X4 FILLER_27_1003 ();
 FILLCELL_X2 FILLER_27_1007 ();
 FILLCELL_X4 FILLER_27_1019 ();
 FILLCELL_X4 FILLER_27_1030 ();
 FILLCELL_X1 FILLER_27_1034 ();
 FILLCELL_X4 FILLER_27_1038 ();
 FILLCELL_X4 FILLER_27_1045 ();
 FILLCELL_X2 FILLER_27_1049 ();
 FILLCELL_X4 FILLER_27_1061 ();
 FILLCELL_X4 FILLER_27_1075 ();
 FILLCELL_X4 FILLER_27_1088 ();
 FILLCELL_X4 FILLER_27_1101 ();
 FILLCELL_X16 FILLER_27_1108 ();
 FILLCELL_X1 FILLER_27_1124 ();
 FILLCELL_X4 FILLER_27_1134 ();
 FILLCELL_X4 FILLER_27_1141 ();
 FILLCELL_X4 FILLER_27_1148 ();
 FILLCELL_X4 FILLER_27_1154 ();
 FILLCELL_X1 FILLER_27_1158 ();
 FILLCELL_X8 FILLER_27_1166 ();
 FILLCELL_X4 FILLER_27_1174 ();
 FILLCELL_X2 FILLER_27_1178 ();
 FILLCELL_X4 FILLER_27_1184 ();
 FILLCELL_X8 FILLER_27_1191 ();
 FILLCELL_X4 FILLER_27_1199 ();
 FILLCELL_X16 FILLER_27_1205 ();
 FILLCELL_X1 FILLER_27_1221 ();
 FILLCELL_X8 FILLER_27_1225 ();
 FILLCELL_X8 FILLER_27_1235 ();
 FILLCELL_X1 FILLER_27_1243 ();
 FILLCELL_X8 FILLER_27_1247 ();
 FILLCELL_X1 FILLER_27_1255 ();
 FILLCELL_X4 FILLER_27_1259 ();
 FILLCELL_X8 FILLER_27_1264 ();
 FILLCELL_X4 FILLER_27_1282 ();
 FILLCELL_X2 FILLER_27_1286 ();
 FILLCELL_X4 FILLER_27_1297 ();
 FILLCELL_X4 FILLER_27_1308 ();
 FILLCELL_X4 FILLER_27_1316 ();
 FILLCELL_X4 FILLER_27_1324 ();
 FILLCELL_X4 FILLER_27_1331 ();
 FILLCELL_X8 FILLER_27_1338 ();
 FILLCELL_X1 FILLER_27_1346 ();
 FILLCELL_X8 FILLER_27_1350 ();
 FILLCELL_X4 FILLER_27_1362 ();
 FILLCELL_X16 FILLER_27_1369 ();
 FILLCELL_X4 FILLER_27_1385 ();
 FILLCELL_X1 FILLER_27_1389 ();
 FILLCELL_X4 FILLER_27_1393 ();
 FILLCELL_X8 FILLER_27_1407 ();
 FILLCELL_X1 FILLER_27_1415 ();
 FILLCELL_X4 FILLER_27_1425 ();
 FILLCELL_X4 FILLER_27_1432 ();
 FILLCELL_X4 FILLER_27_1439 ();
 FILLCELL_X4 FILLER_27_1446 ();
 FILLCELL_X8 FILLER_27_1452 ();
 FILLCELL_X4 FILLER_27_1463 ();
 FILLCELL_X32 FILLER_27_1474 ();
 FILLCELL_X32 FILLER_27_1506 ();
 FILLCELL_X32 FILLER_27_1538 ();
 FILLCELL_X32 FILLER_27_1570 ();
 FILLCELL_X32 FILLER_27_1602 ();
 FILLCELL_X32 FILLER_27_1634 ();
 FILLCELL_X32 FILLER_27_1666 ();
 FILLCELL_X32 FILLER_27_1698 ();
 FILLCELL_X32 FILLER_27_1730 ();
 FILLCELL_X16 FILLER_28_1 ();
 FILLCELL_X4 FILLER_28_26 ();
 FILLCELL_X8 FILLER_28_33 ();
 FILLCELL_X4 FILLER_28_41 ();
 FILLCELL_X1 FILLER_28_45 ();
 FILLCELL_X4 FILLER_28_48 ();
 FILLCELL_X4 FILLER_28_59 ();
 FILLCELL_X1 FILLER_28_63 ();
 FILLCELL_X4 FILLER_28_71 ();
 FILLCELL_X8 FILLER_28_85 ();
 FILLCELL_X1 FILLER_28_93 ();
 FILLCELL_X4 FILLER_28_98 ();
 FILLCELL_X4 FILLER_28_105 ();
 FILLCELL_X1 FILLER_28_109 ();
 FILLCELL_X4 FILLER_28_117 ();
 FILLCELL_X8 FILLER_28_124 ();
 FILLCELL_X2 FILLER_28_132 ();
 FILLCELL_X8 FILLER_28_137 ();
 FILLCELL_X2 FILLER_28_145 ();
 FILLCELL_X1 FILLER_28_147 ();
 FILLCELL_X8 FILLER_28_150 ();
 FILLCELL_X4 FILLER_28_161 ();
 FILLCELL_X2 FILLER_28_165 ();
 FILLCELL_X8 FILLER_28_176 ();
 FILLCELL_X2 FILLER_28_184 ();
 FILLCELL_X1 FILLER_28_186 ();
 FILLCELL_X8 FILLER_28_189 ();
 FILLCELL_X4 FILLER_28_197 ();
 FILLCELL_X2 FILLER_28_201 ();
 FILLCELL_X4 FILLER_28_206 ();
 FILLCELL_X4 FILLER_28_219 ();
 FILLCELL_X2 FILLER_28_223 ();
 FILLCELL_X16 FILLER_28_235 ();
 FILLCELL_X1 FILLER_28_251 ();
 FILLCELL_X8 FILLER_28_256 ();
 FILLCELL_X4 FILLER_28_268 ();
 FILLCELL_X1 FILLER_28_272 ();
 FILLCELL_X4 FILLER_28_277 ();
 FILLCELL_X4 FILLER_28_284 ();
 FILLCELL_X2 FILLER_28_288 ();
 FILLCELL_X1 FILLER_28_290 ();
 FILLCELL_X4 FILLER_28_300 ();
 FILLCELL_X2 FILLER_28_304 ();
 FILLCELL_X16 FILLER_28_309 ();
 FILLCELL_X2 FILLER_28_325 ();
 FILLCELL_X1 FILLER_28_327 ();
 FILLCELL_X4 FILLER_28_331 ();
 FILLCELL_X8 FILLER_28_338 ();
 FILLCELL_X1 FILLER_28_346 ();
 FILLCELL_X4 FILLER_28_350 ();
 FILLCELL_X4 FILLER_28_358 ();
 FILLCELL_X2 FILLER_28_362 ();
 FILLCELL_X1 FILLER_28_364 ();
 FILLCELL_X4 FILLER_28_368 ();
 FILLCELL_X4 FILLER_28_375 ();
 FILLCELL_X2 FILLER_28_379 ();
 FILLCELL_X4 FILLER_28_385 ();
 FILLCELL_X4 FILLER_28_391 ();
 FILLCELL_X1 FILLER_28_395 ();
 FILLCELL_X4 FILLER_28_399 ();
 FILLCELL_X4 FILLER_28_413 ();
 FILLCELL_X1 FILLER_28_417 ();
 FILLCELL_X16 FILLER_28_420 ();
 FILLCELL_X4 FILLER_28_436 ();
 FILLCELL_X2 FILLER_28_440 ();
 FILLCELL_X16 FILLER_28_445 ();
 FILLCELL_X4 FILLER_28_461 ();
 FILLCELL_X2 FILLER_28_465 ();
 FILLCELL_X1 FILLER_28_467 ();
 FILLCELL_X8 FILLER_28_474 ();
 FILLCELL_X4 FILLER_28_482 ();
 FILLCELL_X2 FILLER_28_486 ();
 FILLCELL_X1 FILLER_28_488 ();
 FILLCELL_X4 FILLER_28_493 ();
 FILLCELL_X8 FILLER_28_500 ();
 FILLCELL_X1 FILLER_28_508 ();
 FILLCELL_X4 FILLER_28_511 ();
 FILLCELL_X1 FILLER_28_515 ();
 FILLCELL_X4 FILLER_28_523 ();
 FILLCELL_X8 FILLER_28_532 ();
 FILLCELL_X1 FILLER_28_540 ();
 FILLCELL_X4 FILLER_28_544 ();
 FILLCELL_X4 FILLER_28_552 ();
 FILLCELL_X2 FILLER_28_556 ();
 FILLCELL_X1 FILLER_28_558 ();
 FILLCELL_X4 FILLER_28_563 ();
 FILLCELL_X4 FILLER_28_576 ();
 FILLCELL_X4 FILLER_28_585 ();
 FILLCELL_X2 FILLER_28_589 ();
 FILLCELL_X8 FILLER_28_595 ();
 FILLCELL_X8 FILLER_28_608 ();
 FILLCELL_X4 FILLER_28_616 ();
 FILLCELL_X4 FILLER_28_624 ();
 FILLCELL_X2 FILLER_28_628 ();
 FILLCELL_X1 FILLER_28_630 ();
 FILLCELL_X4 FILLER_28_632 ();
 FILLCELL_X2 FILLER_28_636 ();
 FILLCELL_X1 FILLER_28_638 ();
 FILLCELL_X8 FILLER_28_649 ();
 FILLCELL_X1 FILLER_28_657 ();
 FILLCELL_X4 FILLER_28_662 ();
 FILLCELL_X4 FILLER_28_670 ();
 FILLCELL_X4 FILLER_28_683 ();
 FILLCELL_X2 FILLER_28_687 ();
 FILLCELL_X4 FILLER_28_693 ();
 FILLCELL_X2 FILLER_28_697 ();
 FILLCELL_X4 FILLER_28_702 ();
 FILLCELL_X4 FILLER_28_710 ();
 FILLCELL_X4 FILLER_28_724 ();
 FILLCELL_X4 FILLER_28_730 ();
 FILLCELL_X8 FILLER_28_744 ();
 FILLCELL_X4 FILLER_28_752 ();
 FILLCELL_X2 FILLER_28_756 ();
 FILLCELL_X4 FILLER_28_761 ();
 FILLCELL_X4 FILLER_28_769 ();
 FILLCELL_X4 FILLER_28_782 ();
 FILLCELL_X2 FILLER_28_786 ();
 FILLCELL_X4 FILLER_28_791 ();
 FILLCELL_X4 FILLER_28_798 ();
 FILLCELL_X4 FILLER_28_805 ();
 FILLCELL_X4 FILLER_28_818 ();
 FILLCELL_X8 FILLER_28_824 ();
 FILLCELL_X8 FILLER_28_842 ();
 FILLCELL_X1 FILLER_28_850 ();
 FILLCELL_X4 FILLER_28_855 ();
 FILLCELL_X4 FILLER_28_869 ();
 FILLCELL_X4 FILLER_28_876 ();
 FILLCELL_X4 FILLER_28_887 ();
 FILLCELL_X1 FILLER_28_891 ();
 FILLCELL_X4 FILLER_28_895 ();
 FILLCELL_X4 FILLER_28_902 ();
 FILLCELL_X4 FILLER_28_910 ();
 FILLCELL_X4 FILLER_28_923 ();
 FILLCELL_X16 FILLER_28_931 ();
 FILLCELL_X4 FILLER_28_957 ();
 FILLCELL_X4 FILLER_28_971 ();
 FILLCELL_X1 FILLER_28_975 ();
 FILLCELL_X4 FILLER_28_980 ();
 FILLCELL_X4 FILLER_28_993 ();
 FILLCELL_X4 FILLER_28_1000 ();
 FILLCELL_X4 FILLER_28_1006 ();
 FILLCELL_X2 FILLER_28_1010 ();
 FILLCELL_X4 FILLER_28_1015 ();
 FILLCELL_X4 FILLER_28_1021 ();
 FILLCELL_X4 FILLER_28_1027 ();
 FILLCELL_X4 FILLER_28_1033 ();
 FILLCELL_X2 FILLER_28_1037 ();
 FILLCELL_X1 FILLER_28_1039 ();
 FILLCELL_X4 FILLER_28_1043 ();
 FILLCELL_X4 FILLER_28_1050 ();
 FILLCELL_X8 FILLER_28_1056 ();
 FILLCELL_X16 FILLER_28_1067 ();
 FILLCELL_X8 FILLER_28_1083 ();
 FILLCELL_X2 FILLER_28_1091 ();
 FILLCELL_X1 FILLER_28_1093 ();
 FILLCELL_X8 FILLER_28_1097 ();
 FILLCELL_X1 FILLER_28_1105 ();
 FILLCELL_X4 FILLER_28_1108 ();
 FILLCELL_X8 FILLER_28_1122 ();
 FILLCELL_X4 FILLER_28_1130 ();
 FILLCELL_X2 FILLER_28_1134 ();
 FILLCELL_X4 FILLER_28_1146 ();
 FILLCELL_X2 FILLER_28_1150 ();
 FILLCELL_X1 FILLER_28_1152 ();
 FILLCELL_X4 FILLER_28_1162 ();
 FILLCELL_X4 FILLER_28_1176 ();
 FILLCELL_X16 FILLER_28_1189 ();
 FILLCELL_X8 FILLER_28_1205 ();
 FILLCELL_X2 FILLER_28_1213 ();
 FILLCELL_X4 FILLER_28_1224 ();
 FILLCELL_X8 FILLER_28_1231 ();
 FILLCELL_X8 FILLER_28_1242 ();
 FILLCELL_X4 FILLER_28_1250 ();
 FILLCELL_X4 FILLER_28_1258 ();
 FILLCELL_X4 FILLER_28_1266 ();
 FILLCELL_X4 FILLER_28_1273 ();
 FILLCELL_X8 FILLER_28_1280 ();
 FILLCELL_X4 FILLER_28_1291 ();
 FILLCELL_X4 FILLER_28_1305 ();
 FILLCELL_X4 FILLER_28_1319 ();
 FILLCELL_X4 FILLER_28_1332 ();
 FILLCELL_X4 FILLER_28_1345 ();
 FILLCELL_X2 FILLER_28_1349 ();
 FILLCELL_X4 FILLER_28_1358 ();
 FILLCELL_X4 FILLER_28_1372 ();
 FILLCELL_X2 FILLER_28_1376 ();
 FILLCELL_X1 FILLER_28_1378 ();
 FILLCELL_X4 FILLER_28_1383 ();
 FILLCELL_X4 FILLER_28_1397 ();
 FILLCELL_X4 FILLER_28_1408 ();
 FILLCELL_X1 FILLER_28_1412 ();
 FILLCELL_X4 FILLER_28_1417 ();
 FILLCELL_X8 FILLER_28_1430 ();
 FILLCELL_X1 FILLER_28_1438 ();
 FILLCELL_X4 FILLER_28_1442 ();
 FILLCELL_X2 FILLER_28_1446 ();
 FILLCELL_X4 FILLER_28_1458 ();
 FILLCELL_X4 FILLER_28_1466 ();
 FILLCELL_X32 FILLER_28_1473 ();
 FILLCELL_X32 FILLER_28_1505 ();
 FILLCELL_X32 FILLER_28_1537 ();
 FILLCELL_X32 FILLER_28_1569 ();
 FILLCELL_X32 FILLER_28_1601 ();
 FILLCELL_X32 FILLER_28_1633 ();
 FILLCELL_X32 FILLER_28_1665 ();
 FILLCELL_X32 FILLER_28_1697 ();
 FILLCELL_X32 FILLER_28_1729 ();
 FILLCELL_X1 FILLER_28_1761 ();
 FILLCELL_X8 FILLER_29_1 ();
 FILLCELL_X4 FILLER_29_9 ();
 FILLCELL_X4 FILLER_29_17 ();
 FILLCELL_X4 FILLER_29_30 ();
 FILLCELL_X4 FILLER_29_38 ();
 FILLCELL_X4 FILLER_29_45 ();
 FILLCELL_X1 FILLER_29_49 ();
 FILLCELL_X4 FILLER_29_60 ();
 FILLCELL_X8 FILLER_29_67 ();
 FILLCELL_X1 FILLER_29_75 ();
 FILLCELL_X8 FILLER_29_80 ();
 FILLCELL_X1 FILLER_29_88 ();
 FILLCELL_X4 FILLER_29_98 ();
 FILLCELL_X4 FILLER_29_111 ();
 FILLCELL_X4 FILLER_29_125 ();
 FILLCELL_X1 FILLER_29_129 ();
 FILLCELL_X4 FILLER_29_139 ();
 FILLCELL_X4 FILLER_29_146 ();
 FILLCELL_X2 FILLER_29_150 ();
 FILLCELL_X1 FILLER_29_152 ();
 FILLCELL_X4 FILLER_29_160 ();
 FILLCELL_X8 FILLER_29_174 ();
 FILLCELL_X4 FILLER_29_182 ();
 FILLCELL_X4 FILLER_29_193 ();
 FILLCELL_X1 FILLER_29_197 ();
 FILLCELL_X4 FILLER_29_200 ();
 FILLCELL_X4 FILLER_29_213 ();
 FILLCELL_X1 FILLER_29_217 ();
 FILLCELL_X4 FILLER_29_221 ();
 FILLCELL_X4 FILLER_29_228 ();
 FILLCELL_X8 FILLER_29_235 ();
 FILLCELL_X4 FILLER_29_243 ();
 FILLCELL_X2 FILLER_29_247 ();
 FILLCELL_X4 FILLER_29_258 ();
 FILLCELL_X8 FILLER_29_271 ();
 FILLCELL_X2 FILLER_29_279 ();
 FILLCELL_X4 FILLER_29_285 ();
 FILLCELL_X4 FILLER_29_293 ();
 FILLCELL_X8 FILLER_29_300 ();
 FILLCELL_X4 FILLER_29_308 ();
 FILLCELL_X2 FILLER_29_312 ();
 FILLCELL_X8 FILLER_29_316 ();
 FILLCELL_X2 FILLER_29_324 ();
 FILLCELL_X1 FILLER_29_326 ();
 FILLCELL_X4 FILLER_29_336 ();
 FILLCELL_X16 FILLER_29_345 ();
 FILLCELL_X4 FILLER_29_361 ();
 FILLCELL_X4 FILLER_29_368 ();
 FILLCELL_X4 FILLER_29_382 ();
 FILLCELL_X2 FILLER_29_386 ();
 FILLCELL_X4 FILLER_29_398 ();
 FILLCELL_X1 FILLER_29_402 ();
 FILLCELL_X4 FILLER_29_410 ();
 FILLCELL_X2 FILLER_29_414 ();
 FILLCELL_X1 FILLER_29_416 ();
 FILLCELL_X16 FILLER_29_421 ();
 FILLCELL_X1 FILLER_29_437 ();
 FILLCELL_X4 FILLER_29_440 ();
 FILLCELL_X8 FILLER_29_450 ();
 FILLCELL_X2 FILLER_29_458 ();
 FILLCELL_X4 FILLER_29_464 ();
 FILLCELL_X4 FILLER_29_475 ();
 FILLCELL_X1 FILLER_29_479 ();
 FILLCELL_X4 FILLER_29_486 ();
 FILLCELL_X4 FILLER_29_500 ();
 FILLCELL_X4 FILLER_29_507 ();
 FILLCELL_X2 FILLER_29_511 ();
 FILLCELL_X8 FILLER_29_522 ();
 FILLCELL_X1 FILLER_29_530 ();
 FILLCELL_X8 FILLER_29_538 ();
 FILLCELL_X8 FILLER_29_556 ();
 FILLCELL_X1 FILLER_29_564 ();
 FILLCELL_X4 FILLER_29_574 ();
 FILLCELL_X4 FILLER_29_581 ();
 FILLCELL_X4 FILLER_29_589 ();
 FILLCELL_X8 FILLER_29_602 ();
 FILLCELL_X1 FILLER_29_610 ();
 FILLCELL_X4 FILLER_29_614 ();
 FILLCELL_X4 FILLER_29_627 ();
 FILLCELL_X8 FILLER_29_635 ();
 FILLCELL_X2 FILLER_29_643 ();
 FILLCELL_X1 FILLER_29_645 ();
 FILLCELL_X4 FILLER_29_651 ();
 FILLCELL_X4 FILLER_29_659 ();
 FILLCELL_X4 FILLER_29_672 ();
 FILLCELL_X4 FILLER_29_679 ();
 FILLCELL_X2 FILLER_29_683 ();
 FILLCELL_X4 FILLER_29_689 ();
 FILLCELL_X4 FILLER_29_702 ();
 FILLCELL_X1 FILLER_29_706 ();
 FILLCELL_X4 FILLER_29_710 ();
 FILLCELL_X4 FILLER_29_717 ();
 FILLCELL_X8 FILLER_29_725 ();
 FILLCELL_X4 FILLER_29_737 ();
 FILLCELL_X8 FILLER_29_751 ();
 FILLCELL_X1 FILLER_29_759 ();
 FILLCELL_X4 FILLER_29_763 ();
 FILLCELL_X8 FILLER_29_776 ();
 FILLCELL_X2 FILLER_29_784 ();
 FILLCELL_X4 FILLER_29_789 ();
 FILLCELL_X8 FILLER_29_798 ();
 FILLCELL_X1 FILLER_29_806 ();
 FILLCELL_X4 FILLER_29_813 ();
 FILLCELL_X4 FILLER_29_821 ();
 FILLCELL_X2 FILLER_29_825 ();
 FILLCELL_X1 FILLER_29_827 ();
 FILLCELL_X4 FILLER_29_831 ();
 FILLCELL_X4 FILLER_29_844 ();
 FILLCELL_X1 FILLER_29_848 ();
 FILLCELL_X32 FILLER_29_853 ();
 FILLCELL_X8 FILLER_29_885 ();
 FILLCELL_X2 FILLER_29_893 ();
 FILLCELL_X1 FILLER_29_895 ();
 FILLCELL_X8 FILLER_29_903 ();
 FILLCELL_X4 FILLER_29_914 ();
 FILLCELL_X2 FILLER_29_918 ();
 FILLCELL_X1 FILLER_29_920 ();
 FILLCELL_X4 FILLER_29_924 ();
 FILLCELL_X4 FILLER_29_937 ();
 FILLCELL_X1 FILLER_29_941 ();
 FILLCELL_X4 FILLER_29_944 ();
 FILLCELL_X4 FILLER_29_951 ();
 FILLCELL_X4 FILLER_29_959 ();
 FILLCELL_X8 FILLER_29_965 ();
 FILLCELL_X4 FILLER_29_973 ();
 FILLCELL_X1 FILLER_29_977 ();
 FILLCELL_X4 FILLER_29_987 ();
 FILLCELL_X4 FILLER_29_995 ();
 FILLCELL_X4 FILLER_29_1002 ();
 FILLCELL_X4 FILLER_29_1009 ();
 FILLCELL_X2 FILLER_29_1013 ();
 FILLCELL_X4 FILLER_29_1022 ();
 FILLCELL_X2 FILLER_29_1026 ();
 FILLCELL_X1 FILLER_29_1028 ();
 FILLCELL_X4 FILLER_29_1038 ();
 FILLCELL_X4 FILLER_29_1045 ();
 FILLCELL_X2 FILLER_29_1049 ();
 FILLCELL_X4 FILLER_29_1060 ();
 FILLCELL_X16 FILLER_29_1066 ();
 FILLCELL_X4 FILLER_29_1091 ();
 FILLCELL_X4 FILLER_29_1099 ();
 FILLCELL_X1 FILLER_29_1103 ();
 FILLCELL_X4 FILLER_29_1108 ();
 FILLCELL_X4 FILLER_29_1122 ();
 FILLCELL_X4 FILLER_29_1129 ();
 FILLCELL_X1 FILLER_29_1133 ();
 FILLCELL_X4 FILLER_29_1137 ();
 FILLCELL_X16 FILLER_29_1148 ();
 FILLCELL_X4 FILLER_29_1164 ();
 FILLCELL_X4 FILLER_29_1172 ();
 FILLCELL_X8 FILLER_29_1179 ();
 FILLCELL_X2 FILLER_29_1187 ();
 FILLCELL_X4 FILLER_29_1198 ();
 FILLCELL_X4 FILLER_29_1205 ();
 FILLCELL_X4 FILLER_29_1212 ();
 FILLCELL_X4 FILLER_29_1225 ();
 FILLCELL_X4 FILLER_29_1238 ();
 FILLCELL_X1 FILLER_29_1242 ();
 FILLCELL_X8 FILLER_29_1253 ();
 FILLCELL_X2 FILLER_29_1261 ();
 FILLCELL_X4 FILLER_29_1264 ();
 FILLCELL_X4 FILLER_29_1277 ();
 FILLCELL_X8 FILLER_29_1284 ();
 FILLCELL_X4 FILLER_29_1292 ();
 FILLCELL_X2 FILLER_29_1296 ();
 FILLCELL_X1 FILLER_29_1298 ();
 FILLCELL_X8 FILLER_29_1301 ();
 FILLCELL_X8 FILLER_29_1312 ();
 FILLCELL_X4 FILLER_29_1320 ();
 FILLCELL_X4 FILLER_29_1327 ();
 FILLCELL_X2 FILLER_29_1331 ();
 FILLCELL_X1 FILLER_29_1333 ();
 FILLCELL_X8 FILLER_29_1337 ();
 FILLCELL_X4 FILLER_29_1345 ();
 FILLCELL_X2 FILLER_29_1349 ();
 FILLCELL_X1 FILLER_29_1351 ();
 FILLCELL_X4 FILLER_29_1356 ();
 FILLCELL_X2 FILLER_29_1360 ();
 FILLCELL_X1 FILLER_29_1362 ();
 FILLCELL_X4 FILLER_29_1366 ();
 FILLCELL_X16 FILLER_29_1372 ();
 FILLCELL_X4 FILLER_29_1388 ();
 FILLCELL_X2 FILLER_29_1392 ();
 FILLCELL_X1 FILLER_29_1394 ();
 FILLCELL_X4 FILLER_29_1398 ();
 FILLCELL_X4 FILLER_29_1411 ();
 FILLCELL_X4 FILLER_29_1418 ();
 FILLCELL_X4 FILLER_29_1425 ();
 FILLCELL_X4 FILLER_29_1433 ();
 FILLCELL_X1 FILLER_29_1437 ();
 FILLCELL_X4 FILLER_29_1448 ();
 FILLCELL_X2 FILLER_29_1452 ();
 FILLCELL_X8 FILLER_29_1458 ();
 FILLCELL_X32 FILLER_29_1472 ();
 FILLCELL_X8 FILLER_29_1504 ();
 FILLCELL_X4 FILLER_29_1512 ();
 FILLCELL_X4 FILLER_29_1520 ();
 FILLCELL_X32 FILLER_29_1543 ();
 FILLCELL_X32 FILLER_29_1575 ();
 FILLCELL_X32 FILLER_29_1607 ();
 FILLCELL_X32 FILLER_29_1639 ();
 FILLCELL_X32 FILLER_29_1671 ();
 FILLCELL_X32 FILLER_29_1703 ();
 FILLCELL_X16 FILLER_29_1735 ();
 FILLCELL_X8 FILLER_29_1751 ();
 FILLCELL_X2 FILLER_29_1759 ();
 FILLCELL_X1 FILLER_29_1761 ();
 FILLCELL_X8 FILLER_30_1 ();
 FILLCELL_X4 FILLER_30_9 ();
 FILLCELL_X2 FILLER_30_13 ();
 FILLCELL_X4 FILLER_30_19 ();
 FILLCELL_X4 FILLER_30_27 ();
 FILLCELL_X8 FILLER_30_34 ();
 FILLCELL_X4 FILLER_30_42 ();
 FILLCELL_X8 FILLER_30_55 ();
 FILLCELL_X4 FILLER_30_63 ();
 FILLCELL_X2 FILLER_30_67 ();
 FILLCELL_X16 FILLER_30_71 ();
 FILLCELL_X8 FILLER_30_87 ();
 FILLCELL_X4 FILLER_30_95 ();
 FILLCELL_X4 FILLER_30_102 ();
 FILLCELL_X4 FILLER_30_109 ();
 FILLCELL_X2 FILLER_30_113 ();
 FILLCELL_X8 FILLER_30_119 ();
 FILLCELL_X2 FILLER_30_127 ();
 FILLCELL_X4 FILLER_30_138 ();
 FILLCELL_X4 FILLER_30_152 ();
 FILLCELL_X2 FILLER_30_156 ();
 FILLCELL_X1 FILLER_30_158 ();
 FILLCELL_X8 FILLER_30_169 ();
 FILLCELL_X4 FILLER_30_181 ();
 FILLCELL_X4 FILLER_30_195 ();
 FILLCELL_X8 FILLER_30_202 ();
 FILLCELL_X2 FILLER_30_210 ();
 FILLCELL_X1 FILLER_30_212 ();
 FILLCELL_X4 FILLER_30_216 ();
 FILLCELL_X4 FILLER_30_230 ();
 FILLCELL_X4 FILLER_30_238 ();
 FILLCELL_X2 FILLER_30_242 ();
 FILLCELL_X1 FILLER_30_244 ();
 FILLCELL_X4 FILLER_30_249 ();
 FILLCELL_X4 FILLER_30_256 ();
 FILLCELL_X1 FILLER_30_260 ();
 FILLCELL_X4 FILLER_30_264 ();
 FILLCELL_X2 FILLER_30_268 ();
 FILLCELL_X4 FILLER_30_273 ();
 FILLCELL_X4 FILLER_30_281 ();
 FILLCELL_X8 FILLER_30_294 ();
 FILLCELL_X4 FILLER_30_302 ();
 FILLCELL_X4 FILLER_30_310 ();
 FILLCELL_X1 FILLER_30_314 ();
 FILLCELL_X4 FILLER_30_325 ();
 FILLCELL_X2 FILLER_30_329 ();
 FILLCELL_X4 FILLER_30_334 ();
 FILLCELL_X8 FILLER_30_347 ();
 FILLCELL_X4 FILLER_30_355 ();
 FILLCELL_X2 FILLER_30_359 ();
 FILLCELL_X1 FILLER_30_361 ();
 FILLCELL_X16 FILLER_30_364 ();
 FILLCELL_X8 FILLER_30_380 ();
 FILLCELL_X4 FILLER_30_388 ();
 FILLCELL_X4 FILLER_30_395 ();
 FILLCELL_X4 FILLER_30_402 ();
 FILLCELL_X2 FILLER_30_406 ();
 FILLCELL_X1 FILLER_30_408 ();
 FILLCELL_X4 FILLER_30_412 ();
 FILLCELL_X8 FILLER_30_426 ();
 FILLCELL_X4 FILLER_30_434 ();
 FILLCELL_X8 FILLER_30_445 ();
 FILLCELL_X2 FILLER_30_453 ();
 FILLCELL_X1 FILLER_30_455 ();
 FILLCELL_X4 FILLER_30_465 ();
 FILLCELL_X8 FILLER_30_473 ();
 FILLCELL_X4 FILLER_30_488 ();
 FILLCELL_X8 FILLER_30_501 ();
 FILLCELL_X2 FILLER_30_509 ();
 FILLCELL_X1 FILLER_30_511 ();
 FILLCELL_X4 FILLER_30_515 ();
 FILLCELL_X4 FILLER_30_523 ();
 FILLCELL_X16 FILLER_30_546 ();
 FILLCELL_X8 FILLER_30_562 ();
 FILLCELL_X1 FILLER_30_570 ();
 FILLCELL_X8 FILLER_30_575 ();
 FILLCELL_X4 FILLER_30_583 ();
 FILLCELL_X2 FILLER_30_587 ();
 FILLCELL_X1 FILLER_30_589 ();
 FILLCELL_X4 FILLER_30_599 ();
 FILLCELL_X4 FILLER_30_607 ();
 FILLCELL_X8 FILLER_30_614 ();
 FILLCELL_X2 FILLER_30_622 ();
 FILLCELL_X4 FILLER_30_627 ();
 FILLCELL_X4 FILLER_30_632 ();
 FILLCELL_X4 FILLER_30_646 ();
 FILLCELL_X1 FILLER_30_650 ();
 FILLCELL_X16 FILLER_30_653 ();
 FILLCELL_X2 FILLER_30_669 ();
 FILLCELL_X1 FILLER_30_671 ();
 FILLCELL_X4 FILLER_30_675 ();
 FILLCELL_X2 FILLER_30_679 ();
 FILLCELL_X1 FILLER_30_681 ();
 FILLCELL_X4 FILLER_30_685 ();
 FILLCELL_X8 FILLER_30_692 ();
 FILLCELL_X4 FILLER_30_704 ();
 FILLCELL_X8 FILLER_30_717 ();
 FILLCELL_X2 FILLER_30_725 ();
 FILLCELL_X4 FILLER_30_737 ();
 FILLCELL_X8 FILLER_30_743 ();
 FILLCELL_X4 FILLER_30_751 ();
 FILLCELL_X2 FILLER_30_755 ();
 FILLCELL_X1 FILLER_30_757 ();
 FILLCELL_X4 FILLER_30_761 ();
 FILLCELL_X4 FILLER_30_769 ();
 FILLCELL_X8 FILLER_30_777 ();
 FILLCELL_X1 FILLER_30_785 ();
 FILLCELL_X4 FILLER_30_793 ();
 FILLCELL_X4 FILLER_30_803 ();
 FILLCELL_X1 FILLER_30_807 ();
 FILLCELL_X4 FILLER_30_814 ();
 FILLCELL_X4 FILLER_30_821 ();
 FILLCELL_X1 FILLER_30_825 ();
 FILLCELL_X4 FILLER_30_829 ();
 FILLCELL_X4 FILLER_30_836 ();
 FILLCELL_X1 FILLER_30_840 ();
 FILLCELL_X4 FILLER_30_845 ();
 FILLCELL_X16 FILLER_30_858 ();
 FILLCELL_X8 FILLER_30_874 ();
 FILLCELL_X1 FILLER_30_882 ();
 FILLCELL_X4 FILLER_30_885 ();
 FILLCELL_X8 FILLER_30_899 ();
 FILLCELL_X1 FILLER_30_907 ();
 FILLCELL_X8 FILLER_30_927 ();
 FILLCELL_X2 FILLER_30_935 ();
 FILLCELL_X1 FILLER_30_937 ();
 FILLCELL_X4 FILLER_30_941 ();
 FILLCELL_X8 FILLER_30_948 ();
 FILLCELL_X4 FILLER_30_966 ();
 FILLCELL_X16 FILLER_30_973 ();
 FILLCELL_X4 FILLER_30_989 ();
 FILLCELL_X2 FILLER_30_993 ();
 FILLCELL_X4 FILLER_30_997 ();
 FILLCELL_X4 FILLER_30_1003 ();
 FILLCELL_X4 FILLER_30_1009 ();
 FILLCELL_X4 FILLER_30_1023 ();
 FILLCELL_X2 FILLER_30_1027 ();
 FILLCELL_X1 FILLER_30_1029 ();
 FILLCELL_X4 FILLER_30_1039 ();
 FILLCELL_X4 FILLER_30_1048 ();
 FILLCELL_X1 FILLER_30_1052 ();
 FILLCELL_X4 FILLER_30_1062 ();
 FILLCELL_X4 FILLER_30_1069 ();
 FILLCELL_X8 FILLER_30_1076 ();
 FILLCELL_X2 FILLER_30_1084 ();
 FILLCELL_X1 FILLER_30_1086 ();
 FILLCELL_X4 FILLER_30_1096 ();
 FILLCELL_X4 FILLER_30_1103 ();
 FILLCELL_X4 FILLER_30_1110 ();
 FILLCELL_X8 FILLER_30_1121 ();
 FILLCELL_X4 FILLER_30_1129 ();
 FILLCELL_X2 FILLER_30_1133 ();
 FILLCELL_X1 FILLER_30_1135 ();
 FILLCELL_X8 FILLER_30_1146 ();
 FILLCELL_X1 FILLER_30_1154 ();
 FILLCELL_X4 FILLER_30_1164 ();
 FILLCELL_X8 FILLER_30_1171 ();
 FILLCELL_X4 FILLER_30_1179 ();
 FILLCELL_X4 FILLER_30_1186 ();
 FILLCELL_X4 FILLER_30_1199 ();
 FILLCELL_X1 FILLER_30_1203 ();
 FILLCELL_X4 FILLER_30_1214 ();
 FILLCELL_X1 FILLER_30_1218 ();
 FILLCELL_X4 FILLER_30_1222 ();
 FILLCELL_X4 FILLER_30_1229 ();
 FILLCELL_X2 FILLER_30_1233 ();
 FILLCELL_X4 FILLER_30_1238 ();
 FILLCELL_X2 FILLER_30_1242 ();
 FILLCELL_X1 FILLER_30_1244 ();
 FILLCELL_X8 FILLER_30_1248 ();
 FILLCELL_X4 FILLER_30_1256 ();
 FILLCELL_X1 FILLER_30_1260 ();
 FILLCELL_X4 FILLER_30_1265 ();
 FILLCELL_X8 FILLER_30_1278 ();
 FILLCELL_X4 FILLER_30_1293 ();
 FILLCELL_X16 FILLER_30_1299 ();
 FILLCELL_X1 FILLER_30_1315 ();
 FILLCELL_X4 FILLER_30_1319 ();
 FILLCELL_X8 FILLER_30_1332 ();
 FILLCELL_X4 FILLER_30_1347 ();
 FILLCELL_X4 FILLER_30_1361 ();
 FILLCELL_X4 FILLER_30_1375 ();
 FILLCELL_X2 FILLER_30_1379 ();
 FILLCELL_X16 FILLER_30_1390 ();
 FILLCELL_X8 FILLER_30_1406 ();
 FILLCELL_X4 FILLER_30_1414 ();
 FILLCELL_X1 FILLER_30_1418 ();
 FILLCELL_X4 FILLER_30_1429 ();
 FILLCELL_X8 FILLER_30_1435 ();
 FILLCELL_X4 FILLER_30_1443 ();
 FILLCELL_X4 FILLER_30_1451 ();
 FILLCELL_X4 FILLER_30_1462 ();
 FILLCELL_X32 FILLER_30_1472 ();
 FILLCELL_X32 FILLER_30_1504 ();
 FILLCELL_X32 FILLER_30_1536 ();
 FILLCELL_X32 FILLER_30_1568 ();
 FILLCELL_X32 FILLER_30_1600 ();
 FILLCELL_X32 FILLER_30_1632 ();
 FILLCELL_X32 FILLER_30_1664 ();
 FILLCELL_X32 FILLER_30_1696 ();
 FILLCELL_X16 FILLER_30_1728 ();
 FILLCELL_X8 FILLER_30_1744 ();
 FILLCELL_X2 FILLER_30_1752 ();
 FILLCELL_X1 FILLER_30_1754 ();
 FILLCELL_X4 FILLER_30_1758 ();
 FILLCELL_X8 FILLER_31_1 ();
 FILLCELL_X1 FILLER_31_9 ();
 FILLCELL_X4 FILLER_31_19 ();
 FILLCELL_X2 FILLER_31_23 ();
 FILLCELL_X8 FILLER_31_29 ();
 FILLCELL_X4 FILLER_31_37 ();
 FILLCELL_X1 FILLER_31_41 ();
 FILLCELL_X4 FILLER_31_45 ();
 FILLCELL_X4 FILLER_31_52 ();
 FILLCELL_X1 FILLER_31_56 ();
 FILLCELL_X4 FILLER_31_67 ();
 FILLCELL_X4 FILLER_31_73 ();
 FILLCELL_X4 FILLER_31_87 ();
 FILLCELL_X16 FILLER_31_98 ();
 FILLCELL_X8 FILLER_31_114 ();
 FILLCELL_X4 FILLER_31_122 ();
 FILLCELL_X2 FILLER_31_126 ();
 FILLCELL_X4 FILLER_31_135 ();
 FILLCELL_X8 FILLER_31_142 ();
 FILLCELL_X4 FILLER_31_150 ();
 FILLCELL_X8 FILLER_31_157 ();
 FILLCELL_X4 FILLER_31_165 ();
 FILLCELL_X4 FILLER_31_171 ();
 FILLCELL_X4 FILLER_31_185 ();
 FILLCELL_X4 FILLER_31_192 ();
 FILLCELL_X4 FILLER_31_199 ();
 FILLCELL_X2 FILLER_31_203 ();
 FILLCELL_X1 FILLER_31_205 ();
 FILLCELL_X16 FILLER_31_213 ();
 FILLCELL_X2 FILLER_31_229 ();
 FILLCELL_X4 FILLER_31_240 ();
 FILLCELL_X4 FILLER_31_253 ();
 FILLCELL_X8 FILLER_31_261 ();
 FILLCELL_X1 FILLER_31_269 ();
 FILLCELL_X8 FILLER_31_274 ();
 FILLCELL_X2 FILLER_31_282 ();
 FILLCELL_X4 FILLER_31_287 ();
 FILLCELL_X4 FILLER_31_296 ();
 FILLCELL_X4 FILLER_31_303 ();
 FILLCELL_X4 FILLER_31_317 ();
 FILLCELL_X4 FILLER_31_328 ();
 FILLCELL_X8 FILLER_31_342 ();
 FILLCELL_X4 FILLER_31_360 ();
 FILLCELL_X8 FILLER_31_374 ();
 FILLCELL_X2 FILLER_31_382 ();
 FILLCELL_X1 FILLER_31_384 ();
 FILLCELL_X4 FILLER_31_389 ();
 FILLCELL_X2 FILLER_31_393 ();
 FILLCELL_X4 FILLER_31_399 ();
 FILLCELL_X4 FILLER_31_412 ();
 FILLCELL_X2 FILLER_31_416 ();
 FILLCELL_X8 FILLER_31_422 ();
 FILLCELL_X2 FILLER_31_430 ();
 FILLCELL_X1 FILLER_31_432 ();
 FILLCELL_X8 FILLER_31_458 ();
 FILLCELL_X4 FILLER_31_476 ();
 FILLCELL_X1 FILLER_31_480 ();
 FILLCELL_X4 FILLER_31_483 ();
 FILLCELL_X16 FILLER_31_497 ();
 FILLCELL_X4 FILLER_31_523 ();
 FILLCELL_X4 FILLER_31_530 ();
 FILLCELL_X16 FILLER_31_536 ();
 FILLCELL_X2 FILLER_31_552 ();
 FILLCELL_X1 FILLER_31_554 ();
 FILLCELL_X4 FILLER_31_558 ();
 FILLCELL_X8 FILLER_31_569 ();
 FILLCELL_X8 FILLER_31_587 ();
 FILLCELL_X4 FILLER_31_599 ();
 FILLCELL_X16 FILLER_31_612 ();
 FILLCELL_X4 FILLER_31_628 ();
 FILLCELL_X2 FILLER_31_632 ();
 FILLCELL_X8 FILLER_31_637 ();
 FILLCELL_X2 FILLER_31_645 ();
 FILLCELL_X4 FILLER_31_649 ();
 FILLCELL_X4 FILLER_31_655 ();
 FILLCELL_X4 FILLER_31_666 ();
 FILLCELL_X4 FILLER_31_680 ();
 FILLCELL_X4 FILLER_31_688 ();
 FILLCELL_X2 FILLER_31_692 ();
 FILLCELL_X8 FILLER_31_704 ();
 FILLCELL_X4 FILLER_31_712 ();
 FILLCELL_X1 FILLER_31_716 ();
 FILLCELL_X8 FILLER_31_720 ();
 FILLCELL_X8 FILLER_31_747 ();
 FILLCELL_X4 FILLER_31_755 ();
 FILLCELL_X1 FILLER_31_759 ();
 FILLCELL_X4 FILLER_31_764 ();
 FILLCELL_X8 FILLER_31_773 ();
 FILLCELL_X2 FILLER_31_781 ();
 FILLCELL_X8 FILLER_31_789 ();
 FILLCELL_X4 FILLER_31_801 ();
 FILLCELL_X8 FILLER_31_810 ();
 FILLCELL_X4 FILLER_31_822 ();
 FILLCELL_X8 FILLER_31_835 ();
 FILLCELL_X4 FILLER_31_843 ();
 FILLCELL_X1 FILLER_31_847 ();
 FILLCELL_X16 FILLER_31_852 ();
 FILLCELL_X1 FILLER_31_868 ();
 FILLCELL_X4 FILLER_31_873 ();
 FILLCELL_X4 FILLER_31_881 ();
 FILLCELL_X4 FILLER_31_889 ();
 FILLCELL_X4 FILLER_31_903 ();
 FILLCELL_X8 FILLER_31_910 ();
 FILLCELL_X4 FILLER_31_918 ();
 FILLCELL_X2 FILLER_31_922 ();
 FILLCELL_X4 FILLER_31_926 ();
 FILLCELL_X4 FILLER_31_939 ();
 FILLCELL_X4 FILLER_31_952 ();
 FILLCELL_X4 FILLER_31_963 ();
 FILLCELL_X4 FILLER_31_971 ();
 FILLCELL_X4 FILLER_31_979 ();
 FILLCELL_X2 FILLER_31_983 ();
 FILLCELL_X4 FILLER_31_992 ();
 FILLCELL_X4 FILLER_31_998 ();
 FILLCELL_X8 FILLER_31_1004 ();
 FILLCELL_X4 FILLER_31_1022 ();
 FILLCELL_X8 FILLER_31_1029 ();
 FILLCELL_X1 FILLER_31_1037 ();
 FILLCELL_X4 FILLER_31_1048 ();
 FILLCELL_X4 FILLER_31_1055 ();
 FILLCELL_X2 FILLER_31_1059 ();
 FILLCELL_X1 FILLER_31_1061 ();
 FILLCELL_X4 FILLER_31_1072 ();
 FILLCELL_X4 FILLER_31_1080 ();
 FILLCELL_X2 FILLER_31_1084 ();
 FILLCELL_X1 FILLER_31_1086 ();
 FILLCELL_X4 FILLER_31_1091 ();
 FILLCELL_X4 FILLER_31_1099 ();
 FILLCELL_X8 FILLER_31_1106 ();
 FILLCELL_X4 FILLER_31_1117 ();
 FILLCELL_X8 FILLER_31_1124 ();
 FILLCELL_X2 FILLER_31_1132 ();
 FILLCELL_X4 FILLER_31_1137 ();
 FILLCELL_X8 FILLER_31_1143 ();
 FILLCELL_X4 FILLER_31_1158 ();
 FILLCELL_X4 FILLER_31_1165 ();
 FILLCELL_X4 FILLER_31_1172 ();
 FILLCELL_X4 FILLER_31_1179 ();
 FILLCELL_X2 FILLER_31_1183 ();
 FILLCELL_X4 FILLER_31_1187 ();
 FILLCELL_X8 FILLER_31_1196 ();
 FILLCELL_X4 FILLER_31_1211 ();
 FILLCELL_X4 FILLER_31_1218 ();
 FILLCELL_X1 FILLER_31_1222 ();
 FILLCELL_X4 FILLER_31_1232 ();
 FILLCELL_X4 FILLER_31_1239 ();
 FILLCELL_X8 FILLER_31_1250 ();
 FILLCELL_X4 FILLER_31_1258 ();
 FILLCELL_X1 FILLER_31_1262 ();
 FILLCELL_X8 FILLER_31_1264 ();
 FILLCELL_X1 FILLER_31_1272 ();
 FILLCELL_X4 FILLER_31_1283 ();
 FILLCELL_X4 FILLER_31_1297 ();
 FILLCELL_X8 FILLER_31_1311 ();
 FILLCELL_X4 FILLER_31_1319 ();
 FILLCELL_X4 FILLER_31_1332 ();
 FILLCELL_X2 FILLER_31_1336 ();
 FILLCELL_X1 FILLER_31_1338 ();
 FILLCELL_X4 FILLER_31_1349 ();
 FILLCELL_X16 FILLER_31_1356 ();
 FILLCELL_X4 FILLER_31_1372 ();
 FILLCELL_X4 FILLER_31_1380 ();
 FILLCELL_X4 FILLER_31_1388 ();
 FILLCELL_X16 FILLER_31_1395 ();
 FILLCELL_X4 FILLER_31_1411 ();
 FILLCELL_X8 FILLER_31_1422 ();
 FILLCELL_X32 FILLER_31_1439 ();
 FILLCELL_X32 FILLER_31_1471 ();
 FILLCELL_X32 FILLER_31_1503 ();
 FILLCELL_X32 FILLER_31_1535 ();
 FILLCELL_X32 FILLER_31_1567 ();
 FILLCELL_X32 FILLER_31_1599 ();
 FILLCELL_X32 FILLER_31_1631 ();
 FILLCELL_X32 FILLER_31_1663 ();
 FILLCELL_X32 FILLER_31_1695 ();
 FILLCELL_X32 FILLER_31_1727 ();
 FILLCELL_X2 FILLER_31_1759 ();
 FILLCELL_X1 FILLER_31_1761 ();
 FILLCELL_X8 FILLER_32_1 ();
 FILLCELL_X2 FILLER_32_9 ();
 FILLCELL_X4 FILLER_32_14 ();
 FILLCELL_X4 FILLER_32_27 ();
 FILLCELL_X4 FILLER_32_35 ();
 FILLCELL_X2 FILLER_32_39 ();
 FILLCELL_X16 FILLER_32_44 ();
 FILLCELL_X1 FILLER_32_60 ();
 FILLCELL_X8 FILLER_32_68 ();
 FILLCELL_X4 FILLER_32_76 ();
 FILLCELL_X1 FILLER_32_80 ();
 FILLCELL_X4 FILLER_32_91 ();
 FILLCELL_X4 FILLER_32_105 ();
 FILLCELL_X8 FILLER_32_111 ();
 FILLCELL_X1 FILLER_32_119 ();
 FILLCELL_X4 FILLER_32_122 ();
 FILLCELL_X16 FILLER_32_136 ();
 FILLCELL_X1 FILLER_32_152 ();
 FILLCELL_X4 FILLER_32_156 ();
 FILLCELL_X1 FILLER_32_160 ();
 FILLCELL_X8 FILLER_32_164 ();
 FILLCELL_X8 FILLER_32_181 ();
 FILLCELL_X1 FILLER_32_189 ();
 FILLCELL_X4 FILLER_32_200 ();
 FILLCELL_X4 FILLER_32_206 ();
 FILLCELL_X8 FILLER_32_229 ();
 FILLCELL_X4 FILLER_32_237 ();
 FILLCELL_X4 FILLER_32_245 ();
 FILLCELL_X8 FILLER_32_252 ();
 FILLCELL_X2 FILLER_32_260 ();
 FILLCELL_X1 FILLER_32_262 ();
 FILLCELL_X4 FILLER_32_267 ();
 FILLCELL_X4 FILLER_32_280 ();
 FILLCELL_X16 FILLER_32_289 ();
 FILLCELL_X1 FILLER_32_305 ();
 FILLCELL_X4 FILLER_32_309 ();
 FILLCELL_X16 FILLER_32_316 ();
 FILLCELL_X8 FILLER_32_332 ();
 FILLCELL_X4 FILLER_32_340 ();
 FILLCELL_X2 FILLER_32_344 ();
 FILLCELL_X4 FILLER_32_350 ();
 FILLCELL_X2 FILLER_32_354 ();
 FILLCELL_X4 FILLER_32_363 ();
 FILLCELL_X4 FILLER_32_370 ();
 FILLCELL_X2 FILLER_32_374 ();
 FILLCELL_X4 FILLER_32_385 ();
 FILLCELL_X4 FILLER_32_398 ();
 FILLCELL_X8 FILLER_32_405 ();
 FILLCELL_X4 FILLER_32_413 ();
 FILLCELL_X2 FILLER_32_417 ();
 FILLCELL_X16 FILLER_32_424 ();
 FILLCELL_X2 FILLER_32_440 ();
 FILLCELL_X4 FILLER_32_445 ();
 FILLCELL_X4 FILLER_32_456 ();
 FILLCELL_X32 FILLER_32_463 ();
 FILLCELL_X2 FILLER_32_495 ();
 FILLCELL_X1 FILLER_32_497 ();
 FILLCELL_X4 FILLER_32_507 ();
 FILLCELL_X1 FILLER_32_511 ();
 FILLCELL_X4 FILLER_32_521 ();
 FILLCELL_X8 FILLER_32_535 ();
 FILLCELL_X4 FILLER_32_543 ();
 FILLCELL_X1 FILLER_32_547 ();
 FILLCELL_X4 FILLER_32_558 ();
 FILLCELL_X4 FILLER_32_567 ();
 FILLCELL_X4 FILLER_32_573 ();
 FILLCELL_X2 FILLER_32_577 ();
 FILLCELL_X1 FILLER_32_579 ();
 FILLCELL_X4 FILLER_32_587 ();
 FILLCELL_X8 FILLER_32_594 ();
 FILLCELL_X4 FILLER_32_602 ();
 FILLCELL_X2 FILLER_32_606 ();
 FILLCELL_X4 FILLER_32_627 ();
 FILLCELL_X8 FILLER_32_632 ();
 FILLCELL_X4 FILLER_32_650 ();
 FILLCELL_X2 FILLER_32_654 ();
 FILLCELL_X1 FILLER_32_656 ();
 FILLCELL_X8 FILLER_32_676 ();
 FILLCELL_X4 FILLER_32_684 ();
 FILLCELL_X2 FILLER_32_688 ();
 FILLCELL_X1 FILLER_32_690 ();
 FILLCELL_X16 FILLER_32_695 ();
 FILLCELL_X8 FILLER_32_711 ();
 FILLCELL_X4 FILLER_32_719 ();
 FILLCELL_X2 FILLER_32_723 ();
 FILLCELL_X1 FILLER_32_725 ();
 FILLCELL_X4 FILLER_32_730 ();
 FILLCELL_X4 FILLER_32_753 ();
 FILLCELL_X4 FILLER_32_776 ();
 FILLCELL_X1 FILLER_32_780 ();
 FILLCELL_X8 FILLER_32_784 ();
 FILLCELL_X4 FILLER_32_792 ();
 FILLCELL_X4 FILLER_32_800 ();
 FILLCELL_X4 FILLER_32_811 ();
 FILLCELL_X4 FILLER_32_819 ();
 FILLCELL_X2 FILLER_32_823 ();
 FILLCELL_X1 FILLER_32_825 ();
 FILLCELL_X4 FILLER_32_829 ();
 FILLCELL_X1 FILLER_32_833 ();
 FILLCELL_X4 FILLER_32_837 ();
 FILLCELL_X4 FILLER_32_845 ();
 FILLCELL_X8 FILLER_32_858 ();
 FILLCELL_X4 FILLER_32_869 ();
 FILLCELL_X4 FILLER_32_882 ();
 FILLCELL_X16 FILLER_32_890 ();
 FILLCELL_X8 FILLER_32_906 ();
 FILLCELL_X4 FILLER_32_914 ();
 FILLCELL_X1 FILLER_32_918 ();
 FILLCELL_X16 FILLER_32_929 ();
 FILLCELL_X4 FILLER_32_945 ();
 FILLCELL_X4 FILLER_32_959 ();
 FILLCELL_X8 FILLER_32_965 ();
 FILLCELL_X4 FILLER_32_982 ();
 FILLCELL_X4 FILLER_32_996 ();
 FILLCELL_X4 FILLER_32_1006 ();
 FILLCELL_X4 FILLER_32_1013 ();
 FILLCELL_X4 FILLER_32_1020 ();
 FILLCELL_X1 FILLER_32_1024 ();
 FILLCELL_X4 FILLER_32_1029 ();
 FILLCELL_X2 FILLER_32_1033 ();
 FILLCELL_X8 FILLER_32_1044 ();
 FILLCELL_X1 FILLER_32_1052 ();
 FILLCELL_X4 FILLER_32_1060 ();
 FILLCELL_X4 FILLER_32_1069 ();
 FILLCELL_X4 FILLER_32_1076 ();
 FILLCELL_X4 FILLER_32_1083 ();
 FILLCELL_X2 FILLER_32_1087 ();
 FILLCELL_X1 FILLER_32_1089 ();
 FILLCELL_X4 FILLER_32_1093 ();
 FILLCELL_X4 FILLER_32_1099 ();
 FILLCELL_X4 FILLER_32_1105 ();
 FILLCELL_X2 FILLER_32_1109 ();
 FILLCELL_X1 FILLER_32_1111 ();
 FILLCELL_X4 FILLER_32_1121 ();
 FILLCELL_X4 FILLER_32_1129 ();
 FILLCELL_X4 FILLER_32_1135 ();
 FILLCELL_X8 FILLER_32_1146 ();
 FILLCELL_X2 FILLER_32_1154 ();
 FILLCELL_X1 FILLER_32_1156 ();
 FILLCELL_X8 FILLER_32_1167 ();
 FILLCELL_X4 FILLER_32_1175 ();
 FILLCELL_X4 FILLER_32_1183 ();
 FILLCELL_X4 FILLER_32_1190 ();
 FILLCELL_X8 FILLER_32_1204 ();
 FILLCELL_X4 FILLER_32_1212 ();
 FILLCELL_X8 FILLER_32_1226 ();
 FILLCELL_X4 FILLER_32_1236 ();
 FILLCELL_X4 FILLER_32_1250 ();
 FILLCELL_X4 FILLER_32_1264 ();
 FILLCELL_X8 FILLER_32_1272 ();
 FILLCELL_X4 FILLER_32_1280 ();
 FILLCELL_X2 FILLER_32_1284 ();
 FILLCELL_X1 FILLER_32_1286 ();
 FILLCELL_X4 FILLER_32_1289 ();
 FILLCELL_X4 FILLER_32_1300 ();
 FILLCELL_X4 FILLER_32_1314 ();
 FILLCELL_X4 FILLER_32_1321 ();
 FILLCELL_X2 FILLER_32_1325 ();
 FILLCELL_X1 FILLER_32_1327 ();
 FILLCELL_X8 FILLER_32_1331 ();
 FILLCELL_X4 FILLER_32_1342 ();
 FILLCELL_X16 FILLER_32_1348 ();
 FILLCELL_X4 FILLER_32_1364 ();
 FILLCELL_X1 FILLER_32_1368 ();
 FILLCELL_X4 FILLER_32_1373 ();
 FILLCELL_X4 FILLER_32_1386 ();
 FILLCELL_X4 FILLER_32_1393 ();
 FILLCELL_X4 FILLER_32_1401 ();
 FILLCELL_X4 FILLER_32_1415 ();
 FILLCELL_X8 FILLER_32_1422 ();
 FILLCELL_X1 FILLER_32_1430 ();
 FILLCELL_X4 FILLER_32_1441 ();
 FILLCELL_X32 FILLER_32_1448 ();
 FILLCELL_X32 FILLER_32_1480 ();
 FILLCELL_X32 FILLER_32_1512 ();
 FILLCELL_X32 FILLER_32_1544 ();
 FILLCELL_X32 FILLER_32_1576 ();
 FILLCELL_X32 FILLER_32_1608 ();
 FILLCELL_X32 FILLER_32_1640 ();
 FILLCELL_X32 FILLER_32_1672 ();
 FILLCELL_X32 FILLER_32_1704 ();
 FILLCELL_X16 FILLER_32_1736 ();
 FILLCELL_X8 FILLER_32_1752 ();
 FILLCELL_X2 FILLER_32_1760 ();
 FILLCELL_X4 FILLER_33_1 ();
 FILLCELL_X2 FILLER_33_5 ();
 FILLCELL_X1 FILLER_33_7 ();
 FILLCELL_X4 FILLER_33_11 ();
 FILLCELL_X2 FILLER_33_15 ();
 FILLCELL_X8 FILLER_33_20 ();
 FILLCELL_X4 FILLER_33_28 ();
 FILLCELL_X2 FILLER_33_32 ();
 FILLCELL_X4 FILLER_33_43 ();
 FILLCELL_X8 FILLER_33_56 ();
 FILLCELL_X8 FILLER_33_74 ();
 FILLCELL_X4 FILLER_33_82 ();
 FILLCELL_X1 FILLER_33_86 ();
 FILLCELL_X4 FILLER_33_90 ();
 FILLCELL_X4 FILLER_33_97 ();
 FILLCELL_X4 FILLER_33_108 ();
 FILLCELL_X2 FILLER_33_112 ();
 FILLCELL_X1 FILLER_33_114 ();
 FILLCELL_X4 FILLER_33_118 ();
 FILLCELL_X4 FILLER_33_132 ();
 FILLCELL_X2 FILLER_33_136 ();
 FILLCELL_X4 FILLER_33_142 ();
 FILLCELL_X4 FILLER_33_150 ();
 FILLCELL_X4 FILLER_33_163 ();
 FILLCELL_X8 FILLER_33_171 ();
 FILLCELL_X4 FILLER_33_188 ();
 FILLCELL_X8 FILLER_33_195 ();
 FILLCELL_X4 FILLER_33_203 ();
 FILLCELL_X1 FILLER_33_207 ();
 FILLCELL_X32 FILLER_33_233 ();
 FILLCELL_X4 FILLER_33_265 ();
 FILLCELL_X2 FILLER_33_269 ();
 FILLCELL_X4 FILLER_33_275 ();
 FILLCELL_X8 FILLER_33_282 ();
 FILLCELL_X2 FILLER_33_290 ();
 FILLCELL_X4 FILLER_33_296 ();
 FILLCELL_X8 FILLER_33_309 ();
 FILLCELL_X4 FILLER_33_326 ();
 FILLCELL_X4 FILLER_33_337 ();
 FILLCELL_X4 FILLER_33_343 ();
 FILLCELL_X2 FILLER_33_347 ();
 FILLCELL_X1 FILLER_33_349 ();
 FILLCELL_X4 FILLER_33_353 ();
 FILLCELL_X8 FILLER_33_359 ();
 FILLCELL_X4 FILLER_33_367 ();
 FILLCELL_X4 FILLER_33_374 ();
 FILLCELL_X4 FILLER_33_381 ();
 FILLCELL_X4 FILLER_33_389 ();
 FILLCELL_X8 FILLER_33_396 ();
 FILLCELL_X4 FILLER_33_404 ();
 FILLCELL_X2 FILLER_33_408 ();
 FILLCELL_X1 FILLER_33_410 ();
 FILLCELL_X4 FILLER_33_414 ();
 FILLCELL_X4 FILLER_33_427 ();
 FILLCELL_X1 FILLER_33_431 ();
 FILLCELL_X16 FILLER_33_439 ();
 FILLCELL_X4 FILLER_33_458 ();
 FILLCELL_X1 FILLER_33_462 ();
 FILLCELL_X8 FILLER_33_468 ();
 FILLCELL_X4 FILLER_33_476 ();
 FILLCELL_X2 FILLER_33_480 ();
 FILLCELL_X4 FILLER_33_489 ();
 FILLCELL_X4 FILLER_33_502 ();
 FILLCELL_X4 FILLER_33_509 ();
 FILLCELL_X8 FILLER_33_516 ();
 FILLCELL_X16 FILLER_33_527 ();
 FILLCELL_X8 FILLER_33_543 ();
 FILLCELL_X4 FILLER_33_561 ();
 FILLCELL_X4 FILLER_33_574 ();
 FILLCELL_X4 FILLER_33_580 ();
 FILLCELL_X2 FILLER_33_584 ();
 FILLCELL_X8 FILLER_33_596 ();
 FILLCELL_X2 FILLER_33_604 ();
 FILLCELL_X4 FILLER_33_612 ();
 FILLCELL_X8 FILLER_33_622 ();
 FILLCELL_X2 FILLER_33_630 ();
 FILLCELL_X8 FILLER_33_645 ();
 FILLCELL_X4 FILLER_33_653 ();
 FILLCELL_X2 FILLER_33_657 ();
 FILLCELL_X1 FILLER_33_659 ();
 FILLCELL_X16 FILLER_33_664 ();
 FILLCELL_X4 FILLER_33_699 ();
 FILLCELL_X32 FILLER_33_722 ();
 FILLCELL_X8 FILLER_33_754 ();
 FILLCELL_X4 FILLER_33_762 ();
 FILLCELL_X16 FILLER_33_770 ();
 FILLCELL_X8 FILLER_33_786 ();
 FILLCELL_X1 FILLER_33_794 ();
 FILLCELL_X4 FILLER_33_801 ();
 FILLCELL_X4 FILLER_33_811 ();
 FILLCELL_X2 FILLER_33_815 ();
 FILLCELL_X4 FILLER_33_821 ();
 FILLCELL_X4 FILLER_33_835 ();
 FILLCELL_X4 FILLER_33_841 ();
 FILLCELL_X4 FILLER_33_849 ();
 FILLCELL_X8 FILLER_33_862 ();
 FILLCELL_X4 FILLER_33_873 ();
 FILLCELL_X4 FILLER_33_880 ();
 FILLCELL_X8 FILLER_33_893 ();
 FILLCELL_X2 FILLER_33_901 ();
 FILLCELL_X4 FILLER_33_905 ();
 FILLCELL_X4 FILLER_33_913 ();
 FILLCELL_X4 FILLER_33_927 ();
 FILLCELL_X8 FILLER_33_938 ();
 FILLCELL_X16 FILLER_33_949 ();
 FILLCELL_X1 FILLER_33_965 ();
 FILLCELL_X4 FILLER_33_968 ();
 FILLCELL_X4 FILLER_33_975 ();
 FILLCELL_X1 FILLER_33_979 ();
 FILLCELL_X4 FILLER_33_984 ();
 FILLCELL_X4 FILLER_33_991 ();
 FILLCELL_X4 FILLER_33_998 ();
 FILLCELL_X4 FILLER_33_1005 ();
 FILLCELL_X2 FILLER_33_1009 ();
 FILLCELL_X4 FILLER_33_1017 ();
 FILLCELL_X4 FILLER_33_1025 ();
 FILLCELL_X4 FILLER_33_1033 ();
 FILLCELL_X1 FILLER_33_1037 ();
 FILLCELL_X8 FILLER_33_1048 ();
 FILLCELL_X1 FILLER_33_1056 ();
 FILLCELL_X8 FILLER_33_1061 ();
 FILLCELL_X4 FILLER_33_1072 ();
 FILLCELL_X4 FILLER_33_1082 ();
 FILLCELL_X4 FILLER_33_1090 ();
 FILLCELL_X2 FILLER_33_1094 ();
 FILLCELL_X4 FILLER_33_1098 ();
 FILLCELL_X4 FILLER_33_1106 ();
 FILLCELL_X4 FILLER_33_1119 ();
 FILLCELL_X2 FILLER_33_1123 ();
 FILLCELL_X1 FILLER_33_1125 ();
 FILLCELL_X4 FILLER_33_1136 ();
 FILLCELL_X4 FILLER_33_1150 ();
 FILLCELL_X4 FILLER_33_1158 ();
 FILLCELL_X8 FILLER_33_1165 ();
 FILLCELL_X4 FILLER_33_1173 ();
 FILLCELL_X2 FILLER_33_1177 ();
 FILLCELL_X4 FILLER_33_1189 ();
 FILLCELL_X4 FILLER_33_1200 ();
 FILLCELL_X4 FILLER_33_1206 ();
 FILLCELL_X2 FILLER_33_1210 ();
 FILLCELL_X1 FILLER_33_1212 ();
 FILLCELL_X4 FILLER_33_1216 ();
 FILLCELL_X1 FILLER_33_1220 ();
 FILLCELL_X4 FILLER_33_1228 ();
 FILLCELL_X8 FILLER_33_1234 ();
 FILLCELL_X4 FILLER_33_1242 ();
 FILLCELL_X4 FILLER_33_1249 ();
 FILLCELL_X4 FILLER_33_1256 ();
 FILLCELL_X2 FILLER_33_1260 ();
 FILLCELL_X1 FILLER_33_1262 ();
 FILLCELL_X4 FILLER_33_1264 ();
 FILLCELL_X2 FILLER_33_1268 ();
 FILLCELL_X4 FILLER_33_1274 ();
 FILLCELL_X4 FILLER_33_1282 ();
 FILLCELL_X8 FILLER_33_1289 ();
 FILLCELL_X1 FILLER_33_1297 ();
 FILLCELL_X4 FILLER_33_1301 ();
 FILLCELL_X8 FILLER_33_1309 ();
 FILLCELL_X4 FILLER_33_1317 ();
 FILLCELL_X1 FILLER_33_1321 ();
 FILLCELL_X4 FILLER_33_1331 ();
 FILLCELL_X4 FILLER_33_1339 ();
 FILLCELL_X4 FILLER_33_1347 ();
 FILLCELL_X8 FILLER_33_1360 ();
 FILLCELL_X8 FILLER_33_1371 ();
 FILLCELL_X8 FILLER_33_1382 ();
 FILLCELL_X4 FILLER_33_1390 ();
 FILLCELL_X4 FILLER_33_1398 ();
 FILLCELL_X8 FILLER_33_1411 ();
 FILLCELL_X4 FILLER_33_1419 ();
 FILLCELL_X2 FILLER_33_1423 ();
 FILLCELL_X1 FILLER_33_1425 ();
 FILLCELL_X4 FILLER_33_1429 ();
 FILLCELL_X4 FILLER_33_1440 ();
 FILLCELL_X1 FILLER_33_1444 ();
 FILLCELL_X32 FILLER_33_1449 ();
 FILLCELL_X32 FILLER_33_1481 ();
 FILLCELL_X32 FILLER_33_1513 ();
 FILLCELL_X32 FILLER_33_1545 ();
 FILLCELL_X32 FILLER_33_1577 ();
 FILLCELL_X32 FILLER_33_1609 ();
 FILLCELL_X32 FILLER_33_1641 ();
 FILLCELL_X32 FILLER_33_1673 ();
 FILLCELL_X32 FILLER_33_1705 ();
 FILLCELL_X16 FILLER_33_1737 ();
 FILLCELL_X8 FILLER_33_1753 ();
 FILLCELL_X1 FILLER_33_1761 ();
 FILLCELL_X16 FILLER_34_1 ();
 FILLCELL_X4 FILLER_34_17 ();
 FILLCELL_X8 FILLER_34_31 ();
 FILLCELL_X4 FILLER_34_39 ();
 FILLCELL_X1 FILLER_34_43 ();
 FILLCELL_X4 FILLER_34_47 ();
 FILLCELL_X4 FILLER_34_54 ();
 FILLCELL_X4 FILLER_34_62 ();
 FILLCELL_X8 FILLER_34_69 ();
 FILLCELL_X4 FILLER_34_77 ();
 FILLCELL_X2 FILLER_34_81 ();
 FILLCELL_X4 FILLER_34_87 ();
 FILLCELL_X4 FILLER_34_101 ();
 FILLCELL_X2 FILLER_34_105 ();
 FILLCELL_X8 FILLER_34_114 ();
 FILLCELL_X1 FILLER_34_122 ();
 FILLCELL_X16 FILLER_34_126 ();
 FILLCELL_X2 FILLER_34_142 ();
 FILLCELL_X1 FILLER_34_144 ();
 FILLCELL_X4 FILLER_34_154 ();
 FILLCELL_X1 FILLER_34_158 ();
 FILLCELL_X16 FILLER_34_162 ();
 FILLCELL_X8 FILLER_34_178 ();
 FILLCELL_X4 FILLER_34_186 ();
 FILLCELL_X4 FILLER_34_194 ();
 FILLCELL_X4 FILLER_34_202 ();
 FILLCELL_X16 FILLER_34_210 ();
 FILLCELL_X4 FILLER_34_226 ();
 FILLCELL_X2 FILLER_34_230 ();
 FILLCELL_X1 FILLER_34_232 ();
 FILLCELL_X4 FILLER_34_237 ();
 FILLCELL_X8 FILLER_34_244 ();
 FILLCELL_X4 FILLER_34_252 ();
 FILLCELL_X4 FILLER_34_260 ();
 FILLCELL_X4 FILLER_34_267 ();
 FILLCELL_X2 FILLER_34_271 ();
 FILLCELL_X4 FILLER_34_282 ();
 FILLCELL_X1 FILLER_34_286 ();
 FILLCELL_X4 FILLER_34_291 ();
 FILLCELL_X8 FILLER_34_304 ();
 FILLCELL_X4 FILLER_34_315 ();
 FILLCELL_X4 FILLER_34_324 ();
 FILLCELL_X4 FILLER_34_337 ();
 FILLCELL_X4 FILLER_34_351 ();
 FILLCELL_X4 FILLER_34_365 ();
 FILLCELL_X8 FILLER_34_378 ();
 FILLCELL_X1 FILLER_34_386 ();
 FILLCELL_X4 FILLER_34_391 ();
 FILLCELL_X4 FILLER_34_399 ();
 FILLCELL_X4 FILLER_34_407 ();
 FILLCELL_X1 FILLER_34_411 ();
 FILLCELL_X4 FILLER_34_415 ();
 FILLCELL_X4 FILLER_34_429 ();
 FILLCELL_X4 FILLER_34_443 ();
 FILLCELL_X4 FILLER_34_451 ();
 FILLCELL_X4 FILLER_34_464 ();
 FILLCELL_X2 FILLER_34_468 ();
 FILLCELL_X4 FILLER_34_480 ();
 FILLCELL_X8 FILLER_34_494 ();
 FILLCELL_X4 FILLER_34_502 ();
 FILLCELL_X4 FILLER_34_509 ();
 FILLCELL_X2 FILLER_34_513 ();
 FILLCELL_X4 FILLER_34_520 ();
 FILLCELL_X4 FILLER_34_527 ();
 FILLCELL_X16 FILLER_34_534 ();
 FILLCELL_X1 FILLER_34_550 ();
 FILLCELL_X8 FILLER_34_564 ();
 FILLCELL_X1 FILLER_34_572 ();
 FILLCELL_X16 FILLER_34_583 ();
 FILLCELL_X4 FILLER_34_618 ();
 FILLCELL_X1 FILLER_34_622 ();
 FILLCELL_X4 FILLER_34_627 ();
 FILLCELL_X4 FILLER_34_632 ();
 FILLCELL_X8 FILLER_34_639 ();
 FILLCELL_X4 FILLER_34_666 ();
 FILLCELL_X2 FILLER_34_670 ();
 FILLCELL_X1 FILLER_34_672 ();
 FILLCELL_X8 FILLER_34_692 ();
 FILLCELL_X4 FILLER_34_700 ();
 FILLCELL_X1 FILLER_34_704 ();
 FILLCELL_X4 FILLER_34_709 ();
 FILLCELL_X2 FILLER_34_713 ();
 FILLCELL_X1 FILLER_34_715 ();
 FILLCELL_X8 FILLER_34_735 ();
 FILLCELL_X4 FILLER_34_743 ();
 FILLCELL_X2 FILLER_34_747 ();
 FILLCELL_X4 FILLER_34_753 ();
 FILLCELL_X4 FILLER_34_776 ();
 FILLCELL_X8 FILLER_34_799 ();
 FILLCELL_X8 FILLER_34_811 ();
 FILLCELL_X4 FILLER_34_819 ();
 FILLCELL_X1 FILLER_34_823 ();
 FILLCELL_X4 FILLER_34_828 ();
 FILLCELL_X2 FILLER_34_832 ();
 FILLCELL_X1 FILLER_34_834 ();
 FILLCELL_X4 FILLER_34_838 ();
 FILLCELL_X16 FILLER_34_845 ();
 FILLCELL_X2 FILLER_34_861 ();
 FILLCELL_X8 FILLER_34_866 ();
 FILLCELL_X16 FILLER_34_876 ();
 FILLCELL_X2 FILLER_34_892 ();
 FILLCELL_X1 FILLER_34_894 ();
 FILLCELL_X16 FILLER_34_899 ();
 FILLCELL_X4 FILLER_34_915 ();
 FILLCELL_X4 FILLER_34_922 ();
 FILLCELL_X2 FILLER_34_926 ();
 FILLCELL_X4 FILLER_34_937 ();
 FILLCELL_X1 FILLER_34_941 ();
 FILLCELL_X4 FILLER_34_951 ();
 FILLCELL_X8 FILLER_34_958 ();
 FILLCELL_X8 FILLER_34_970 ();
 FILLCELL_X1 FILLER_34_978 ();
 FILLCELL_X4 FILLER_34_983 ();
 FILLCELL_X4 FILLER_34_990 ();
 FILLCELL_X2 FILLER_34_994 ();
 FILLCELL_X1 FILLER_34_996 ();
 FILLCELL_X4 FILLER_34_1001 ();
 FILLCELL_X4 FILLER_34_1009 ();
 FILLCELL_X1 FILLER_34_1013 ();
 FILLCELL_X4 FILLER_34_1019 ();
 FILLCELL_X8 FILLER_34_1027 ();
 FILLCELL_X4 FILLER_34_1039 ();
 FILLCELL_X1 FILLER_34_1043 ();
 FILLCELL_X4 FILLER_34_1051 ();
 FILLCELL_X4 FILLER_34_1065 ();
 FILLCELL_X4 FILLER_34_1072 ();
 FILLCELL_X4 FILLER_34_1078 ();
 FILLCELL_X1 FILLER_34_1082 ();
 FILLCELL_X4 FILLER_34_1089 ();
 FILLCELL_X8 FILLER_34_1097 ();
 FILLCELL_X4 FILLER_34_1105 ();
 FILLCELL_X4 FILLER_34_1113 ();
 FILLCELL_X4 FILLER_34_1120 ();
 FILLCELL_X4 FILLER_34_1128 ();
 FILLCELL_X4 FILLER_34_1134 ();
 FILLCELL_X16 FILLER_34_1140 ();
 FILLCELL_X2 FILLER_34_1156 ();
 FILLCELL_X4 FILLER_34_1167 ();
 FILLCELL_X8 FILLER_34_1181 ();
 FILLCELL_X4 FILLER_34_1193 ();
 FILLCELL_X4 FILLER_34_1199 ();
 FILLCELL_X1 FILLER_34_1203 ();
 FILLCELL_X8 FILLER_34_1211 ();
 FILLCELL_X4 FILLER_34_1229 ();
 FILLCELL_X4 FILLER_34_1236 ();
 FILLCELL_X4 FILLER_34_1243 ();
 FILLCELL_X4 FILLER_34_1256 ();
 FILLCELL_X4 FILLER_34_1263 ();
 FILLCELL_X1 FILLER_34_1267 ();
 FILLCELL_X4 FILLER_34_1277 ();
 FILLCELL_X4 FILLER_34_1290 ();
 FILLCELL_X4 FILLER_34_1303 ();
 FILLCELL_X4 FILLER_34_1311 ();
 FILLCELL_X4 FILLER_34_1318 ();
 FILLCELL_X4 FILLER_34_1331 ();
 FILLCELL_X4 FILLER_34_1339 ();
 FILLCELL_X1 FILLER_34_1343 ();
 FILLCELL_X4 FILLER_34_1348 ();
 FILLCELL_X4 FILLER_34_1361 ();
 FILLCELL_X8 FILLER_34_1368 ();
 FILLCELL_X2 FILLER_34_1376 ();
 FILLCELL_X4 FILLER_34_1383 ();
 FILLCELL_X8 FILLER_34_1389 ();
 FILLCELL_X2 FILLER_34_1397 ();
 FILLCELL_X1 FILLER_34_1399 ();
 FILLCELL_X4 FILLER_34_1403 ();
 FILLCELL_X8 FILLER_34_1410 ();
 FILLCELL_X2 FILLER_34_1418 ();
 FILLCELL_X4 FILLER_34_1424 ();
 FILLCELL_X4 FILLER_34_1441 ();
 FILLCELL_X2 FILLER_34_1445 ();
 FILLCELL_X1 FILLER_34_1447 ();
 FILLCELL_X32 FILLER_34_1467 ();
 FILLCELL_X32 FILLER_34_1499 ();
 FILLCELL_X32 FILLER_34_1531 ();
 FILLCELL_X32 FILLER_34_1563 ();
 FILLCELL_X32 FILLER_34_1595 ();
 FILLCELL_X32 FILLER_34_1627 ();
 FILLCELL_X32 FILLER_34_1659 ();
 FILLCELL_X32 FILLER_34_1691 ();
 FILLCELL_X32 FILLER_34_1723 ();
 FILLCELL_X4 FILLER_34_1755 ();
 FILLCELL_X2 FILLER_34_1759 ();
 FILLCELL_X1 FILLER_34_1761 ();
 FILLCELL_X4 FILLER_35_1 ();
 FILLCELL_X8 FILLER_35_8 ();
 FILLCELL_X4 FILLER_35_16 ();
 FILLCELL_X8 FILLER_35_22 ();
 FILLCELL_X2 FILLER_35_30 ();
 FILLCELL_X1 FILLER_35_32 ();
 FILLCELL_X4 FILLER_35_35 ();
 FILLCELL_X4 FILLER_35_48 ();
 FILLCELL_X8 FILLER_35_55 ();
 FILLCELL_X2 FILLER_35_63 ();
 FILLCELL_X8 FILLER_35_74 ();
 FILLCELL_X4 FILLER_35_82 ();
 FILLCELL_X1 FILLER_35_86 ();
 FILLCELL_X4 FILLER_35_96 ();
 FILLCELL_X4 FILLER_35_104 ();
 FILLCELL_X4 FILLER_35_118 ();
 FILLCELL_X4 FILLER_35_131 ();
 FILLCELL_X8 FILLER_35_138 ();
 FILLCELL_X1 FILLER_35_146 ();
 FILLCELL_X4 FILLER_35_151 ();
 FILLCELL_X2 FILLER_35_155 ();
 FILLCELL_X1 FILLER_35_157 ();
 FILLCELL_X4 FILLER_35_161 ();
 FILLCELL_X8 FILLER_35_168 ();
 FILLCELL_X4 FILLER_35_176 ();
 FILLCELL_X8 FILLER_35_185 ();
 FILLCELL_X8 FILLER_35_212 ();
 FILLCELL_X4 FILLER_35_220 ();
 FILLCELL_X2 FILLER_35_224 ();
 FILLCELL_X4 FILLER_35_230 ();
 FILLCELL_X4 FILLER_35_243 ();
 FILLCELL_X4 FILLER_35_252 ();
 FILLCELL_X1 FILLER_35_256 ();
 FILLCELL_X4 FILLER_35_266 ();
 FILLCELL_X16 FILLER_35_274 ();
 FILLCELL_X2 FILLER_35_290 ();
 FILLCELL_X8 FILLER_35_296 ();
 FILLCELL_X2 FILLER_35_304 ();
 FILLCELL_X4 FILLER_35_311 ();
 FILLCELL_X4 FILLER_35_318 ();
 FILLCELL_X4 FILLER_35_325 ();
 FILLCELL_X8 FILLER_35_339 ();
 FILLCELL_X4 FILLER_35_347 ();
 FILLCELL_X2 FILLER_35_351 ();
 FILLCELL_X4 FILLER_35_360 ();
 FILLCELL_X1 FILLER_35_364 ();
 FILLCELL_X4 FILLER_35_368 ();
 FILLCELL_X4 FILLER_35_376 ();
 FILLCELL_X8 FILLER_35_383 ();
 FILLCELL_X4 FILLER_35_391 ();
 FILLCELL_X2 FILLER_35_395 ();
 FILLCELL_X4 FILLER_35_406 ();
 FILLCELL_X4 FILLER_35_419 ();
 FILLCELL_X2 FILLER_35_423 ();
 FILLCELL_X1 FILLER_35_425 ();
 FILLCELL_X4 FILLER_35_429 ();
 FILLCELL_X8 FILLER_35_435 ();
 FILLCELL_X4 FILLER_35_443 ();
 FILLCELL_X8 FILLER_35_456 ();
 FILLCELL_X2 FILLER_35_464 ();
 FILLCELL_X4 FILLER_35_470 ();
 FILLCELL_X4 FILLER_35_478 ();
 FILLCELL_X8 FILLER_35_485 ();
 FILLCELL_X1 FILLER_35_493 ();
 FILLCELL_X4 FILLER_35_503 ();
 FILLCELL_X4 FILLER_35_516 ();
 FILLCELL_X4 FILLER_35_529 ();
 FILLCELL_X4 FILLER_35_543 ();
 FILLCELL_X4 FILLER_35_549 ();
 FILLCELL_X1 FILLER_35_553 ();
 FILLCELL_X4 FILLER_35_557 ();
 FILLCELL_X2 FILLER_35_561 ();
 FILLCELL_X4 FILLER_35_566 ();
 FILLCELL_X8 FILLER_35_580 ();
 FILLCELL_X2 FILLER_35_588 ();
 FILLCELL_X1 FILLER_35_590 ();
 FILLCELL_X4 FILLER_35_610 ();
 FILLCELL_X8 FILLER_35_618 ();
 FILLCELL_X4 FILLER_35_626 ();
 FILLCELL_X2 FILLER_35_630 ();
 FILLCELL_X1 FILLER_35_632 ();
 FILLCELL_X8 FILLER_35_637 ();
 FILLCELL_X4 FILLER_35_645 ();
 FILLCELL_X2 FILLER_35_649 ();
 FILLCELL_X1 FILLER_35_651 ();
 FILLCELL_X16 FILLER_35_656 ();
 FILLCELL_X16 FILLER_35_676 ();
 FILLCELL_X8 FILLER_35_692 ();
 FILLCELL_X8 FILLER_35_705 ();
 FILLCELL_X4 FILLER_35_713 ();
 FILLCELL_X2 FILLER_35_717 ();
 FILLCELL_X4 FILLER_35_723 ();
 FILLCELL_X4 FILLER_35_746 ();
 FILLCELL_X8 FILLER_35_769 ();
 FILLCELL_X4 FILLER_35_777 ();
 FILLCELL_X1 FILLER_35_781 ();
 FILLCELL_X32 FILLER_35_786 ();
 FILLCELL_X16 FILLER_35_818 ();
 FILLCELL_X8 FILLER_35_844 ();
 FILLCELL_X2 FILLER_35_852 ();
 FILLCELL_X4 FILLER_35_858 ();
 FILLCELL_X8 FILLER_35_872 ();
 FILLCELL_X1 FILLER_35_880 ();
 FILLCELL_X4 FILLER_35_885 ();
 FILLCELL_X4 FILLER_35_899 ();
 FILLCELL_X8 FILLER_35_913 ();
 FILLCELL_X4 FILLER_35_921 ();
 FILLCELL_X2 FILLER_35_925 ();
 FILLCELL_X4 FILLER_35_930 ();
 FILLCELL_X8 FILLER_35_937 ();
 FILLCELL_X1 FILLER_35_945 ();
 FILLCELL_X4 FILLER_35_953 ();
 FILLCELL_X2 FILLER_35_957 ();
 FILLCELL_X1 FILLER_35_959 ();
 FILLCELL_X4 FILLER_35_964 ();
 FILLCELL_X8 FILLER_35_977 ();
 FILLCELL_X1 FILLER_35_985 ();
 FILLCELL_X4 FILLER_35_993 ();
 FILLCELL_X4 FILLER_35_1003 ();
 FILLCELL_X4 FILLER_35_1013 ();
 FILLCELL_X4 FILLER_35_1023 ();
 FILLCELL_X4 FILLER_35_1033 ();
 FILLCELL_X4 FILLER_35_1041 ();
 FILLCELL_X4 FILLER_35_1049 ();
 FILLCELL_X8 FILLER_35_1055 ();
 FILLCELL_X1 FILLER_35_1063 ();
 FILLCELL_X4 FILLER_35_1067 ();
 FILLCELL_X4 FILLER_35_1073 ();
 FILLCELL_X4 FILLER_35_1079 ();
 FILLCELL_X4 FILLER_35_1087 ();
 FILLCELL_X1 FILLER_35_1091 ();
 FILLCELL_X4 FILLER_35_1109 ();
 FILLCELL_X4 FILLER_35_1115 ();
 FILLCELL_X2 FILLER_35_1119 ();
 FILLCELL_X1 FILLER_35_1121 ();
 FILLCELL_X8 FILLER_35_1131 ();
 FILLCELL_X4 FILLER_35_1139 ();
 FILLCELL_X4 FILLER_35_1147 ();
 FILLCELL_X4 FILLER_35_1154 ();
 FILLCELL_X2 FILLER_35_1158 ();
 FILLCELL_X1 FILLER_35_1160 ();
 FILLCELL_X4 FILLER_35_1170 ();
 FILLCELL_X4 FILLER_35_1177 ();
 FILLCELL_X8 FILLER_35_1184 ();
 FILLCELL_X8 FILLER_35_1202 ();
 FILLCELL_X2 FILLER_35_1210 ();
 FILLCELL_X1 FILLER_35_1212 ();
 FILLCELL_X4 FILLER_35_1223 ();
 FILLCELL_X8 FILLER_35_1231 ();
 FILLCELL_X4 FILLER_35_1239 ();
 FILLCELL_X2 FILLER_35_1243 ();
 FILLCELL_X8 FILLER_35_1254 ();
 FILLCELL_X1 FILLER_35_1262 ();
 FILLCELL_X8 FILLER_35_1264 ();
 FILLCELL_X2 FILLER_35_1272 ();
 FILLCELL_X1 FILLER_35_1274 ();
 FILLCELL_X4 FILLER_35_1279 ();
 FILLCELL_X4 FILLER_35_1286 ();
 FILLCELL_X4 FILLER_35_1293 ();
 FILLCELL_X2 FILLER_35_1297 ();
 FILLCELL_X16 FILLER_35_1302 ();
 FILLCELL_X4 FILLER_35_1318 ();
 FILLCELL_X16 FILLER_35_1329 ();
 FILLCELL_X4 FILLER_35_1345 ();
 FILLCELL_X2 FILLER_35_1349 ();
 FILLCELL_X8 FILLER_35_1355 ();
 FILLCELL_X2 FILLER_35_1363 ();
 FILLCELL_X4 FILLER_35_1369 ();
 FILLCELL_X4 FILLER_35_1380 ();
 FILLCELL_X4 FILLER_35_1401 ();
 FILLCELL_X4 FILLER_35_1414 ();
 FILLCELL_X4 FILLER_35_1422 ();
 FILLCELL_X2 FILLER_35_1426 ();
 FILLCELL_X4 FILLER_35_1434 ();
 FILLCELL_X32 FILLER_35_1444 ();
 FILLCELL_X32 FILLER_35_1476 ();
 FILLCELL_X32 FILLER_35_1508 ();
 FILLCELL_X32 FILLER_35_1540 ();
 FILLCELL_X32 FILLER_35_1572 ();
 FILLCELL_X32 FILLER_35_1604 ();
 FILLCELL_X32 FILLER_35_1636 ();
 FILLCELL_X32 FILLER_35_1668 ();
 FILLCELL_X32 FILLER_35_1700 ();
 FILLCELL_X16 FILLER_35_1732 ();
 FILLCELL_X8 FILLER_35_1748 ();
 FILLCELL_X4 FILLER_35_1756 ();
 FILLCELL_X2 FILLER_35_1760 ();
 FILLCELL_X16 FILLER_36_1 ();
 FILLCELL_X4 FILLER_36_17 ();
 FILLCELL_X2 FILLER_36_21 ();
 FILLCELL_X4 FILLER_36_30 ();
 FILLCELL_X2 FILLER_36_34 ();
 FILLCELL_X1 FILLER_36_36 ();
 FILLCELL_X8 FILLER_36_47 ();
 FILLCELL_X2 FILLER_36_55 ();
 FILLCELL_X1 FILLER_36_57 ();
 FILLCELL_X4 FILLER_36_61 ();
 FILLCELL_X4 FILLER_36_69 ();
 FILLCELL_X1 FILLER_36_73 ();
 FILLCELL_X8 FILLER_36_77 ();
 FILLCELL_X4 FILLER_36_85 ();
 FILLCELL_X1 FILLER_36_89 ();
 FILLCELL_X4 FILLER_36_100 ();
 FILLCELL_X4 FILLER_36_106 ();
 FILLCELL_X1 FILLER_36_110 ();
 FILLCELL_X8 FILLER_36_114 ();
 FILLCELL_X8 FILLER_36_125 ();
 FILLCELL_X4 FILLER_36_133 ();
 FILLCELL_X2 FILLER_36_137 ();
 FILLCELL_X4 FILLER_36_143 ();
 FILLCELL_X4 FILLER_36_156 ();
 FILLCELL_X2 FILLER_36_160 ();
 FILLCELL_X1 FILLER_36_162 ();
 FILLCELL_X4 FILLER_36_166 ();
 FILLCELL_X2 FILLER_36_170 ();
 FILLCELL_X4 FILLER_36_174 ();
 FILLCELL_X32 FILLER_36_195 ();
 FILLCELL_X8 FILLER_36_227 ();
 FILLCELL_X1 FILLER_36_235 ();
 FILLCELL_X8 FILLER_36_240 ();
 FILLCELL_X1 FILLER_36_248 ();
 FILLCELL_X4 FILLER_36_253 ();
 FILLCELL_X4 FILLER_36_266 ();
 FILLCELL_X4 FILLER_36_273 ();
 FILLCELL_X8 FILLER_36_281 ();
 FILLCELL_X2 FILLER_36_289 ();
 FILLCELL_X4 FILLER_36_295 ();
 FILLCELL_X1 FILLER_36_299 ();
 FILLCELL_X4 FILLER_36_309 ();
 FILLCELL_X8 FILLER_36_318 ();
 FILLCELL_X2 FILLER_36_326 ();
 FILLCELL_X32 FILLER_36_332 ();
 FILLCELL_X2 FILLER_36_364 ();
 FILLCELL_X4 FILLER_36_370 ();
 FILLCELL_X4 FILLER_36_383 ();
 FILLCELL_X4 FILLER_36_392 ();
 FILLCELL_X16 FILLER_36_399 ();
 FILLCELL_X1 FILLER_36_415 ();
 FILLCELL_X16 FILLER_36_418 ();
 FILLCELL_X16 FILLER_36_438 ();
 FILLCELL_X8 FILLER_36_454 ();
 FILLCELL_X1 FILLER_36_462 ();
 FILLCELL_X4 FILLER_36_467 ();
 FILLCELL_X8 FILLER_36_474 ();
 FILLCELL_X4 FILLER_36_482 ();
 FILLCELL_X1 FILLER_36_486 ();
 FILLCELL_X16 FILLER_36_489 ();
 FILLCELL_X8 FILLER_36_505 ();
 FILLCELL_X4 FILLER_36_513 ();
 FILLCELL_X8 FILLER_36_520 ();
 FILLCELL_X1 FILLER_36_528 ();
 FILLCELL_X16 FILLER_36_532 ();
 FILLCELL_X1 FILLER_36_548 ();
 FILLCELL_X4 FILLER_36_552 ();
 FILLCELL_X8 FILLER_36_560 ();
 FILLCELL_X4 FILLER_36_568 ();
 FILLCELL_X2 FILLER_36_572 ();
 FILLCELL_X1 FILLER_36_574 ();
 FILLCELL_X4 FILLER_36_594 ();
 FILLCELL_X16 FILLER_36_602 ();
 FILLCELL_X8 FILLER_36_618 ();
 FILLCELL_X4 FILLER_36_626 ();
 FILLCELL_X1 FILLER_36_630 ();
 FILLCELL_X4 FILLER_36_632 ();
 FILLCELL_X16 FILLER_36_655 ();
 FILLCELL_X2 FILLER_36_671 ();
 FILLCELL_X8 FILLER_36_692 ();
 FILLCELL_X1 FILLER_36_700 ();
 FILLCELL_X8 FILLER_36_720 ();
 FILLCELL_X4 FILLER_36_728 ();
 FILLCELL_X1 FILLER_36_732 ();
 FILLCELL_X32 FILLER_36_737 ();
 FILLCELL_X4 FILLER_36_769 ();
 FILLCELL_X8 FILLER_36_792 ();
 FILLCELL_X2 FILLER_36_800 ();
 FILLCELL_X16 FILLER_36_821 ();
 FILLCELL_X1 FILLER_36_837 ();
 FILLCELL_X4 FILLER_36_841 ();
 FILLCELL_X4 FILLER_36_852 ();
 FILLCELL_X4 FILLER_36_859 ();
 FILLCELL_X4 FILLER_36_870 ();
 FILLCELL_X4 FILLER_36_880 ();
 FILLCELL_X1 FILLER_36_884 ();
 FILLCELL_X4 FILLER_36_891 ();
 FILLCELL_X4 FILLER_36_898 ();
 FILLCELL_X4 FILLER_36_904 ();
 FILLCELL_X2 FILLER_36_908 ();
 FILLCELL_X4 FILLER_36_914 ();
 FILLCELL_X4 FILLER_36_927 ();
 FILLCELL_X4 FILLER_36_934 ();
 FILLCELL_X2 FILLER_36_938 ();
 FILLCELL_X1 FILLER_36_940 ();
 FILLCELL_X8 FILLER_36_951 ();
 FILLCELL_X1 FILLER_36_959 ();
 FILLCELL_X4 FILLER_36_969 ();
 FILLCELL_X8 FILLER_36_977 ();
 FILLCELL_X1 FILLER_36_985 ();
 FILLCELL_X4 FILLER_36_989 ();
 FILLCELL_X1 FILLER_36_993 ();
 FILLCELL_X4 FILLER_36_1000 ();
 FILLCELL_X4 FILLER_36_1006 ();
 FILLCELL_X4 FILLER_36_1012 ();
 FILLCELL_X4 FILLER_36_1018 ();
 FILLCELL_X1 FILLER_36_1022 ();
 FILLCELL_X4 FILLER_36_1025 ();
 FILLCELL_X4 FILLER_36_1035 ();
 FILLCELL_X4 FILLER_36_1043 ();
 FILLCELL_X2 FILLER_36_1047 ();
 FILLCELL_X1 FILLER_36_1049 ();
 FILLCELL_X8 FILLER_36_1069 ();
 FILLCELL_X2 FILLER_36_1077 ();
 FILLCELL_X4 FILLER_36_1088 ();
 FILLCELL_X4 FILLER_36_1097 ();
 FILLCELL_X8 FILLER_36_1105 ();
 FILLCELL_X1 FILLER_36_1113 ();
 FILLCELL_X4 FILLER_36_1121 ();
 FILLCELL_X4 FILLER_36_1142 ();
 FILLCELL_X4 FILLER_36_1155 ();
 FILLCELL_X4 FILLER_36_1162 ();
 FILLCELL_X16 FILLER_36_1169 ();
 FILLCELL_X8 FILLER_36_1185 ();
 FILLCELL_X16 FILLER_36_1196 ();
 FILLCELL_X4 FILLER_36_1212 ();
 FILLCELL_X4 FILLER_36_1220 ();
 FILLCELL_X2 FILLER_36_1224 ();
 FILLCELL_X4 FILLER_36_1235 ();
 FILLCELL_X4 FILLER_36_1242 ();
 FILLCELL_X8 FILLER_36_1249 ();
 FILLCELL_X2 FILLER_36_1257 ();
 FILLCELL_X1 FILLER_36_1259 ();
 FILLCELL_X4 FILLER_36_1264 ();
 FILLCELL_X4 FILLER_36_1275 ();
 FILLCELL_X1 FILLER_36_1279 ();
 FILLCELL_X8 FILLER_36_1284 ();
 FILLCELL_X4 FILLER_36_1292 ();
 FILLCELL_X2 FILLER_36_1296 ();
 FILLCELL_X4 FILLER_36_1307 ();
 FILLCELL_X4 FILLER_36_1314 ();
 FILLCELL_X2 FILLER_36_1318 ();
 FILLCELL_X1 FILLER_36_1320 ();
 FILLCELL_X4 FILLER_36_1331 ();
 FILLCELL_X8 FILLER_36_1337 ();
 FILLCELL_X2 FILLER_36_1345 ();
 FILLCELL_X4 FILLER_36_1350 ();
 FILLCELL_X4 FILLER_36_1357 ();
 FILLCELL_X4 FILLER_36_1364 ();
 FILLCELL_X8 FILLER_36_1372 ();
 FILLCELL_X2 FILLER_36_1380 ();
 FILLCELL_X8 FILLER_36_1387 ();
 FILLCELL_X4 FILLER_36_1395 ();
 FILLCELL_X4 FILLER_36_1403 ();
 FILLCELL_X8 FILLER_36_1410 ();
 FILLCELL_X2 FILLER_36_1418 ();
 FILLCELL_X1 FILLER_36_1420 ();
 FILLCELL_X4 FILLER_36_1426 ();
 FILLCELL_X32 FILLER_36_1434 ();
 FILLCELL_X32 FILLER_36_1466 ();
 FILLCELL_X32 FILLER_36_1498 ();
 FILLCELL_X32 FILLER_36_1530 ();
 FILLCELL_X32 FILLER_36_1562 ();
 FILLCELL_X32 FILLER_36_1594 ();
 FILLCELL_X32 FILLER_36_1626 ();
 FILLCELL_X32 FILLER_36_1658 ();
 FILLCELL_X32 FILLER_36_1690 ();
 FILLCELL_X32 FILLER_36_1722 ();
 FILLCELL_X8 FILLER_36_1754 ();
 FILLCELL_X16 FILLER_37_1 ();
 FILLCELL_X2 FILLER_37_17 ();
 FILLCELL_X4 FILLER_37_29 ();
 FILLCELL_X4 FILLER_37_36 ();
 FILLCELL_X2 FILLER_37_40 ();
 FILLCELL_X1 FILLER_37_42 ();
 FILLCELL_X8 FILLER_37_50 ();
 FILLCELL_X4 FILLER_37_62 ();
 FILLCELL_X4 FILLER_37_75 ();
 FILLCELL_X4 FILLER_37_83 ();
 FILLCELL_X2 FILLER_37_87 ();
 FILLCELL_X4 FILLER_37_92 ();
 FILLCELL_X8 FILLER_37_99 ();
 FILLCELL_X1 FILLER_37_107 ();
 FILLCELL_X8 FILLER_37_110 ();
 FILLCELL_X1 FILLER_37_118 ();
 FILLCELL_X4 FILLER_37_128 ();
 FILLCELL_X4 FILLER_37_135 ();
 FILLCELL_X2 FILLER_37_139 ();
 FILLCELL_X4 FILLER_37_150 ();
 FILLCELL_X4 FILLER_37_158 ();
 FILLCELL_X4 FILLER_37_165 ();
 FILLCELL_X4 FILLER_37_173 ();
 FILLCELL_X4 FILLER_37_184 ();
 FILLCELL_X4 FILLER_37_193 ();
 FILLCELL_X1 FILLER_37_197 ();
 FILLCELL_X16 FILLER_37_217 ();
 FILLCELL_X1 FILLER_37_233 ();
 FILLCELL_X4 FILLER_37_243 ();
 FILLCELL_X8 FILLER_37_250 ();
 FILLCELL_X2 FILLER_37_258 ();
 FILLCELL_X1 FILLER_37_260 ();
 FILLCELL_X4 FILLER_37_264 ();
 FILLCELL_X4 FILLER_37_271 ();
 FILLCELL_X8 FILLER_37_285 ();
 FILLCELL_X2 FILLER_37_293 ();
 FILLCELL_X4 FILLER_37_299 ();
 FILLCELL_X4 FILLER_37_312 ();
 FILLCELL_X8 FILLER_37_319 ();
 FILLCELL_X4 FILLER_37_329 ();
 FILLCELL_X4 FILLER_37_340 ();
 FILLCELL_X4 FILLER_37_354 ();
 FILLCELL_X8 FILLER_37_361 ();
 FILLCELL_X4 FILLER_37_372 ();
 FILLCELL_X8 FILLER_37_379 ();
 FILLCELL_X2 FILLER_37_387 ();
 FILLCELL_X4 FILLER_37_392 ();
 FILLCELL_X1 FILLER_37_396 ();
 FILLCELL_X4 FILLER_37_400 ();
 FILLCELL_X4 FILLER_37_414 ();
 FILLCELL_X2 FILLER_37_418 ();
 FILLCELL_X1 FILLER_37_420 ();
 FILLCELL_X4 FILLER_37_428 ();
 FILLCELL_X8 FILLER_37_442 ();
 FILLCELL_X2 FILLER_37_450 ();
 FILLCELL_X1 FILLER_37_452 ();
 FILLCELL_X8 FILLER_37_459 ();
 FILLCELL_X2 FILLER_37_467 ();
 FILLCELL_X4 FILLER_37_486 ();
 FILLCELL_X4 FILLER_37_497 ();
 FILLCELL_X4 FILLER_37_510 ();
 FILLCELL_X4 FILLER_37_524 ();
 FILLCELL_X2 FILLER_37_528 ();
 FILLCELL_X4 FILLER_37_532 ();
 FILLCELL_X4 FILLER_37_540 ();
 FILLCELL_X4 FILLER_37_548 ();
 FILLCELL_X16 FILLER_37_557 ();
 FILLCELL_X8 FILLER_37_573 ();
 FILLCELL_X1 FILLER_37_581 ();
 FILLCELL_X32 FILLER_37_586 ();
 FILLCELL_X1 FILLER_37_618 ();
 FILLCELL_X8 FILLER_37_638 ();
 FILLCELL_X4 FILLER_37_646 ();
 FILLCELL_X4 FILLER_37_669 ();
 FILLCELL_X2 FILLER_37_673 ();
 FILLCELL_X1 FILLER_37_675 ();
 FILLCELL_X8 FILLER_37_695 ();
 FILLCELL_X4 FILLER_37_707 ();
 FILLCELL_X4 FILLER_37_730 ();
 FILLCELL_X4 FILLER_37_753 ();
 FILLCELL_X4 FILLER_37_776 ();
 FILLCELL_X4 FILLER_37_799 ();
 FILLCELL_X4 FILLER_37_822 ();
 FILLCELL_X4 FILLER_37_845 ();
 FILLCELL_X1 FILLER_37_849 ();
 FILLCELL_X4 FILLER_37_856 ();
 FILLCELL_X8 FILLER_37_866 ();
 FILLCELL_X1 FILLER_37_874 ();
 FILLCELL_X4 FILLER_37_879 ();
 FILLCELL_X4 FILLER_37_893 ();
 FILLCELL_X4 FILLER_37_904 ();
 FILLCELL_X1 FILLER_37_908 ();
 FILLCELL_X4 FILLER_37_913 ();
 FILLCELL_X4 FILLER_37_926 ();
 FILLCELL_X4 FILLER_37_933 ();
 FILLCELL_X2 FILLER_37_937 ();
 FILLCELL_X1 FILLER_37_939 ();
 FILLCELL_X4 FILLER_37_944 ();
 FILLCELL_X4 FILLER_37_958 ();
 FILLCELL_X16 FILLER_37_965 ();
 FILLCELL_X8 FILLER_37_981 ();
 FILLCELL_X2 FILLER_37_989 ();
 FILLCELL_X1 FILLER_37_991 ();
 FILLCELL_X4 FILLER_37_994 ();
 FILLCELL_X1 FILLER_37_998 ();
 FILLCELL_X16 FILLER_37_1003 ();
 FILLCELL_X8 FILLER_37_1019 ();
 FILLCELL_X4 FILLER_37_1027 ();
 FILLCELL_X2 FILLER_37_1031 ();
 FILLCELL_X4 FILLER_37_1039 ();
 FILLCELL_X8 FILLER_37_1062 ();
 FILLCELL_X2 FILLER_37_1070 ();
 FILLCELL_X1 FILLER_37_1072 ();
 FILLCELL_X4 FILLER_37_1092 ();
 FILLCELL_X1 FILLER_37_1096 ();
 FILLCELL_X4 FILLER_37_1102 ();
 FILLCELL_X4 FILLER_37_1113 ();
 FILLCELL_X16 FILLER_37_1126 ();
 FILLCELL_X2 FILLER_37_1142 ();
 FILLCELL_X1 FILLER_37_1144 ();
 FILLCELL_X4 FILLER_37_1154 ();
 FILLCELL_X8 FILLER_37_1161 ();
 FILLCELL_X1 FILLER_37_1169 ();
 FILLCELL_X4 FILLER_37_1174 ();
 FILLCELL_X4 FILLER_37_1182 ();
 FILLCELL_X4 FILLER_37_1195 ();
 FILLCELL_X2 FILLER_37_1199 ();
 FILLCELL_X4 FILLER_37_1210 ();
 FILLCELL_X8 FILLER_37_1217 ();
 FILLCELL_X2 FILLER_37_1225 ();
 FILLCELL_X1 FILLER_37_1227 ();
 FILLCELL_X4 FILLER_37_1231 ();
 FILLCELL_X4 FILLER_37_1244 ();
 FILLCELL_X1 FILLER_37_1248 ();
 FILLCELL_X4 FILLER_37_1259 ();
 FILLCELL_X4 FILLER_37_1264 ();
 FILLCELL_X4 FILLER_37_1278 ();
 FILLCELL_X4 FILLER_37_1291 ();
 FILLCELL_X4 FILLER_37_1298 ();
 FILLCELL_X1 FILLER_37_1302 ();
 FILLCELL_X4 FILLER_37_1307 ();
 FILLCELL_X4 FILLER_37_1314 ();
 FILLCELL_X4 FILLER_37_1321 ();
 FILLCELL_X4 FILLER_37_1335 ();
 FILLCELL_X1 FILLER_37_1339 ();
 FILLCELL_X4 FILLER_37_1344 ();
 FILLCELL_X4 FILLER_37_1357 ();
 FILLCELL_X8 FILLER_37_1365 ();
 FILLCELL_X1 FILLER_37_1373 ();
 FILLCELL_X32 FILLER_37_1378 ();
 FILLCELL_X2 FILLER_37_1410 ();
 FILLCELL_X1 FILLER_37_1412 ();
 FILLCELL_X4 FILLER_37_1420 ();
 FILLCELL_X32 FILLER_37_1441 ();
 FILLCELL_X32 FILLER_37_1473 ();
 FILLCELL_X32 FILLER_37_1505 ();
 FILLCELL_X32 FILLER_37_1537 ();
 FILLCELL_X32 FILLER_37_1569 ();
 FILLCELL_X32 FILLER_37_1601 ();
 FILLCELL_X32 FILLER_37_1633 ();
 FILLCELL_X32 FILLER_37_1665 ();
 FILLCELL_X32 FILLER_37_1697 ();
 FILLCELL_X32 FILLER_37_1729 ();
 FILLCELL_X1 FILLER_37_1761 ();
 FILLCELL_X16 FILLER_38_1 ();
 FILLCELL_X4 FILLER_38_17 ();
 FILLCELL_X4 FILLER_38_25 ();
 FILLCELL_X2 FILLER_38_29 ();
 FILLCELL_X8 FILLER_38_34 ();
 FILLCELL_X4 FILLER_38_42 ();
 FILLCELL_X1 FILLER_38_46 ();
 FILLCELL_X4 FILLER_38_57 ();
 FILLCELL_X4 FILLER_38_64 ();
 FILLCELL_X2 FILLER_38_68 ();
 FILLCELL_X8 FILLER_38_73 ();
 FILLCELL_X4 FILLER_38_81 ();
 FILLCELL_X2 FILLER_38_85 ();
 FILLCELL_X1 FILLER_38_87 ();
 FILLCELL_X4 FILLER_38_97 ();
 FILLCELL_X4 FILLER_38_104 ();
 FILLCELL_X2 FILLER_38_108 ();
 FILLCELL_X4 FILLER_38_114 ();
 FILLCELL_X4 FILLER_38_125 ();
 FILLCELL_X16 FILLER_38_139 ();
 FILLCELL_X4 FILLER_38_155 ();
 FILLCELL_X1 FILLER_38_159 ();
 FILLCELL_X4 FILLER_38_164 ();
 FILLCELL_X2 FILLER_38_168 ();
 FILLCELL_X1 FILLER_38_170 ();
 FILLCELL_X4 FILLER_38_174 ();
 FILLCELL_X4 FILLER_38_182 ();
 FILLCELL_X4 FILLER_38_190 ();
 FILLCELL_X1 FILLER_38_194 ();
 FILLCELL_X4 FILLER_38_199 ();
 FILLCELL_X4 FILLER_38_222 ();
 FILLCELL_X8 FILLER_38_229 ();
 FILLCELL_X8 FILLER_38_240 ();
 FILLCELL_X4 FILLER_38_252 ();
 FILLCELL_X16 FILLER_38_260 ();
 FILLCELL_X2 FILLER_38_276 ();
 FILLCELL_X1 FILLER_38_278 ();
 FILLCELL_X16 FILLER_38_286 ();
 FILLCELL_X4 FILLER_38_306 ();
 FILLCELL_X8 FILLER_38_313 ();
 FILLCELL_X4 FILLER_38_321 ();
 FILLCELL_X2 FILLER_38_325 ();
 FILLCELL_X4 FILLER_38_337 ();
 FILLCELL_X2 FILLER_38_341 ();
 FILLCELL_X4 FILLER_38_347 ();
 FILLCELL_X8 FILLER_38_361 ();
 FILLCELL_X2 FILLER_38_369 ();
 FILLCELL_X1 FILLER_38_371 ();
 FILLCELL_X4 FILLER_38_381 ();
 FILLCELL_X4 FILLER_38_389 ();
 FILLCELL_X1 FILLER_38_393 ();
 FILLCELL_X4 FILLER_38_403 ();
 FILLCELL_X16 FILLER_38_409 ();
 FILLCELL_X4 FILLER_38_425 ();
 FILLCELL_X4 FILLER_38_433 ();
 FILLCELL_X4 FILLER_38_440 ();
 FILLCELL_X2 FILLER_38_444 ();
 FILLCELL_X1 FILLER_38_446 ();
 FILLCELL_X4 FILLER_38_453 ();
 FILLCELL_X4 FILLER_38_470 ();
 FILLCELL_X1 FILLER_38_474 ();
 FILLCELL_X8 FILLER_38_481 ();
 FILLCELL_X4 FILLER_38_499 ();
 FILLCELL_X2 FILLER_38_503 ();
 FILLCELL_X8 FILLER_38_515 ();
 FILLCELL_X4 FILLER_38_527 ();
 FILLCELL_X4 FILLER_38_540 ();
 FILLCELL_X8 FILLER_38_553 ();
 FILLCELL_X1 FILLER_38_561 ();
 FILLCELL_X4 FILLER_38_581 ();
 FILLCELL_X4 FILLER_38_604 ();
 FILLCELL_X4 FILLER_38_627 ();
 FILLCELL_X8 FILLER_38_632 ();
 FILLCELL_X4 FILLER_38_640 ();
 FILLCELL_X8 FILLER_38_663 ();
 FILLCELL_X1 FILLER_38_671 ();
 FILLCELL_X4 FILLER_38_676 ();
 FILLCELL_X8 FILLER_38_684 ();
 FILLCELL_X2 FILLER_38_692 ();
 FILLCELL_X4 FILLER_38_713 ();
 FILLCELL_X4 FILLER_38_721 ();
 FILLCELL_X8 FILLER_38_729 ();
 FILLCELL_X4 FILLER_38_737 ();
 FILLCELL_X2 FILLER_38_741 ();
 FILLCELL_X8 FILLER_38_747 ();
 FILLCELL_X4 FILLER_38_755 ();
 FILLCELL_X8 FILLER_38_763 ();
 FILLCELL_X2 FILLER_38_771 ();
 FILLCELL_X1 FILLER_38_773 ();
 FILLCELL_X8 FILLER_38_778 ();
 FILLCELL_X2 FILLER_38_786 ();
 FILLCELL_X1 FILLER_38_788 ();
 FILLCELL_X8 FILLER_38_793 ();
 FILLCELL_X4 FILLER_38_805 ();
 FILLCELL_X4 FILLER_38_813 ();
 FILLCELL_X2 FILLER_38_817 ();
 FILLCELL_X1 FILLER_38_819 ();
 FILLCELL_X32 FILLER_38_824 ();
 FILLCELL_X16 FILLER_38_856 ();
 FILLCELL_X8 FILLER_38_872 ();
 FILLCELL_X4 FILLER_38_880 ();
 FILLCELL_X2 FILLER_38_884 ();
 FILLCELL_X1 FILLER_38_886 ();
 FILLCELL_X16 FILLER_38_891 ();
 FILLCELL_X8 FILLER_38_907 ();
 FILLCELL_X2 FILLER_38_915 ();
 FILLCELL_X16 FILLER_38_921 ();
 FILLCELL_X1 FILLER_38_937 ();
 FILLCELL_X16 FILLER_38_940 ();
 FILLCELL_X8 FILLER_38_956 ();
 FILLCELL_X4 FILLER_38_968 ();
 FILLCELL_X1 FILLER_38_972 ();
 FILLCELL_X4 FILLER_38_992 ();
 FILLCELL_X2 FILLER_38_996 ();
 FILLCELL_X1 FILLER_38_998 ();
 FILLCELL_X32 FILLER_38_1018 ();
 FILLCELL_X8 FILLER_38_1050 ();
 FILLCELL_X4 FILLER_38_1058 ();
 FILLCELL_X2 FILLER_38_1062 ();
 FILLCELL_X1 FILLER_38_1064 ();
 FILLCELL_X16 FILLER_38_1069 ();
 FILLCELL_X8 FILLER_38_1085 ();
 FILLCELL_X1 FILLER_38_1093 ();
 FILLCELL_X16 FILLER_38_1097 ();
 FILLCELL_X1 FILLER_38_1113 ();
 FILLCELL_X16 FILLER_38_1119 ();
 FILLCELL_X8 FILLER_38_1135 ();
 FILLCELL_X2 FILLER_38_1143 ();
 FILLCELL_X4 FILLER_38_1149 ();
 FILLCELL_X8 FILLER_38_1157 ();
 FILLCELL_X2 FILLER_38_1165 ();
 FILLCELL_X1 FILLER_38_1167 ();
 FILLCELL_X8 FILLER_38_1187 ();
 FILLCELL_X2 FILLER_38_1195 ();
 FILLCELL_X4 FILLER_38_1200 ();
 FILLCELL_X1 FILLER_38_1204 ();
 FILLCELL_X4 FILLER_38_1209 ();
 FILLCELL_X16 FILLER_38_1217 ();
 FILLCELL_X4 FILLER_38_1233 ();
 FILLCELL_X4 FILLER_38_1241 ();
 FILLCELL_X8 FILLER_38_1249 ();
 FILLCELL_X2 FILLER_38_1257 ();
 FILLCELL_X8 FILLER_38_1261 ();
 FILLCELL_X2 FILLER_38_1269 ();
 FILLCELL_X16 FILLER_38_1274 ();
 FILLCELL_X2 FILLER_38_1290 ();
 FILLCELL_X1 FILLER_38_1292 ();
 FILLCELL_X4 FILLER_38_1296 ();
 FILLCELL_X4 FILLER_38_1309 ();
 FILLCELL_X8 FILLER_38_1317 ();
 FILLCELL_X8 FILLER_38_1329 ();
 FILLCELL_X2 FILLER_38_1337 ();
 FILLCELL_X1 FILLER_38_1339 ();
 FILLCELL_X4 FILLER_38_1349 ();
 FILLCELL_X4 FILLER_38_1356 ();
 FILLCELL_X1 FILLER_38_1360 ();
 FILLCELL_X4 FILLER_38_1365 ();
 FILLCELL_X8 FILLER_38_1388 ();
 FILLCELL_X4 FILLER_38_1396 ();
 FILLCELL_X1 FILLER_38_1400 ();
 FILLCELL_X4 FILLER_38_1405 ();
 FILLCELL_X4 FILLER_38_1413 ();
 FILLCELL_X4 FILLER_38_1422 ();
 FILLCELL_X32 FILLER_38_1428 ();
 FILLCELL_X32 FILLER_38_1460 ();
 FILLCELL_X32 FILLER_38_1492 ();
 FILLCELL_X32 FILLER_38_1524 ();
 FILLCELL_X32 FILLER_38_1556 ();
 FILLCELL_X32 FILLER_38_1588 ();
 FILLCELL_X32 FILLER_38_1620 ();
 FILLCELL_X32 FILLER_38_1652 ();
 FILLCELL_X32 FILLER_38_1684 ();
 FILLCELL_X32 FILLER_38_1716 ();
 FILLCELL_X8 FILLER_38_1748 ();
 FILLCELL_X4 FILLER_38_1756 ();
 FILLCELL_X2 FILLER_38_1760 ();
 FILLCELL_X16 FILLER_39_1 ();
 FILLCELL_X4 FILLER_39_17 ();
 FILLCELL_X2 FILLER_39_21 ();
 FILLCELL_X1 FILLER_39_23 ();
 FILLCELL_X4 FILLER_39_33 ();
 FILLCELL_X2 FILLER_39_37 ();
 FILLCELL_X16 FILLER_39_42 ();
 FILLCELL_X1 FILLER_39_58 ();
 FILLCELL_X8 FILLER_39_68 ();
 FILLCELL_X4 FILLER_39_76 ();
 FILLCELL_X2 FILLER_39_80 ();
 FILLCELL_X1 FILLER_39_82 ();
 FILLCELL_X4 FILLER_39_93 ();
 FILLCELL_X4 FILLER_39_107 ();
 FILLCELL_X8 FILLER_39_118 ();
 FILLCELL_X4 FILLER_39_126 ();
 FILLCELL_X1 FILLER_39_130 ();
 FILLCELL_X16 FILLER_39_135 ();
 FILLCELL_X2 FILLER_39_151 ();
 FILLCELL_X4 FILLER_39_157 ();
 FILLCELL_X4 FILLER_39_170 ();
 FILLCELL_X2 FILLER_39_174 ();
 FILLCELL_X1 FILLER_39_176 ();
 FILLCELL_X8 FILLER_39_180 ();
 FILLCELL_X16 FILLER_39_192 ();
 FILLCELL_X4 FILLER_39_208 ();
 FILLCELL_X4 FILLER_39_216 ();
 FILLCELL_X4 FILLER_39_229 ();
 FILLCELL_X4 FILLER_39_237 ();
 FILLCELL_X2 FILLER_39_241 ();
 FILLCELL_X1 FILLER_39_243 ();
 FILLCELL_X8 FILLER_39_261 ();
 FILLCELL_X4 FILLER_39_269 ();
 FILLCELL_X4 FILLER_39_283 ();
 FILLCELL_X8 FILLER_39_289 ();
 FILLCELL_X4 FILLER_39_297 ();
 FILLCELL_X4 FILLER_39_305 ();
 FILLCELL_X4 FILLER_39_312 ();
 FILLCELL_X2 FILLER_39_316 ();
 FILLCELL_X1 FILLER_39_318 ();
 FILLCELL_X4 FILLER_39_323 ();
 FILLCELL_X16 FILLER_39_336 ();
 FILLCELL_X4 FILLER_39_352 ();
 FILLCELL_X2 FILLER_39_356 ();
 FILLCELL_X1 FILLER_39_358 ();
 FILLCELL_X4 FILLER_39_361 ();
 FILLCELL_X4 FILLER_39_372 ();
 FILLCELL_X1 FILLER_39_376 ();
 FILLCELL_X4 FILLER_39_380 ();
 FILLCELL_X8 FILLER_39_393 ();
 FILLCELL_X4 FILLER_39_411 ();
 FILLCELL_X4 FILLER_39_422 ();
 FILLCELL_X1 FILLER_39_426 ();
 FILLCELL_X4 FILLER_39_437 ();
 FILLCELL_X8 FILLER_39_444 ();
 FILLCELL_X2 FILLER_39_452 ();
 FILLCELL_X4 FILLER_39_458 ();
 FILLCELL_X4 FILLER_39_466 ();
 FILLCELL_X2 FILLER_39_470 ();
 FILLCELL_X4 FILLER_39_474 ();
 FILLCELL_X4 FILLER_39_480 ();
 FILLCELL_X4 FILLER_39_487 ();
 FILLCELL_X1 FILLER_39_491 ();
 FILLCELL_X8 FILLER_39_496 ();
 FILLCELL_X2 FILLER_39_504 ();
 FILLCELL_X32 FILLER_39_509 ();
 FILLCELL_X16 FILLER_39_544 ();
 FILLCELL_X8 FILLER_39_560 ();
 FILLCELL_X2 FILLER_39_568 ();
 FILLCELL_X1 FILLER_39_570 ();
 FILLCELL_X16 FILLER_39_575 ();
 FILLCELL_X2 FILLER_39_591 ();
 FILLCELL_X16 FILLER_39_597 ();
 FILLCELL_X1 FILLER_39_613 ();
 FILLCELL_X4 FILLER_39_618 ();
 FILLCELL_X1 FILLER_39_622 ();
 FILLCELL_X4 FILLER_39_627 ();
 FILLCELL_X8 FILLER_39_632 ();
 FILLCELL_X2 FILLER_39_640 ();
 FILLCELL_X4 FILLER_39_646 ();
 FILLCELL_X32 FILLER_39_654 ();
 FILLCELL_X8 FILLER_39_686 ();
 FILLCELL_X4 FILLER_39_694 ();
 FILLCELL_X1 FILLER_39_698 ();
 FILLCELL_X32 FILLER_39_704 ();
 FILLCELL_X32 FILLER_39_736 ();
 FILLCELL_X4 FILLER_39_768 ();
 FILLCELL_X1 FILLER_39_772 ();
 FILLCELL_X32 FILLER_39_778 ();
 FILLCELL_X32 FILLER_39_810 ();
 FILLCELL_X4 FILLER_39_842 ();
 FILLCELL_X1 FILLER_39_846 ();
 FILLCELL_X32 FILLER_39_852 ();
 FILLCELL_X2 FILLER_39_884 ();
 FILLCELL_X1 FILLER_39_886 ();
 FILLCELL_X32 FILLER_39_890 ();
 FILLCELL_X32 FILLER_39_922 ();
 FILLCELL_X32 FILLER_39_954 ();
 FILLCELL_X32 FILLER_39_986 ();
 FILLCELL_X32 FILLER_39_1018 ();
 FILLCELL_X32 FILLER_39_1050 ();
 FILLCELL_X32 FILLER_39_1082 ();
 FILLCELL_X32 FILLER_39_1114 ();
 FILLCELL_X32 FILLER_39_1146 ();
 FILLCELL_X32 FILLER_39_1178 ();
 FILLCELL_X32 FILLER_39_1210 ();
 FILLCELL_X16 FILLER_39_1242 ();
 FILLCELL_X4 FILLER_39_1258 ();
 FILLCELL_X32 FILLER_39_1263 ();
 FILLCELL_X32 FILLER_39_1295 ();
 FILLCELL_X4 FILLER_39_1327 ();
 FILLCELL_X2 FILLER_39_1331 ();
 FILLCELL_X1 FILLER_39_1333 ();
 FILLCELL_X32 FILLER_39_1338 ();
 FILLCELL_X16 FILLER_39_1370 ();
 FILLCELL_X4 FILLER_39_1386 ();
 FILLCELL_X1 FILLER_39_1390 ();
 FILLCELL_X4 FILLER_39_1396 ();
 FILLCELL_X8 FILLER_39_1403 ();
 FILLCELL_X2 FILLER_39_1411 ();
 FILLCELL_X1 FILLER_39_1413 ();
 FILLCELL_X4 FILLER_39_1418 ();
 FILLCELL_X2 FILLER_39_1422 ();
 FILLCELL_X32 FILLER_39_1427 ();
 FILLCELL_X32 FILLER_39_1459 ();
 FILLCELL_X32 FILLER_39_1491 ();
 FILLCELL_X32 FILLER_39_1523 ();
 FILLCELL_X32 FILLER_39_1555 ();
 FILLCELL_X32 FILLER_39_1587 ();
 FILLCELL_X32 FILLER_39_1619 ();
 FILLCELL_X32 FILLER_39_1651 ();
 FILLCELL_X32 FILLER_39_1683 ();
 FILLCELL_X32 FILLER_39_1715 ();
 FILLCELL_X8 FILLER_39_1747 ();
 FILLCELL_X4 FILLER_39_1755 ();
 FILLCELL_X2 FILLER_39_1759 ();
 FILLCELL_X1 FILLER_39_1761 ();
 FILLCELL_X8 FILLER_40_1 ();
 FILLCELL_X4 FILLER_40_9 ();
 FILLCELL_X2 FILLER_40_13 ();
 FILLCELL_X4 FILLER_40_19 ();
 FILLCELL_X4 FILLER_40_27 ();
 FILLCELL_X4 FILLER_40_40 ();
 FILLCELL_X4 FILLER_40_47 ();
 FILLCELL_X4 FILLER_40_55 ();
 FILLCELL_X4 FILLER_40_68 ();
 FILLCELL_X4 FILLER_40_76 ();
 FILLCELL_X8 FILLER_40_83 ();
 FILLCELL_X1 FILLER_40_91 ();
 FILLCELL_X16 FILLER_40_94 ();
 FILLCELL_X2 FILLER_40_110 ();
 FILLCELL_X4 FILLER_40_122 ();
 FILLCELL_X4 FILLER_40_130 ();
 FILLCELL_X1 FILLER_40_134 ();
 FILLCELL_X4 FILLER_40_144 ();
 FILLCELL_X4 FILLER_40_152 ();
 FILLCELL_X1 FILLER_40_156 ();
 FILLCELL_X4 FILLER_40_166 ();
 FILLCELL_X8 FILLER_40_174 ();
 FILLCELL_X4 FILLER_40_186 ();
 FILLCELL_X8 FILLER_40_199 ();
 FILLCELL_X4 FILLER_40_207 ();
 FILLCELL_X2 FILLER_40_211 ();
 FILLCELL_X1 FILLER_40_213 ();
 FILLCELL_X4 FILLER_40_218 ();
 FILLCELL_X4 FILLER_40_231 ();
 FILLCELL_X8 FILLER_40_238 ();
 FILLCELL_X4 FILLER_40_246 ();
 FILLCELL_X4 FILLER_40_260 ();
 FILLCELL_X4 FILLER_40_267 ();
 FILLCELL_X2 FILLER_40_271 ();
 FILLCELL_X8 FILLER_40_276 ();
 FILLCELL_X2 FILLER_40_284 ();
 FILLCELL_X4 FILLER_40_293 ();
 FILLCELL_X4 FILLER_40_307 ();
 FILLCELL_X4 FILLER_40_316 ();
 FILLCELL_X4 FILLER_40_323 ();
 FILLCELL_X4 FILLER_40_331 ();
 FILLCELL_X8 FILLER_40_338 ();
 FILLCELL_X4 FILLER_40_346 ();
 FILLCELL_X4 FILLER_40_360 ();
 FILLCELL_X4 FILLER_40_374 ();
 FILLCELL_X2 FILLER_40_378 ();
 FILLCELL_X32 FILLER_40_1518 ();
 FILLCELL_X32 FILLER_40_1550 ();
 FILLCELL_X32 FILLER_40_1582 ();
 FILLCELL_X32 FILLER_40_1614 ();
 FILLCELL_X32 FILLER_40_1646 ();
 FILLCELL_X32 FILLER_40_1678 ();
 FILLCELL_X32 FILLER_40_1710 ();
 FILLCELL_X16 FILLER_40_1742 ();
 FILLCELL_X4 FILLER_40_1758 ();
 FILLCELL_X16 FILLER_41_1 ();
 FILLCELL_X8 FILLER_41_17 ();
 FILLCELL_X4 FILLER_41_25 ();
 FILLCELL_X2 FILLER_41_29 ();
 FILLCELL_X1 FILLER_41_31 ();
 FILLCELL_X16 FILLER_41_36 ();
 FILLCELL_X4 FILLER_41_52 ();
 FILLCELL_X8 FILLER_41_60 ();
 FILLCELL_X4 FILLER_41_71 ();
 FILLCELL_X8 FILLER_41_78 ();
 FILLCELL_X2 FILLER_41_86 ();
 FILLCELL_X1 FILLER_41_88 ();
 FILLCELL_X16 FILLER_41_98 ();
 FILLCELL_X1 FILLER_41_114 ();
 FILLCELL_X4 FILLER_41_118 ();
 FILLCELL_X4 FILLER_41_124 ();
 FILLCELL_X2 FILLER_41_128 ();
 FILLCELL_X4 FILLER_41_134 ();
 FILLCELL_X1 FILLER_41_138 ();
 FILLCELL_X4 FILLER_41_142 ();
 FILLCELL_X32 FILLER_41_149 ();
 FILLCELL_X4 FILLER_41_181 ();
 FILLCELL_X4 FILLER_41_189 ();
 FILLCELL_X4 FILLER_41_202 ();
 FILLCELL_X8 FILLER_41_209 ();
 FILLCELL_X4 FILLER_41_217 ();
 FILLCELL_X1 FILLER_41_221 ();
 FILLCELL_X8 FILLER_41_225 ();
 FILLCELL_X4 FILLER_41_233 ();
 FILLCELL_X2 FILLER_41_237 ();
 FILLCELL_X4 FILLER_41_241 ();
 FILLCELL_X4 FILLER_41_247 ();
 FILLCELL_X4 FILLER_41_258 ();
 FILLCELL_X4 FILLER_41_271 ();
 FILLCELL_X8 FILLER_41_285 ();
 FILLCELL_X1 FILLER_41_293 ();
 FILLCELL_X8 FILLER_41_303 ();
 FILLCELL_X1 FILLER_41_311 ();
 FILLCELL_X4 FILLER_41_315 ();
 FILLCELL_X4 FILLER_41_323 ();
 FILLCELL_X4 FILLER_41_336 ();
 FILLCELL_X4 FILLER_41_343 ();
 FILLCELL_X8 FILLER_41_351 ();
 FILLCELL_X2 FILLER_41_359 ();
 FILLCELL_X8 FILLER_41_365 ();
 FILLCELL_X4 FILLER_41_376 ();
 FILLCELL_X32 FILLER_41_1518 ();
 FILLCELL_X32 FILLER_41_1550 ();
 FILLCELL_X32 FILLER_41_1582 ();
 FILLCELL_X32 FILLER_41_1614 ();
 FILLCELL_X32 FILLER_41_1646 ();
 FILLCELL_X32 FILLER_41_1678 ();
 FILLCELL_X32 FILLER_41_1710 ();
 FILLCELL_X16 FILLER_41_1742 ();
 FILLCELL_X4 FILLER_41_1758 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X16 FILLER_42_33 ();
 FILLCELL_X8 FILLER_42_49 ();
 FILLCELL_X4 FILLER_42_57 ();
 FILLCELL_X2 FILLER_42_61 ();
 FILLCELL_X4 FILLER_42_67 ();
 FILLCELL_X4 FILLER_42_74 ();
 FILLCELL_X4 FILLER_42_82 ();
 FILLCELL_X4 FILLER_42_90 ();
 FILLCELL_X4 FILLER_42_103 ();
 FILLCELL_X8 FILLER_42_112 ();
 FILLCELL_X1 FILLER_42_120 ();
 FILLCELL_X4 FILLER_42_128 ();
 FILLCELL_X4 FILLER_42_137 ();
 FILLCELL_X2 FILLER_42_141 ();
 FILLCELL_X1 FILLER_42_143 ();
 FILLCELL_X4 FILLER_42_148 ();
 FILLCELL_X1 FILLER_42_152 ();
 FILLCELL_X4 FILLER_42_157 ();
 FILLCELL_X1 FILLER_42_161 ();
 FILLCELL_X4 FILLER_42_166 ();
 FILLCELL_X16 FILLER_42_173 ();
 FILLCELL_X4 FILLER_42_189 ();
 FILLCELL_X4 FILLER_42_196 ();
 FILLCELL_X8 FILLER_42_203 ();
 FILLCELL_X1 FILLER_42_211 ();
 FILLCELL_X4 FILLER_42_216 ();
 FILLCELL_X4 FILLER_42_230 ();
 FILLCELL_X4 FILLER_42_241 ();
 FILLCELL_X4 FILLER_42_255 ();
 FILLCELL_X8 FILLER_42_262 ();
 FILLCELL_X1 FILLER_42_270 ();
 FILLCELL_X8 FILLER_42_274 ();
 FILLCELL_X4 FILLER_42_282 ();
 FILLCELL_X1 FILLER_42_286 ();
 FILLCELL_X8 FILLER_42_289 ();
 FILLCELL_X1 FILLER_42_297 ();
 FILLCELL_X4 FILLER_42_307 ();
 FILLCELL_X8 FILLER_42_314 ();
 FILLCELL_X4 FILLER_42_322 ();
 FILLCELL_X2 FILLER_42_326 ();
 FILLCELL_X4 FILLER_42_331 ();
 FILLCELL_X4 FILLER_42_338 ();
 FILLCELL_X4 FILLER_42_351 ();
 FILLCELL_X4 FILLER_42_364 ();
 FILLCELL_X2 FILLER_42_368 ();
 FILLCELL_X1 FILLER_42_370 ();
 FILLCELL_X4 FILLER_42_376 ();
 FILLCELL_X32 FILLER_42_1518 ();
 FILLCELL_X32 FILLER_42_1550 ();
 FILLCELL_X32 FILLER_42_1582 ();
 FILLCELL_X32 FILLER_42_1614 ();
 FILLCELL_X32 FILLER_42_1646 ();
 FILLCELL_X32 FILLER_42_1678 ();
 FILLCELL_X32 FILLER_42_1710 ();
 FILLCELL_X16 FILLER_42_1742 ();
 FILLCELL_X4 FILLER_42_1758 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X16 FILLER_43_33 ();
 FILLCELL_X4 FILLER_43_49 ();
 FILLCELL_X2 FILLER_43_53 ();
 FILLCELL_X1 FILLER_43_55 ();
 FILLCELL_X4 FILLER_43_60 ();
 FILLCELL_X4 FILLER_43_73 ();
 FILLCELL_X8 FILLER_43_80 ();
 FILLCELL_X2 FILLER_43_88 ();
 FILLCELL_X1 FILLER_43_90 ();
 FILLCELL_X4 FILLER_43_94 ();
 FILLCELL_X8 FILLER_43_101 ();
 FILLCELL_X4 FILLER_43_109 ();
 FILLCELL_X8 FILLER_43_130 ();
 FILLCELL_X4 FILLER_43_138 ();
 FILLCELL_X4 FILLER_43_151 ();
 FILLCELL_X2 FILLER_43_155 ();
 FILLCELL_X4 FILLER_43_161 ();
 FILLCELL_X4 FILLER_43_174 ();
 FILLCELL_X4 FILLER_43_181 ();
 FILLCELL_X4 FILLER_43_187 ();
 FILLCELL_X2 FILLER_43_191 ();
 FILLCELL_X1 FILLER_43_193 ();
 FILLCELL_X16 FILLER_43_198 ();
 FILLCELL_X1 FILLER_43_214 ();
 FILLCELL_X4 FILLER_43_217 ();
 FILLCELL_X8 FILLER_43_231 ();
 FILLCELL_X1 FILLER_43_239 ();
 FILLCELL_X4 FILLER_43_244 ();
 FILLCELL_X16 FILLER_43_257 ();
 FILLCELL_X4 FILLER_43_282 ();
 FILLCELL_X4 FILLER_43_291 ();
 FILLCELL_X4 FILLER_43_298 ();
 FILLCELL_X4 FILLER_43_306 ();
 FILLCELL_X2 FILLER_43_310 ();
 FILLCELL_X4 FILLER_43_314 ();
 FILLCELL_X4 FILLER_43_321 ();
 FILLCELL_X4 FILLER_43_335 ();
 FILLCELL_X1 FILLER_43_339 ();
 FILLCELL_X4 FILLER_43_343 ();
 FILLCELL_X8 FILLER_43_351 ();
 FILLCELL_X8 FILLER_43_363 ();
 FILLCELL_X4 FILLER_43_375 ();
 FILLCELL_X1 FILLER_43_379 ();
 FILLCELL_X32 FILLER_43_1518 ();
 FILLCELL_X32 FILLER_43_1550 ();
 FILLCELL_X32 FILLER_43_1582 ();
 FILLCELL_X32 FILLER_43_1614 ();
 FILLCELL_X32 FILLER_43_1646 ();
 FILLCELL_X32 FILLER_43_1678 ();
 FILLCELL_X32 FILLER_43_1710 ();
 FILLCELL_X16 FILLER_43_1742 ();
 FILLCELL_X4 FILLER_43_1758 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X8 FILLER_44_33 ();
 FILLCELL_X4 FILLER_44_41 ();
 FILLCELL_X1 FILLER_44_45 ();
 FILLCELL_X8 FILLER_44_50 ();
 FILLCELL_X2 FILLER_44_58 ();
 FILLCELL_X4 FILLER_44_64 ();
 FILLCELL_X4 FILLER_44_77 ();
 FILLCELL_X16 FILLER_44_84 ();
 FILLCELL_X8 FILLER_44_100 ();
 FILLCELL_X4 FILLER_44_108 ();
 FILLCELL_X2 FILLER_44_112 ();
 FILLCELL_X4 FILLER_44_118 ();
 FILLCELL_X4 FILLER_44_127 ();
 FILLCELL_X8 FILLER_44_135 ();
 FILLCELL_X1 FILLER_44_143 ();
 FILLCELL_X8 FILLER_44_147 ();
 FILLCELL_X2 FILLER_44_155 ();
 FILLCELL_X4 FILLER_44_160 ();
 FILLCELL_X4 FILLER_44_168 ();
 FILLCELL_X4 FILLER_44_181 ();
 FILLCELL_X2 FILLER_44_185 ();
 FILLCELL_X4 FILLER_44_190 ();
 FILLCELL_X4 FILLER_44_204 ();
 FILLCELL_X16 FILLER_44_215 ();
 FILLCELL_X8 FILLER_44_231 ();
 FILLCELL_X2 FILLER_44_239 ();
 FILLCELL_X4 FILLER_44_244 ();
 FILLCELL_X1 FILLER_44_248 ();
 FILLCELL_X4 FILLER_44_251 ();
 FILLCELL_X2 FILLER_44_255 ();
 FILLCELL_X1 FILLER_44_257 ();
 FILLCELL_X4 FILLER_44_261 ();
 FILLCELL_X4 FILLER_44_268 ();
 FILLCELL_X4 FILLER_44_281 ();
 FILLCELL_X8 FILLER_44_289 ();
 FILLCELL_X1 FILLER_44_297 ();
 FILLCELL_X4 FILLER_44_308 ();
 FILLCELL_X4 FILLER_44_322 ();
 FILLCELL_X4 FILLER_44_333 ();
 FILLCELL_X8 FILLER_44_341 ();
 FILLCELL_X4 FILLER_44_352 ();
 FILLCELL_X4 FILLER_44_359 ();
 FILLCELL_X4 FILLER_44_366 ();
 FILLCELL_X1 FILLER_44_370 ();
 FILLCELL_X4 FILLER_44_376 ();
 FILLCELL_X32 FILLER_44_1518 ();
 FILLCELL_X32 FILLER_44_1550 ();
 FILLCELL_X32 FILLER_44_1582 ();
 FILLCELL_X32 FILLER_44_1614 ();
 FILLCELL_X32 FILLER_44_1646 ();
 FILLCELL_X32 FILLER_44_1678 ();
 FILLCELL_X32 FILLER_44_1710 ();
 FILLCELL_X16 FILLER_44_1742 ();
 FILLCELL_X4 FILLER_44_1758 ();
 FILLCELL_X4 FILLER_45_1 ();
 FILLCELL_X32 FILLER_45_8 ();
 FILLCELL_X16 FILLER_45_40 ();
 FILLCELL_X8 FILLER_45_56 ();
 FILLCELL_X2 FILLER_45_64 ();
 FILLCELL_X1 FILLER_45_66 ();
 FILLCELL_X4 FILLER_45_70 ();
 FILLCELL_X8 FILLER_45_84 ();
 FILLCELL_X2 FILLER_45_92 ();
 FILLCELL_X1 FILLER_45_94 ();
 FILLCELL_X4 FILLER_45_99 ();
 FILLCELL_X4 FILLER_45_107 ();
 FILLCELL_X4 FILLER_45_114 ();
 FILLCELL_X1 FILLER_45_118 ();
 FILLCELL_X8 FILLER_45_123 ();
 FILLCELL_X4 FILLER_45_131 ();
 FILLCELL_X2 FILLER_45_135 ();
 FILLCELL_X1 FILLER_45_137 ();
 FILLCELL_X4 FILLER_45_142 ();
 FILLCELL_X8 FILLER_45_150 ();
 FILLCELL_X4 FILLER_45_162 ();
 FILLCELL_X8 FILLER_45_185 ();
 FILLCELL_X1 FILLER_45_193 ();
 FILLCELL_X8 FILLER_45_204 ();
 FILLCELL_X4 FILLER_45_222 ();
 FILLCELL_X4 FILLER_45_229 ();
 FILLCELL_X4 FILLER_45_242 ();
 FILLCELL_X1 FILLER_45_246 ();
 FILLCELL_X4 FILLER_45_257 ();
 FILLCELL_X2 FILLER_45_261 ();
 FILLCELL_X4 FILLER_45_268 ();
 FILLCELL_X4 FILLER_45_279 ();
 FILLCELL_X8 FILLER_45_293 ();
 FILLCELL_X2 FILLER_45_301 ();
 FILLCELL_X4 FILLER_45_306 ();
 FILLCELL_X2 FILLER_45_310 ();
 FILLCELL_X8 FILLER_45_315 ();
 FILLCELL_X1 FILLER_45_323 ();
 FILLCELL_X4 FILLER_45_329 ();
 FILLCELL_X2 FILLER_45_333 ();
 FILLCELL_X1 FILLER_45_335 ();
 FILLCELL_X4 FILLER_45_345 ();
 FILLCELL_X2 FILLER_45_349 ();
 FILLCELL_X1 FILLER_45_351 ();
 FILLCELL_X4 FILLER_45_355 ();
 FILLCELL_X4 FILLER_45_363 ();
 FILLCELL_X4 FILLER_45_376 ();
 FILLCELL_X32 FILLER_45_1518 ();
 FILLCELL_X32 FILLER_45_1550 ();
 FILLCELL_X32 FILLER_45_1582 ();
 FILLCELL_X32 FILLER_45_1614 ();
 FILLCELL_X32 FILLER_45_1646 ();
 FILLCELL_X32 FILLER_45_1678 ();
 FILLCELL_X32 FILLER_45_1710 ();
 FILLCELL_X16 FILLER_45_1742 ();
 FILLCELL_X4 FILLER_45_1758 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X16 FILLER_46_33 ();
 FILLCELL_X2 FILLER_46_49 ();
 FILLCELL_X4 FILLER_46_54 ();
 FILLCELL_X4 FILLER_46_61 ();
 FILLCELL_X8 FILLER_46_68 ();
 FILLCELL_X16 FILLER_46_80 ();
 FILLCELL_X1 FILLER_46_96 ();
 FILLCELL_X8 FILLER_46_106 ();
 FILLCELL_X1 FILLER_46_114 ();
 FILLCELL_X8 FILLER_46_134 ();
 FILLCELL_X2 FILLER_46_142 ();
 FILLCELL_X4 FILLER_46_153 ();
 FILLCELL_X32 FILLER_46_161 ();
 FILLCELL_X8 FILLER_46_193 ();
 FILLCELL_X4 FILLER_46_203 ();
 FILLCELL_X4 FILLER_46_211 ();
 FILLCELL_X4 FILLER_46_225 ();
 FILLCELL_X8 FILLER_46_238 ();
 FILLCELL_X4 FILLER_46_249 ();
 FILLCELL_X4 FILLER_46_262 ();
 FILLCELL_X4 FILLER_46_269 ();
 FILLCELL_X8 FILLER_46_275 ();
 FILLCELL_X2 FILLER_46_283 ();
 FILLCELL_X4 FILLER_46_288 ();
 FILLCELL_X1 FILLER_46_292 ();
 FILLCELL_X4 FILLER_46_295 ();
 FILLCELL_X4 FILLER_46_306 ();
 FILLCELL_X4 FILLER_46_319 ();
 FILLCELL_X8 FILLER_46_326 ();
 FILLCELL_X4 FILLER_46_334 ();
 FILLCELL_X2 FILLER_46_338 ();
 FILLCELL_X4 FILLER_46_344 ();
 FILLCELL_X8 FILLER_46_357 ();
 FILLCELL_X2 FILLER_46_365 ();
 FILLCELL_X4 FILLER_46_376 ();
 FILLCELL_X32 FILLER_46_1518 ();
 FILLCELL_X32 FILLER_46_1550 ();
 FILLCELL_X32 FILLER_46_1582 ();
 FILLCELL_X32 FILLER_46_1614 ();
 FILLCELL_X32 FILLER_46_1646 ();
 FILLCELL_X32 FILLER_46_1678 ();
 FILLCELL_X32 FILLER_46_1710 ();
 FILLCELL_X16 FILLER_46_1742 ();
 FILLCELL_X4 FILLER_46_1758 ();
 FILLCELL_X32 FILLER_47_1 ();
 FILLCELL_X4 FILLER_47_33 ();
 FILLCELL_X2 FILLER_47_37 ();
 FILLCELL_X4 FILLER_47_43 ();
 FILLCELL_X4 FILLER_47_56 ();
 FILLCELL_X4 FILLER_47_62 ();
 FILLCELL_X4 FILLER_47_73 ();
 FILLCELL_X8 FILLER_47_87 ();
 FILLCELL_X4 FILLER_47_104 ();
 FILLCELL_X8 FILLER_47_112 ();
 FILLCELL_X1 FILLER_47_120 ();
 FILLCELL_X4 FILLER_47_125 ();
 FILLCELL_X2 FILLER_47_129 ();
 FILLCELL_X1 FILLER_47_131 ();
 FILLCELL_X4 FILLER_47_135 ();
 FILLCELL_X8 FILLER_47_148 ();
 FILLCELL_X1 FILLER_47_156 ();
 FILLCELL_X4 FILLER_47_160 ();
 FILLCELL_X2 FILLER_47_164 ();
 FILLCELL_X8 FILLER_47_170 ();
 FILLCELL_X4 FILLER_47_187 ();
 FILLCELL_X16 FILLER_47_194 ();
 FILLCELL_X4 FILLER_47_210 ();
 FILLCELL_X2 FILLER_47_214 ();
 FILLCELL_X8 FILLER_47_223 ();
 FILLCELL_X4 FILLER_47_234 ();
 FILLCELL_X8 FILLER_47_241 ();
 FILLCELL_X1 FILLER_47_249 ();
 FILLCELL_X16 FILLER_47_259 ();
 FILLCELL_X8 FILLER_47_275 ();
 FILLCELL_X1 FILLER_47_283 ();
 FILLCELL_X8 FILLER_47_291 ();
 FILLCELL_X16 FILLER_47_309 ();
 FILLCELL_X8 FILLER_47_334 ();
 FILLCELL_X4 FILLER_47_342 ();
 FILLCELL_X1 FILLER_47_346 ();
 FILLCELL_X8 FILLER_47_350 ();
 FILLCELL_X4 FILLER_47_358 ();
 FILLCELL_X4 FILLER_47_366 ();
 FILLCELL_X4 FILLER_47_374 ();
 FILLCELL_X2 FILLER_47_378 ();
 FILLCELL_X4 FILLER_47_1518 ();
 FILLCELL_X32 FILLER_47_1541 ();
 FILLCELL_X32 FILLER_47_1573 ();
 FILLCELL_X32 FILLER_47_1605 ();
 FILLCELL_X32 FILLER_47_1637 ();
 FILLCELL_X32 FILLER_47_1669 ();
 FILLCELL_X32 FILLER_47_1701 ();
 FILLCELL_X16 FILLER_47_1733 ();
 FILLCELL_X8 FILLER_47_1749 ();
 FILLCELL_X4 FILLER_47_1757 ();
 FILLCELL_X1 FILLER_47_1761 ();
 FILLCELL_X32 FILLER_48_1 ();
 FILLCELL_X8 FILLER_48_33 ();
 FILLCELL_X1 FILLER_48_41 ();
 FILLCELL_X4 FILLER_48_46 ();
 FILLCELL_X8 FILLER_48_59 ();
 FILLCELL_X4 FILLER_48_67 ();
 FILLCELL_X16 FILLER_48_75 ();
 FILLCELL_X8 FILLER_48_91 ();
 FILLCELL_X4 FILLER_48_102 ();
 FILLCELL_X4 FILLER_48_108 ();
 FILLCELL_X4 FILLER_48_115 ();
 FILLCELL_X1 FILLER_48_119 ();
 FILLCELL_X4 FILLER_48_130 ();
 FILLCELL_X8 FILLER_48_137 ();
 FILLCELL_X1 FILLER_48_145 ();
 FILLCELL_X4 FILLER_48_149 ();
 FILLCELL_X1 FILLER_48_153 ();
 FILLCELL_X4 FILLER_48_157 ();
 FILLCELL_X4 FILLER_48_166 ();
 FILLCELL_X4 FILLER_48_174 ();
 FILLCELL_X4 FILLER_48_187 ();
 FILLCELL_X4 FILLER_48_194 ();
 FILLCELL_X1 FILLER_48_198 ();
 FILLCELL_X4 FILLER_48_203 ();
 FILLCELL_X8 FILLER_48_211 ();
 FILLCELL_X4 FILLER_48_219 ();
 FILLCELL_X1 FILLER_48_223 ();
 FILLCELL_X4 FILLER_48_228 ();
 FILLCELL_X4 FILLER_48_239 ();
 FILLCELL_X4 FILLER_48_246 ();
 FILLCELL_X8 FILLER_48_252 ();
 FILLCELL_X4 FILLER_48_264 ();
 FILLCELL_X2 FILLER_48_268 ();
 FILLCELL_X4 FILLER_48_280 ();
 FILLCELL_X4 FILLER_48_294 ();
 FILLCELL_X1 FILLER_48_298 ();
 FILLCELL_X4 FILLER_48_302 ();
 FILLCELL_X4 FILLER_48_309 ();
 FILLCELL_X8 FILLER_48_318 ();
 FILLCELL_X4 FILLER_48_326 ();
 FILLCELL_X4 FILLER_48_332 ();
 FILLCELL_X4 FILLER_48_339 ();
 FILLCELL_X4 FILLER_48_347 ();
 FILLCELL_X1 FILLER_48_351 ();
 FILLCELL_X4 FILLER_48_355 ();
 FILLCELL_X4 FILLER_48_369 ();
 FILLCELL_X4 FILLER_48_376 ();
 FILLCELL_X32 FILLER_48_1518 ();
 FILLCELL_X32 FILLER_48_1550 ();
 FILLCELL_X32 FILLER_48_1582 ();
 FILLCELL_X32 FILLER_48_1614 ();
 FILLCELL_X32 FILLER_48_1646 ();
 FILLCELL_X32 FILLER_48_1678 ();
 FILLCELL_X32 FILLER_48_1710 ();
 FILLCELL_X16 FILLER_48_1742 ();
 FILLCELL_X4 FILLER_48_1758 ();
 FILLCELL_X32 FILLER_49_1 ();
 FILLCELL_X16 FILLER_49_33 ();
 FILLCELL_X8 FILLER_49_49 ();
 FILLCELL_X4 FILLER_49_57 ();
 FILLCELL_X1 FILLER_49_61 ();
 FILLCELL_X4 FILLER_49_66 ();
 FILLCELL_X4 FILLER_49_79 ();
 FILLCELL_X16 FILLER_49_86 ();
 FILLCELL_X4 FILLER_49_102 ();
 FILLCELL_X1 FILLER_49_106 ();
 FILLCELL_X4 FILLER_49_117 ();
 FILLCELL_X8 FILLER_49_125 ();
 FILLCELL_X4 FILLER_49_133 ();
 FILLCELL_X4 FILLER_49_141 ();
 FILLCELL_X4 FILLER_49_149 ();
 FILLCELL_X4 FILLER_49_157 ();
 FILLCELL_X8 FILLER_49_164 ();
 FILLCELL_X4 FILLER_49_172 ();
 FILLCELL_X1 FILLER_49_176 ();
 FILLCELL_X4 FILLER_49_181 ();
 FILLCELL_X4 FILLER_49_188 ();
 FILLCELL_X2 FILLER_49_192 ();
 FILLCELL_X1 FILLER_49_194 ();
 FILLCELL_X4 FILLER_49_198 ();
 FILLCELL_X4 FILLER_49_211 ();
 FILLCELL_X4 FILLER_49_218 ();
 FILLCELL_X2 FILLER_49_222 ();
 FILLCELL_X1 FILLER_49_224 ();
 FILLCELL_X4 FILLER_49_227 ();
 FILLCELL_X4 FILLER_49_241 ();
 FILLCELL_X1 FILLER_49_245 ();
 FILLCELL_X4 FILLER_49_253 ();
 FILLCELL_X4 FILLER_49_267 ();
 FILLCELL_X4 FILLER_49_274 ();
 FILLCELL_X2 FILLER_49_278 ();
 FILLCELL_X4 FILLER_49_283 ();
 FILLCELL_X8 FILLER_49_289 ();
 FILLCELL_X4 FILLER_49_297 ();
 FILLCELL_X1 FILLER_49_301 ();
 FILLCELL_X8 FILLER_49_311 ();
 FILLCELL_X2 FILLER_49_319 ();
 FILLCELL_X4 FILLER_49_331 ();
 FILLCELL_X1 FILLER_49_335 ();
 FILLCELL_X4 FILLER_49_346 ();
 FILLCELL_X8 FILLER_49_357 ();
 FILLCELL_X1 FILLER_49_365 ();
 FILLCELL_X4 FILLER_49_376 ();
 FILLCELL_X32 FILLER_49_1518 ();
 FILLCELL_X32 FILLER_49_1550 ();
 FILLCELL_X32 FILLER_49_1582 ();
 FILLCELL_X32 FILLER_49_1614 ();
 FILLCELL_X32 FILLER_49_1646 ();
 FILLCELL_X32 FILLER_49_1678 ();
 FILLCELL_X32 FILLER_49_1710 ();
 FILLCELL_X16 FILLER_49_1742 ();
 FILLCELL_X4 FILLER_49_1758 ();
 FILLCELL_X16 FILLER_50_1 ();
 FILLCELL_X8 FILLER_50_17 ();
 FILLCELL_X2 FILLER_50_25 ();
 FILLCELL_X1 FILLER_50_27 ();
 FILLCELL_X4 FILLER_50_32 ();
 FILLCELL_X4 FILLER_50_40 ();
 FILLCELL_X1 FILLER_50_44 ();
 FILLCELL_X16 FILLER_50_49 ();
 FILLCELL_X1 FILLER_50_65 ();
 FILLCELL_X4 FILLER_50_75 ();
 FILLCELL_X8 FILLER_50_84 ();
 FILLCELL_X1 FILLER_50_92 ();
 FILLCELL_X4 FILLER_50_102 ();
 FILLCELL_X16 FILLER_50_109 ();
 FILLCELL_X8 FILLER_50_125 ();
 FILLCELL_X1 FILLER_50_133 ();
 FILLCELL_X4 FILLER_50_137 ();
 FILLCELL_X1 FILLER_50_141 ();
 FILLCELL_X4 FILLER_50_151 ();
 FILLCELL_X4 FILLER_50_164 ();
 FILLCELL_X4 FILLER_50_171 ();
 FILLCELL_X2 FILLER_50_175 ();
 FILLCELL_X4 FILLER_50_179 ();
 FILLCELL_X8 FILLER_50_185 ();
 FILLCELL_X4 FILLER_50_193 ();
 FILLCELL_X4 FILLER_50_201 ();
 FILLCELL_X4 FILLER_50_214 ();
 FILLCELL_X2 FILLER_50_218 ();
 FILLCELL_X4 FILLER_50_230 ();
 FILLCELL_X8 FILLER_50_244 ();
 FILLCELL_X1 FILLER_50_252 ();
 FILLCELL_X4 FILLER_50_257 ();
 FILLCELL_X4 FILLER_50_271 ();
 FILLCELL_X4 FILLER_50_278 ();
 FILLCELL_X2 FILLER_50_282 ();
 FILLCELL_X4 FILLER_50_288 ();
 FILLCELL_X8 FILLER_50_295 ();
 FILLCELL_X4 FILLER_50_303 ();
 FILLCELL_X2 FILLER_50_307 ();
 FILLCELL_X16 FILLER_50_318 ();
 FILLCELL_X1 FILLER_50_334 ();
 FILLCELL_X8 FILLER_50_337 ();
 FILLCELL_X4 FILLER_50_345 ();
 FILLCELL_X2 FILLER_50_349 ();
 FILLCELL_X1 FILLER_50_351 ();
 FILLCELL_X4 FILLER_50_355 ();
 FILLCELL_X4 FILLER_50_362 ();
 FILLCELL_X4 FILLER_50_368 ();
 FILLCELL_X1 FILLER_50_372 ();
 FILLCELL_X4 FILLER_50_375 ();
 FILLCELL_X1 FILLER_50_379 ();
 FILLCELL_X32 FILLER_50_1518 ();
 FILLCELL_X32 FILLER_50_1550 ();
 FILLCELL_X32 FILLER_50_1582 ();
 FILLCELL_X32 FILLER_50_1614 ();
 FILLCELL_X32 FILLER_50_1646 ();
 FILLCELL_X32 FILLER_50_1678 ();
 FILLCELL_X32 FILLER_50_1710 ();
 FILLCELL_X8 FILLER_50_1742 ();
 FILLCELL_X4 FILLER_50_1750 ();
 FILLCELL_X1 FILLER_50_1754 ();
 FILLCELL_X4 FILLER_50_1758 ();
 FILLCELL_X32 FILLER_51_1 ();
 FILLCELL_X4 FILLER_51_42 ();
 FILLCELL_X8 FILLER_51_49 ();
 FILLCELL_X4 FILLER_51_57 ();
 FILLCELL_X2 FILLER_51_61 ();
 FILLCELL_X1 FILLER_51_63 ();
 FILLCELL_X4 FILLER_51_68 ();
 FILLCELL_X8 FILLER_51_75 ();
 FILLCELL_X4 FILLER_51_83 ();
 FILLCELL_X2 FILLER_51_87 ();
 FILLCELL_X8 FILLER_51_98 ();
 FILLCELL_X4 FILLER_51_109 ();
 FILLCELL_X4 FILLER_51_116 ();
 FILLCELL_X2 FILLER_51_120 ();
 FILLCELL_X4 FILLER_51_132 ();
 FILLCELL_X2 FILLER_51_136 ();
 FILLCELL_X8 FILLER_51_141 ();
 FILLCELL_X4 FILLER_51_149 ();
 FILLCELL_X1 FILLER_51_153 ();
 FILLCELL_X8 FILLER_51_157 ();
 FILLCELL_X4 FILLER_51_165 ();
 FILLCELL_X2 FILLER_51_169 ();
 FILLCELL_X1 FILLER_51_171 ();
 FILLCELL_X4 FILLER_51_176 ();
 FILLCELL_X4 FILLER_51_190 ();
 FILLCELL_X8 FILLER_51_197 ();
 FILLCELL_X8 FILLER_51_208 ();
 FILLCELL_X4 FILLER_51_216 ();
 FILLCELL_X1 FILLER_51_220 ();
 FILLCELL_X16 FILLER_51_224 ();
 FILLCELL_X2 FILLER_51_240 ();
 FILLCELL_X1 FILLER_51_242 ();
 FILLCELL_X4 FILLER_51_245 ();
 FILLCELL_X4 FILLER_51_259 ();
 FILLCELL_X4 FILLER_51_270 ();
 FILLCELL_X2 FILLER_51_274 ();
 FILLCELL_X4 FILLER_51_285 ();
 FILLCELL_X4 FILLER_51_298 ();
 FILLCELL_X4 FILLER_51_306 ();
 FILLCELL_X4 FILLER_51_320 ();
 FILLCELL_X8 FILLER_51_327 ();
 FILLCELL_X1 FILLER_51_335 ();
 FILLCELL_X4 FILLER_51_346 ();
 FILLCELL_X4 FILLER_51_359 ();
 FILLCELL_X2 FILLER_51_363 ();
 FILLCELL_X1 FILLER_51_365 ();
 FILLCELL_X4 FILLER_51_376 ();
 FILLCELL_X32 FILLER_51_1518 ();
 FILLCELL_X32 FILLER_51_1550 ();
 FILLCELL_X32 FILLER_51_1582 ();
 FILLCELL_X32 FILLER_51_1614 ();
 FILLCELL_X32 FILLER_51_1646 ();
 FILLCELL_X32 FILLER_51_1678 ();
 FILLCELL_X32 FILLER_51_1710 ();
 FILLCELL_X16 FILLER_51_1742 ();
 FILLCELL_X4 FILLER_51_1758 ();
 FILLCELL_X16 FILLER_52_1 ();
 FILLCELL_X1 FILLER_52_17 ();
 FILLCELL_X4 FILLER_52_22 ();
 FILLCELL_X4 FILLER_52_35 ();
 FILLCELL_X4 FILLER_52_42 ();
 FILLCELL_X4 FILLER_52_50 ();
 FILLCELL_X4 FILLER_52_56 ();
 FILLCELL_X4 FILLER_52_63 ();
 FILLCELL_X4 FILLER_52_77 ();
 FILLCELL_X4 FILLER_52_88 ();
 FILLCELL_X2 FILLER_52_92 ();
 FILLCELL_X1 FILLER_52_94 ();
 FILLCELL_X4 FILLER_52_99 ();
 FILLCELL_X4 FILLER_52_107 ();
 FILLCELL_X1 FILLER_52_111 ();
 FILLCELL_X4 FILLER_52_114 ();
 FILLCELL_X4 FILLER_52_120 ();
 FILLCELL_X8 FILLER_52_131 ();
 FILLCELL_X4 FILLER_52_146 ();
 FILLCELL_X8 FILLER_52_153 ();
 FILLCELL_X4 FILLER_52_161 ();
 FILLCELL_X1 FILLER_52_165 ();
 FILLCELL_X4 FILLER_52_170 ();
 FILLCELL_X4 FILLER_52_177 ();
 FILLCELL_X2 FILLER_52_181 ();
 FILLCELL_X4 FILLER_52_193 ();
 FILLCELL_X2 FILLER_52_197 ();
 FILLCELL_X1 FILLER_52_199 ();
 FILLCELL_X8 FILLER_52_209 ();
 FILLCELL_X1 FILLER_52_217 ();
 FILLCELL_X4 FILLER_52_228 ();
 FILLCELL_X2 FILLER_52_232 ();
 FILLCELL_X4 FILLER_52_237 ();
 FILLCELL_X8 FILLER_52_243 ();
 FILLCELL_X4 FILLER_52_251 ();
 FILLCELL_X2 FILLER_52_255 ();
 FILLCELL_X1 FILLER_52_257 ();
 FILLCELL_X4 FILLER_52_261 ();
 FILLCELL_X1 FILLER_52_265 ();
 FILLCELL_X4 FILLER_52_269 ();
 FILLCELL_X8 FILLER_52_276 ();
 FILLCELL_X4 FILLER_52_287 ();
 FILLCELL_X16 FILLER_52_295 ();
 FILLCELL_X8 FILLER_52_311 ();
 FILLCELL_X4 FILLER_52_319 ();
 FILLCELL_X2 FILLER_52_323 ();
 FILLCELL_X4 FILLER_52_334 ();
 FILLCELL_X4 FILLER_52_341 ();
 FILLCELL_X2 FILLER_52_345 ();
 FILLCELL_X4 FILLER_52_350 ();
 FILLCELL_X8 FILLER_52_358 ();
 FILLCELL_X1 FILLER_52_366 ();
 FILLCELL_X8 FILLER_52_371 ();
 FILLCELL_X1 FILLER_52_379 ();
 FILLCELL_X32 FILLER_52_1518 ();
 FILLCELL_X32 FILLER_52_1550 ();
 FILLCELL_X32 FILLER_52_1582 ();
 FILLCELL_X32 FILLER_52_1614 ();
 FILLCELL_X32 FILLER_52_1646 ();
 FILLCELL_X32 FILLER_52_1678 ();
 FILLCELL_X32 FILLER_52_1710 ();
 FILLCELL_X16 FILLER_52_1742 ();
 FILLCELL_X4 FILLER_52_1758 ();
 FILLCELL_X16 FILLER_53_1 ();
 FILLCELL_X8 FILLER_53_17 ();
 FILLCELL_X4 FILLER_53_25 ();
 FILLCELL_X2 FILLER_53_29 ();
 FILLCELL_X1 FILLER_53_31 ();
 FILLCELL_X8 FILLER_53_35 ();
 FILLCELL_X4 FILLER_53_52 ();
 FILLCELL_X8 FILLER_53_59 ();
 FILLCELL_X4 FILLER_53_67 ();
 FILLCELL_X4 FILLER_53_81 ();
 FILLCELL_X2 FILLER_53_85 ();
 FILLCELL_X4 FILLER_53_91 ();
 FILLCELL_X8 FILLER_53_104 ();
 FILLCELL_X1 FILLER_53_112 ();
 FILLCELL_X4 FILLER_53_123 ();
 FILLCELL_X1 FILLER_53_127 ();
 FILLCELL_X4 FILLER_53_137 ();
 FILLCELL_X2 FILLER_53_141 ();
 FILLCELL_X4 FILLER_53_145 ();
 FILLCELL_X4 FILLER_53_159 ();
 FILLCELL_X1 FILLER_53_163 ();
 FILLCELL_X4 FILLER_53_174 ();
 FILLCELL_X4 FILLER_53_180 ();
 FILLCELL_X1 FILLER_53_184 ();
 FILLCELL_X8 FILLER_53_192 ();
 FILLCELL_X4 FILLER_53_200 ();
 FILLCELL_X4 FILLER_53_206 ();
 FILLCELL_X4 FILLER_53_213 ();
 FILLCELL_X4 FILLER_53_224 ();
 FILLCELL_X2 FILLER_53_228 ();
 FILLCELL_X4 FILLER_53_239 ();
 FILLCELL_X1 FILLER_53_243 ();
 FILLCELL_X4 FILLER_53_251 ();
 FILLCELL_X8 FILLER_53_264 ();
 FILLCELL_X1 FILLER_53_272 ();
 FILLCELL_X4 FILLER_53_276 ();
 FILLCELL_X16 FILLER_53_282 ();
 FILLCELL_X4 FILLER_53_298 ();
 FILLCELL_X4 FILLER_53_306 ();
 FILLCELL_X8 FILLER_53_317 ();
 FILLCELL_X4 FILLER_53_325 ();
 FILLCELL_X2 FILLER_53_329 ();
 FILLCELL_X1 FILLER_53_331 ();
 FILLCELL_X4 FILLER_53_342 ();
 FILLCELL_X8 FILLER_53_356 ();
 FILLCELL_X4 FILLER_53_374 ();
 FILLCELL_X2 FILLER_53_378 ();
 FILLCELL_X32 FILLER_53_1518 ();
 FILLCELL_X32 FILLER_53_1550 ();
 FILLCELL_X32 FILLER_53_1582 ();
 FILLCELL_X32 FILLER_53_1614 ();
 FILLCELL_X32 FILLER_53_1646 ();
 FILLCELL_X32 FILLER_53_1678 ();
 FILLCELL_X32 FILLER_53_1710 ();
 FILLCELL_X16 FILLER_53_1742 ();
 FILLCELL_X4 FILLER_53_1758 ();
 FILLCELL_X4 FILLER_54_1 ();
 FILLCELL_X16 FILLER_54_8 ();
 FILLCELL_X8 FILLER_54_24 ();
 FILLCELL_X1 FILLER_54_32 ();
 FILLCELL_X4 FILLER_54_37 ();
 FILLCELL_X4 FILLER_54_45 ();
 FILLCELL_X8 FILLER_54_52 ();
 FILLCELL_X1 FILLER_54_60 ();
 FILLCELL_X4 FILLER_54_65 ();
 FILLCELL_X16 FILLER_54_71 ();
 FILLCELL_X1 FILLER_54_87 ();
 FILLCELL_X4 FILLER_54_92 ();
 FILLCELL_X2 FILLER_54_96 ();
 FILLCELL_X4 FILLER_54_101 ();
 FILLCELL_X4 FILLER_54_114 ();
 FILLCELL_X4 FILLER_54_128 ();
 FILLCELL_X1 FILLER_54_132 ();
 FILLCELL_X4 FILLER_54_136 ();
 FILLCELL_X8 FILLER_54_149 ();
 FILLCELL_X4 FILLER_54_157 ();
 FILLCELL_X2 FILLER_54_161 ();
 FILLCELL_X8 FILLER_54_167 ();
 FILLCELL_X4 FILLER_54_175 ();
 FILLCELL_X2 FILLER_54_179 ();
 FILLCELL_X1 FILLER_54_181 ();
 FILLCELL_X8 FILLER_54_186 ();
 FILLCELL_X1 FILLER_54_194 ();
 FILLCELL_X4 FILLER_54_198 ();
 FILLCELL_X8 FILLER_54_212 ();
 FILLCELL_X1 FILLER_54_220 ();
 FILLCELL_X8 FILLER_54_225 ();
 FILLCELL_X4 FILLER_54_236 ();
 FILLCELL_X8 FILLER_54_250 ();
 FILLCELL_X4 FILLER_54_267 ();
 FILLCELL_X4 FILLER_54_281 ();
 FILLCELL_X4 FILLER_54_292 ();
 FILLCELL_X1 FILLER_54_296 ();
 FILLCELL_X4 FILLER_54_299 ();
 FILLCELL_X4 FILLER_54_305 ();
 FILLCELL_X4 FILLER_54_319 ();
 FILLCELL_X2 FILLER_54_323 ();
 FILLCELL_X4 FILLER_54_328 ();
 FILLCELL_X2 FILLER_54_332 ();
 FILLCELL_X1 FILLER_54_334 ();
 FILLCELL_X4 FILLER_54_339 ();
 FILLCELL_X4 FILLER_54_345 ();
 FILLCELL_X2 FILLER_54_349 ();
 FILLCELL_X4 FILLER_54_354 ();
 FILLCELL_X8 FILLER_54_367 ();
 FILLCELL_X4 FILLER_54_375 ();
 FILLCELL_X1 FILLER_54_379 ();
 FILLCELL_X32 FILLER_54_1518 ();
 FILLCELL_X32 FILLER_54_1550 ();
 FILLCELL_X32 FILLER_54_1582 ();
 FILLCELL_X32 FILLER_54_1614 ();
 FILLCELL_X32 FILLER_54_1646 ();
 FILLCELL_X32 FILLER_54_1678 ();
 FILLCELL_X32 FILLER_54_1710 ();
 FILLCELL_X16 FILLER_54_1742 ();
 FILLCELL_X4 FILLER_54_1758 ();
 FILLCELL_X16 FILLER_55_1 ();
 FILLCELL_X8 FILLER_55_17 ();
 FILLCELL_X4 FILLER_55_25 ();
 FILLCELL_X1 FILLER_55_29 ();
 FILLCELL_X4 FILLER_55_34 ();
 FILLCELL_X4 FILLER_55_47 ();
 FILLCELL_X1 FILLER_55_51 ();
 FILLCELL_X4 FILLER_55_55 ();
 FILLCELL_X16 FILLER_55_69 ();
 FILLCELL_X1 FILLER_55_85 ();
 FILLCELL_X8 FILLER_55_96 ();
 FILLCELL_X1 FILLER_55_104 ();
 FILLCELL_X4 FILLER_55_114 ();
 FILLCELL_X2 FILLER_55_118 ();
 FILLCELL_X1 FILLER_55_120 ();
 FILLCELL_X4 FILLER_55_124 ();
 FILLCELL_X2 FILLER_55_128 ();
 FILLCELL_X16 FILLER_55_133 ();
 FILLCELL_X4 FILLER_55_149 ();
 FILLCELL_X2 FILLER_55_153 ();
 FILLCELL_X4 FILLER_55_174 ();
 FILLCELL_X4 FILLER_55_188 ();
 FILLCELL_X1 FILLER_55_192 ();
 FILLCELL_X4 FILLER_55_202 ();
 FILLCELL_X8 FILLER_55_209 ();
 FILLCELL_X4 FILLER_55_226 ();
 FILLCELL_X4 FILLER_55_234 ();
 FILLCELL_X2 FILLER_55_238 ();
 FILLCELL_X1 FILLER_55_240 ();
 FILLCELL_X4 FILLER_55_251 ();
 FILLCELL_X16 FILLER_55_258 ();
 FILLCELL_X4 FILLER_55_274 ();
 FILLCELL_X8 FILLER_55_288 ();
 FILLCELL_X8 FILLER_55_306 ();
 FILLCELL_X1 FILLER_55_314 ();
 FILLCELL_X4 FILLER_55_319 ();
 FILLCELL_X4 FILLER_55_333 ();
 FILLCELL_X8 FILLER_55_342 ();
 FILLCELL_X4 FILLER_55_350 ();
 FILLCELL_X2 FILLER_55_354 ();
 FILLCELL_X4 FILLER_55_359 ();
 FILLCELL_X8 FILLER_55_366 ();
 FILLCELL_X4 FILLER_55_374 ();
 FILLCELL_X2 FILLER_55_378 ();
 FILLCELL_X32 FILLER_55_1518 ();
 FILLCELL_X32 FILLER_55_1550 ();
 FILLCELL_X32 FILLER_55_1582 ();
 FILLCELL_X32 FILLER_55_1614 ();
 FILLCELL_X32 FILLER_55_1646 ();
 FILLCELL_X32 FILLER_55_1678 ();
 FILLCELL_X32 FILLER_55_1710 ();
 FILLCELL_X16 FILLER_55_1742 ();
 FILLCELL_X4 FILLER_55_1758 ();
 FILLCELL_X32 FILLER_56_1 ();
 FILLCELL_X8 FILLER_56_33 ();
 FILLCELL_X8 FILLER_56_44 ();
 FILLCELL_X4 FILLER_56_56 ();
 FILLCELL_X4 FILLER_56_70 ();
 FILLCELL_X2 FILLER_56_74 ();
 FILLCELL_X4 FILLER_56_86 ();
 FILLCELL_X8 FILLER_56_97 ();
 FILLCELL_X4 FILLER_56_105 ();
 FILLCELL_X1 FILLER_56_109 ();
 FILLCELL_X4 FILLER_56_113 ();
 FILLCELL_X4 FILLER_56_120 ();
 FILLCELL_X4 FILLER_56_127 ();
 FILLCELL_X1 FILLER_56_131 ();
 FILLCELL_X8 FILLER_56_134 ();
 FILLCELL_X2 FILLER_56_142 ();
 FILLCELL_X4 FILLER_56_147 ();
 FILLCELL_X8 FILLER_56_161 ();
 FILLCELL_X4 FILLER_56_169 ();
 FILLCELL_X2 FILLER_56_173 ();
 FILLCELL_X4 FILLER_56_179 ();
 FILLCELL_X4 FILLER_56_193 ();
 FILLCELL_X4 FILLER_56_204 ();
 FILLCELL_X8 FILLER_56_211 ();
 FILLCELL_X1 FILLER_56_219 ();
 FILLCELL_X4 FILLER_56_224 ();
 FILLCELL_X2 FILLER_56_228 ();
 FILLCELL_X16 FILLER_56_233 ();
 FILLCELL_X2 FILLER_56_249 ();
 FILLCELL_X1 FILLER_56_251 ();
 FILLCELL_X4 FILLER_56_255 ();
 FILLCELL_X16 FILLER_56_262 ();
 FILLCELL_X4 FILLER_56_278 ();
 FILLCELL_X1 FILLER_56_282 ();
 FILLCELL_X8 FILLER_56_292 ();
 FILLCELL_X1 FILLER_56_300 ();
 FILLCELL_X4 FILLER_56_311 ();
 FILLCELL_X8 FILLER_56_318 ();
 FILLCELL_X1 FILLER_56_326 ();
 FILLCELL_X4 FILLER_56_330 ();
 FILLCELL_X4 FILLER_56_336 ();
 FILLCELL_X4 FILLER_56_350 ();
 FILLCELL_X4 FILLER_56_363 ();
 FILLCELL_X4 FILLER_56_373 ();
 FILLCELL_X2 FILLER_56_377 ();
 FILLCELL_X1 FILLER_56_379 ();
 FILLCELL_X32 FILLER_56_1518 ();
 FILLCELL_X32 FILLER_56_1550 ();
 FILLCELL_X32 FILLER_56_1582 ();
 FILLCELL_X32 FILLER_56_1614 ();
 FILLCELL_X32 FILLER_56_1646 ();
 FILLCELL_X32 FILLER_56_1678 ();
 FILLCELL_X32 FILLER_56_1710 ();
 FILLCELL_X16 FILLER_56_1742 ();
 FILLCELL_X4 FILLER_56_1758 ();
 FILLCELL_X8 FILLER_57_1 ();
 FILLCELL_X4 FILLER_57_9 ();
 FILLCELL_X2 FILLER_57_13 ();
 FILLCELL_X4 FILLER_57_19 ();
 FILLCELL_X4 FILLER_57_33 ();
 FILLCELL_X8 FILLER_57_40 ();
 FILLCELL_X1 FILLER_57_48 ();
 FILLCELL_X4 FILLER_57_59 ();
 FILLCELL_X8 FILLER_57_66 ();
 FILLCELL_X4 FILLER_57_74 ();
 FILLCELL_X4 FILLER_57_81 ();
 FILLCELL_X4 FILLER_57_87 ();
 FILLCELL_X1 FILLER_57_91 ();
 FILLCELL_X8 FILLER_57_96 ();
 FILLCELL_X2 FILLER_57_104 ();
 FILLCELL_X4 FILLER_57_115 ();
 FILLCELL_X2 FILLER_57_119 ();
 FILLCELL_X1 FILLER_57_121 ();
 FILLCELL_X4 FILLER_57_125 ();
 FILLCELL_X1 FILLER_57_129 ();
 FILLCELL_X4 FILLER_57_140 ();
 FILLCELL_X4 FILLER_57_148 ();
 FILLCELL_X2 FILLER_57_152 ();
 FILLCELL_X4 FILLER_57_163 ();
 FILLCELL_X1 FILLER_57_167 ();
 FILLCELL_X8 FILLER_57_171 ();
 FILLCELL_X4 FILLER_57_179 ();
 FILLCELL_X2 FILLER_57_183 ();
 FILLCELL_X4 FILLER_57_188 ();
 FILLCELL_X8 FILLER_57_201 ();
 FILLCELL_X1 FILLER_57_209 ();
 FILLCELL_X4 FILLER_57_219 ();
 FILLCELL_X8 FILLER_57_226 ();
 FILLCELL_X2 FILLER_57_234 ();
 FILLCELL_X4 FILLER_57_245 ();
 FILLCELL_X4 FILLER_57_258 ();
 FILLCELL_X8 FILLER_57_265 ();
 FILLCELL_X1 FILLER_57_273 ();
 FILLCELL_X4 FILLER_57_278 ();
 FILLCELL_X4 FILLER_57_285 ();
 FILLCELL_X4 FILLER_57_292 ();
 FILLCELL_X16 FILLER_57_299 ();
 FILLCELL_X4 FILLER_57_315 ();
 FILLCELL_X2 FILLER_57_319 ();
 FILLCELL_X8 FILLER_57_324 ();
 FILLCELL_X4 FILLER_57_342 ();
 FILLCELL_X4 FILLER_57_353 ();
 FILLCELL_X4 FILLER_57_360 ();
 FILLCELL_X2 FILLER_57_364 ();
 FILLCELL_X8 FILLER_57_372 ();
 FILLCELL_X32 FILLER_57_1518 ();
 FILLCELL_X32 FILLER_57_1550 ();
 FILLCELL_X32 FILLER_57_1582 ();
 FILLCELL_X32 FILLER_57_1614 ();
 FILLCELL_X32 FILLER_57_1646 ();
 FILLCELL_X32 FILLER_57_1678 ();
 FILLCELL_X32 FILLER_57_1710 ();
 FILLCELL_X16 FILLER_57_1742 ();
 FILLCELL_X4 FILLER_57_1758 ();
 FILLCELL_X32 FILLER_58_1 ();
 FILLCELL_X8 FILLER_58_33 ();
 FILLCELL_X4 FILLER_58_41 ();
 FILLCELL_X2 FILLER_58_45 ();
 FILLCELL_X1 FILLER_58_47 ();
 FILLCELL_X4 FILLER_58_55 ();
 FILLCELL_X1 FILLER_58_59 ();
 FILLCELL_X4 FILLER_58_63 ();
 FILLCELL_X4 FILLER_58_76 ();
 FILLCELL_X1 FILLER_58_80 ();
 FILLCELL_X4 FILLER_58_84 ();
 FILLCELL_X4 FILLER_58_97 ();
 FILLCELL_X16 FILLER_58_105 ();
 FILLCELL_X8 FILLER_58_121 ();
 FILLCELL_X4 FILLER_58_129 ();
 FILLCELL_X1 FILLER_58_133 ();
 FILLCELL_X4 FILLER_58_144 ();
 FILLCELL_X8 FILLER_58_151 ();
 FILLCELL_X4 FILLER_58_159 ();
 FILLCELL_X2 FILLER_58_163 ();
 FILLCELL_X4 FILLER_58_168 ();
 FILLCELL_X16 FILLER_58_175 ();
 FILLCELL_X1 FILLER_58_191 ();
 FILLCELL_X4 FILLER_58_202 ();
 FILLCELL_X4 FILLER_58_209 ();
 FILLCELL_X2 FILLER_58_213 ();
 FILLCELL_X4 FILLER_58_218 ();
 FILLCELL_X32 FILLER_58_225 ();
 FILLCELL_X1 FILLER_58_257 ();
 FILLCELL_X4 FILLER_58_262 ();
 FILLCELL_X4 FILLER_58_270 ();
 FILLCELL_X4 FILLER_58_283 ();
 FILLCELL_X8 FILLER_58_290 ();
 FILLCELL_X1 FILLER_58_298 ();
 FILLCELL_X8 FILLER_58_303 ();
 FILLCELL_X2 FILLER_58_311 ();
 FILLCELL_X4 FILLER_58_315 ();
 FILLCELL_X16 FILLER_58_329 ();
 FILLCELL_X8 FILLER_58_345 ();
 FILLCELL_X4 FILLER_58_353 ();
 FILLCELL_X2 FILLER_58_357 ();
 FILLCELL_X1 FILLER_58_359 ();
 FILLCELL_X4 FILLER_58_364 ();
 FILLCELL_X4 FILLER_58_375 ();
 FILLCELL_X1 FILLER_58_379 ();
 FILLCELL_X32 FILLER_58_1518 ();
 FILLCELL_X32 FILLER_58_1550 ();
 FILLCELL_X32 FILLER_58_1582 ();
 FILLCELL_X32 FILLER_58_1614 ();
 FILLCELL_X32 FILLER_58_1646 ();
 FILLCELL_X32 FILLER_58_1678 ();
 FILLCELL_X32 FILLER_58_1710 ();
 FILLCELL_X16 FILLER_58_1742 ();
 FILLCELL_X4 FILLER_58_1758 ();
 FILLCELL_X16 FILLER_59_1 ();
 FILLCELL_X2 FILLER_59_17 ();
 FILLCELL_X1 FILLER_59_19 ();
 FILLCELL_X4 FILLER_59_22 ();
 FILLCELL_X4 FILLER_59_33 ();
 FILLCELL_X2 FILLER_59_37 ();
 FILLCELL_X1 FILLER_59_39 ();
 FILLCELL_X4 FILLER_59_50 ();
 FILLCELL_X4 FILLER_59_63 ();
 FILLCELL_X4 FILLER_59_70 ();
 FILLCELL_X8 FILLER_59_76 ();
 FILLCELL_X4 FILLER_59_84 ();
 FILLCELL_X1 FILLER_59_88 ();
 FILLCELL_X4 FILLER_59_93 ();
 FILLCELL_X8 FILLER_59_100 ();
 FILLCELL_X1 FILLER_59_108 ();
 FILLCELL_X16 FILLER_59_113 ();
 FILLCELL_X1 FILLER_59_129 ();
 FILLCELL_X4 FILLER_59_132 ();
 FILLCELL_X8 FILLER_59_143 ();
 FILLCELL_X4 FILLER_59_151 ();
 FILLCELL_X2 FILLER_59_155 ();
 FILLCELL_X1 FILLER_59_157 ();
 FILLCELL_X4 FILLER_59_164 ();
 FILLCELL_X4 FILLER_59_181 ();
 FILLCELL_X8 FILLER_59_188 ();
 FILLCELL_X2 FILLER_59_196 ();
 FILLCELL_X1 FILLER_59_198 ();
 FILLCELL_X4 FILLER_59_201 ();
 FILLCELL_X4 FILLER_59_209 ();
 FILLCELL_X4 FILLER_59_223 ();
 FILLCELL_X4 FILLER_59_236 ();
 FILLCELL_X1 FILLER_59_240 ();
 FILLCELL_X4 FILLER_59_251 ();
 FILLCELL_X8 FILLER_59_262 ();
 FILLCELL_X4 FILLER_59_279 ();
 FILLCELL_X8 FILLER_59_286 ();
 FILLCELL_X4 FILLER_59_297 ();
 FILLCELL_X8 FILLER_59_311 ();
 FILLCELL_X4 FILLER_59_328 ();
 FILLCELL_X1 FILLER_59_332 ();
 FILLCELL_X4 FILLER_59_336 ();
 FILLCELL_X8 FILLER_59_349 ();
 FILLCELL_X4 FILLER_59_357 ();
 FILLCELL_X2 FILLER_59_361 ();
 FILLCELL_X8 FILLER_59_369 ();
 FILLCELL_X2 FILLER_59_377 ();
 FILLCELL_X1 FILLER_59_379 ();
 FILLCELL_X32 FILLER_59_1518 ();
 FILLCELL_X32 FILLER_59_1550 ();
 FILLCELL_X32 FILLER_59_1582 ();
 FILLCELL_X32 FILLER_59_1614 ();
 FILLCELL_X32 FILLER_59_1646 ();
 FILLCELL_X32 FILLER_59_1678 ();
 FILLCELL_X32 FILLER_59_1710 ();
 FILLCELL_X8 FILLER_59_1742 ();
 FILLCELL_X4 FILLER_59_1750 ();
 FILLCELL_X1 FILLER_59_1754 ();
 FILLCELL_X4 FILLER_59_1758 ();
 FILLCELL_X8 FILLER_60_1 ();
 FILLCELL_X1 FILLER_60_9 ();
 FILLCELL_X4 FILLER_60_14 ();
 FILLCELL_X2 FILLER_60_18 ();
 FILLCELL_X1 FILLER_60_20 ();
 FILLCELL_X4 FILLER_60_31 ();
 FILLCELL_X8 FILLER_60_38 ();
 FILLCELL_X4 FILLER_60_48 ();
 FILLCELL_X4 FILLER_60_55 ();
 FILLCELL_X4 FILLER_60_68 ();
 FILLCELL_X8 FILLER_60_75 ();
 FILLCELL_X1 FILLER_60_83 ();
 FILLCELL_X8 FILLER_60_93 ();
 FILLCELL_X1 FILLER_60_101 ();
 FILLCELL_X4 FILLER_60_106 ();
 FILLCELL_X4 FILLER_60_123 ();
 FILLCELL_X8 FILLER_60_133 ();
 FILLCELL_X4 FILLER_60_141 ();
 FILLCELL_X1 FILLER_60_145 ();
 FILLCELL_X4 FILLER_60_148 ();
 FILLCELL_X2 FILLER_60_152 ();
 FILLCELL_X4 FILLER_60_161 ();
 FILLCELL_X8 FILLER_60_171 ();
 FILLCELL_X2 FILLER_60_179 ();
 FILLCELL_X16 FILLER_60_200 ();
 FILLCELL_X2 FILLER_60_216 ();
 FILLCELL_X8 FILLER_60_225 ();
 FILLCELL_X1 FILLER_60_233 ();
 FILLCELL_X4 FILLER_60_236 ();
 FILLCELL_X4 FILLER_60_250 ();
 FILLCELL_X4 FILLER_60_257 ();
 FILLCELL_X1 FILLER_60_261 ();
 FILLCELL_X32 FILLER_60_266 ();
 FILLCELL_X4 FILLER_60_305 ();
 FILLCELL_X2 FILLER_60_309 ();
 FILLCELL_X1 FILLER_60_311 ();
 FILLCELL_X8 FILLER_60_319 ();
 FILLCELL_X1 FILLER_60_327 ();
 FILLCELL_X4 FILLER_60_331 ();
 FILLCELL_X4 FILLER_60_344 ();
 FILLCELL_X2 FILLER_60_348 ();
 FILLCELL_X4 FILLER_60_360 ();
 FILLCELL_X1 FILLER_60_364 ();
 FILLCELL_X4 FILLER_60_367 ();
 FILLCELL_X4 FILLER_60_375 ();
 FILLCELL_X1 FILLER_60_379 ();
 FILLCELL_X32 FILLER_60_1518 ();
 FILLCELL_X32 FILLER_60_1550 ();
 FILLCELL_X32 FILLER_60_1582 ();
 FILLCELL_X32 FILLER_60_1614 ();
 FILLCELL_X32 FILLER_60_1646 ();
 FILLCELL_X32 FILLER_60_1678 ();
 FILLCELL_X32 FILLER_60_1710 ();
 FILLCELL_X16 FILLER_60_1742 ();
 FILLCELL_X4 FILLER_60_1758 ();
 FILLCELL_X4 FILLER_61_1 ();
 FILLCELL_X8 FILLER_61_22 ();
 FILLCELL_X4 FILLER_61_39 ();
 FILLCELL_X8 FILLER_61_46 ();
 FILLCELL_X1 FILLER_61_54 ();
 FILLCELL_X4 FILLER_61_58 ();
 FILLCELL_X4 FILLER_61_72 ();
 FILLCELL_X2 FILLER_61_76 ();
 FILLCELL_X4 FILLER_61_88 ();
 FILLCELL_X1 FILLER_61_92 ();
 FILLCELL_X4 FILLER_61_99 ();
 FILLCELL_X8 FILLER_61_109 ();
 FILLCELL_X4 FILLER_61_120 ();
 FILLCELL_X4 FILLER_61_133 ();
 FILLCELL_X4 FILLER_61_147 ();
 FILLCELL_X2 FILLER_61_151 ();
 FILLCELL_X1 FILLER_61_153 ();
 FILLCELL_X8 FILLER_61_164 ();
 FILLCELL_X2 FILLER_61_172 ();
 FILLCELL_X8 FILLER_61_178 ();
 FILLCELL_X1 FILLER_61_186 ();
 FILLCELL_X4 FILLER_61_197 ();
 FILLCELL_X8 FILLER_61_204 ();
 FILLCELL_X1 FILLER_61_212 ();
 FILLCELL_X4 FILLER_61_223 ();
 FILLCELL_X16 FILLER_61_229 ();
 FILLCELL_X4 FILLER_61_245 ();
 FILLCELL_X4 FILLER_61_256 ();
 FILLCELL_X8 FILLER_61_270 ();
 FILLCELL_X4 FILLER_61_278 ();
 FILLCELL_X1 FILLER_61_282 ();
 FILLCELL_X4 FILLER_61_285 ();
 FILLCELL_X4 FILLER_61_293 ();
 FILLCELL_X4 FILLER_61_307 ();
 FILLCELL_X2 FILLER_61_311 ();
 FILLCELL_X4 FILLER_61_322 ();
 FILLCELL_X1 FILLER_61_326 ();
 FILLCELL_X4 FILLER_61_337 ();
 FILLCELL_X2 FILLER_61_341 ();
 FILLCELL_X4 FILLER_61_346 ();
 FILLCELL_X2 FILLER_61_350 ();
 FILLCELL_X8 FILLER_61_354 ();
 FILLCELL_X1 FILLER_61_362 ();
 FILLCELL_X8 FILLER_61_370 ();
 FILLCELL_X2 FILLER_61_378 ();
 FILLCELL_X32 FILLER_61_1518 ();
 FILLCELL_X32 FILLER_61_1550 ();
 FILLCELL_X32 FILLER_61_1582 ();
 FILLCELL_X32 FILLER_61_1614 ();
 FILLCELL_X32 FILLER_61_1646 ();
 FILLCELL_X32 FILLER_61_1678 ();
 FILLCELL_X32 FILLER_61_1710 ();
 FILLCELL_X16 FILLER_61_1742 ();
 FILLCELL_X4 FILLER_61_1758 ();
 FILLCELL_X4 FILLER_62_1 ();
 FILLCELL_X4 FILLER_62_9 ();
 FILLCELL_X2 FILLER_62_13 ();
 FILLCELL_X8 FILLER_62_18 ();
 FILLCELL_X2 FILLER_62_26 ();
 FILLCELL_X4 FILLER_62_37 ();
 FILLCELL_X2 FILLER_62_41 ();
 FILLCELL_X4 FILLER_62_47 ();
 FILLCELL_X8 FILLER_62_54 ();
 FILLCELL_X4 FILLER_62_62 ();
 FILLCELL_X2 FILLER_62_66 ();
 FILLCELL_X1 FILLER_62_68 ();
 FILLCELL_X4 FILLER_62_76 ();
 FILLCELL_X4 FILLER_62_83 ();
 FILLCELL_X4 FILLER_62_89 ();
 FILLCELL_X2 FILLER_62_93 ();
 FILLCELL_X8 FILLER_62_105 ();
 FILLCELL_X4 FILLER_62_113 ();
 FILLCELL_X2 FILLER_62_117 ();
 FILLCELL_X8 FILLER_62_122 ();
 FILLCELL_X4 FILLER_62_133 ();
 FILLCELL_X2 FILLER_62_137 ();
 FILLCELL_X4 FILLER_62_142 ();
 FILLCELL_X8 FILLER_62_155 ();
 FILLCELL_X2 FILLER_62_163 ();
 FILLCELL_X1 FILLER_62_165 ();
 FILLCELL_X8 FILLER_62_169 ();
 FILLCELL_X1 FILLER_62_177 ();
 FILLCELL_X8 FILLER_62_185 ();
 FILLCELL_X2 FILLER_62_193 ();
 FILLCELL_X4 FILLER_62_198 ();
 FILLCELL_X4 FILLER_62_206 ();
 FILLCELL_X8 FILLER_62_214 ();
 FILLCELL_X4 FILLER_62_222 ();
 FILLCELL_X2 FILLER_62_226 ();
 FILLCELL_X1 FILLER_62_228 ();
 FILLCELL_X4 FILLER_62_232 ();
 FILLCELL_X8 FILLER_62_239 ();
 FILLCELL_X1 FILLER_62_247 ();
 FILLCELL_X4 FILLER_62_258 ();
 FILLCELL_X4 FILLER_62_265 ();
 FILLCELL_X4 FILLER_62_273 ();
 FILLCELL_X4 FILLER_62_286 ();
 FILLCELL_X4 FILLER_62_300 ();
 FILLCELL_X4 FILLER_62_307 ();
 FILLCELL_X4 FILLER_62_314 ();
 FILLCELL_X4 FILLER_62_321 ();
 FILLCELL_X16 FILLER_62_332 ();
 FILLCELL_X2 FILLER_62_348 ();
 FILLCELL_X1 FILLER_62_350 ();
 FILLCELL_X4 FILLER_62_355 ();
 FILLCELL_X2 FILLER_62_359 ();
 FILLCELL_X8 FILLER_62_371 ();
 FILLCELL_X1 FILLER_62_379 ();
 FILLCELL_X32 FILLER_62_1518 ();
 FILLCELL_X32 FILLER_62_1550 ();
 FILLCELL_X32 FILLER_62_1582 ();
 FILLCELL_X32 FILLER_62_1614 ();
 FILLCELL_X32 FILLER_62_1646 ();
 FILLCELL_X32 FILLER_62_1678 ();
 FILLCELL_X32 FILLER_62_1710 ();
 FILLCELL_X16 FILLER_62_1742 ();
 FILLCELL_X4 FILLER_62_1758 ();
 FILLCELL_X4 FILLER_63_1 ();
 FILLCELL_X4 FILLER_63_12 ();
 FILLCELL_X4 FILLER_63_20 ();
 FILLCELL_X4 FILLER_63_27 ();
 FILLCELL_X2 FILLER_63_31 ();
 FILLCELL_X1 FILLER_63_33 ();
 FILLCELL_X4 FILLER_63_37 ();
 FILLCELL_X16 FILLER_63_51 ();
 FILLCELL_X4 FILLER_63_67 ();
 FILLCELL_X1 FILLER_63_71 ();
 FILLCELL_X8 FILLER_63_82 ();
 FILLCELL_X4 FILLER_63_94 ();
 FILLCELL_X4 FILLER_63_101 ();
 FILLCELL_X2 FILLER_63_105 ();
 FILLCELL_X8 FILLER_63_116 ();
 FILLCELL_X2 FILLER_63_124 ();
 FILLCELL_X8 FILLER_63_130 ();
 FILLCELL_X1 FILLER_63_138 ();
 FILLCELL_X4 FILLER_63_148 ();
 FILLCELL_X4 FILLER_63_156 ();
 FILLCELL_X8 FILLER_63_163 ();
 FILLCELL_X2 FILLER_63_171 ();
 FILLCELL_X4 FILLER_63_183 ();
 FILLCELL_X4 FILLER_63_189 ();
 FILLCELL_X2 FILLER_63_193 ();
 FILLCELL_X1 FILLER_63_195 ();
 FILLCELL_X4 FILLER_63_199 ();
 FILLCELL_X8 FILLER_63_212 ();
 FILLCELL_X2 FILLER_63_220 ();
 FILLCELL_X4 FILLER_63_226 ();
 FILLCELL_X4 FILLER_63_239 ();
 FILLCELL_X4 FILLER_63_247 ();
 FILLCELL_X4 FILLER_63_253 ();
 FILLCELL_X8 FILLER_63_260 ();
 FILLCELL_X2 FILLER_63_268 ();
 FILLCELL_X4 FILLER_63_274 ();
 FILLCELL_X32 FILLER_63_281 ();
 FILLCELL_X8 FILLER_63_313 ();
 FILLCELL_X1 FILLER_63_321 ();
 FILLCELL_X8 FILLER_63_324 ();
 FILLCELL_X4 FILLER_63_335 ();
 FILLCELL_X4 FILLER_63_342 ();
 FILLCELL_X4 FILLER_63_356 ();
 FILLCELL_X2 FILLER_63_360 ();
 FILLCELL_X8 FILLER_63_365 ();
 FILLCELL_X4 FILLER_63_373 ();
 FILLCELL_X2 FILLER_63_377 ();
 FILLCELL_X1 FILLER_63_379 ();
 FILLCELL_X32 FILLER_63_1518 ();
 FILLCELL_X32 FILLER_63_1550 ();
 FILLCELL_X32 FILLER_63_1582 ();
 FILLCELL_X32 FILLER_63_1614 ();
 FILLCELL_X32 FILLER_63_1646 ();
 FILLCELL_X32 FILLER_63_1678 ();
 FILLCELL_X32 FILLER_63_1710 ();
 FILLCELL_X16 FILLER_63_1742 ();
 FILLCELL_X4 FILLER_63_1758 ();
 FILLCELL_X8 FILLER_64_1 ();
 FILLCELL_X2 FILLER_64_9 ();
 FILLCELL_X4 FILLER_64_20 ();
 FILLCELL_X8 FILLER_64_28 ();
 FILLCELL_X4 FILLER_64_36 ();
 FILLCELL_X2 FILLER_64_40 ();
 FILLCELL_X1 FILLER_64_42 ();
 FILLCELL_X16 FILLER_64_45 ();
 FILLCELL_X4 FILLER_64_61 ();
 FILLCELL_X2 FILLER_64_65 ();
 FILLCELL_X1 FILLER_64_67 ();
 FILLCELL_X8 FILLER_64_71 ();
 FILLCELL_X4 FILLER_64_79 ();
 FILLCELL_X2 FILLER_64_83 ();
 FILLCELL_X4 FILLER_64_89 ();
 FILLCELL_X4 FILLER_64_103 ();
 FILLCELL_X4 FILLER_64_110 ();
 FILLCELL_X1 FILLER_64_114 ();
 FILLCELL_X4 FILLER_64_122 ();
 FILLCELL_X8 FILLER_64_136 ();
 FILLCELL_X4 FILLER_64_144 ();
 FILLCELL_X2 FILLER_64_148 ();
 FILLCELL_X4 FILLER_64_159 ();
 FILLCELL_X8 FILLER_64_167 ();
 FILLCELL_X2 FILLER_64_175 ();
 FILLCELL_X1 FILLER_64_177 ();
 FILLCELL_X4 FILLER_64_181 ();
 FILLCELL_X4 FILLER_64_187 ();
 FILLCELL_X2 FILLER_64_191 ();
 FILLCELL_X4 FILLER_64_197 ();
 FILLCELL_X16 FILLER_64_210 ();
 FILLCELL_X4 FILLER_64_235 ();
 FILLCELL_X8 FILLER_64_243 ();
 FILLCELL_X8 FILLER_64_255 ();
 FILLCELL_X2 FILLER_64_263 ();
 FILLCELL_X4 FILLER_64_269 ();
 FILLCELL_X4 FILLER_64_282 ();
 FILLCELL_X8 FILLER_64_289 ();
 FILLCELL_X2 FILLER_64_297 ();
 FILLCELL_X4 FILLER_64_303 ();
 FILLCELL_X4 FILLER_64_316 ();
 FILLCELL_X2 FILLER_64_320 ();
 FILLCELL_X1 FILLER_64_322 ();
 FILLCELL_X4 FILLER_64_327 ();
 FILLCELL_X8 FILLER_64_341 ();
 FILLCELL_X1 FILLER_64_349 ();
 FILLCELL_X16 FILLER_64_359 ();
 FILLCELL_X4 FILLER_64_375 ();
 FILLCELL_X1 FILLER_64_379 ();
 FILLCELL_X32 FILLER_64_1518 ();
 FILLCELL_X32 FILLER_64_1550 ();
 FILLCELL_X32 FILLER_64_1582 ();
 FILLCELL_X32 FILLER_64_1614 ();
 FILLCELL_X32 FILLER_64_1646 ();
 FILLCELL_X32 FILLER_64_1678 ();
 FILLCELL_X32 FILLER_64_1710 ();
 FILLCELL_X16 FILLER_64_1742 ();
 FILLCELL_X4 FILLER_64_1758 ();
 FILLCELL_X4 FILLER_65_1 ();
 FILLCELL_X2 FILLER_65_5 ();
 FILLCELL_X1 FILLER_65_7 ();
 FILLCELL_X4 FILLER_65_17 ();
 FILLCELL_X4 FILLER_65_24 ();
 FILLCELL_X2 FILLER_65_28 ();
 FILLCELL_X4 FILLER_65_33 ();
 FILLCELL_X4 FILLER_65_41 ();
 FILLCELL_X4 FILLER_65_52 ();
 FILLCELL_X2 FILLER_65_56 ();
 FILLCELL_X1 FILLER_65_58 ();
 FILLCELL_X4 FILLER_65_61 ();
 FILLCELL_X4 FILLER_65_75 ();
 FILLCELL_X4 FILLER_65_86 ();
 FILLCELL_X16 FILLER_65_92 ();
 FILLCELL_X4 FILLER_65_108 ();
 FILLCELL_X2 FILLER_65_112 ();
 FILLCELL_X1 FILLER_65_114 ();
 FILLCELL_X4 FILLER_65_117 ();
 FILLCELL_X4 FILLER_65_128 ();
 FILLCELL_X8 FILLER_65_135 ();
 FILLCELL_X1 FILLER_65_143 ();
 FILLCELL_X4 FILLER_65_147 ();
 FILLCELL_X8 FILLER_65_155 ();
 FILLCELL_X2 FILLER_65_163 ();
 FILLCELL_X4 FILLER_65_174 ();
 FILLCELL_X8 FILLER_65_188 ();
 FILLCELL_X1 FILLER_65_196 ();
 FILLCELL_X4 FILLER_65_204 ();
 FILLCELL_X16 FILLER_65_211 ();
 FILLCELL_X2 FILLER_65_227 ();
 FILLCELL_X8 FILLER_65_232 ();
 FILLCELL_X2 FILLER_65_240 ();
 FILLCELL_X4 FILLER_65_246 ();
 FILLCELL_X4 FILLER_65_259 ();
 FILLCELL_X8 FILLER_65_266 ();
 FILLCELL_X1 FILLER_65_274 ();
 FILLCELL_X8 FILLER_65_278 ();
 FILLCELL_X2 FILLER_65_286 ();
 FILLCELL_X4 FILLER_65_292 ();
 FILLCELL_X4 FILLER_65_305 ();
 FILLCELL_X2 FILLER_65_309 ();
 FILLCELL_X16 FILLER_65_321 ();
 FILLCELL_X2 FILLER_65_337 ();
 FILLCELL_X4 FILLER_65_342 ();
 FILLCELL_X4 FILLER_65_349 ();
 FILLCELL_X4 FILLER_65_356 ();
 FILLCELL_X8 FILLER_65_369 ();
 FILLCELL_X2 FILLER_65_377 ();
 FILLCELL_X1 FILLER_65_379 ();
 FILLCELL_X32 FILLER_65_1518 ();
 FILLCELL_X32 FILLER_65_1550 ();
 FILLCELL_X32 FILLER_65_1582 ();
 FILLCELL_X32 FILLER_65_1614 ();
 FILLCELL_X32 FILLER_65_1646 ();
 FILLCELL_X32 FILLER_65_1678 ();
 FILLCELL_X32 FILLER_65_1710 ();
 FILLCELL_X16 FILLER_65_1742 ();
 FILLCELL_X4 FILLER_65_1758 ();
 FILLCELL_X8 FILLER_66_1 ();
 FILLCELL_X8 FILLER_66_12 ();
 FILLCELL_X4 FILLER_66_20 ();
 FILLCELL_X2 FILLER_66_24 ();
 FILLCELL_X4 FILLER_66_29 ();
 FILLCELL_X4 FILLER_66_42 ();
 FILLCELL_X4 FILLER_66_56 ();
 FILLCELL_X2 FILLER_66_60 ();
 FILLCELL_X1 FILLER_66_62 ();
 FILLCELL_X4 FILLER_66_73 ();
 FILLCELL_X4 FILLER_66_80 ();
 FILLCELL_X2 FILLER_66_84 ();
 FILLCELL_X8 FILLER_66_96 ();
 FILLCELL_X4 FILLER_66_104 ();
 FILLCELL_X2 FILLER_66_108 ();
 FILLCELL_X4 FILLER_66_113 ();
 FILLCELL_X2 FILLER_66_117 ();
 FILLCELL_X1 FILLER_66_119 ();
 FILLCELL_X16 FILLER_66_130 ();
 FILLCELL_X8 FILLER_66_146 ();
 FILLCELL_X4 FILLER_66_154 ();
 FILLCELL_X1 FILLER_66_158 ();
 FILLCELL_X8 FILLER_66_162 ();
 FILLCELL_X2 FILLER_66_170 ();
 FILLCELL_X1 FILLER_66_172 ();
 FILLCELL_X4 FILLER_66_182 ();
 FILLCELL_X8 FILLER_66_189 ();
 FILLCELL_X4 FILLER_66_207 ();
 FILLCELL_X4 FILLER_66_214 ();
 FILLCELL_X2 FILLER_66_218 ();
 FILLCELL_X1 FILLER_66_220 ();
 FILLCELL_X4 FILLER_66_230 ();
 FILLCELL_X8 FILLER_66_237 ();
 FILLCELL_X4 FILLER_66_245 ();
 FILLCELL_X4 FILLER_66_253 ();
 FILLCELL_X8 FILLER_66_260 ();
 FILLCELL_X4 FILLER_66_268 ();
 FILLCELL_X1 FILLER_66_272 ();
 FILLCELL_X4 FILLER_66_277 ();
 FILLCELL_X4 FILLER_66_290 ();
 FILLCELL_X1 FILLER_66_294 ();
 FILLCELL_X4 FILLER_66_298 ();
 FILLCELL_X4 FILLER_66_305 ();
 FILLCELL_X4 FILLER_66_312 ();
 FILLCELL_X4 FILLER_66_318 ();
 FILLCELL_X1 FILLER_66_322 ();
 FILLCELL_X4 FILLER_66_325 ();
 FILLCELL_X4 FILLER_66_339 ();
 FILLCELL_X4 FILLER_66_352 ();
 FILLCELL_X4 FILLER_66_360 ();
 FILLCELL_X4 FILLER_66_373 ();
 FILLCELL_X2 FILLER_66_377 ();
 FILLCELL_X1 FILLER_66_379 ();
 FILLCELL_X32 FILLER_66_1518 ();
 FILLCELL_X32 FILLER_66_1550 ();
 FILLCELL_X32 FILLER_66_1582 ();
 FILLCELL_X32 FILLER_66_1614 ();
 FILLCELL_X32 FILLER_66_1646 ();
 FILLCELL_X32 FILLER_66_1678 ();
 FILLCELL_X32 FILLER_66_1710 ();
 FILLCELL_X16 FILLER_66_1742 ();
 FILLCELL_X4 FILLER_66_1758 ();
 FILLCELL_X4 FILLER_67_1 ();
 FILLCELL_X2 FILLER_67_5 ();
 FILLCELL_X4 FILLER_67_17 ();
 FILLCELL_X4 FILLER_67_25 ();
 FILLCELL_X4 FILLER_67_32 ();
 FILLCELL_X2 FILLER_67_36 ();
 FILLCELL_X1 FILLER_67_38 ();
 FILLCELL_X4 FILLER_67_43 ();
 FILLCELL_X8 FILLER_67_50 ();
 FILLCELL_X4 FILLER_67_58 ();
 FILLCELL_X1 FILLER_67_62 ();
 FILLCELL_X4 FILLER_67_72 ();
 FILLCELL_X4 FILLER_67_79 ();
 FILLCELL_X1 FILLER_67_83 ();
 FILLCELL_X4 FILLER_67_93 ();
 FILLCELL_X4 FILLER_67_106 ();
 FILLCELL_X4 FILLER_67_120 ();
 FILLCELL_X4 FILLER_67_126 ();
 FILLCELL_X1 FILLER_67_130 ();
 FILLCELL_X4 FILLER_67_134 ();
 FILLCELL_X8 FILLER_67_148 ();
 FILLCELL_X2 FILLER_67_156 ();
 FILLCELL_X1 FILLER_67_158 ();
 FILLCELL_X16 FILLER_67_163 ();
 FILLCELL_X8 FILLER_67_179 ();
 FILLCELL_X4 FILLER_67_187 ();
 FILLCELL_X2 FILLER_67_191 ();
 FILLCELL_X4 FILLER_67_195 ();
 FILLCELL_X4 FILLER_67_203 ();
 FILLCELL_X4 FILLER_67_210 ();
 FILLCELL_X4 FILLER_67_223 ();
 FILLCELL_X4 FILLER_67_230 ();
 FILLCELL_X2 FILLER_67_234 ();
 FILLCELL_X1 FILLER_67_236 ();
 FILLCELL_X4 FILLER_67_244 ();
 FILLCELL_X8 FILLER_67_257 ();
 FILLCELL_X1 FILLER_67_265 ();
 FILLCELL_X4 FILLER_67_270 ();
 FILLCELL_X4 FILLER_67_283 ();
 FILLCELL_X8 FILLER_67_290 ();
 FILLCELL_X4 FILLER_67_298 ();
 FILLCELL_X4 FILLER_67_305 ();
 FILLCELL_X4 FILLER_67_313 ();
 FILLCELL_X2 FILLER_67_317 ();
 FILLCELL_X1 FILLER_67_319 ();
 FILLCELL_X4 FILLER_67_330 ();
 FILLCELL_X4 FILLER_67_341 ();
 FILLCELL_X8 FILLER_67_348 ();
 FILLCELL_X4 FILLER_67_359 ();
 FILLCELL_X4 FILLER_67_367 ();
 FILLCELL_X4 FILLER_67_375 ();
 FILLCELL_X1 FILLER_67_379 ();
 FILLCELL_X32 FILLER_67_1518 ();
 FILLCELL_X32 FILLER_67_1550 ();
 FILLCELL_X32 FILLER_67_1582 ();
 FILLCELL_X32 FILLER_67_1614 ();
 FILLCELL_X32 FILLER_67_1646 ();
 FILLCELL_X32 FILLER_67_1678 ();
 FILLCELL_X32 FILLER_67_1710 ();
 FILLCELL_X16 FILLER_67_1742 ();
 FILLCELL_X4 FILLER_67_1758 ();
 FILLCELL_X16 FILLER_68_1 ();
 FILLCELL_X2 FILLER_68_17 ();
 FILLCELL_X1 FILLER_68_19 ();
 FILLCELL_X4 FILLER_68_30 ();
 FILLCELL_X4 FILLER_68_43 ();
 FILLCELL_X4 FILLER_68_56 ();
 FILLCELL_X8 FILLER_68_63 ();
 FILLCELL_X2 FILLER_68_71 ();
 FILLCELL_X4 FILLER_68_76 ();
 FILLCELL_X4 FILLER_68_83 ();
 FILLCELL_X8 FILLER_68_97 ();
 FILLCELL_X1 FILLER_68_105 ();
 FILLCELL_X4 FILLER_68_109 ();
 FILLCELL_X4 FILLER_68_116 ();
 FILLCELL_X1 FILLER_68_120 ();
 FILLCELL_X8 FILLER_68_124 ();
 FILLCELL_X2 FILLER_68_132 ();
 FILLCELL_X1 FILLER_68_134 ();
 FILLCELL_X8 FILLER_68_139 ();
 FILLCELL_X4 FILLER_68_154 ();
 FILLCELL_X4 FILLER_68_168 ();
 FILLCELL_X4 FILLER_68_175 ();
 FILLCELL_X2 FILLER_68_179 ();
 FILLCELL_X8 FILLER_68_184 ();
 FILLCELL_X4 FILLER_68_202 ();
 FILLCELL_X2 FILLER_68_206 ();
 FILLCELL_X1 FILLER_68_208 ();
 FILLCELL_X4 FILLER_68_216 ();
 FILLCELL_X4 FILLER_68_223 ();
 FILLCELL_X1 FILLER_68_227 ();
 FILLCELL_X4 FILLER_68_238 ();
 FILLCELL_X4 FILLER_68_252 ();
 FILLCELL_X8 FILLER_68_259 ();
 FILLCELL_X4 FILLER_68_267 ();
 FILLCELL_X8 FILLER_68_275 ();
 FILLCELL_X2 FILLER_68_283 ();
 FILLCELL_X4 FILLER_68_288 ();
 FILLCELL_X4 FILLER_68_296 ();
 FILLCELL_X8 FILLER_68_310 ();
 FILLCELL_X4 FILLER_68_318 ();
 FILLCELL_X1 FILLER_68_322 ();
 FILLCELL_X16 FILLER_68_326 ();
 FILLCELL_X4 FILLER_68_351 ();
 FILLCELL_X4 FILLER_68_358 ();
 FILLCELL_X2 FILLER_68_362 ();
 FILLCELL_X8 FILLER_68_367 ();
 FILLCELL_X4 FILLER_68_375 ();
 FILLCELL_X1 FILLER_68_379 ();
 FILLCELL_X32 FILLER_68_1518 ();
 FILLCELL_X32 FILLER_68_1550 ();
 FILLCELL_X32 FILLER_68_1582 ();
 FILLCELL_X32 FILLER_68_1614 ();
 FILLCELL_X32 FILLER_68_1646 ();
 FILLCELL_X32 FILLER_68_1678 ();
 FILLCELL_X32 FILLER_68_1710 ();
 FILLCELL_X16 FILLER_68_1742 ();
 FILLCELL_X4 FILLER_68_1758 ();
 FILLCELL_X4 FILLER_69_1 ();
 FILLCELL_X1 FILLER_69_5 ();
 FILLCELL_X4 FILLER_69_9 ();
 FILLCELL_X4 FILLER_69_23 ();
 FILLCELL_X4 FILLER_69_34 ();
 FILLCELL_X8 FILLER_69_41 ();
 FILLCELL_X2 FILLER_69_49 ();
 FILLCELL_X1 FILLER_69_51 ();
 FILLCELL_X16 FILLER_69_55 ();
 FILLCELL_X8 FILLER_69_74 ();
 FILLCELL_X4 FILLER_69_82 ();
 FILLCELL_X2 FILLER_69_86 ();
 FILLCELL_X8 FILLER_69_95 ();
 FILLCELL_X2 FILLER_69_103 ();
 FILLCELL_X4 FILLER_69_114 ();
 FILLCELL_X4 FILLER_69_120 ();
 FILLCELL_X4 FILLER_69_127 ();
 FILLCELL_X4 FILLER_69_135 ();
 FILLCELL_X8 FILLER_69_143 ();
 FILLCELL_X1 FILLER_69_151 ();
 FILLCELL_X4 FILLER_69_162 ();
 FILLCELL_X4 FILLER_69_168 ();
 FILLCELL_X1 FILLER_69_172 ();
 FILLCELL_X4 FILLER_69_182 ();
 FILLCELL_X4 FILLER_69_190 ();
 FILLCELL_X4 FILLER_69_197 ();
 FILLCELL_X2 FILLER_69_201 ();
 FILLCELL_X1 FILLER_69_203 ();
 FILLCELL_X4 FILLER_69_208 ();
 FILLCELL_X8 FILLER_69_222 ();
 FILLCELL_X4 FILLER_69_230 ();
 FILLCELL_X2 FILLER_69_234 ();
 FILLCELL_X4 FILLER_69_238 ();
 FILLCELL_X2 FILLER_69_242 ();
 FILLCELL_X16 FILLER_69_248 ();
 FILLCELL_X4 FILLER_69_264 ();
 FILLCELL_X1 FILLER_69_268 ();
 FILLCELL_X4 FILLER_69_278 ();
 FILLCELL_X8 FILLER_69_285 ();
 FILLCELL_X4 FILLER_69_293 ();
 FILLCELL_X2 FILLER_69_297 ();
 FILLCELL_X16 FILLER_69_309 ();
 FILLCELL_X4 FILLER_69_325 ();
 FILLCELL_X2 FILLER_69_329 ();
 FILLCELL_X1 FILLER_69_331 ();
 FILLCELL_X4 FILLER_69_342 ();
 FILLCELL_X4 FILLER_69_355 ();
 FILLCELL_X2 FILLER_69_359 ();
 FILLCELL_X4 FILLER_69_368 ();
 FILLCELL_X4 FILLER_69_376 ();
 FILLCELL_X32 FILLER_69_1518 ();
 FILLCELL_X32 FILLER_69_1550 ();
 FILLCELL_X32 FILLER_69_1582 ();
 FILLCELL_X32 FILLER_69_1614 ();
 FILLCELL_X32 FILLER_69_1646 ();
 FILLCELL_X32 FILLER_69_1678 ();
 FILLCELL_X32 FILLER_69_1710 ();
 FILLCELL_X8 FILLER_69_1742 ();
 FILLCELL_X4 FILLER_69_1750 ();
 FILLCELL_X1 FILLER_69_1754 ();
 FILLCELL_X4 FILLER_69_1758 ();
 FILLCELL_X4 FILLER_70_1 ();
 FILLCELL_X1 FILLER_70_5 ();
 FILLCELL_X8 FILLER_70_9 ();
 FILLCELL_X4 FILLER_70_21 ();
 FILLCELL_X4 FILLER_70_27 ();
 FILLCELL_X2 FILLER_70_31 ();
 FILLCELL_X1 FILLER_70_33 ();
 FILLCELL_X4 FILLER_70_44 ();
 FILLCELL_X4 FILLER_70_57 ();
 FILLCELL_X4 FILLER_70_64 ();
 FILLCELL_X2 FILLER_70_68 ();
 FILLCELL_X1 FILLER_70_70 ();
 FILLCELL_X4 FILLER_70_80 ();
 FILLCELL_X4 FILLER_70_87 ();
 FILLCELL_X2 FILLER_70_91 ();
 FILLCELL_X1 FILLER_70_93 ();
 FILLCELL_X4 FILLER_70_98 ();
 FILLCELL_X4 FILLER_70_104 ();
 FILLCELL_X2 FILLER_70_108 ();
 FILLCELL_X4 FILLER_70_114 ();
 FILLCELL_X2 FILLER_70_118 ();
 FILLCELL_X1 FILLER_70_120 ();
 FILLCELL_X4 FILLER_70_130 ();
 FILLCELL_X16 FILLER_70_143 ();
 FILLCELL_X2 FILLER_70_159 ();
 FILLCELL_X8 FILLER_70_164 ();
 FILLCELL_X4 FILLER_70_176 ();
 FILLCELL_X4 FILLER_70_189 ();
 FILLCELL_X8 FILLER_70_196 ();
 FILLCELL_X8 FILLER_70_208 ();
 FILLCELL_X8 FILLER_70_219 ();
 FILLCELL_X2 FILLER_70_227 ();
 FILLCELL_X8 FILLER_70_232 ();
 FILLCELL_X4 FILLER_70_240 ();
 FILLCELL_X2 FILLER_70_244 ();
 FILLCELL_X4 FILLER_70_250 ();
 FILLCELL_X4 FILLER_70_258 ();
 FILLCELL_X4 FILLER_70_266 ();
 FILLCELL_X4 FILLER_70_274 ();
 FILLCELL_X16 FILLER_70_280 ();
 FILLCELL_X1 FILLER_70_296 ();
 FILLCELL_X8 FILLER_70_299 ();
 FILLCELL_X4 FILLER_70_307 ();
 FILLCELL_X4 FILLER_70_314 ();
 FILLCELL_X4 FILLER_70_327 ();
 FILLCELL_X8 FILLER_70_333 ();
 FILLCELL_X4 FILLER_70_344 ();
 FILLCELL_X8 FILLER_70_351 ();
 FILLCELL_X4 FILLER_70_369 ();
 FILLCELL_X4 FILLER_70_375 ();
 FILLCELL_X1 FILLER_70_379 ();
 FILLCELL_X32 FILLER_70_1518 ();
 FILLCELL_X32 FILLER_70_1550 ();
 FILLCELL_X32 FILLER_70_1582 ();
 FILLCELL_X32 FILLER_70_1614 ();
 FILLCELL_X32 FILLER_70_1646 ();
 FILLCELL_X32 FILLER_70_1678 ();
 FILLCELL_X32 FILLER_70_1710 ();
 FILLCELL_X16 FILLER_70_1742 ();
 FILLCELL_X4 FILLER_70_1758 ();
 FILLCELL_X4 FILLER_71_1 ();
 FILLCELL_X4 FILLER_71_7 ();
 FILLCELL_X4 FILLER_71_18 ();
 FILLCELL_X4 FILLER_71_25 ();
 FILLCELL_X8 FILLER_71_31 ();
 FILLCELL_X1 FILLER_71_39 ();
 FILLCELL_X8 FILLER_71_43 ();
 FILLCELL_X4 FILLER_71_54 ();
 FILLCELL_X4 FILLER_71_61 ();
 FILLCELL_X8 FILLER_71_74 ();
 FILLCELL_X4 FILLER_71_92 ();
 FILLCELL_X4 FILLER_71_98 ();
 FILLCELL_X4 FILLER_71_109 ();
 FILLCELL_X8 FILLER_71_123 ();
 FILLCELL_X16 FILLER_71_134 ();
 FILLCELL_X4 FILLER_71_150 ();
 FILLCELL_X1 FILLER_71_154 ();
 FILLCELL_X8 FILLER_71_159 ();
 FILLCELL_X8 FILLER_71_171 ();
 FILLCELL_X1 FILLER_71_179 ();
 FILLCELL_X8 FILLER_71_184 ();
 FILLCELL_X1 FILLER_71_192 ();
 FILLCELL_X4 FILLER_71_200 ();
 FILLCELL_X8 FILLER_71_214 ();
 FILLCELL_X2 FILLER_71_222 ();
 FILLCELL_X4 FILLER_71_228 ();
 FILLCELL_X4 FILLER_71_236 ();
 FILLCELL_X4 FILLER_71_243 ();
 FILLCELL_X8 FILLER_71_266 ();
 FILLCELL_X1 FILLER_71_274 ();
 FILLCELL_X4 FILLER_71_279 ();
 FILLCELL_X8 FILLER_71_292 ();
 FILLCELL_X2 FILLER_71_300 ();
 FILLCELL_X4 FILLER_71_309 ();
 FILLCELL_X2 FILLER_71_313 ();
 FILLCELL_X4 FILLER_71_324 ();
 FILLCELL_X1 FILLER_71_328 ();
 FILLCELL_X8 FILLER_71_336 ();
 FILLCELL_X8 FILLER_71_348 ();
 FILLCELL_X4 FILLER_71_359 ();
 FILLCELL_X4 FILLER_71_373 ();
 FILLCELL_X2 FILLER_71_377 ();
 FILLCELL_X1 FILLER_71_379 ();
 FILLCELL_X32 FILLER_71_1518 ();
 FILLCELL_X32 FILLER_71_1550 ();
 FILLCELL_X32 FILLER_71_1582 ();
 FILLCELL_X32 FILLER_71_1614 ();
 FILLCELL_X32 FILLER_71_1646 ();
 FILLCELL_X32 FILLER_71_1678 ();
 FILLCELL_X32 FILLER_71_1710 ();
 FILLCELL_X16 FILLER_71_1742 ();
 FILLCELL_X4 FILLER_71_1758 ();
 FILLCELL_X4 FILLER_72_1 ();
 FILLCELL_X2 FILLER_72_5 ();
 FILLCELL_X8 FILLER_72_17 ();
 FILLCELL_X1 FILLER_72_25 ();
 FILLCELL_X4 FILLER_72_33 ();
 FILLCELL_X4 FILLER_72_46 ();
 FILLCELL_X4 FILLER_72_53 ();
 FILLCELL_X2 FILLER_72_57 ();
 FILLCELL_X1 FILLER_72_59 ();
 FILLCELL_X4 FILLER_72_67 ();
 FILLCELL_X4 FILLER_72_74 ();
 FILLCELL_X1 FILLER_72_78 ();
 FILLCELL_X8 FILLER_72_86 ();
 FILLCELL_X4 FILLER_72_97 ();
 FILLCELL_X4 FILLER_72_111 ();
 FILLCELL_X8 FILLER_72_118 ();
 FILLCELL_X4 FILLER_72_126 ();
 FILLCELL_X4 FILLER_72_137 ();
 FILLCELL_X4 FILLER_72_144 ();
 FILLCELL_X2 FILLER_72_148 ();
 FILLCELL_X1 FILLER_72_150 ();
 FILLCELL_X4 FILLER_72_160 ();
 FILLCELL_X4 FILLER_72_173 ();
 FILLCELL_X16 FILLER_72_181 ();
 FILLCELL_X4 FILLER_72_207 ();
 FILLCELL_X4 FILLER_72_213 ();
 FILLCELL_X1 FILLER_72_217 ();
 FILLCELL_X4 FILLER_72_227 ();
 FILLCELL_X4 FILLER_72_240 ();
 FILLCELL_X16 FILLER_72_247 ();
 FILLCELL_X4 FILLER_72_263 ();
 FILLCELL_X4 FILLER_72_270 ();
 FILLCELL_X4 FILLER_72_283 ();
 FILLCELL_X2 FILLER_72_287 ();
 FILLCELL_X1 FILLER_72_289 ();
 FILLCELL_X4 FILLER_72_294 ();
 FILLCELL_X8 FILLER_72_308 ();
 FILLCELL_X2 FILLER_72_316 ();
 FILLCELL_X4 FILLER_72_321 ();
 FILLCELL_X4 FILLER_72_328 ();
 FILLCELL_X8 FILLER_72_342 ();
 FILLCELL_X1 FILLER_72_350 ();
 FILLCELL_X16 FILLER_72_355 ();
 FILLCELL_X1 FILLER_72_371 ();
 FILLCELL_X4 FILLER_72_376 ();
 FILLCELL_X32 FILLER_72_1518 ();
 FILLCELL_X32 FILLER_72_1550 ();
 FILLCELL_X32 FILLER_72_1582 ();
 FILLCELL_X32 FILLER_72_1614 ();
 FILLCELL_X32 FILLER_72_1646 ();
 FILLCELL_X32 FILLER_72_1678 ();
 FILLCELL_X32 FILLER_72_1710 ();
 FILLCELL_X16 FILLER_72_1742 ();
 FILLCELL_X4 FILLER_72_1758 ();
 FILLCELL_X8 FILLER_73_1 ();
 FILLCELL_X1 FILLER_73_9 ();
 FILLCELL_X4 FILLER_73_20 ();
 FILLCELL_X8 FILLER_73_34 ();
 FILLCELL_X4 FILLER_73_42 ();
 FILLCELL_X4 FILLER_73_55 ();
 FILLCELL_X4 FILLER_73_62 ();
 FILLCELL_X2 FILLER_73_66 ();
 FILLCELL_X1 FILLER_73_68 ();
 FILLCELL_X4 FILLER_73_79 ();
 FILLCELL_X8 FILLER_73_85 ();
 FILLCELL_X4 FILLER_73_93 ();
 FILLCELL_X1 FILLER_73_97 ();
 FILLCELL_X8 FILLER_73_105 ();
 FILLCELL_X2 FILLER_73_113 ();
 FILLCELL_X8 FILLER_73_125 ();
 FILLCELL_X4 FILLER_73_133 ();
 FILLCELL_X2 FILLER_73_137 ();
 FILLCELL_X4 FILLER_73_149 ();
 FILLCELL_X8 FILLER_73_157 ();
 FILLCELL_X8 FILLER_73_168 ();
 FILLCELL_X4 FILLER_73_176 ();
 FILLCELL_X2 FILLER_73_180 ();
 FILLCELL_X16 FILLER_73_186 ();
 FILLCELL_X4 FILLER_73_202 ();
 FILLCELL_X2 FILLER_73_206 ();
 FILLCELL_X16 FILLER_73_211 ();
 FILLCELL_X4 FILLER_73_227 ();
 FILLCELL_X1 FILLER_73_231 ();
 FILLCELL_X16 FILLER_73_236 ();
 FILLCELL_X8 FILLER_73_252 ();
 FILLCELL_X1 FILLER_73_260 ();
 FILLCELL_X4 FILLER_73_265 ();
 FILLCELL_X2 FILLER_73_269 ();
 FILLCELL_X4 FILLER_73_281 ();
 FILLCELL_X1 FILLER_73_285 ();
 FILLCELL_X4 FILLER_73_289 ();
 FILLCELL_X4 FILLER_73_296 ();
 FILLCELL_X1 FILLER_73_300 ();
 FILLCELL_X8 FILLER_73_304 ();
 FILLCELL_X2 FILLER_73_312 ();
 FILLCELL_X4 FILLER_73_317 ();
 FILLCELL_X16 FILLER_73_325 ();
 FILLCELL_X1 FILLER_73_341 ();
 FILLCELL_X4 FILLER_73_345 ();
 FILLCELL_X8 FILLER_73_353 ();
 FILLCELL_X1 FILLER_73_361 ();
 FILLCELL_X8 FILLER_73_371 ();
 FILLCELL_X1 FILLER_73_379 ();
 FILLCELL_X32 FILLER_73_1518 ();
 FILLCELL_X32 FILLER_73_1550 ();
 FILLCELL_X32 FILLER_73_1582 ();
 FILLCELL_X32 FILLER_73_1614 ();
 FILLCELL_X32 FILLER_73_1646 ();
 FILLCELL_X32 FILLER_73_1678 ();
 FILLCELL_X32 FILLER_73_1710 ();
 FILLCELL_X16 FILLER_73_1742 ();
 FILLCELL_X4 FILLER_73_1758 ();
 FILLCELL_X8 FILLER_74_1 ();
 FILLCELL_X2 FILLER_74_9 ();
 FILLCELL_X4 FILLER_74_20 ();
 FILLCELL_X8 FILLER_74_27 ();
 FILLCELL_X4 FILLER_74_35 ();
 FILLCELL_X2 FILLER_74_39 ();
 FILLCELL_X8 FILLER_74_51 ();
 FILLCELL_X1 FILLER_74_59 ();
 FILLCELL_X8 FILLER_74_70 ();
 FILLCELL_X8 FILLER_74_88 ();
 FILLCELL_X1 FILLER_74_96 ();
 FILLCELL_X4 FILLER_74_107 ();
 FILLCELL_X4 FILLER_74_113 ();
 FILLCELL_X2 FILLER_74_117 ();
 FILLCELL_X8 FILLER_74_122 ();
 FILLCELL_X1 FILLER_74_130 ();
 FILLCELL_X4 FILLER_74_141 ();
 FILLCELL_X8 FILLER_74_147 ();
 FILLCELL_X2 FILLER_74_155 ();
 FILLCELL_X8 FILLER_74_160 ();
 FILLCELL_X1 FILLER_74_168 ();
 FILLCELL_X4 FILLER_74_176 ();
 FILLCELL_X8 FILLER_74_190 ();
 FILLCELL_X4 FILLER_74_201 ();
 FILLCELL_X4 FILLER_74_209 ();
 FILLCELL_X2 FILLER_74_213 ();
 FILLCELL_X8 FILLER_74_219 ();
 FILLCELL_X4 FILLER_74_227 ();
 FILLCELL_X2 FILLER_74_231 ();
 FILLCELL_X1 FILLER_74_233 ();
 FILLCELL_X4 FILLER_74_238 ();
 FILLCELL_X4 FILLER_74_246 ();
 FILLCELL_X8 FILLER_74_259 ();
 FILLCELL_X4 FILLER_74_277 ();
 FILLCELL_X8 FILLER_74_284 ();
 FILLCELL_X4 FILLER_74_292 ();
 FILLCELL_X8 FILLER_74_305 ();
 FILLCELL_X4 FILLER_74_313 ();
 FILLCELL_X4 FILLER_74_321 ();
 FILLCELL_X8 FILLER_74_334 ();
 FILLCELL_X8 FILLER_74_347 ();
 FILLCELL_X4 FILLER_74_364 ();
 FILLCELL_X8 FILLER_74_371 ();
 FILLCELL_X1 FILLER_74_379 ();
 FILLCELL_X32 FILLER_74_1518 ();
 FILLCELL_X32 FILLER_74_1550 ();
 FILLCELL_X32 FILLER_74_1582 ();
 FILLCELL_X32 FILLER_74_1614 ();
 FILLCELL_X32 FILLER_74_1646 ();
 FILLCELL_X32 FILLER_74_1678 ();
 FILLCELL_X32 FILLER_74_1710 ();
 FILLCELL_X16 FILLER_74_1742 ();
 FILLCELL_X4 FILLER_74_1758 ();
 FILLCELL_X4 FILLER_75_1 ();
 FILLCELL_X4 FILLER_75_8 ();
 FILLCELL_X8 FILLER_75_21 ();
 FILLCELL_X4 FILLER_75_29 ();
 FILLCELL_X4 FILLER_75_35 ();
 FILLCELL_X1 FILLER_75_39 ();
 FILLCELL_X4 FILLER_75_47 ();
 FILLCELL_X8 FILLER_75_54 ();
 FILLCELL_X4 FILLER_75_66 ();
 FILLCELL_X2 FILLER_75_70 ();
 FILLCELL_X8 FILLER_75_74 ();
 FILLCELL_X2 FILLER_75_82 ();
 FILLCELL_X1 FILLER_75_84 ();
 FILLCELL_X4 FILLER_75_88 ();
 FILLCELL_X8 FILLER_75_96 ();
 FILLCELL_X4 FILLER_75_107 ();
 FILLCELL_X4 FILLER_75_114 ();
 FILLCELL_X8 FILLER_75_127 ();
 FILLCELL_X4 FILLER_75_135 ();
 FILLCELL_X2 FILLER_75_139 ();
 FILLCELL_X1 FILLER_75_141 ();
 FILLCELL_X8 FILLER_75_145 ();
 FILLCELL_X1 FILLER_75_153 ();
 FILLCELL_X8 FILLER_75_158 ();
 FILLCELL_X1 FILLER_75_166 ();
 FILLCELL_X4 FILLER_75_177 ();
 FILLCELL_X1 FILLER_75_181 ();
 FILLCELL_X8 FILLER_75_185 ();
 FILLCELL_X4 FILLER_75_193 ();
 FILLCELL_X2 FILLER_75_197 ();
 FILLCELL_X4 FILLER_75_208 ();
 FILLCELL_X4 FILLER_75_221 ();
 FILLCELL_X4 FILLER_75_229 ();
 FILLCELL_X4 FILLER_75_237 ();
 FILLCELL_X4 FILLER_75_250 ();
 FILLCELL_X2 FILLER_75_254 ();
 FILLCELL_X1 FILLER_75_256 ();
 FILLCELL_X4 FILLER_75_260 ();
 FILLCELL_X8 FILLER_75_267 ();
 FILLCELL_X8 FILLER_75_282 ();
 FILLCELL_X4 FILLER_75_294 ();
 FILLCELL_X4 FILLER_75_302 ();
 FILLCELL_X4 FILLER_75_309 ();
 FILLCELL_X4 FILLER_75_317 ();
 FILLCELL_X4 FILLER_75_330 ();
 FILLCELL_X4 FILLER_75_337 ();
 FILLCELL_X4 FILLER_75_351 ();
 FILLCELL_X8 FILLER_75_358 ();
 FILLCELL_X4 FILLER_75_366 ();
 FILLCELL_X2 FILLER_75_370 ();
 FILLCELL_X1 FILLER_75_372 ();
 FILLCELL_X4 FILLER_75_376 ();
 FILLCELL_X32 FILLER_75_1518 ();
 FILLCELL_X32 FILLER_75_1550 ();
 FILLCELL_X32 FILLER_75_1582 ();
 FILLCELL_X32 FILLER_75_1614 ();
 FILLCELL_X32 FILLER_75_1646 ();
 FILLCELL_X32 FILLER_75_1678 ();
 FILLCELL_X32 FILLER_75_1710 ();
 FILLCELL_X16 FILLER_75_1742 ();
 FILLCELL_X4 FILLER_75_1758 ();
 FILLCELL_X8 FILLER_76_1 ();
 FILLCELL_X4 FILLER_76_18 ();
 FILLCELL_X2 FILLER_76_22 ();
 FILLCELL_X4 FILLER_76_34 ();
 FILLCELL_X2 FILLER_76_38 ();
 FILLCELL_X1 FILLER_76_40 ();
 FILLCELL_X8 FILLER_76_45 ();
 FILLCELL_X8 FILLER_76_56 ();
 FILLCELL_X16 FILLER_76_67 ();
 FILLCELL_X4 FILLER_76_86 ();
 FILLCELL_X4 FILLER_76_99 ();
 FILLCELL_X4 FILLER_76_107 ();
 FILLCELL_X2 FILLER_76_111 ();
 FILLCELL_X1 FILLER_76_113 ();
 FILLCELL_X8 FILLER_76_123 ();
 FILLCELL_X2 FILLER_76_131 ();
 FILLCELL_X4 FILLER_76_136 ();
 FILLCELL_X4 FILLER_76_144 ();
 FILLCELL_X4 FILLER_76_157 ();
 FILLCELL_X4 FILLER_76_165 ();
 FILLCELL_X2 FILLER_76_169 ();
 FILLCELL_X1 FILLER_76_171 ();
 FILLCELL_X4 FILLER_76_174 ();
 FILLCELL_X4 FILLER_76_181 ();
 FILLCELL_X2 FILLER_76_185 ();
 FILLCELL_X16 FILLER_76_191 ();
 FILLCELL_X4 FILLER_76_207 ();
 FILLCELL_X2 FILLER_76_211 ();
 FILLCELL_X1 FILLER_76_213 ();
 FILLCELL_X16 FILLER_76_217 ();
 FILLCELL_X8 FILLER_76_233 ();
 FILLCELL_X4 FILLER_76_244 ();
 FILLCELL_X4 FILLER_76_252 ();
 FILLCELL_X8 FILLER_76_259 ();
 FILLCELL_X2 FILLER_76_267 ();
 FILLCELL_X4 FILLER_76_271 ();
 FILLCELL_X8 FILLER_76_277 ();
 FILLCELL_X4 FILLER_76_285 ();
 FILLCELL_X1 FILLER_76_289 ();
 FILLCELL_X4 FILLER_76_294 ();
 FILLCELL_X4 FILLER_76_307 ();
 FILLCELL_X8 FILLER_76_314 ();
 FILLCELL_X1 FILLER_76_322 ();
 FILLCELL_X4 FILLER_76_326 ();
 FILLCELL_X8 FILLER_76_333 ();
 FILLCELL_X2 FILLER_76_341 ();
 FILLCELL_X16 FILLER_76_345 ();
 FILLCELL_X2 FILLER_76_361 ();
 FILLCELL_X1 FILLER_76_363 ();
 FILLCELL_X8 FILLER_76_370 ();
 FILLCELL_X2 FILLER_76_378 ();
 FILLCELL_X32 FILLER_76_1518 ();
 FILLCELL_X32 FILLER_76_1550 ();
 FILLCELL_X32 FILLER_76_1582 ();
 FILLCELL_X32 FILLER_76_1614 ();
 FILLCELL_X32 FILLER_76_1646 ();
 FILLCELL_X32 FILLER_76_1678 ();
 FILLCELL_X32 FILLER_76_1710 ();
 FILLCELL_X16 FILLER_76_1742 ();
 FILLCELL_X4 FILLER_76_1758 ();
 FILLCELL_X8 FILLER_77_1 ();
 FILLCELL_X1 FILLER_77_9 ();
 FILLCELL_X4 FILLER_77_20 ();
 FILLCELL_X4 FILLER_77_26 ();
 FILLCELL_X4 FILLER_77_34 ();
 FILLCELL_X4 FILLER_77_48 ();
 FILLCELL_X2 FILLER_77_52 ();
 FILLCELL_X1 FILLER_77_54 ();
 FILLCELL_X4 FILLER_77_59 ();
 FILLCELL_X8 FILLER_77_72 ();
 FILLCELL_X4 FILLER_77_80 ();
 FILLCELL_X4 FILLER_77_87 ();
 FILLCELL_X4 FILLER_77_100 ();
 FILLCELL_X8 FILLER_77_108 ();
 FILLCELL_X2 FILLER_77_116 ();
 FILLCELL_X16 FILLER_77_122 ();
 FILLCELL_X2 FILLER_77_138 ();
 FILLCELL_X1 FILLER_77_140 ();
 FILLCELL_X4 FILLER_77_150 ();
 FILLCELL_X8 FILLER_77_157 ();
 FILLCELL_X4 FILLER_77_165 ();
 FILLCELL_X4 FILLER_77_172 ();
 FILLCELL_X4 FILLER_77_179 ();
 FILLCELL_X4 FILLER_77_192 ();
 FILLCELL_X4 FILLER_77_200 ();
 FILLCELL_X16 FILLER_77_208 ();
 FILLCELL_X1 FILLER_77_224 ();
 FILLCELL_X4 FILLER_77_229 ();
 FILLCELL_X4 FILLER_77_237 ();
 FILLCELL_X2 FILLER_77_241 ();
 FILLCELL_X1 FILLER_77_243 ();
 FILLCELL_X4 FILLER_77_248 ();
 FILLCELL_X4 FILLER_77_254 ();
 FILLCELL_X4 FILLER_77_262 ();
 FILLCELL_X4 FILLER_77_270 ();
 FILLCELL_X4 FILLER_77_284 ();
 FILLCELL_X8 FILLER_77_291 ();
 FILLCELL_X2 FILLER_77_299 ();
 FILLCELL_X4 FILLER_77_304 ();
 FILLCELL_X16 FILLER_77_310 ();
 FILLCELL_X2 FILLER_77_326 ();
 FILLCELL_X1 FILLER_77_328 ();
 FILLCELL_X4 FILLER_77_332 ();
 FILLCELL_X2 FILLER_77_336 ();
 FILLCELL_X1 FILLER_77_338 ();
 FILLCELL_X4 FILLER_77_343 ();
 FILLCELL_X4 FILLER_77_350 ();
 FILLCELL_X4 FILLER_77_364 ();
 FILLCELL_X4 FILLER_77_375 ();
 FILLCELL_X1 FILLER_77_379 ();
 FILLCELL_X32 FILLER_77_1518 ();
 FILLCELL_X32 FILLER_77_1550 ();
 FILLCELL_X32 FILLER_77_1582 ();
 FILLCELL_X32 FILLER_77_1614 ();
 FILLCELL_X32 FILLER_77_1646 ();
 FILLCELL_X32 FILLER_77_1678 ();
 FILLCELL_X32 FILLER_77_1710 ();
 FILLCELL_X16 FILLER_77_1742 ();
 FILLCELL_X4 FILLER_77_1758 ();
 FILLCELL_X4 FILLER_78_1 ();
 FILLCELL_X4 FILLER_78_8 ();
 FILLCELL_X4 FILLER_78_15 ();
 FILLCELL_X4 FILLER_78_22 ();
 FILLCELL_X8 FILLER_78_29 ();
 FILLCELL_X2 FILLER_78_37 ();
 FILLCELL_X1 FILLER_78_39 ();
 FILLCELL_X8 FILLER_78_47 ();
 FILLCELL_X1 FILLER_78_55 ();
 FILLCELL_X4 FILLER_78_60 ();
 FILLCELL_X4 FILLER_78_73 ();
 FILLCELL_X8 FILLER_78_80 ();
 FILLCELL_X4 FILLER_78_88 ();
 FILLCELL_X1 FILLER_78_92 ();
 FILLCELL_X8 FILLER_78_96 ();
 FILLCELL_X4 FILLER_78_104 ();
 FILLCELL_X2 FILLER_78_108 ();
 FILLCELL_X1 FILLER_78_110 ();
 FILLCELL_X4 FILLER_78_115 ();
 FILLCELL_X4 FILLER_78_128 ();
 FILLCELL_X4 FILLER_78_135 ();
 FILLCELL_X8 FILLER_78_143 ();
 FILLCELL_X1 FILLER_78_151 ();
 FILLCELL_X4 FILLER_78_155 ();
 FILLCELL_X4 FILLER_78_163 ();
 FILLCELL_X1 FILLER_78_167 ();
 FILLCELL_X4 FILLER_78_172 ();
 FILLCELL_X8 FILLER_78_185 ();
 FILLCELL_X2 FILLER_78_193 ();
 FILLCELL_X1 FILLER_78_195 ();
 FILLCELL_X4 FILLER_78_200 ();
 FILLCELL_X4 FILLER_78_213 ();
 FILLCELL_X8 FILLER_78_220 ();
 FILLCELL_X4 FILLER_78_237 ();
 FILLCELL_X4 FILLER_78_244 ();
 FILLCELL_X4 FILLER_78_257 ();
 FILLCELL_X4 FILLER_78_270 ();
 FILLCELL_X2 FILLER_78_274 ();
 FILLCELL_X1 FILLER_78_276 ();
 FILLCELL_X4 FILLER_78_287 ();
 FILLCELL_X8 FILLER_78_298 ();
 FILLCELL_X1 FILLER_78_306 ();
 FILLCELL_X4 FILLER_78_311 ();
 FILLCELL_X8 FILLER_78_325 ();
 FILLCELL_X4 FILLER_78_343 ();
 FILLCELL_X4 FILLER_78_357 ();
 FILLCELL_X1 FILLER_78_361 ();
 FILLCELL_X4 FILLER_78_368 ();
 FILLCELL_X4 FILLER_78_375 ();
 FILLCELL_X1 FILLER_78_379 ();
 FILLCELL_X32 FILLER_78_1518 ();
 FILLCELL_X32 FILLER_78_1550 ();
 FILLCELL_X32 FILLER_78_1582 ();
 FILLCELL_X32 FILLER_78_1614 ();
 FILLCELL_X32 FILLER_78_1646 ();
 FILLCELL_X32 FILLER_78_1678 ();
 FILLCELL_X32 FILLER_78_1710 ();
 FILLCELL_X8 FILLER_78_1742 ();
 FILLCELL_X4 FILLER_78_1750 ();
 FILLCELL_X1 FILLER_78_1754 ();
 FILLCELL_X4 FILLER_78_1758 ();
 FILLCELL_X4 FILLER_79_1 ();
 FILLCELL_X1 FILLER_79_5 ();
 FILLCELL_X4 FILLER_79_9 ();
 FILLCELL_X8 FILLER_79_17 ();
 FILLCELL_X1 FILLER_79_25 ();
 FILLCELL_X4 FILLER_79_29 ();
 FILLCELL_X4 FILLER_79_36 ();
 FILLCELL_X4 FILLER_79_43 ();
 FILLCELL_X8 FILLER_79_57 ();
 FILLCELL_X8 FILLER_79_69 ();
 FILLCELL_X4 FILLER_79_77 ();
 FILLCELL_X2 FILLER_79_81 ();
 FILLCELL_X1 FILLER_79_83 ();
 FILLCELL_X4 FILLER_79_88 ();
 FILLCELL_X8 FILLER_79_102 ();
 FILLCELL_X1 FILLER_79_110 ();
 FILLCELL_X4 FILLER_79_114 ();
 FILLCELL_X4 FILLER_79_122 ();
 FILLCELL_X4 FILLER_79_135 ();
 FILLCELL_X2 FILLER_79_139 ();
 FILLCELL_X4 FILLER_79_148 ();
 FILLCELL_X2 FILLER_79_152 ();
 FILLCELL_X1 FILLER_79_154 ();
 FILLCELL_X4 FILLER_79_159 ();
 FILLCELL_X4 FILLER_79_172 ();
 FILLCELL_X16 FILLER_79_180 ();
 FILLCELL_X2 FILLER_79_196 ();
 FILLCELL_X4 FILLER_79_201 ();
 FILLCELL_X8 FILLER_79_209 ();
 FILLCELL_X2 FILLER_79_217 ();
 FILLCELL_X4 FILLER_79_222 ();
 FILLCELL_X4 FILLER_79_230 ();
 FILLCELL_X8 FILLER_79_243 ();
 FILLCELL_X1 FILLER_79_251 ();
 FILLCELL_X4 FILLER_79_255 ();
 FILLCELL_X16 FILLER_79_262 ();
 FILLCELL_X1 FILLER_79_278 ();
 FILLCELL_X8 FILLER_79_282 ();
 FILLCELL_X2 FILLER_79_290 ();
 FILLCELL_X4 FILLER_79_301 ();
 FILLCELL_X2 FILLER_79_305 ();
 FILLCELL_X4 FILLER_79_317 ();
 FILLCELL_X8 FILLER_79_325 ();
 FILLCELL_X4 FILLER_79_333 ();
 FILLCELL_X8 FILLER_79_346 ();
 FILLCELL_X4 FILLER_79_358 ();
 FILLCELL_X16 FILLER_79_364 ();
 FILLCELL_X32 FILLER_79_1518 ();
 FILLCELL_X32 FILLER_79_1550 ();
 FILLCELL_X32 FILLER_79_1582 ();
 FILLCELL_X32 FILLER_79_1614 ();
 FILLCELL_X32 FILLER_79_1646 ();
 FILLCELL_X32 FILLER_79_1678 ();
 FILLCELL_X32 FILLER_79_1710 ();
 FILLCELL_X16 FILLER_79_1742 ();
 FILLCELL_X4 FILLER_79_1758 ();
 FILLCELL_X4 FILLER_80_1 ();
 FILLCELL_X2 FILLER_80_5 ();
 FILLCELL_X1 FILLER_80_7 ();
 FILLCELL_X4 FILLER_80_17 ();
 FILLCELL_X1 FILLER_80_21 ();
 FILLCELL_X4 FILLER_80_31 ();
 FILLCELL_X4 FILLER_80_44 ();
 FILLCELL_X1 FILLER_80_48 ();
 FILLCELL_X4 FILLER_80_51 ();
 FILLCELL_X2 FILLER_80_55 ();
 FILLCELL_X1 FILLER_80_57 ();
 FILLCELL_X4 FILLER_80_61 ();
 FILLCELL_X8 FILLER_80_75 ();
 FILLCELL_X1 FILLER_80_83 ();
 FILLCELL_X4 FILLER_80_86 ();
 FILLCELL_X4 FILLER_80_97 ();
 FILLCELL_X8 FILLER_80_105 ();
 FILLCELL_X4 FILLER_80_113 ();
 FILLCELL_X8 FILLER_80_120 ();
 FILLCELL_X4 FILLER_80_128 ();
 FILLCELL_X4 FILLER_80_135 ();
 FILLCELL_X4 FILLER_80_149 ();
 FILLCELL_X4 FILLER_80_155 ();
 FILLCELL_X1 FILLER_80_159 ();
 FILLCELL_X4 FILLER_80_163 ();
 FILLCELL_X1 FILLER_80_167 ();
 FILLCELL_X4 FILLER_80_171 ();
 FILLCELL_X8 FILLER_80_184 ();
 FILLCELL_X4 FILLER_80_195 ();
 FILLCELL_X2 FILLER_80_199 ();
 FILLCELL_X4 FILLER_80_204 ();
 FILLCELL_X16 FILLER_80_217 ();
 FILLCELL_X8 FILLER_80_236 ();
 FILLCELL_X4 FILLER_80_244 ();
 FILLCELL_X16 FILLER_80_251 ();
 FILLCELL_X4 FILLER_80_267 ();
 FILLCELL_X8 FILLER_80_275 ();
 FILLCELL_X1 FILLER_80_283 ();
 FILLCELL_X4 FILLER_80_293 ();
 FILLCELL_X4 FILLER_80_300 ();
 FILLCELL_X2 FILLER_80_304 ();
 FILLCELL_X1 FILLER_80_306 ();
 FILLCELL_X4 FILLER_80_310 ();
 FILLCELL_X1 FILLER_80_314 ();
 FILLCELL_X4 FILLER_80_318 ();
 FILLCELL_X8 FILLER_80_324 ();
 FILLCELL_X2 FILLER_80_332 ();
 FILLCELL_X1 FILLER_80_334 ();
 FILLCELL_X4 FILLER_80_338 ();
 FILLCELL_X16 FILLER_80_345 ();
 FILLCELL_X2 FILLER_80_361 ();
 FILLCELL_X8 FILLER_80_367 ();
 FILLCELL_X4 FILLER_80_375 ();
 FILLCELL_X1 FILLER_80_379 ();
 FILLCELL_X32 FILLER_80_1518 ();
 FILLCELL_X32 FILLER_80_1550 ();
 FILLCELL_X32 FILLER_80_1582 ();
 FILLCELL_X32 FILLER_80_1614 ();
 FILLCELL_X32 FILLER_80_1646 ();
 FILLCELL_X32 FILLER_80_1678 ();
 FILLCELL_X32 FILLER_80_1710 ();
 FILLCELL_X16 FILLER_80_1742 ();
 FILLCELL_X4 FILLER_80_1758 ();
 FILLCELL_X8 FILLER_81_1 ();
 FILLCELL_X1 FILLER_81_9 ();
 FILLCELL_X4 FILLER_81_14 ();
 FILLCELL_X4 FILLER_81_22 ();
 FILLCELL_X4 FILLER_81_30 ();
 FILLCELL_X16 FILLER_81_37 ();
 FILLCELL_X2 FILLER_81_53 ();
 FILLCELL_X1 FILLER_81_55 ();
 FILLCELL_X4 FILLER_81_58 ();
 FILLCELL_X4 FILLER_81_69 ();
 FILLCELL_X8 FILLER_81_83 ();
 FILLCELL_X2 FILLER_81_91 ();
 FILLCELL_X4 FILLER_81_103 ();
 FILLCELL_X1 FILLER_81_107 ();
 FILLCELL_X8 FILLER_81_111 ();
 FILLCELL_X2 FILLER_81_119 ();
 FILLCELL_X16 FILLER_81_125 ();
 FILLCELL_X8 FILLER_81_141 ();
 FILLCELL_X1 FILLER_81_149 ();
 FILLCELL_X16 FILLER_81_160 ();
 FILLCELL_X4 FILLER_81_176 ();
 FILLCELL_X2 FILLER_81_180 ();
 FILLCELL_X1 FILLER_81_182 ();
 FILLCELL_X4 FILLER_81_187 ();
 FILLCELL_X8 FILLER_81_201 ();
 FILLCELL_X4 FILLER_81_209 ();
 FILLCELL_X1 FILLER_81_213 ();
 FILLCELL_X4 FILLER_81_218 ();
 FILLCELL_X8 FILLER_81_229 ();
 FILLCELL_X1 FILLER_81_237 ();
 FILLCELL_X4 FILLER_81_242 ();
 FILLCELL_X8 FILLER_81_256 ();
 FILLCELL_X2 FILLER_81_264 ();
 FILLCELL_X1 FILLER_81_266 ();
 FILLCELL_X4 FILLER_81_271 ();
 FILLCELL_X8 FILLER_81_284 ();
 FILLCELL_X8 FILLER_81_295 ();
 FILLCELL_X2 FILLER_81_303 ();
 FILLCELL_X1 FILLER_81_305 ();
 FILLCELL_X4 FILLER_81_316 ();
 FILLCELL_X4 FILLER_81_330 ();
 FILLCELL_X4 FILLER_81_343 ();
 FILLCELL_X4 FILLER_81_350 ();
 FILLCELL_X2 FILLER_81_354 ();
 FILLCELL_X1 FILLER_81_356 ();
 FILLCELL_X4 FILLER_81_376 ();
 FILLCELL_X32 FILLER_81_1518 ();
 FILLCELL_X32 FILLER_81_1550 ();
 FILLCELL_X32 FILLER_81_1582 ();
 FILLCELL_X32 FILLER_81_1614 ();
 FILLCELL_X32 FILLER_81_1646 ();
 FILLCELL_X32 FILLER_81_1678 ();
 FILLCELL_X32 FILLER_81_1710 ();
 FILLCELL_X16 FILLER_81_1742 ();
 FILLCELL_X4 FILLER_81_1758 ();
 FILLCELL_X4 FILLER_82_1 ();
 FILLCELL_X2 FILLER_82_5 ();
 FILLCELL_X8 FILLER_82_16 ();
 FILLCELL_X4 FILLER_82_34 ();
 FILLCELL_X2 FILLER_82_38 ();
 FILLCELL_X1 FILLER_82_40 ();
 FILLCELL_X16 FILLER_82_45 ();
 FILLCELL_X4 FILLER_82_64 ();
 FILLCELL_X8 FILLER_82_71 ();
 FILLCELL_X2 FILLER_82_79 ();
 FILLCELL_X1 FILLER_82_81 ();
 FILLCELL_X4 FILLER_82_85 ();
 FILLCELL_X4 FILLER_82_93 ();
 FILLCELL_X4 FILLER_82_106 ();
 FILLCELL_X1 FILLER_82_110 ();
 FILLCELL_X4 FILLER_82_115 ();
 FILLCELL_X4 FILLER_82_128 ();
 FILLCELL_X4 FILLER_82_136 ();
 FILLCELL_X2 FILLER_82_140 ();
 FILLCELL_X1 FILLER_82_142 ();
 FILLCELL_X4 FILLER_82_146 ();
 FILLCELL_X2 FILLER_82_150 ();
 FILLCELL_X1 FILLER_82_152 ();
 FILLCELL_X4 FILLER_82_157 ();
 FILLCELL_X4 FILLER_82_164 ();
 FILLCELL_X4 FILLER_82_178 ();
 FILLCELL_X4 FILLER_82_186 ();
 FILLCELL_X1 FILLER_82_190 ();
 FILLCELL_X4 FILLER_82_198 ();
 FILLCELL_X4 FILLER_82_212 ();
 FILLCELL_X4 FILLER_82_226 ();
 FILLCELL_X4 FILLER_82_240 ();
 FILLCELL_X4 FILLER_82_251 ();
 FILLCELL_X8 FILLER_82_265 ();
 FILLCELL_X2 FILLER_82_273 ();
 FILLCELL_X4 FILLER_82_279 ();
 FILLCELL_X4 FILLER_82_285 ();
 FILLCELL_X1 FILLER_82_289 ();
 FILLCELL_X4 FILLER_82_293 ();
 FILLCELL_X16 FILLER_82_304 ();
 FILLCELL_X8 FILLER_82_327 ();
 FILLCELL_X4 FILLER_82_344 ();
 FILLCELL_X4 FILLER_82_358 ();
 FILLCELL_X16 FILLER_82_364 ();
 FILLCELL_X32 FILLER_82_1518 ();
 FILLCELL_X32 FILLER_82_1550 ();
 FILLCELL_X32 FILLER_82_1582 ();
 FILLCELL_X32 FILLER_82_1614 ();
 FILLCELL_X32 FILLER_82_1646 ();
 FILLCELL_X32 FILLER_82_1678 ();
 FILLCELL_X32 FILLER_82_1710 ();
 FILLCELL_X16 FILLER_82_1742 ();
 FILLCELL_X4 FILLER_82_1758 ();
 FILLCELL_X4 FILLER_83_1 ();
 FILLCELL_X16 FILLER_83_8 ();
 FILLCELL_X4 FILLER_83_31 ();
 FILLCELL_X1 FILLER_83_35 ();
 FILLCELL_X4 FILLER_83_39 ();
 FILLCELL_X8 FILLER_83_52 ();
 FILLCELL_X1 FILLER_83_60 ();
 FILLCELL_X4 FILLER_83_70 ();
 FILLCELL_X4 FILLER_83_77 ();
 FILLCELL_X2 FILLER_83_81 ();
 FILLCELL_X1 FILLER_83_83 ();
 FILLCELL_X4 FILLER_83_87 ();
 FILLCELL_X4 FILLER_83_100 ();
 FILLCELL_X16 FILLER_83_108 ();
 FILLCELL_X4 FILLER_83_124 ();
 FILLCELL_X2 FILLER_83_128 ();
 FILLCELL_X4 FILLER_83_137 ();
 FILLCELL_X8 FILLER_83_151 ();
 FILLCELL_X2 FILLER_83_159 ();
 FILLCELL_X1 FILLER_83_161 ();
 FILLCELL_X4 FILLER_83_169 ();
 FILLCELL_X16 FILLER_83_175 ();
 FILLCELL_X8 FILLER_83_191 ();
 FILLCELL_X16 FILLER_83_201 ();
 FILLCELL_X4 FILLER_83_217 ();
 FILLCELL_X4 FILLER_83_224 ();
 FILLCELL_X16 FILLER_83_230 ();
 FILLCELL_X4 FILLER_83_246 ();
 FILLCELL_X2 FILLER_83_250 ();
 FILLCELL_X1 FILLER_83_252 ();
 FILLCELL_X4 FILLER_83_255 ();
 FILLCELL_X4 FILLER_83_262 ();
 FILLCELL_X4 FILLER_83_269 ();
 FILLCELL_X4 FILLER_83_282 ();
 FILLCELL_X4 FILLER_83_296 ();
 FILLCELL_X4 FILLER_83_310 ();
 FILLCELL_X16 FILLER_83_323 ();
 FILLCELL_X2 FILLER_83_339 ();
 FILLCELL_X4 FILLER_83_344 ();
 FILLCELL_X4 FILLER_83_350 ();
 FILLCELL_X16 FILLER_83_361 ();
 FILLCELL_X2 FILLER_83_377 ();
 FILLCELL_X1 FILLER_83_379 ();
 FILLCELL_X32 FILLER_83_1518 ();
 FILLCELL_X32 FILLER_83_1550 ();
 FILLCELL_X32 FILLER_83_1582 ();
 FILLCELL_X32 FILLER_83_1614 ();
 FILLCELL_X32 FILLER_83_1646 ();
 FILLCELL_X32 FILLER_83_1678 ();
 FILLCELL_X32 FILLER_83_1710 ();
 FILLCELL_X16 FILLER_83_1742 ();
 FILLCELL_X4 FILLER_83_1758 ();
 FILLCELL_X8 FILLER_84_1 ();
 FILLCELL_X4 FILLER_84_12 ();
 FILLCELL_X2 FILLER_84_16 ();
 FILLCELL_X1 FILLER_84_18 ();
 FILLCELL_X4 FILLER_84_21 ();
 FILLCELL_X4 FILLER_84_35 ();
 FILLCELL_X1 FILLER_84_39 ();
 FILLCELL_X4 FILLER_84_43 ();
 FILLCELL_X8 FILLER_84_50 ();
 FILLCELL_X4 FILLER_84_58 ();
 FILLCELL_X1 FILLER_84_62 ();
 FILLCELL_X4 FILLER_84_72 ();
 FILLCELL_X8 FILLER_84_79 ();
 FILLCELL_X4 FILLER_84_87 ();
 FILLCELL_X2 FILLER_84_91 ();
 FILLCELL_X16 FILLER_84_97 ();
 FILLCELL_X4 FILLER_84_113 ();
 FILLCELL_X1 FILLER_84_117 ();
 FILLCELL_X8 FILLER_84_121 ();
 FILLCELL_X2 FILLER_84_129 ();
 FILLCELL_X1 FILLER_84_131 ();
 FILLCELL_X4 FILLER_84_142 ();
 FILLCELL_X8 FILLER_84_148 ();
 FILLCELL_X2 FILLER_84_156 ();
 FILLCELL_X4 FILLER_84_168 ();
 FILLCELL_X4 FILLER_84_175 ();
 FILLCELL_X4 FILLER_84_183 ();
 FILLCELL_X4 FILLER_84_191 ();
 FILLCELL_X1 FILLER_84_195 ();
 FILLCELL_X8 FILLER_84_200 ();
 FILLCELL_X4 FILLER_84_208 ();
 FILLCELL_X2 FILLER_84_212 ();
 FILLCELL_X4 FILLER_84_218 ();
 FILLCELL_X16 FILLER_84_226 ();
 FILLCELL_X2 FILLER_84_242 ();
 FILLCELL_X4 FILLER_84_248 ();
 FILLCELL_X2 FILLER_84_252 ();
 FILLCELL_X4 FILLER_84_257 ();
 FILLCELL_X4 FILLER_84_266 ();
 FILLCELL_X4 FILLER_84_279 ();
 FILLCELL_X8 FILLER_84_288 ();
 FILLCELL_X1 FILLER_84_296 ();
 FILLCELL_X32 FILLER_84_299 ();
 FILLCELL_X2 FILLER_84_331 ();
 FILLCELL_X1 FILLER_84_333 ();
 FILLCELL_X8 FILLER_84_344 ();
 FILLCELL_X1 FILLER_84_352 ();
 FILLCELL_X4 FILLER_84_356 ();
 FILLCELL_X8 FILLER_84_370 ();
 FILLCELL_X2 FILLER_84_378 ();
 FILLCELL_X32 FILLER_84_1518 ();
 FILLCELL_X32 FILLER_84_1550 ();
 FILLCELL_X32 FILLER_84_1582 ();
 FILLCELL_X32 FILLER_84_1614 ();
 FILLCELL_X32 FILLER_84_1646 ();
 FILLCELL_X32 FILLER_84_1678 ();
 FILLCELL_X32 FILLER_84_1710 ();
 FILLCELL_X16 FILLER_84_1742 ();
 FILLCELL_X4 FILLER_84_1758 ();
 FILLCELL_X4 FILLER_85_1 ();
 FILLCELL_X2 FILLER_85_5 ();
 FILLCELL_X4 FILLER_85_17 ();
 FILLCELL_X8 FILLER_85_25 ();
 FILLCELL_X1 FILLER_85_33 ();
 FILLCELL_X4 FILLER_85_38 ();
 FILLCELL_X8 FILLER_85_51 ();
 FILLCELL_X4 FILLER_85_69 ();
 FILLCELL_X8 FILLER_85_83 ();
 FILLCELL_X2 FILLER_85_91 ();
 FILLCELL_X1 FILLER_85_93 ();
 FILLCELL_X8 FILLER_85_98 ();
 FILLCELL_X4 FILLER_85_109 ();
 FILLCELL_X4 FILLER_85_122 ();
 FILLCELL_X8 FILLER_85_135 ();
 FILLCELL_X4 FILLER_85_143 ();
 FILLCELL_X16 FILLER_85_150 ();
 FILLCELL_X2 FILLER_85_166 ();
 FILLCELL_X4 FILLER_85_171 ();
 FILLCELL_X8 FILLER_85_184 ();
 FILLCELL_X4 FILLER_85_192 ();
 FILLCELL_X4 FILLER_85_200 ();
 FILLCELL_X2 FILLER_85_204 ();
 FILLCELL_X4 FILLER_85_210 ();
 FILLCELL_X2 FILLER_85_214 ();
 FILLCELL_X1 FILLER_85_216 ();
 FILLCELL_X4 FILLER_85_226 ();
 FILLCELL_X4 FILLER_85_233 ();
 FILLCELL_X1 FILLER_85_237 ();
 FILLCELL_X4 FILLER_85_242 ();
 FILLCELL_X4 FILLER_85_255 ();
 FILLCELL_X2 FILLER_85_259 ();
 FILLCELL_X1 FILLER_85_261 ();
 FILLCELL_X4 FILLER_85_265 ();
 FILLCELL_X4 FILLER_85_279 ();
 FILLCELL_X16 FILLER_85_286 ();
 FILLCELL_X4 FILLER_85_302 ();
 FILLCELL_X1 FILLER_85_306 ();
 FILLCELL_X4 FILLER_85_309 ();
 FILLCELL_X1 FILLER_85_313 ();
 FILLCELL_X4 FILLER_85_317 ();
 FILLCELL_X4 FILLER_85_324 ();
 FILLCELL_X4 FILLER_85_338 ();
 FILLCELL_X4 FILLER_85_349 ();
 FILLCELL_X4 FILLER_85_356 ();
 FILLCELL_X2 FILLER_85_360 ();
 FILLCELL_X8 FILLER_85_366 ();
 FILLCELL_X4 FILLER_85_374 ();
 FILLCELL_X2 FILLER_85_378 ();
 FILLCELL_X32 FILLER_85_1518 ();
 FILLCELL_X32 FILLER_85_1550 ();
 FILLCELL_X32 FILLER_85_1582 ();
 FILLCELL_X32 FILLER_85_1614 ();
 FILLCELL_X32 FILLER_85_1646 ();
 FILLCELL_X32 FILLER_85_1678 ();
 FILLCELL_X32 FILLER_85_1710 ();
 FILLCELL_X16 FILLER_85_1742 ();
 FILLCELL_X4 FILLER_85_1758 ();
 FILLCELL_X8 FILLER_86_1 ();
 FILLCELL_X2 FILLER_86_9 ();
 FILLCELL_X4 FILLER_86_18 ();
 FILLCELL_X4 FILLER_86_31 ();
 FILLCELL_X16 FILLER_86_38 ();
 FILLCELL_X4 FILLER_86_54 ();
 FILLCELL_X2 FILLER_86_58 ();
 FILLCELL_X1 FILLER_86_60 ();
 FILLCELL_X4 FILLER_86_64 ();
 FILLCELL_X4 FILLER_86_75 ();
 FILLCELL_X4 FILLER_86_81 ();
 FILLCELL_X1 FILLER_86_85 ();
 FILLCELL_X4 FILLER_86_89 ();
 FILLCELL_X4 FILLER_86_102 ();
 FILLCELL_X8 FILLER_86_110 ();
 FILLCELL_X2 FILLER_86_118 ();
 FILLCELL_X1 FILLER_86_120 ();
 FILLCELL_X8 FILLER_86_124 ();
 FILLCELL_X1 FILLER_86_132 ();
 FILLCELL_X4 FILLER_86_136 ();
 FILLCELL_X4 FILLER_86_144 ();
 FILLCELL_X2 FILLER_86_148 ();
 FILLCELL_X4 FILLER_86_154 ();
 FILLCELL_X8 FILLER_86_162 ();
 FILLCELL_X2 FILLER_86_170 ();
 FILLCELL_X1 FILLER_86_172 ();
 FILLCELL_X4 FILLER_86_177 ();
 FILLCELL_X4 FILLER_86_184 ();
 FILLCELL_X4 FILLER_86_191 ();
 FILLCELL_X8 FILLER_86_204 ();
 FILLCELL_X2 FILLER_86_212 ();
 FILLCELL_X4 FILLER_86_218 ();
 FILLCELL_X4 FILLER_86_231 ();
 FILLCELL_X2 FILLER_86_235 ();
 FILLCELL_X1 FILLER_86_237 ();
 FILLCELL_X4 FILLER_86_241 ();
 FILLCELL_X4 FILLER_86_249 ();
 FILLCELL_X4 FILLER_86_262 ();
 FILLCELL_X1 FILLER_86_266 ();
 FILLCELL_X16 FILLER_86_271 ();
 FILLCELL_X8 FILLER_86_287 ();
 FILLCELL_X4 FILLER_86_295 ();
 FILLCELL_X2 FILLER_86_299 ();
 FILLCELL_X4 FILLER_86_305 ();
 FILLCELL_X2 FILLER_86_309 ();
 FILLCELL_X4 FILLER_86_321 ();
 FILLCELL_X2 FILLER_86_325 ();
 FILLCELL_X1 FILLER_86_327 ();
 FILLCELL_X4 FILLER_86_331 ();
 FILLCELL_X8 FILLER_86_344 ();
 FILLCELL_X4 FILLER_86_356 ();
 FILLCELL_X8 FILLER_86_369 ();
 FILLCELL_X2 FILLER_86_377 ();
 FILLCELL_X1 FILLER_86_379 ();
 FILLCELL_X32 FILLER_86_1518 ();
 FILLCELL_X32 FILLER_86_1550 ();
 FILLCELL_X32 FILLER_86_1582 ();
 FILLCELL_X32 FILLER_86_1614 ();
 FILLCELL_X32 FILLER_86_1646 ();
 FILLCELL_X32 FILLER_86_1678 ();
 FILLCELL_X32 FILLER_86_1710 ();
 FILLCELL_X16 FILLER_86_1742 ();
 FILLCELL_X4 FILLER_86_1758 ();
 FILLCELL_X4 FILLER_87_1 ();
 FILLCELL_X1 FILLER_87_5 ();
 FILLCELL_X4 FILLER_87_9 ();
 FILLCELL_X8 FILLER_87_15 ();
 FILLCELL_X4 FILLER_87_26 ();
 FILLCELL_X1 FILLER_87_30 ();
 FILLCELL_X4 FILLER_87_34 ();
 FILLCELL_X8 FILLER_87_47 ();
 FILLCELL_X4 FILLER_87_62 ();
 FILLCELL_X8 FILLER_87_76 ();
 FILLCELL_X2 FILLER_87_84 ();
 FILLCELL_X1 FILLER_87_86 ();
 FILLCELL_X8 FILLER_87_91 ();
 FILLCELL_X4 FILLER_87_108 ();
 FILLCELL_X4 FILLER_87_115 ();
 FILLCELL_X2 FILLER_87_119 ();
 FILLCELL_X1 FILLER_87_121 ();
 FILLCELL_X4 FILLER_87_126 ();
 FILLCELL_X2 FILLER_87_130 ();
 FILLCELL_X4 FILLER_87_141 ();
 FILLCELL_X8 FILLER_87_154 ();
 FILLCELL_X4 FILLER_87_162 ();
 FILLCELL_X1 FILLER_87_166 ();
 FILLCELL_X8 FILLER_87_176 ();
 FILLCELL_X1 FILLER_87_184 ();
 FILLCELL_X4 FILLER_87_188 ();
 FILLCELL_X4 FILLER_87_195 ();
 FILLCELL_X8 FILLER_87_208 ();
 FILLCELL_X4 FILLER_87_219 ();
 FILLCELL_X4 FILLER_87_226 ();
 FILLCELL_X8 FILLER_87_233 ();
 FILLCELL_X4 FILLER_87_241 ();
 FILLCELL_X4 FILLER_87_248 ();
 FILLCELL_X1 FILLER_87_252 ();
 FILLCELL_X4 FILLER_87_256 ();
 FILLCELL_X4 FILLER_87_270 ();
 FILLCELL_X4 FILLER_87_299 ();
 FILLCELL_X1 FILLER_87_303 ();
 FILLCELL_X4 FILLER_87_314 ();
 FILLCELL_X4 FILLER_87_327 ();
 FILLCELL_X16 FILLER_87_334 ();
 FILLCELL_X1 FILLER_87_350 ();
 FILLCELL_X4 FILLER_87_355 ();
 FILLCELL_X4 FILLER_87_368 ();
 FILLCELL_X4 FILLER_87_375 ();
 FILLCELL_X1 FILLER_87_379 ();
 FILLCELL_X32 FILLER_87_1518 ();
 FILLCELL_X32 FILLER_87_1550 ();
 FILLCELL_X32 FILLER_87_1582 ();
 FILLCELL_X32 FILLER_87_1614 ();
 FILLCELL_X32 FILLER_87_1646 ();
 FILLCELL_X32 FILLER_87_1678 ();
 FILLCELL_X32 FILLER_87_1710 ();
 FILLCELL_X16 FILLER_87_1742 ();
 FILLCELL_X4 FILLER_87_1758 ();
 FILLCELL_X8 FILLER_88_1 ();
 FILLCELL_X2 FILLER_88_9 ();
 FILLCELL_X4 FILLER_88_21 ();
 FILLCELL_X16 FILLER_88_28 ();
 FILLCELL_X1 FILLER_88_44 ();
 FILLCELL_X8 FILLER_88_48 ();
 FILLCELL_X2 FILLER_88_56 ();
 FILLCELL_X1 FILLER_88_58 ();
 FILLCELL_X4 FILLER_88_61 ();
 FILLCELL_X1 FILLER_88_65 ();
 FILLCELL_X8 FILLER_88_69 ();
 FILLCELL_X1 FILLER_88_77 ();
 FILLCELL_X4 FILLER_88_81 ();
 FILLCELL_X2 FILLER_88_85 ();
 FILLCELL_X4 FILLER_88_90 ();
 FILLCELL_X4 FILLER_88_97 ();
 FILLCELL_X1 FILLER_88_101 ();
 FILLCELL_X8 FILLER_88_109 ();
 FILLCELL_X4 FILLER_88_120 ();
 FILLCELL_X4 FILLER_88_127 ();
 FILLCELL_X4 FILLER_88_133 ();
 FILLCELL_X2 FILLER_88_137 ();
 FILLCELL_X1 FILLER_88_139 ();
 FILLCELL_X8 FILLER_88_143 ();
 FILLCELL_X4 FILLER_88_151 ();
 FILLCELL_X2 FILLER_88_155 ();
 FILLCELL_X4 FILLER_88_160 ();
 FILLCELL_X2 FILLER_88_164 ();
 FILLCELL_X8 FILLER_88_170 ();
 FILLCELL_X1 FILLER_88_178 ();
 FILLCELL_X4 FILLER_88_183 ();
 FILLCELL_X4 FILLER_88_191 ();
 FILLCELL_X8 FILLER_88_198 ();
 FILLCELL_X1 FILLER_88_206 ();
 FILLCELL_X8 FILLER_88_211 ();
 FILLCELL_X2 FILLER_88_219 ();
 FILLCELL_X4 FILLER_88_225 ();
 FILLCELL_X4 FILLER_88_239 ();
 FILLCELL_X2 FILLER_88_243 ();
 FILLCELL_X4 FILLER_88_247 ();
 FILLCELL_X8 FILLER_88_253 ();
 FILLCELL_X2 FILLER_88_261 ();
 FILLCELL_X1 FILLER_88_263 ();
 FILLCELL_X4 FILLER_88_266 ();
 FILLCELL_X16 FILLER_88_274 ();
 FILLCELL_X4 FILLER_88_293 ();
 FILLCELL_X8 FILLER_88_301 ();
 FILLCELL_X1 FILLER_88_309 ();
 FILLCELL_X4 FILLER_88_317 ();
 FILLCELL_X2 FILLER_88_321 ();
 FILLCELL_X1 FILLER_88_323 ();
 FILLCELL_X4 FILLER_88_327 ();
 FILLCELL_X4 FILLER_88_333 ();
 FILLCELL_X4 FILLER_88_347 ();
 FILLCELL_X1 FILLER_88_351 ();
 FILLCELL_X4 FILLER_88_355 ();
 FILLCELL_X4 FILLER_88_363 ();
 FILLCELL_X8 FILLER_88_370 ();
 FILLCELL_X2 FILLER_88_378 ();
 FILLCELL_X32 FILLER_88_1518 ();
 FILLCELL_X32 FILLER_88_1550 ();
 FILLCELL_X32 FILLER_88_1582 ();
 FILLCELL_X32 FILLER_88_1614 ();
 FILLCELL_X32 FILLER_88_1646 ();
 FILLCELL_X32 FILLER_88_1678 ();
 FILLCELL_X32 FILLER_88_1710 ();
 FILLCELL_X8 FILLER_88_1742 ();
 FILLCELL_X4 FILLER_88_1750 ();
 FILLCELL_X1 FILLER_88_1754 ();
 FILLCELL_X4 FILLER_88_1758 ();
 FILLCELL_X4 FILLER_89_1 ();
 FILLCELL_X2 FILLER_89_5 ();
 FILLCELL_X4 FILLER_89_16 ();
 FILLCELL_X1 FILLER_89_20 ();
 FILLCELL_X4 FILLER_89_24 ();
 FILLCELL_X4 FILLER_89_37 ();
 FILLCELL_X4 FILLER_89_51 ();
 FILLCELL_X4 FILLER_89_65 ();
 FILLCELL_X8 FILLER_89_78 ();
 FILLCELL_X4 FILLER_89_96 ();
 FILLCELL_X2 FILLER_89_100 ();
 FILLCELL_X1 FILLER_89_102 ();
 FILLCELL_X4 FILLER_89_105 ();
 FILLCELL_X4 FILLER_89_119 ();
 FILLCELL_X4 FILLER_89_133 ();
 FILLCELL_X4 FILLER_89_141 ();
 FILLCELL_X2 FILLER_89_145 ();
 FILLCELL_X1 FILLER_89_147 ();
 FILLCELL_X4 FILLER_89_150 ();
 FILLCELL_X4 FILLER_89_164 ();
 FILLCELL_X4 FILLER_89_171 ();
 FILLCELL_X8 FILLER_89_184 ();
 FILLCELL_X4 FILLER_89_192 ();
 FILLCELL_X2 FILLER_89_196 ();
 FILLCELL_X1 FILLER_89_198 ();
 FILLCELL_X4 FILLER_89_202 ();
 FILLCELL_X4 FILLER_89_216 ();
 FILLCELL_X1 FILLER_89_220 ();
 FILLCELL_X4 FILLER_89_223 ();
 FILLCELL_X4 FILLER_89_234 ();
 FILLCELL_X4 FILLER_89_248 ();
 FILLCELL_X8 FILLER_89_255 ();
 FILLCELL_X2 FILLER_89_263 ();
 FILLCELL_X4 FILLER_89_268 ();
 FILLCELL_X16 FILLER_89_279 ();
 FILLCELL_X4 FILLER_89_295 ();
 FILLCELL_X1 FILLER_89_299 ();
 FILLCELL_X4 FILLER_89_309 ();
 FILLCELL_X8 FILLER_89_316 ();
 FILLCELL_X2 FILLER_89_324 ();
 FILLCELL_X4 FILLER_89_330 ();
 FILLCELL_X32 FILLER_89_341 ();
 FILLCELL_X4 FILLER_89_373 ();
 FILLCELL_X2 FILLER_89_377 ();
 FILLCELL_X1 FILLER_89_379 ();
 FILLCELL_X32 FILLER_89_1518 ();
 FILLCELL_X32 FILLER_89_1550 ();
 FILLCELL_X32 FILLER_89_1582 ();
 FILLCELL_X32 FILLER_89_1614 ();
 FILLCELL_X32 FILLER_89_1646 ();
 FILLCELL_X32 FILLER_89_1678 ();
 FILLCELL_X32 FILLER_89_1710 ();
 FILLCELL_X16 FILLER_89_1742 ();
 FILLCELL_X4 FILLER_89_1758 ();
 FILLCELL_X8 FILLER_90_1 ();
 FILLCELL_X4 FILLER_90_9 ();
 FILLCELL_X2 FILLER_90_13 ();
 FILLCELL_X8 FILLER_90_25 ();
 FILLCELL_X2 FILLER_90_33 ();
 FILLCELL_X4 FILLER_90_38 ();
 FILLCELL_X8 FILLER_90_49 ();
 FILLCELL_X4 FILLER_90_57 ();
 FILLCELL_X2 FILLER_90_61 ();
 FILLCELL_X1 FILLER_90_63 ();
 FILLCELL_X4 FILLER_90_67 ();
 FILLCELL_X4 FILLER_90_80 ();
 FILLCELL_X4 FILLER_90_86 ();
 FILLCELL_X4 FILLER_90_100 ();
 FILLCELL_X16 FILLER_90_106 ();
 FILLCELL_X8 FILLER_90_122 ();
 FILLCELL_X4 FILLER_90_130 ();
 FILLCELL_X8 FILLER_90_136 ();
 FILLCELL_X1 FILLER_90_144 ();
 FILLCELL_X4 FILLER_90_155 ();
 FILLCELL_X4 FILLER_90_166 ();
 FILLCELL_X2 FILLER_90_170 ();
 FILLCELL_X4 FILLER_90_176 ();
 FILLCELL_X2 FILLER_90_180 ();
 FILLCELL_X1 FILLER_90_182 ();
 FILLCELL_X4 FILLER_90_187 ();
 FILLCELL_X4 FILLER_90_195 ();
 FILLCELL_X4 FILLER_90_206 ();
 FILLCELL_X8 FILLER_90_220 ();
 FILLCELL_X4 FILLER_90_232 ();
 FILLCELL_X4 FILLER_90_245 ();
 FILLCELL_X4 FILLER_90_258 ();
 FILLCELL_X4 FILLER_90_272 ();
 FILLCELL_X4 FILLER_90_286 ();
 FILLCELL_X4 FILLER_90_294 ();
 FILLCELL_X4 FILLER_90_307 ();
 FILLCELL_X4 FILLER_90_315 ();
 FILLCELL_X8 FILLER_90_324 ();
 FILLCELL_X2 FILLER_90_332 ();
 FILLCELL_X8 FILLER_90_344 ();
 FILLCELL_X1 FILLER_90_352 ();
 FILLCELL_X4 FILLER_90_359 ();
 FILLCELL_X4 FILLER_90_373 ();
 FILLCELL_X2 FILLER_90_377 ();
 FILLCELL_X1 FILLER_90_379 ();
 FILLCELL_X4 FILLER_90_1518 ();
 FILLCELL_X2 FILLER_90_1522 ();
 FILLCELL_X1 FILLER_90_1524 ();
 FILLCELL_X32 FILLER_90_1529 ();
 FILLCELL_X32 FILLER_90_1561 ();
 FILLCELL_X32 FILLER_90_1593 ();
 FILLCELL_X32 FILLER_90_1625 ();
 FILLCELL_X32 FILLER_90_1657 ();
 FILLCELL_X32 FILLER_90_1689 ();
 FILLCELL_X32 FILLER_90_1721 ();
 FILLCELL_X8 FILLER_90_1753 ();
 FILLCELL_X1 FILLER_90_1761 ();
 FILLCELL_X8 FILLER_91_1 ();
 FILLCELL_X1 FILLER_91_9 ();
 FILLCELL_X4 FILLER_91_12 ();
 FILLCELL_X4 FILLER_91_20 ();
 FILLCELL_X4 FILLER_91_34 ();
 FILLCELL_X4 FILLER_91_41 ();
 FILLCELL_X1 FILLER_91_45 ();
 FILLCELL_X16 FILLER_91_55 ();
 FILLCELL_X8 FILLER_91_71 ();
 FILLCELL_X4 FILLER_91_79 ();
 FILLCELL_X1 FILLER_91_83 ();
 FILLCELL_X8 FILLER_91_91 ();
 FILLCELL_X1 FILLER_91_99 ();
 FILLCELL_X4 FILLER_91_103 ();
 FILLCELL_X2 FILLER_91_107 ();
 FILLCELL_X4 FILLER_91_119 ();
 FILLCELL_X1 FILLER_91_123 ();
 FILLCELL_X4 FILLER_91_131 ();
 FILLCELL_X8 FILLER_91_145 ();
 FILLCELL_X4 FILLER_91_153 ();
 FILLCELL_X2 FILLER_91_157 ();
 FILLCELL_X1 FILLER_91_159 ();
 FILLCELL_X4 FILLER_91_163 ();
 FILLCELL_X4 FILLER_91_176 ();
 FILLCELL_X2 FILLER_91_180 ();
 FILLCELL_X4 FILLER_91_185 ();
 FILLCELL_X8 FILLER_91_198 ();
 FILLCELL_X4 FILLER_91_206 ();
 FILLCELL_X1 FILLER_91_210 ();
 FILLCELL_X8 FILLER_91_213 ();
 FILLCELL_X2 FILLER_91_221 ();
 FILLCELL_X1 FILLER_91_223 ();
 FILLCELL_X4 FILLER_91_228 ();
 FILLCELL_X4 FILLER_91_241 ();
 FILLCELL_X2 FILLER_91_245 ();
 FILLCELL_X1 FILLER_91_247 ();
 FILLCELL_X16 FILLER_91_251 ();
 FILLCELL_X4 FILLER_91_267 ();
 FILLCELL_X2 FILLER_91_271 ();
 FILLCELL_X8 FILLER_91_275 ();
 FILLCELL_X4 FILLER_91_283 ();
 FILLCELL_X2 FILLER_91_287 ();
 FILLCELL_X4 FILLER_91_292 ();
 FILLCELL_X8 FILLER_91_300 ();
 FILLCELL_X4 FILLER_91_311 ();
 FILLCELL_X4 FILLER_91_334 ();
 FILLCELL_X4 FILLER_91_341 ();
 FILLCELL_X1 FILLER_91_345 ();
 FILLCELL_X4 FILLER_91_348 ();
 FILLCELL_X4 FILLER_91_356 ();
 FILLCELL_X8 FILLER_91_367 ();
 FILLCELL_X4 FILLER_91_375 ();
 FILLCELL_X1 FILLER_91_379 ();
 FILLCELL_X4 FILLER_91_1518 ();
 FILLCELL_X2 FILLER_91_1522 ();
 FILLCELL_X1 FILLER_91_1524 ();
 FILLCELL_X32 FILLER_91_1544 ();
 FILLCELL_X32 FILLER_91_1576 ();
 FILLCELL_X32 FILLER_91_1608 ();
 FILLCELL_X32 FILLER_91_1640 ();
 FILLCELL_X32 FILLER_91_1672 ();
 FILLCELL_X32 FILLER_91_1704 ();
 FILLCELL_X16 FILLER_91_1736 ();
 FILLCELL_X8 FILLER_91_1752 ();
 FILLCELL_X2 FILLER_91_1760 ();
 FILLCELL_X4 FILLER_92_1 ();
 FILLCELL_X2 FILLER_92_5 ();
 FILLCELL_X1 FILLER_92_7 ();
 FILLCELL_X4 FILLER_92_18 ();
 FILLCELL_X16 FILLER_92_25 ();
 FILLCELL_X1 FILLER_92_41 ();
 FILLCELL_X4 FILLER_92_52 ();
 FILLCELL_X8 FILLER_92_58 ();
 FILLCELL_X1 FILLER_92_66 ();
 FILLCELL_X4 FILLER_92_70 ();
 FILLCELL_X4 FILLER_92_84 ();
 FILLCELL_X4 FILLER_92_90 ();
 FILLCELL_X4 FILLER_92_103 ();
 FILLCELL_X16 FILLER_92_116 ();
 FILLCELL_X4 FILLER_92_132 ();
 FILLCELL_X2 FILLER_92_136 ();
 FILLCELL_X1 FILLER_92_138 ();
 FILLCELL_X16 FILLER_92_143 ();
 FILLCELL_X4 FILLER_92_161 ();
 FILLCELL_X4 FILLER_92_169 ();
 FILLCELL_X2 FILLER_92_173 ();
 FILLCELL_X4 FILLER_92_178 ();
 FILLCELL_X2 FILLER_92_182 ();
 FILLCELL_X8 FILLER_92_188 ();
 FILLCELL_X2 FILLER_92_196 ();
 FILLCELL_X4 FILLER_92_202 ();
 FILLCELL_X8 FILLER_92_209 ();
 FILLCELL_X1 FILLER_92_217 ();
 FILLCELL_X8 FILLER_92_221 ();
 FILLCELL_X2 FILLER_92_229 ();
 FILLCELL_X8 FILLER_92_235 ();
 FILLCELL_X4 FILLER_92_246 ();
 FILLCELL_X2 FILLER_92_250 ();
 FILLCELL_X1 FILLER_92_252 ();
 FILLCELL_X8 FILLER_92_257 ();
 FILLCELL_X4 FILLER_92_265 ();
 FILLCELL_X4 FILLER_92_273 ();
 FILLCELL_X2 FILLER_92_277 ();
 FILLCELL_X8 FILLER_92_283 ();
 FILLCELL_X4 FILLER_92_291 ();
 FILLCELL_X2 FILLER_92_295 ();
 FILLCELL_X8 FILLER_92_301 ();
 FILLCELL_X1 FILLER_92_309 ();
 FILLCELL_X16 FILLER_92_313 ();
 FILLCELL_X8 FILLER_92_329 ();
 FILLCELL_X4 FILLER_92_343 ();
 FILLCELL_X4 FILLER_92_354 ();
 FILLCELL_X16 FILLER_92_362 ();
 FILLCELL_X2 FILLER_92_378 ();
 FILLCELL_X32 FILLER_92_1518 ();
 FILLCELL_X32 FILLER_92_1550 ();
 FILLCELL_X32 FILLER_92_1582 ();
 FILLCELL_X32 FILLER_92_1614 ();
 FILLCELL_X32 FILLER_92_1646 ();
 FILLCELL_X32 FILLER_92_1678 ();
 FILLCELL_X32 FILLER_92_1710 ();
 FILLCELL_X16 FILLER_92_1742 ();
 FILLCELL_X4 FILLER_92_1758 ();
 FILLCELL_X4 FILLER_93_1 ();
 FILLCELL_X4 FILLER_93_8 ();
 FILLCELL_X4 FILLER_93_16 ();
 FILLCELL_X4 FILLER_93_22 ();
 FILLCELL_X2 FILLER_93_26 ();
 FILLCELL_X1 FILLER_93_28 ();
 FILLCELL_X4 FILLER_93_32 ();
 FILLCELL_X4 FILLER_93_45 ();
 FILLCELL_X1 FILLER_93_49 ();
 FILLCELL_X4 FILLER_93_53 ();
 FILLCELL_X4 FILLER_93_67 ();
 FILLCELL_X2 FILLER_93_71 ();
 FILLCELL_X8 FILLER_93_80 ();
 FILLCELL_X4 FILLER_93_91 ();
 FILLCELL_X8 FILLER_93_105 ();
 FILLCELL_X4 FILLER_93_116 ();
 FILLCELL_X4 FILLER_93_123 ();
 FILLCELL_X8 FILLER_93_136 ();
 FILLCELL_X1 FILLER_93_144 ();
 FILLCELL_X4 FILLER_93_149 ();
 FILLCELL_X4 FILLER_93_157 ();
 FILLCELL_X2 FILLER_93_161 ();
 FILLCELL_X4 FILLER_93_173 ();
 FILLCELL_X2 FILLER_93_177 ();
 FILLCELL_X1 FILLER_93_179 ();
 FILLCELL_X4 FILLER_93_183 ();
 FILLCELL_X8 FILLER_93_196 ();
 FILLCELL_X4 FILLER_93_213 ();
 FILLCELL_X4 FILLER_93_226 ();
 FILLCELL_X1 FILLER_93_230 ();
 FILLCELL_X8 FILLER_93_238 ();
 FILLCELL_X4 FILLER_93_246 ();
 FILLCELL_X8 FILLER_93_267 ();
 FILLCELL_X4 FILLER_93_279 ();
 FILLCELL_X1 FILLER_93_283 ();
 FILLCELL_X4 FILLER_93_293 ();
 FILLCELL_X1 FILLER_93_297 ();
 FILLCELL_X4 FILLER_93_308 ();
 FILLCELL_X2 FILLER_93_312 ();
 FILLCELL_X1 FILLER_93_314 ();
 FILLCELL_X4 FILLER_93_319 ();
 FILLCELL_X4 FILLER_93_332 ();
 FILLCELL_X4 FILLER_93_346 ();
 FILLCELL_X4 FILLER_93_375 ();
 FILLCELL_X1 FILLER_93_379 ();
 FILLCELL_X32 FILLER_93_1518 ();
 FILLCELL_X32 FILLER_93_1550 ();
 FILLCELL_X32 FILLER_93_1582 ();
 FILLCELL_X32 FILLER_93_1614 ();
 FILLCELL_X32 FILLER_93_1646 ();
 FILLCELL_X32 FILLER_93_1678 ();
 FILLCELL_X32 FILLER_93_1710 ();
 FILLCELL_X16 FILLER_93_1742 ();
 FILLCELL_X4 FILLER_93_1758 ();
 FILLCELL_X4 FILLER_94_1 ();
 FILLCELL_X1 FILLER_94_5 ();
 FILLCELL_X4 FILLER_94_10 ();
 FILLCELL_X2 FILLER_94_14 ();
 FILLCELL_X8 FILLER_94_26 ();
 FILLCELL_X2 FILLER_94_34 ();
 FILLCELL_X4 FILLER_94_39 ();
 FILLCELL_X8 FILLER_94_46 ();
 FILLCELL_X4 FILLER_94_57 ();
 FILLCELL_X1 FILLER_94_61 ();
 FILLCELL_X8 FILLER_94_65 ();
 FILLCELL_X2 FILLER_94_73 ();
 FILLCELL_X4 FILLER_94_85 ();
 FILLCELL_X2 FILLER_94_89 ();
 FILLCELL_X1 FILLER_94_91 ();
 FILLCELL_X4 FILLER_94_99 ();
 FILLCELL_X4 FILLER_94_106 ();
 FILLCELL_X4 FILLER_94_113 ();
 FILLCELL_X4 FILLER_94_120 ();
 FILLCELL_X8 FILLER_94_133 ();
 FILLCELL_X1 FILLER_94_141 ();
 FILLCELL_X8 FILLER_94_151 ();
 FILLCELL_X1 FILLER_94_159 ();
 FILLCELL_X8 FILLER_94_170 ();
 FILLCELL_X1 FILLER_94_178 ();
 FILLCELL_X4 FILLER_94_181 ();
 FILLCELL_X4 FILLER_94_188 ();
 FILLCELL_X4 FILLER_94_202 ();
 FILLCELL_X4 FILLER_94_216 ();
 FILLCELL_X2 FILLER_94_220 ();
 FILLCELL_X1 FILLER_94_222 ();
 FILLCELL_X4 FILLER_94_233 ();
 FILLCELL_X16 FILLER_94_247 ();
 FILLCELL_X4 FILLER_94_263 ();
 FILLCELL_X2 FILLER_94_267 ();
 FILLCELL_X4 FILLER_94_273 ();
 FILLCELL_X8 FILLER_94_286 ();
 FILLCELL_X4 FILLER_94_301 ();
 FILLCELL_X8 FILLER_94_315 ();
 FILLCELL_X4 FILLER_94_323 ();
 FILLCELL_X4 FILLER_94_331 ();
 FILLCELL_X4 FILLER_94_338 ();
 FILLCELL_X1 FILLER_94_342 ();
 FILLCELL_X32 FILLER_94_346 ();
 FILLCELL_X2 FILLER_94_378 ();
 FILLCELL_X4 FILLER_94_1518 ();
 FILLCELL_X32 FILLER_94_1526 ();
 FILLCELL_X32 FILLER_94_1558 ();
 FILLCELL_X32 FILLER_94_1590 ();
 FILLCELL_X32 FILLER_94_1622 ();
 FILLCELL_X32 FILLER_94_1654 ();
 FILLCELL_X32 FILLER_94_1686 ();
 FILLCELL_X32 FILLER_94_1718 ();
 FILLCELL_X8 FILLER_94_1750 ();
 FILLCELL_X4 FILLER_94_1758 ();
 FILLCELL_X8 FILLER_95_1 ();
 FILLCELL_X1 FILLER_95_9 ();
 FILLCELL_X4 FILLER_95_14 ();
 FILLCELL_X8 FILLER_95_31 ();
 FILLCELL_X2 FILLER_95_39 ();
 FILLCELL_X4 FILLER_95_45 ();
 FILLCELL_X4 FILLER_95_52 ();
 FILLCELL_X1 FILLER_95_56 ();
 FILLCELL_X4 FILLER_95_60 ();
 FILLCELL_X2 FILLER_95_64 ();
 FILLCELL_X4 FILLER_95_75 ();
 FILLCELL_X4 FILLER_95_82 ();
 FILLCELL_X4 FILLER_95_88 ();
 FILLCELL_X32 FILLER_95_102 ();
 FILLCELL_X8 FILLER_95_134 ();
 FILLCELL_X4 FILLER_95_142 ();
 FILLCELL_X4 FILLER_95_155 ();
 FILLCELL_X1 FILLER_95_159 ();
 FILLCELL_X4 FILLER_95_167 ();
 FILLCELL_X16 FILLER_95_173 ();
 FILLCELL_X4 FILLER_95_189 ();
 FILLCELL_X1 FILLER_95_193 ();
 FILLCELL_X8 FILLER_95_201 ();
 FILLCELL_X2 FILLER_95_209 ();
 FILLCELL_X4 FILLER_95_214 ();
 FILLCELL_X8 FILLER_95_221 ();
 FILLCELL_X1 FILLER_95_229 ();
 FILLCELL_X4 FILLER_95_233 ();
 FILLCELL_X4 FILLER_95_239 ();
 FILLCELL_X2 FILLER_95_243 ();
 FILLCELL_X8 FILLER_95_249 ();
 FILLCELL_X4 FILLER_95_257 ();
 FILLCELL_X1 FILLER_95_261 ();
 FILLCELL_X8 FILLER_95_265 ();
 FILLCELL_X1 FILLER_95_273 ();
 FILLCELL_X4 FILLER_95_277 ();
 FILLCELL_X4 FILLER_95_284 ();
 FILLCELL_X8 FILLER_95_291 ();
 FILLCELL_X2 FILLER_95_299 ();
 FILLCELL_X1 FILLER_95_301 ();
 FILLCELL_X8 FILLER_95_304 ();
 FILLCELL_X4 FILLER_95_315 ();
 FILLCELL_X4 FILLER_95_323 ();
 FILLCELL_X8 FILLER_95_336 ();
 FILLCELL_X4 FILLER_95_344 ();
 FILLCELL_X2 FILLER_95_348 ();
 FILLCELL_X1 FILLER_95_350 ();
 FILLCELL_X16 FILLER_95_358 ();
 FILLCELL_X4 FILLER_95_374 ();
 FILLCELL_X2 FILLER_95_378 ();
 FILLCELL_X8 FILLER_95_1518 ();
 FILLCELL_X32 FILLER_95_1545 ();
 FILLCELL_X32 FILLER_95_1577 ();
 FILLCELL_X32 FILLER_95_1609 ();
 FILLCELL_X32 FILLER_95_1641 ();
 FILLCELL_X32 FILLER_95_1673 ();
 FILLCELL_X32 FILLER_95_1705 ();
 FILLCELL_X16 FILLER_95_1737 ();
 FILLCELL_X8 FILLER_95_1753 ();
 FILLCELL_X1 FILLER_95_1761 ();
 FILLCELL_X4 FILLER_96_1 ();
 FILLCELL_X2 FILLER_96_5 ();
 FILLCELL_X4 FILLER_96_13 ();
 FILLCELL_X8 FILLER_96_20 ();
 FILLCELL_X2 FILLER_96_28 ();
 FILLCELL_X1 FILLER_96_30 ();
 FILLCELL_X4 FILLER_96_40 ();
 FILLCELL_X4 FILLER_96_54 ();
 FILLCELL_X8 FILLER_96_67 ();
 FILLCELL_X1 FILLER_96_75 ();
 FILLCELL_X8 FILLER_96_86 ();
 FILLCELL_X2 FILLER_96_94 ();
 FILLCELL_X1 FILLER_96_96 ();
 FILLCELL_X4 FILLER_96_100 ();
 FILLCELL_X8 FILLER_96_114 ();
 FILLCELL_X4 FILLER_96_122 ();
 FILLCELL_X4 FILLER_96_129 ();
 FILLCELL_X4 FILLER_96_136 ();
 FILLCELL_X4 FILLER_96_143 ();
 FILLCELL_X8 FILLER_96_156 ();
 FILLCELL_X1 FILLER_96_164 ();
 FILLCELL_X8 FILLER_96_172 ();
 FILLCELL_X4 FILLER_96_180 ();
 FILLCELL_X4 FILLER_96_187 ();
 FILLCELL_X4 FILLER_96_200 ();
 FILLCELL_X32 FILLER_96_207 ();
 FILLCELL_X1 FILLER_96_239 ();
 FILLCELL_X4 FILLER_96_244 ();
 FILLCELL_X4 FILLER_96_257 ();
 FILLCELL_X4 FILLER_96_271 ();
 FILLCELL_X8 FILLER_96_277 ();
 FILLCELL_X4 FILLER_96_285 ();
 FILLCELL_X4 FILLER_96_293 ();
 FILLCELL_X1 FILLER_96_297 ();
 FILLCELL_X4 FILLER_96_305 ();
 FILLCELL_X8 FILLER_96_311 ();
 FILLCELL_X4 FILLER_96_328 ();
 FILLCELL_X4 FILLER_96_335 ();
 FILLCELL_X1 FILLER_96_339 ();
 FILLCELL_X4 FILLER_96_343 ();
 FILLCELL_X4 FILLER_96_356 ();
 FILLCELL_X8 FILLER_96_370 ();
 FILLCELL_X2 FILLER_96_378 ();
 FILLCELL_X32 FILLER_96_1518 ();
 FILLCELL_X32 FILLER_96_1550 ();
 FILLCELL_X32 FILLER_96_1582 ();
 FILLCELL_X32 FILLER_96_1614 ();
 FILLCELL_X32 FILLER_96_1646 ();
 FILLCELL_X32 FILLER_96_1678 ();
 FILLCELL_X32 FILLER_96_1710 ();
 FILLCELL_X16 FILLER_96_1742 ();
 FILLCELL_X4 FILLER_96_1758 ();
 FILLCELL_X4 FILLER_97_1 ();
 FILLCELL_X2 FILLER_97_5 ();
 FILLCELL_X8 FILLER_97_13 ();
 FILLCELL_X2 FILLER_97_21 ();
 FILLCELL_X16 FILLER_97_26 ();
 FILLCELL_X8 FILLER_97_42 ();
 FILLCELL_X16 FILLER_97_57 ();
 FILLCELL_X1 FILLER_97_73 ();
 FILLCELL_X16 FILLER_97_81 ();
 FILLCELL_X4 FILLER_97_97 ();
 FILLCELL_X2 FILLER_97_101 ();
 FILLCELL_X4 FILLER_97_110 ();
 FILLCELL_X4 FILLER_97_124 ();
 FILLCELL_X4 FILLER_97_138 ();
 FILLCELL_X2 FILLER_97_142 ();
 FILLCELL_X4 FILLER_97_147 ();
 FILLCELL_X4 FILLER_97_154 ();
 FILLCELL_X4 FILLER_97_168 ();
 FILLCELL_X4 FILLER_97_182 ();
 FILLCELL_X4 FILLER_97_195 ();
 FILLCELL_X8 FILLER_97_203 ();
 FILLCELL_X4 FILLER_97_214 ();
 FILLCELL_X4 FILLER_97_227 ();
 FILLCELL_X2 FILLER_97_231 ();
 FILLCELL_X4 FILLER_97_237 ();
 FILLCELL_X4 FILLER_97_250 ();
 FILLCELL_X2 FILLER_97_254 ();
 FILLCELL_X1 FILLER_97_256 ();
 FILLCELL_X4 FILLER_97_264 ();
 FILLCELL_X4 FILLER_97_278 ();
 FILLCELL_X2 FILLER_97_282 ();
 FILLCELL_X4 FILLER_97_287 ();
 FILLCELL_X4 FILLER_97_301 ();
 FILLCELL_X2 FILLER_97_305 ();
 FILLCELL_X1 FILLER_97_307 ();
 FILLCELL_X4 FILLER_97_318 ();
 FILLCELL_X4 FILLER_97_325 ();
 FILLCELL_X8 FILLER_97_338 ();
 FILLCELL_X4 FILLER_97_346 ();
 FILLCELL_X2 FILLER_97_350 ();
 FILLCELL_X16 FILLER_97_355 ();
 FILLCELL_X8 FILLER_97_371 ();
 FILLCELL_X1 FILLER_97_379 ();
 FILLCELL_X32 FILLER_97_1518 ();
 FILLCELL_X32 FILLER_97_1550 ();
 FILLCELL_X32 FILLER_97_1582 ();
 FILLCELL_X32 FILLER_97_1614 ();
 FILLCELL_X32 FILLER_97_1646 ();
 FILLCELL_X32 FILLER_97_1678 ();
 FILLCELL_X32 FILLER_97_1710 ();
 FILLCELL_X16 FILLER_97_1742 ();
 FILLCELL_X4 FILLER_97_1758 ();
 FILLCELL_X4 FILLER_98_1 ();
 FILLCELL_X2 FILLER_98_5 ();
 FILLCELL_X1 FILLER_98_7 ();
 FILLCELL_X4 FILLER_98_12 ();
 FILLCELL_X2 FILLER_98_16 ();
 FILLCELL_X4 FILLER_98_22 ();
 FILLCELL_X2 FILLER_98_26 ();
 FILLCELL_X8 FILLER_98_32 ();
 FILLCELL_X2 FILLER_98_40 ();
 FILLCELL_X1 FILLER_98_42 ();
 FILLCELL_X4 FILLER_98_47 ();
 FILLCELL_X8 FILLER_98_53 ();
 FILLCELL_X1 FILLER_98_61 ();
 FILLCELL_X4 FILLER_98_64 ();
 FILLCELL_X4 FILLER_98_75 ();
 FILLCELL_X16 FILLER_98_82 ();
 FILLCELL_X2 FILLER_98_98 ();
 FILLCELL_X8 FILLER_98_104 ();
 FILLCELL_X1 FILLER_98_112 ();
 FILLCELL_X4 FILLER_98_115 ();
 FILLCELL_X2 FILLER_98_119 ();
 FILLCELL_X1 FILLER_98_121 ();
 FILLCELL_X4 FILLER_98_124 ();
 FILLCELL_X16 FILLER_98_138 ();
 FILLCELL_X8 FILLER_98_154 ();
 FILLCELL_X2 FILLER_98_162 ();
 FILLCELL_X1 FILLER_98_164 ();
 FILLCELL_X4 FILLER_98_168 ();
 FILLCELL_X8 FILLER_98_174 ();
 FILLCELL_X4 FILLER_98_182 ();
 FILLCELL_X2 FILLER_98_186 ();
 FILLCELL_X1 FILLER_98_188 ();
 FILLCELL_X8 FILLER_98_192 ();
 FILLCELL_X4 FILLER_98_200 ();
 FILLCELL_X4 FILLER_98_207 ();
 FILLCELL_X4 FILLER_98_215 ();
 FILLCELL_X4 FILLER_98_228 ();
 FILLCELL_X2 FILLER_98_232 ();
 FILLCELL_X1 FILLER_98_234 ();
 FILLCELL_X4 FILLER_98_238 ();
 FILLCELL_X4 FILLER_98_245 ();
 FILLCELL_X2 FILLER_98_249 ();
 FILLCELL_X1 FILLER_98_251 ();
 FILLCELL_X16 FILLER_98_255 ();
 FILLCELL_X4 FILLER_98_275 ();
 FILLCELL_X8 FILLER_98_288 ();
 FILLCELL_X2 FILLER_98_296 ();
 FILLCELL_X16 FILLER_98_307 ();
 FILLCELL_X4 FILLER_98_323 ();
 FILLCELL_X2 FILLER_98_327 ();
 FILLCELL_X8 FILLER_98_332 ();
 FILLCELL_X4 FILLER_98_340 ();
 FILLCELL_X1 FILLER_98_344 ();
 FILLCELL_X4 FILLER_98_355 ();
 FILLCELL_X16 FILLER_98_361 ();
 FILLCELL_X2 FILLER_98_377 ();
 FILLCELL_X1 FILLER_98_379 ();
 FILLCELL_X32 FILLER_98_1518 ();
 FILLCELL_X32 FILLER_98_1550 ();
 FILLCELL_X32 FILLER_98_1582 ();
 FILLCELL_X32 FILLER_98_1614 ();
 FILLCELL_X32 FILLER_98_1646 ();
 FILLCELL_X32 FILLER_98_1678 ();
 FILLCELL_X32 FILLER_98_1710 ();
 FILLCELL_X8 FILLER_98_1742 ();
 FILLCELL_X4 FILLER_98_1750 ();
 FILLCELL_X1 FILLER_98_1754 ();
 FILLCELL_X4 FILLER_98_1758 ();
 FILLCELL_X4 FILLER_99_1 ();
 FILLCELL_X1 FILLER_99_5 ();
 FILLCELL_X4 FILLER_99_10 ();
 FILLCELL_X4 FILLER_99_23 ();
 FILLCELL_X4 FILLER_99_36 ();
 FILLCELL_X2 FILLER_99_40 ();
 FILLCELL_X4 FILLER_99_46 ();
 FILLCELL_X1 FILLER_99_50 ();
 FILLCELL_X4 FILLER_99_61 ();
 FILLCELL_X2 FILLER_99_65 ();
 FILLCELL_X8 FILLER_99_77 ();
 FILLCELL_X1 FILLER_99_85 ();
 FILLCELL_X4 FILLER_99_89 ();
 FILLCELL_X4 FILLER_99_96 ();
 FILLCELL_X4 FILLER_99_104 ();
 FILLCELL_X4 FILLER_99_112 ();
 FILLCELL_X8 FILLER_99_119 ();
 FILLCELL_X8 FILLER_99_134 ();
 FILLCELL_X1 FILLER_99_142 ();
 FILLCELL_X4 FILLER_99_147 ();
 FILLCELL_X4 FILLER_99_155 ();
 FILLCELL_X8 FILLER_99_163 ();
 FILLCELL_X1 FILLER_99_171 ();
 FILLCELL_X4 FILLER_99_175 ();
 FILLCELL_X8 FILLER_99_183 ();
 FILLCELL_X4 FILLER_99_191 ();
 FILLCELL_X4 FILLER_99_198 ();
 FILLCELL_X2 FILLER_99_202 ();
 FILLCELL_X8 FILLER_99_206 ();
 FILLCELL_X2 FILLER_99_214 ();
 FILLCELL_X1 FILLER_99_216 ();
 FILLCELL_X16 FILLER_99_220 ();
 FILLCELL_X8 FILLER_99_236 ();
 FILLCELL_X4 FILLER_99_244 ();
 FILLCELL_X8 FILLER_99_251 ();
 FILLCELL_X4 FILLER_99_259 ();
 FILLCELL_X1 FILLER_99_263 ();
 FILLCELL_X8 FILLER_99_267 ();
 FILLCELL_X4 FILLER_99_279 ();
 FILLCELL_X8 FILLER_99_286 ();
 FILLCELL_X4 FILLER_99_297 ();
 FILLCELL_X8 FILLER_99_310 ();
 FILLCELL_X4 FILLER_99_318 ();
 FILLCELL_X2 FILLER_99_322 ();
 FILLCELL_X4 FILLER_99_327 ();
 FILLCELL_X8 FILLER_99_340 ();
 FILLCELL_X4 FILLER_99_348 ();
 FILLCELL_X4 FILLER_99_362 ();
 FILLCELL_X8 FILLER_99_370 ();
 FILLCELL_X2 FILLER_99_378 ();
 FILLCELL_X32 FILLER_99_1518 ();
 FILLCELL_X32 FILLER_99_1550 ();
 FILLCELL_X32 FILLER_99_1582 ();
 FILLCELL_X32 FILLER_99_1614 ();
 FILLCELL_X32 FILLER_99_1646 ();
 FILLCELL_X32 FILLER_99_1678 ();
 FILLCELL_X32 FILLER_99_1710 ();
 FILLCELL_X16 FILLER_99_1742 ();
 FILLCELL_X4 FILLER_99_1758 ();
 FILLCELL_X4 FILLER_100_1 ();
 FILLCELL_X4 FILLER_100_24 ();
 FILLCELL_X4 FILLER_100_31 ();
 FILLCELL_X4 FILLER_100_38 ();
 FILLCELL_X4 FILLER_100_51 ();
 FILLCELL_X4 FILLER_100_58 ();
 FILLCELL_X2 FILLER_100_62 ();
 FILLCELL_X4 FILLER_100_67 ();
 FILLCELL_X8 FILLER_100_81 ();
 FILLCELL_X4 FILLER_100_93 ();
 FILLCELL_X8 FILLER_100_106 ();
 FILLCELL_X2 FILLER_100_114 ();
 FILLCELL_X4 FILLER_100_120 ();
 FILLCELL_X4 FILLER_100_128 ();
 FILLCELL_X2 FILLER_100_132 ();
 FILLCELL_X8 FILLER_100_138 ();
 FILLCELL_X2 FILLER_100_146 ();
 FILLCELL_X4 FILLER_100_157 ();
 FILLCELL_X4 FILLER_100_170 ();
 FILLCELL_X2 FILLER_100_174 ();
 FILLCELL_X4 FILLER_100_186 ();
 FILLCELL_X4 FILLER_100_200 ();
 FILLCELL_X16 FILLER_100_214 ();
 FILLCELL_X2 FILLER_100_230 ();
 FILLCELL_X1 FILLER_100_232 ();
 FILLCELL_X4 FILLER_100_237 ();
 FILLCELL_X4 FILLER_100_245 ();
 FILLCELL_X8 FILLER_100_258 ();
 FILLCELL_X1 FILLER_100_266 ();
 FILLCELL_X4 FILLER_100_271 ();
 FILLCELL_X4 FILLER_100_284 ();
 FILLCELL_X1 FILLER_100_288 ();
 FILLCELL_X4 FILLER_100_292 ();
 FILLCELL_X4 FILLER_100_299 ();
 FILLCELL_X4 FILLER_100_313 ();
 FILLCELL_X8 FILLER_100_319 ();
 FILLCELL_X2 FILLER_100_327 ();
 FILLCELL_X8 FILLER_100_332 ();
 FILLCELL_X2 FILLER_100_340 ();
 FILLCELL_X1 FILLER_100_342 ();
 FILLCELL_X4 FILLER_100_350 ();
 FILLCELL_X16 FILLER_100_357 ();
 FILLCELL_X4 FILLER_100_373 ();
 FILLCELL_X2 FILLER_100_377 ();
 FILLCELL_X1 FILLER_100_379 ();
 FILLCELL_X32 FILLER_100_1518 ();
 FILLCELL_X32 FILLER_100_1550 ();
 FILLCELL_X32 FILLER_100_1582 ();
 FILLCELL_X32 FILLER_100_1614 ();
 FILLCELL_X32 FILLER_100_1646 ();
 FILLCELL_X32 FILLER_100_1678 ();
 FILLCELL_X32 FILLER_100_1710 ();
 FILLCELL_X16 FILLER_100_1742 ();
 FILLCELL_X4 FILLER_100_1758 ();
 FILLCELL_X4 FILLER_101_1 ();
 FILLCELL_X8 FILLER_101_8 ();
 FILLCELL_X4 FILLER_101_16 ();
 FILLCELL_X4 FILLER_101_23 ();
 FILLCELL_X8 FILLER_101_30 ();
 FILLCELL_X1 FILLER_101_38 ();
 FILLCELL_X4 FILLER_101_43 ();
 FILLCELL_X4 FILLER_101_50 ();
 FILLCELL_X2 FILLER_101_54 ();
 FILLCELL_X4 FILLER_101_58 ();
 FILLCELL_X4 FILLER_101_65 ();
 FILLCELL_X16 FILLER_101_78 ();
 FILLCELL_X8 FILLER_101_94 ();
 FILLCELL_X4 FILLER_101_111 ();
 FILLCELL_X2 FILLER_101_115 ();
 FILLCELL_X1 FILLER_101_117 ();
 FILLCELL_X4 FILLER_101_122 ();
 FILLCELL_X1 FILLER_101_126 ();
 FILLCELL_X4 FILLER_101_136 ();
 FILLCELL_X8 FILLER_101_143 ();
 FILLCELL_X2 FILLER_101_151 ();
 FILLCELL_X4 FILLER_101_157 ();
 FILLCELL_X2 FILLER_101_161 ();
 FILLCELL_X1 FILLER_101_163 ();
 FILLCELL_X4 FILLER_101_167 ();
 FILLCELL_X1 FILLER_101_171 ();
 FILLCELL_X4 FILLER_101_174 ();
 FILLCELL_X8 FILLER_101_188 ();
 FILLCELL_X2 FILLER_101_196 ();
 FILLCELL_X4 FILLER_101_205 ();
 FILLCELL_X4 FILLER_101_213 ();
 FILLCELL_X4 FILLER_101_221 ();
 FILLCELL_X8 FILLER_101_234 ();
 FILLCELL_X2 FILLER_101_242 ();
 FILLCELL_X1 FILLER_101_244 ();
 FILLCELL_X4 FILLER_101_248 ();
 FILLCELL_X4 FILLER_101_256 ();
 FILLCELL_X4 FILLER_101_269 ();
 FILLCELL_X2 FILLER_101_273 ();
 FILLCELL_X8 FILLER_101_278 ();
 FILLCELL_X2 FILLER_101_286 ();
 FILLCELL_X16 FILLER_101_291 ();
 FILLCELL_X4 FILLER_101_314 ();
 FILLCELL_X4 FILLER_101_328 ();
 FILLCELL_X8 FILLER_101_341 ();
 FILLCELL_X4 FILLER_101_349 ();
 FILLCELL_X4 FILLER_101_362 ();
 FILLCELL_X8 FILLER_101_370 ();
 FILLCELL_X2 FILLER_101_378 ();
 FILLCELL_X32 FILLER_101_1518 ();
 FILLCELL_X32 FILLER_101_1550 ();
 FILLCELL_X32 FILLER_101_1582 ();
 FILLCELL_X32 FILLER_101_1614 ();
 FILLCELL_X32 FILLER_101_1646 ();
 FILLCELL_X32 FILLER_101_1678 ();
 FILLCELL_X32 FILLER_101_1710 ();
 FILLCELL_X16 FILLER_101_1742 ();
 FILLCELL_X4 FILLER_101_1758 ();
 FILLCELL_X8 FILLER_102_1 ();
 FILLCELL_X1 FILLER_102_9 ();
 FILLCELL_X4 FILLER_102_14 ();
 FILLCELL_X1 FILLER_102_18 ();
 FILLCELL_X4 FILLER_102_26 ();
 FILLCELL_X8 FILLER_102_36 ();
 FILLCELL_X1 FILLER_102_44 ();
 FILLCELL_X4 FILLER_102_54 ();
 FILLCELL_X8 FILLER_102_62 ();
 FILLCELL_X1 FILLER_102_70 ();
 FILLCELL_X4 FILLER_102_74 ();
 FILLCELL_X16 FILLER_102_87 ();
 FILLCELL_X1 FILLER_102_103 ();
 FILLCELL_X4 FILLER_102_107 ();
 FILLCELL_X1 FILLER_102_111 ();
 FILLCELL_X4 FILLER_102_117 ();
 FILLCELL_X4 FILLER_102_124 ();
 FILLCELL_X4 FILLER_102_131 ();
 FILLCELL_X8 FILLER_102_144 ();
 FILLCELL_X4 FILLER_102_152 ();
 FILLCELL_X2 FILLER_102_156 ();
 FILLCELL_X1 FILLER_102_158 ();
 FILLCELL_X8 FILLER_102_162 ();
 FILLCELL_X4 FILLER_102_170 ();
 FILLCELL_X2 FILLER_102_174 ();
 FILLCELL_X1 FILLER_102_176 ();
 FILLCELL_X4 FILLER_102_184 ();
 FILLCELL_X2 FILLER_102_188 ();
 FILLCELL_X8 FILLER_102_194 ();
 FILLCELL_X4 FILLER_102_202 ();
 FILLCELL_X1 FILLER_102_206 ();
 FILLCELL_X4 FILLER_102_211 ();
 FILLCELL_X8 FILLER_102_224 ();
 FILLCELL_X2 FILLER_102_232 ();
 FILLCELL_X4 FILLER_102_237 ();
 FILLCELL_X4 FILLER_102_251 ();
 FILLCELL_X4 FILLER_102_258 ();
 FILLCELL_X16 FILLER_102_264 ();
 FILLCELL_X4 FILLER_102_280 ();
 FILLCELL_X1 FILLER_102_284 ();
 FILLCELL_X16 FILLER_102_289 ();
 FILLCELL_X8 FILLER_102_305 ();
 FILLCELL_X4 FILLER_102_313 ();
 FILLCELL_X2 FILLER_102_317 ();
 FILLCELL_X4 FILLER_102_321 ();
 FILLCELL_X4 FILLER_102_328 ();
 FILLCELL_X4 FILLER_102_335 ();
 FILLCELL_X4 FILLER_102_342 ();
 FILLCELL_X4 FILLER_102_350 ();
 FILLCELL_X4 FILLER_102_363 ();
 FILLCELL_X8 FILLER_102_370 ();
 FILLCELL_X2 FILLER_102_378 ();
 FILLCELL_X32 FILLER_102_1518 ();
 FILLCELL_X32 FILLER_102_1550 ();
 FILLCELL_X32 FILLER_102_1582 ();
 FILLCELL_X32 FILLER_102_1614 ();
 FILLCELL_X32 FILLER_102_1646 ();
 FILLCELL_X32 FILLER_102_1678 ();
 FILLCELL_X32 FILLER_102_1710 ();
 FILLCELL_X16 FILLER_102_1742 ();
 FILLCELL_X4 FILLER_102_1758 ();
 FILLCELL_X4 FILLER_103_1 ();
 FILLCELL_X4 FILLER_103_24 ();
 FILLCELL_X8 FILLER_103_34 ();
 FILLCELL_X2 FILLER_103_42 ();
 FILLCELL_X4 FILLER_103_54 ();
 FILLCELL_X4 FILLER_103_61 ();
 FILLCELL_X1 FILLER_103_65 ();
 FILLCELL_X4 FILLER_103_76 ();
 FILLCELL_X8 FILLER_103_82 ();
 FILLCELL_X8 FILLER_103_93 ();
 FILLCELL_X4 FILLER_103_104 ();
 FILLCELL_X1 FILLER_103_108 ();
 FILLCELL_X4 FILLER_103_119 ();
 FILLCELL_X8 FILLER_103_125 ();
 FILLCELL_X4 FILLER_103_133 ();
 FILLCELL_X4 FILLER_103_140 ();
 FILLCELL_X8 FILLER_103_154 ();
 FILLCELL_X4 FILLER_103_162 ();
 FILLCELL_X4 FILLER_103_175 ();
 FILLCELL_X4 FILLER_103_183 ();
 FILLCELL_X4 FILLER_103_191 ();
 FILLCELL_X8 FILLER_103_198 ();
 FILLCELL_X2 FILLER_103_206 ();
 FILLCELL_X1 FILLER_103_208 ();
 FILLCELL_X4 FILLER_103_212 ();
 FILLCELL_X8 FILLER_103_219 ();
 FILLCELL_X4 FILLER_103_230 ();
 FILLCELL_X8 FILLER_103_237 ();
 FILLCELL_X4 FILLER_103_245 ();
 FILLCELL_X2 FILLER_103_249 ();
 FILLCELL_X4 FILLER_103_258 ();
 FILLCELL_X4 FILLER_103_272 ();
 FILLCELL_X4 FILLER_103_279 ();
 FILLCELL_X8 FILLER_103_293 ();
 FILLCELL_X4 FILLER_103_301 ();
 FILLCELL_X4 FILLER_103_315 ();
 FILLCELL_X4 FILLER_103_329 ();
 FILLCELL_X4 FILLER_103_343 ();
 FILLCELL_X4 FILLER_103_350 ();
 FILLCELL_X16 FILLER_103_358 ();
 FILLCELL_X4 FILLER_103_374 ();
 FILLCELL_X2 FILLER_103_378 ();
 FILLCELL_X32 FILLER_103_1518 ();
 FILLCELL_X32 FILLER_103_1550 ();
 FILLCELL_X32 FILLER_103_1582 ();
 FILLCELL_X32 FILLER_103_1614 ();
 FILLCELL_X32 FILLER_103_1646 ();
 FILLCELL_X32 FILLER_103_1678 ();
 FILLCELL_X32 FILLER_103_1710 ();
 FILLCELL_X16 FILLER_103_1742 ();
 FILLCELL_X4 FILLER_103_1758 ();
 FILLCELL_X16 FILLER_104_1 ();
 FILLCELL_X8 FILLER_104_17 ();
 FILLCELL_X2 FILLER_104_25 ();
 FILLCELL_X1 FILLER_104_27 ();
 FILLCELL_X8 FILLER_104_32 ();
 FILLCELL_X2 FILLER_104_40 ();
 FILLCELL_X16 FILLER_104_49 ();
 FILLCELL_X2 FILLER_104_65 ();
 FILLCELL_X1 FILLER_104_67 ();
 FILLCELL_X4 FILLER_104_71 ();
 FILLCELL_X1 FILLER_104_75 ();
 FILLCELL_X4 FILLER_104_86 ();
 FILLCELL_X4 FILLER_104_99 ();
 FILLCELL_X1 FILLER_104_103 ();
 FILLCELL_X4 FILLER_104_111 ();
 FILLCELL_X4 FILLER_104_125 ();
 FILLCELL_X4 FILLER_104_133 ();
 FILLCELL_X2 FILLER_104_137 ();
 FILLCELL_X1 FILLER_104_139 ();
 FILLCELL_X4 FILLER_104_147 ();
 FILLCELL_X16 FILLER_104_161 ();
 FILLCELL_X4 FILLER_104_186 ();
 FILLCELL_X1 FILLER_104_190 ();
 FILLCELL_X4 FILLER_104_201 ();
 FILLCELL_X8 FILLER_104_207 ();
 FILLCELL_X2 FILLER_104_215 ();
 FILLCELL_X1 FILLER_104_217 ();
 FILLCELL_X4 FILLER_104_222 ();
 FILLCELL_X4 FILLER_104_236 ();
 FILLCELL_X2 FILLER_104_240 ();
 FILLCELL_X1 FILLER_104_242 ();
 FILLCELL_X16 FILLER_104_245 ();
 FILLCELL_X4 FILLER_104_261 ();
 FILLCELL_X1 FILLER_104_265 ();
 FILLCELL_X4 FILLER_104_269 ();
 FILLCELL_X8 FILLER_104_282 ();
 FILLCELL_X2 FILLER_104_290 ();
 FILLCELL_X1 FILLER_104_292 ();
 FILLCELL_X4 FILLER_104_303 ();
 FILLCELL_X4 FILLER_104_316 ();
 FILLCELL_X4 FILLER_104_323 ();
 FILLCELL_X4 FILLER_104_331 ();
 FILLCELL_X32 FILLER_104_339 ();
 FILLCELL_X8 FILLER_104_371 ();
 FILLCELL_X1 FILLER_104_379 ();
 FILLCELL_X4 FILLER_104_1518 ();
 FILLCELL_X32 FILLER_104_1526 ();
 FILLCELL_X32 FILLER_104_1558 ();
 FILLCELL_X32 FILLER_104_1590 ();
 FILLCELL_X32 FILLER_104_1622 ();
 FILLCELL_X32 FILLER_104_1654 ();
 FILLCELL_X32 FILLER_104_1686 ();
 FILLCELL_X32 FILLER_104_1718 ();
 FILLCELL_X8 FILLER_104_1750 ();
 FILLCELL_X4 FILLER_104_1758 ();
 FILLCELL_X4 FILLER_105_1 ();
 FILLCELL_X2 FILLER_105_5 ();
 FILLCELL_X1 FILLER_105_7 ();
 FILLCELL_X4 FILLER_105_12 ();
 FILLCELL_X2 FILLER_105_16 ();
 FILLCELL_X4 FILLER_105_22 ();
 FILLCELL_X4 FILLER_105_35 ();
 FILLCELL_X4 FILLER_105_43 ();
 FILLCELL_X1 FILLER_105_47 ();
 FILLCELL_X4 FILLER_105_52 ();
 FILLCELL_X8 FILLER_105_66 ();
 FILLCELL_X8 FILLER_105_77 ();
 FILLCELL_X2 FILLER_105_85 ();
 FILLCELL_X1 FILLER_105_87 ();
 FILLCELL_X4 FILLER_105_91 ();
 FILLCELL_X2 FILLER_105_95 ();
 FILLCELL_X4 FILLER_105_106 ();
 FILLCELL_X2 FILLER_105_110 ();
 FILLCELL_X8 FILLER_105_115 ();
 FILLCELL_X1 FILLER_105_123 ();
 FILLCELL_X8 FILLER_105_127 ();
 FILLCELL_X4 FILLER_105_137 ();
 FILLCELL_X8 FILLER_105_148 ();
 FILLCELL_X4 FILLER_105_159 ();
 FILLCELL_X4 FILLER_105_166 ();
 FILLCELL_X4 FILLER_105_174 ();
 FILLCELL_X8 FILLER_105_181 ();
 FILLCELL_X1 FILLER_105_189 ();
 FILLCELL_X4 FILLER_105_197 ();
 FILLCELL_X8 FILLER_105_211 ();
 FILLCELL_X1 FILLER_105_219 ();
 FILLCELL_X4 FILLER_105_227 ();
 FILLCELL_X4 FILLER_105_241 ();
 FILLCELL_X2 FILLER_105_245 ();
 FILLCELL_X4 FILLER_105_250 ();
 FILLCELL_X8 FILLER_105_263 ();
 FILLCELL_X2 FILLER_105_271 ();
 FILLCELL_X1 FILLER_105_273 ();
 FILLCELL_X4 FILLER_105_277 ();
 FILLCELL_X2 FILLER_105_281 ();
 FILLCELL_X1 FILLER_105_283 ();
 FILLCELL_X4 FILLER_105_291 ();
 FILLCELL_X4 FILLER_105_298 ();
 FILLCELL_X8 FILLER_105_304 ();
 FILLCELL_X4 FILLER_105_315 ();
 FILLCELL_X4 FILLER_105_329 ();
 FILLCELL_X32 FILLER_105_335 ();
 FILLCELL_X8 FILLER_105_367 ();
 FILLCELL_X4 FILLER_105_375 ();
 FILLCELL_X1 FILLER_105_379 ();
 FILLCELL_X8 FILLER_105_1518 ();
 FILLCELL_X1 FILLER_105_1526 ();
 FILLCELL_X32 FILLER_105_1546 ();
 FILLCELL_X32 FILLER_105_1578 ();
 FILLCELL_X32 FILLER_105_1610 ();
 FILLCELL_X32 FILLER_105_1642 ();
 FILLCELL_X32 FILLER_105_1674 ();
 FILLCELL_X32 FILLER_105_1706 ();
 FILLCELL_X16 FILLER_105_1738 ();
 FILLCELL_X8 FILLER_105_1754 ();
 FILLCELL_X4 FILLER_106_1 ();
 FILLCELL_X8 FILLER_106_24 ();
 FILLCELL_X4 FILLER_106_32 ();
 FILLCELL_X1 FILLER_106_36 ();
 FILLCELL_X4 FILLER_106_46 ();
 FILLCELL_X4 FILLER_106_53 ();
 FILLCELL_X4 FILLER_106_59 ();
 FILLCELL_X4 FILLER_106_70 ();
 FILLCELL_X8 FILLER_106_83 ();
 FILLCELL_X4 FILLER_106_91 ();
 FILLCELL_X4 FILLER_106_98 ();
 FILLCELL_X8 FILLER_106_112 ();
 FILLCELL_X1 FILLER_106_120 ();
 FILLCELL_X4 FILLER_106_124 ();
 FILLCELL_X1 FILLER_106_128 ();
 FILLCELL_X4 FILLER_106_139 ();
 FILLCELL_X1 FILLER_106_143 ();
 FILLCELL_X4 FILLER_106_146 ();
 FILLCELL_X32 FILLER_106_160 ();
 FILLCELL_X8 FILLER_106_192 ();
 FILLCELL_X4 FILLER_106_200 ();
 FILLCELL_X4 FILLER_106_207 ();
 FILLCELL_X4 FILLER_106_220 ();
 FILLCELL_X4 FILLER_106_227 ();
 FILLCELL_X8 FILLER_106_240 ();
 FILLCELL_X2 FILLER_106_248 ();
 FILLCELL_X4 FILLER_106_253 ();
 FILLCELL_X1 FILLER_106_257 ();
 FILLCELL_X4 FILLER_106_261 ();
 FILLCELL_X4 FILLER_106_274 ();
 FILLCELL_X4 FILLER_106_281 ();
 FILLCELL_X8 FILLER_106_287 ();
 FILLCELL_X4 FILLER_106_295 ();
 FILLCELL_X2 FILLER_106_299 ();
 FILLCELL_X1 FILLER_106_301 ();
 FILLCELL_X32 FILLER_106_305 ();
 FILLCELL_X32 FILLER_106_337 ();
 FILLCELL_X8 FILLER_106_369 ();
 FILLCELL_X2 FILLER_106_377 ();
 FILLCELL_X1 FILLER_106_379 ();
 FILLCELL_X32 FILLER_106_1518 ();
 FILLCELL_X32 FILLER_106_1550 ();
 FILLCELL_X32 FILLER_106_1582 ();
 FILLCELL_X32 FILLER_106_1614 ();
 FILLCELL_X32 FILLER_106_1646 ();
 FILLCELL_X32 FILLER_106_1678 ();
 FILLCELL_X32 FILLER_106_1710 ();
 FILLCELL_X16 FILLER_106_1742 ();
 FILLCELL_X4 FILLER_106_1758 ();
 FILLCELL_X16 FILLER_107_1 ();
 FILLCELL_X8 FILLER_107_17 ();
 FILLCELL_X4 FILLER_107_25 ();
 FILLCELL_X1 FILLER_107_29 ();
 FILLCELL_X4 FILLER_107_33 ();
 FILLCELL_X1 FILLER_107_37 ();
 FILLCELL_X8 FILLER_107_41 ();
 FILLCELL_X4 FILLER_107_49 ();
 FILLCELL_X4 FILLER_107_55 ();
 FILLCELL_X2 FILLER_107_59 ();
 FILLCELL_X4 FILLER_107_71 ();
 FILLCELL_X2 FILLER_107_75 ();
 FILLCELL_X1 FILLER_107_77 ();
 FILLCELL_X8 FILLER_107_81 ();
 FILLCELL_X8 FILLER_107_92 ();
 FILLCELL_X1 FILLER_107_100 ();
 FILLCELL_X8 FILLER_107_108 ();
 FILLCELL_X1 FILLER_107_116 ();
 FILLCELL_X8 FILLER_107_126 ();
 FILLCELL_X1 FILLER_107_134 ();
 FILLCELL_X4 FILLER_107_138 ();
 FILLCELL_X4 FILLER_107_151 ();
 FILLCELL_X1 FILLER_107_155 ();
 FILLCELL_X4 FILLER_107_159 ();
 FILLCELL_X8 FILLER_107_172 ();
 FILLCELL_X4 FILLER_107_180 ();
 FILLCELL_X2 FILLER_107_184 ();
 FILLCELL_X1 FILLER_107_186 ();
 FILLCELL_X4 FILLER_107_190 ();
 FILLCELL_X8 FILLER_107_203 ();
 FILLCELL_X8 FILLER_107_214 ();
 FILLCELL_X1 FILLER_107_222 ();
 FILLCELL_X8 FILLER_107_226 ();
 FILLCELL_X4 FILLER_107_234 ();
 FILLCELL_X4 FILLER_107_241 ();
 FILLCELL_X4 FILLER_107_255 ();
 FILLCELL_X1 FILLER_107_259 ();
 FILLCELL_X4 FILLER_107_270 ();
 FILLCELL_X4 FILLER_107_284 ();
 FILLCELL_X8 FILLER_107_298 ();
 FILLCELL_X1 FILLER_107_306 ();
 FILLCELL_X32 FILLER_107_316 ();
 FILLCELL_X32 FILLER_107_348 ();
 FILLCELL_X32 FILLER_107_1518 ();
 FILLCELL_X32 FILLER_107_1550 ();
 FILLCELL_X32 FILLER_107_1582 ();
 FILLCELL_X32 FILLER_107_1614 ();
 FILLCELL_X32 FILLER_107_1646 ();
 FILLCELL_X32 FILLER_107_1678 ();
 FILLCELL_X32 FILLER_107_1710 ();
 FILLCELL_X8 FILLER_107_1742 ();
 FILLCELL_X4 FILLER_107_1750 ();
 FILLCELL_X1 FILLER_107_1754 ();
 FILLCELL_X4 FILLER_107_1758 ();
 FILLCELL_X4 FILLER_108_1 ();
 FILLCELL_X2 FILLER_108_5 ();
 FILLCELL_X1 FILLER_108_7 ();
 FILLCELL_X16 FILLER_108_12 ();
 FILLCELL_X2 FILLER_108_28 ();
 FILLCELL_X16 FILLER_108_34 ();
 FILLCELL_X2 FILLER_108_50 ();
 FILLCELL_X8 FILLER_108_58 ();
 FILLCELL_X1 FILLER_108_66 ();
 FILLCELL_X4 FILLER_108_70 ();
 FILLCELL_X4 FILLER_108_83 ();
 FILLCELL_X4 FILLER_108_97 ();
 FILLCELL_X4 FILLER_108_103 ();
 FILLCELL_X8 FILLER_108_117 ();
 FILLCELL_X1 FILLER_108_125 ();
 FILLCELL_X4 FILLER_108_135 ();
 FILLCELL_X4 FILLER_108_142 ();
 FILLCELL_X4 FILLER_108_149 ();
 FILLCELL_X8 FILLER_108_162 ();
 FILLCELL_X1 FILLER_108_170 ();
 FILLCELL_X4 FILLER_108_180 ();
 FILLCELL_X4 FILLER_108_194 ();
 FILLCELL_X2 FILLER_108_198 ();
 FILLCELL_X4 FILLER_108_203 ();
 FILLCELL_X4 FILLER_108_216 ();
 FILLCELL_X2 FILLER_108_220 ();
 FILLCELL_X16 FILLER_108_232 ();
 FILLCELL_X4 FILLER_108_248 ();
 FILLCELL_X2 FILLER_108_252 ();
 FILLCELL_X1 FILLER_108_254 ();
 FILLCELL_X4 FILLER_108_259 ();
 FILLCELL_X8 FILLER_108_265 ();
 FILLCELL_X2 FILLER_108_273 ();
 FILLCELL_X1 FILLER_108_275 ();
 FILLCELL_X4 FILLER_108_283 ();
 FILLCELL_X2 FILLER_108_287 ();
 FILLCELL_X4 FILLER_108_292 ();
 FILLCELL_X32 FILLER_108_305 ();
 FILLCELL_X32 FILLER_108_337 ();
 FILLCELL_X8 FILLER_108_369 ();
 FILLCELL_X2 FILLER_108_377 ();
 FILLCELL_X1 FILLER_108_379 ();
 FILLCELL_X32 FILLER_108_1518 ();
 FILLCELL_X32 FILLER_108_1550 ();
 FILLCELL_X32 FILLER_108_1582 ();
 FILLCELL_X32 FILLER_108_1614 ();
 FILLCELL_X32 FILLER_108_1646 ();
 FILLCELL_X32 FILLER_108_1678 ();
 FILLCELL_X32 FILLER_108_1710 ();
 FILLCELL_X16 FILLER_108_1742 ();
 FILLCELL_X4 FILLER_108_1758 ();
 FILLCELL_X4 FILLER_109_1 ();
 FILLCELL_X4 FILLER_109_24 ();
 FILLCELL_X2 FILLER_109_28 ();
 FILLCELL_X8 FILLER_109_49 ();
 FILLCELL_X4 FILLER_109_57 ();
 FILLCELL_X8 FILLER_109_65 ();
 FILLCELL_X4 FILLER_109_73 ();
 FILLCELL_X8 FILLER_109_80 ();
 FILLCELL_X2 FILLER_109_88 ();
 FILLCELL_X1 FILLER_109_90 ();
 FILLCELL_X4 FILLER_109_95 ();
 FILLCELL_X2 FILLER_109_99 ();
 FILLCELL_X4 FILLER_109_111 ();
 FILLCELL_X8 FILLER_109_118 ();
 FILLCELL_X2 FILLER_109_126 ();
 FILLCELL_X16 FILLER_109_131 ();
 FILLCELL_X8 FILLER_109_147 ();
 FILLCELL_X4 FILLER_109_155 ();
 FILLCELL_X2 FILLER_109_159 ();
 FILLCELL_X4 FILLER_109_164 ();
 FILLCELL_X8 FILLER_109_171 ();
 FILLCELL_X4 FILLER_109_179 ();
 FILLCELL_X2 FILLER_109_183 ();
 FILLCELL_X1 FILLER_109_185 ();
 FILLCELL_X4 FILLER_109_189 ();
 FILLCELL_X2 FILLER_109_193 ();
 FILLCELL_X1 FILLER_109_195 ();
 FILLCELL_X4 FILLER_109_199 ();
 FILLCELL_X2 FILLER_109_203 ();
 FILLCELL_X8 FILLER_109_215 ();
 FILLCELL_X4 FILLER_109_223 ();
 FILLCELL_X2 FILLER_109_227 ();
 FILLCELL_X4 FILLER_109_239 ();
 FILLCELL_X4 FILLER_109_246 ();
 FILLCELL_X8 FILLER_109_252 ();
 FILLCELL_X1 FILLER_109_260 ();
 FILLCELL_X8 FILLER_109_264 ();
 FILLCELL_X16 FILLER_109_274 ();
 FILLCELL_X4 FILLER_109_290 ();
 FILLCELL_X1 FILLER_109_294 ();
 FILLCELL_X32 FILLER_109_298 ();
 FILLCELL_X32 FILLER_109_330 ();
 FILLCELL_X16 FILLER_109_362 ();
 FILLCELL_X2 FILLER_109_378 ();
 FILLCELL_X32 FILLER_109_1518 ();
 FILLCELL_X32 FILLER_109_1550 ();
 FILLCELL_X32 FILLER_109_1582 ();
 FILLCELL_X32 FILLER_109_1614 ();
 FILLCELL_X32 FILLER_109_1646 ();
 FILLCELL_X32 FILLER_109_1678 ();
 FILLCELL_X32 FILLER_109_1710 ();
 FILLCELL_X16 FILLER_109_1742 ();
 FILLCELL_X4 FILLER_109_1758 ();
 FILLCELL_X32 FILLER_110_1 ();
 FILLCELL_X16 FILLER_110_33 ();
 FILLCELL_X2 FILLER_110_49 ();
 FILLCELL_X1 FILLER_110_51 ();
 FILLCELL_X4 FILLER_110_56 ();
 FILLCELL_X4 FILLER_110_67 ();
 FILLCELL_X4 FILLER_110_77 ();
 FILLCELL_X1 FILLER_110_81 ();
 FILLCELL_X4 FILLER_110_92 ();
 FILLCELL_X1 FILLER_110_96 ();
 FILLCELL_X8 FILLER_110_99 ();
 FILLCELL_X4 FILLER_110_110 ();
 FILLCELL_X4 FILLER_110_117 ();
 FILLCELL_X2 FILLER_110_121 ();
 FILLCELL_X4 FILLER_110_126 ();
 FILLCELL_X2 FILLER_110_130 ();
 FILLCELL_X1 FILLER_110_132 ();
 FILLCELL_X4 FILLER_110_143 ();
 FILLCELL_X4 FILLER_110_149 ();
 FILLCELL_X2 FILLER_110_153 ();
 FILLCELL_X1 FILLER_110_155 ();
 FILLCELL_X4 FILLER_110_159 ();
 FILLCELL_X4 FILLER_110_173 ();
 FILLCELL_X16 FILLER_110_179 ();
 FILLCELL_X2 FILLER_110_195 ();
 FILLCELL_X4 FILLER_110_204 ();
 FILLCELL_X8 FILLER_110_210 ();
 FILLCELL_X2 FILLER_110_218 ();
 FILLCELL_X4 FILLER_110_227 ();
 FILLCELL_X1 FILLER_110_231 ();
 FILLCELL_X4 FILLER_110_241 ();
 FILLCELL_X2 FILLER_110_245 ();
 FILLCELL_X4 FILLER_110_256 ();
 FILLCELL_X4 FILLER_110_270 ();
 FILLCELL_X1 FILLER_110_274 ();
 FILLCELL_X4 FILLER_110_281 ();
 FILLCELL_X4 FILLER_110_289 ();
 FILLCELL_X32 FILLER_110_299 ();
 FILLCELL_X32 FILLER_110_331 ();
 FILLCELL_X16 FILLER_110_363 ();
 FILLCELL_X1 FILLER_110_379 ();
 FILLCELL_X32 FILLER_110_1518 ();
 FILLCELL_X32 FILLER_110_1550 ();
 FILLCELL_X32 FILLER_110_1582 ();
 FILLCELL_X32 FILLER_110_1614 ();
 FILLCELL_X32 FILLER_110_1646 ();
 FILLCELL_X32 FILLER_110_1678 ();
 FILLCELL_X32 FILLER_110_1710 ();
 FILLCELL_X16 FILLER_110_1742 ();
 FILLCELL_X4 FILLER_110_1758 ();
 FILLCELL_X32 FILLER_111_1 ();
 FILLCELL_X16 FILLER_111_33 ();
 FILLCELL_X8 FILLER_111_49 ();
 FILLCELL_X4 FILLER_111_57 ();
 FILLCELL_X8 FILLER_111_67 ();
 FILLCELL_X4 FILLER_111_75 ();
 FILLCELL_X2 FILLER_111_79 ();
 FILLCELL_X4 FILLER_111_85 ();
 FILLCELL_X8 FILLER_111_91 ();
 FILLCELL_X4 FILLER_111_99 ();
 FILLCELL_X2 FILLER_111_103 ();
 FILLCELL_X4 FILLER_111_108 ();
 FILLCELL_X4 FILLER_111_121 ();
 FILLCELL_X2 FILLER_111_125 ();
 FILLCELL_X1 FILLER_111_127 ();
 FILLCELL_X4 FILLER_111_137 ();
 FILLCELL_X4 FILLER_111_145 ();
 FILLCELL_X1 FILLER_111_149 ();
 FILLCELL_X4 FILLER_111_160 ();
 FILLCELL_X1 FILLER_111_164 ();
 FILLCELL_X4 FILLER_111_168 ();
 FILLCELL_X4 FILLER_111_182 ();
 FILLCELL_X8 FILLER_111_189 ();
 FILLCELL_X4 FILLER_111_197 ();
 FILLCELL_X1 FILLER_111_201 ();
 FILLCELL_X4 FILLER_111_205 ();
 FILLCELL_X2 FILLER_111_209 ();
 FILLCELL_X1 FILLER_111_211 ();
 FILLCELL_X8 FILLER_111_216 ();
 FILLCELL_X1 FILLER_111_224 ();
 FILLCELL_X4 FILLER_111_228 ();
 FILLCELL_X4 FILLER_111_235 ();
 FILLCELL_X8 FILLER_111_242 ();
 FILLCELL_X8 FILLER_111_256 ();
 FILLCELL_X4 FILLER_111_271 ();
 FILLCELL_X1 FILLER_111_275 ();
 FILLCELL_X4 FILLER_111_280 ();
 FILLCELL_X4 FILLER_111_291 ();
 FILLCELL_X2 FILLER_111_295 ();
 FILLCELL_X1 FILLER_111_297 ();
 FILLCELL_X32 FILLER_111_317 ();
 FILLCELL_X16 FILLER_111_349 ();
 FILLCELL_X8 FILLER_111_365 ();
 FILLCELL_X4 FILLER_111_373 ();
 FILLCELL_X2 FILLER_111_377 ();
 FILLCELL_X1 FILLER_111_379 ();
 FILLCELL_X32 FILLER_111_1518 ();
 FILLCELL_X32 FILLER_111_1550 ();
 FILLCELL_X32 FILLER_111_1582 ();
 FILLCELL_X32 FILLER_111_1614 ();
 FILLCELL_X32 FILLER_111_1646 ();
 FILLCELL_X32 FILLER_111_1678 ();
 FILLCELL_X32 FILLER_111_1710 ();
 FILLCELL_X16 FILLER_111_1742 ();
 FILLCELL_X4 FILLER_111_1758 ();
 FILLCELL_X4 FILLER_112_1 ();
 FILLCELL_X32 FILLER_112_8 ();
 FILLCELL_X16 FILLER_112_40 ();
 FILLCELL_X8 FILLER_112_56 ();
 FILLCELL_X16 FILLER_112_68 ();
 FILLCELL_X4 FILLER_112_84 ();
 FILLCELL_X2 FILLER_112_88 ();
 FILLCELL_X4 FILLER_112_100 ();
 FILLCELL_X1 FILLER_112_104 ();
 FILLCELL_X4 FILLER_112_112 ();
 FILLCELL_X8 FILLER_112_119 ();
 FILLCELL_X4 FILLER_112_127 ();
 FILLCELL_X2 FILLER_112_131 ();
 FILLCELL_X1 FILLER_112_133 ();
 FILLCELL_X4 FILLER_112_137 ();
 FILLCELL_X4 FILLER_112_151 ();
 FILLCELL_X4 FILLER_112_157 ();
 FILLCELL_X2 FILLER_112_161 ();
 FILLCELL_X4 FILLER_112_170 ();
 FILLCELL_X4 FILLER_112_183 ();
 FILLCELL_X4 FILLER_112_196 ();
 FILLCELL_X4 FILLER_112_210 ();
 FILLCELL_X4 FILLER_112_220 ();
 FILLCELL_X2 FILLER_112_224 ();
 FILLCELL_X1 FILLER_112_226 ();
 FILLCELL_X4 FILLER_112_237 ();
 FILLCELL_X2 FILLER_112_241 ();
 FILLCELL_X1 FILLER_112_243 ();
 FILLCELL_X4 FILLER_112_251 ();
 FILLCELL_X16 FILLER_112_261 ();
 FILLCELL_X2 FILLER_112_277 ();
 FILLCELL_X1 FILLER_112_279 ();
 FILLCELL_X4 FILLER_112_283 ();
 FILLCELL_X1 FILLER_112_287 ();
 FILLCELL_X4 FILLER_112_294 ();
 FILLCELL_X32 FILLER_112_302 ();
 FILLCELL_X32 FILLER_112_334 ();
 FILLCELL_X8 FILLER_112_366 ();
 FILLCELL_X4 FILLER_112_374 ();
 FILLCELL_X2 FILLER_112_378 ();
 FILLCELL_X32 FILLER_112_1518 ();
 FILLCELL_X32 FILLER_112_1550 ();
 FILLCELL_X32 FILLER_112_1582 ();
 FILLCELL_X32 FILLER_112_1614 ();
 FILLCELL_X32 FILLER_112_1646 ();
 FILLCELL_X32 FILLER_112_1678 ();
 FILLCELL_X32 FILLER_112_1710 ();
 FILLCELL_X16 FILLER_112_1742 ();
 FILLCELL_X4 FILLER_112_1758 ();
 FILLCELL_X32 FILLER_113_1 ();
 FILLCELL_X16 FILLER_113_33 ();
 FILLCELL_X8 FILLER_113_49 ();
 FILLCELL_X4 FILLER_113_57 ();
 FILLCELL_X1 FILLER_113_61 ();
 FILLCELL_X16 FILLER_113_81 ();
 FILLCELL_X2 FILLER_113_97 ();
 FILLCELL_X1 FILLER_113_99 ();
 FILLCELL_X4 FILLER_113_106 ();
 FILLCELL_X16 FILLER_113_116 ();
 FILLCELL_X8 FILLER_113_132 ();
 FILLCELL_X2 FILLER_113_140 ();
 FILLCELL_X1 FILLER_113_142 ();
 FILLCELL_X4 FILLER_113_150 ();
 FILLCELL_X2 FILLER_113_154 ();
 FILLCELL_X4 FILLER_113_166 ();
 FILLCELL_X2 FILLER_113_170 ();
 FILLCELL_X1 FILLER_113_172 ();
 FILLCELL_X16 FILLER_113_176 ();
 FILLCELL_X4 FILLER_113_192 ();
 FILLCELL_X1 FILLER_113_196 ();
 FILLCELL_X4 FILLER_113_201 ();
 FILLCELL_X4 FILLER_113_212 ();
 FILLCELL_X1 FILLER_113_216 ();
 FILLCELL_X4 FILLER_113_219 ();
 FILLCELL_X8 FILLER_113_233 ();
 FILLCELL_X4 FILLER_113_241 ();
 FILLCELL_X1 FILLER_113_245 ();
 FILLCELL_X16 FILLER_113_249 ();
 FILLCELL_X2 FILLER_113_265 ();
 FILLCELL_X1 FILLER_113_267 ();
 FILLCELL_X4 FILLER_113_271 ();
 FILLCELL_X4 FILLER_113_278 ();
 FILLCELL_X4 FILLER_113_285 ();
 FILLCELL_X4 FILLER_113_292 ();
 FILLCELL_X2 FILLER_113_296 ();
 FILLCELL_X4 FILLER_113_300 ();
 FILLCELL_X2 FILLER_113_304 ();
 FILLCELL_X4 FILLER_113_309 ();
 FILLCELL_X8 FILLER_113_318 ();
 FILLCELL_X4 FILLER_113_326 ();
 FILLCELL_X2 FILLER_113_330 ();
 FILLCELL_X32 FILLER_113_335 ();
 FILLCELL_X8 FILLER_113_367 ();
 FILLCELL_X4 FILLER_113_375 ();
 FILLCELL_X1 FILLER_113_379 ();
 FILLCELL_X32 FILLER_113_1518 ();
 FILLCELL_X32 FILLER_113_1550 ();
 FILLCELL_X32 FILLER_113_1582 ();
 FILLCELL_X32 FILLER_113_1614 ();
 FILLCELL_X32 FILLER_113_1646 ();
 FILLCELL_X32 FILLER_113_1678 ();
 FILLCELL_X32 FILLER_113_1710 ();
 FILLCELL_X16 FILLER_113_1742 ();
 FILLCELL_X4 FILLER_113_1758 ();
 FILLCELL_X32 FILLER_114_1 ();
 FILLCELL_X32 FILLER_114_33 ();
 FILLCELL_X32 FILLER_114_65 ();
 FILLCELL_X16 FILLER_114_97 ();
 FILLCELL_X1 FILLER_114_113 ();
 FILLCELL_X32 FILLER_114_118 ();
 FILLCELL_X32 FILLER_114_150 ();
 FILLCELL_X16 FILLER_114_182 ();
 FILLCELL_X4 FILLER_114_198 ();
 FILLCELL_X2 FILLER_114_202 ();
 FILLCELL_X1 FILLER_114_204 ();
 FILLCELL_X32 FILLER_114_209 ();
 FILLCELL_X16 FILLER_114_241 ();
 FILLCELL_X4 FILLER_114_257 ();
 FILLCELL_X2 FILLER_114_261 ();
 FILLCELL_X1 FILLER_114_263 ();
 FILLCELL_X4 FILLER_114_267 ();
 FILLCELL_X4 FILLER_114_288 ();
 FILLCELL_X8 FILLER_114_311 ();
 FILLCELL_X2 FILLER_114_319 ();
 FILLCELL_X4 FILLER_114_326 ();
 FILLCELL_X8 FILLER_114_333 ();
 FILLCELL_X2 FILLER_114_341 ();
 FILLCELL_X4 FILLER_114_349 ();
 FILLCELL_X8 FILLER_114_356 ();
 FILLCELL_X2 FILLER_114_364 ();
 FILLCELL_X4 FILLER_114_369 ();
 FILLCELL_X4 FILLER_114_376 ();
 FILLCELL_X32 FILLER_114_1518 ();
 FILLCELL_X32 FILLER_114_1550 ();
 FILLCELL_X32 FILLER_114_1582 ();
 FILLCELL_X32 FILLER_114_1614 ();
 FILLCELL_X32 FILLER_114_1646 ();
 FILLCELL_X32 FILLER_114_1678 ();
 FILLCELL_X32 FILLER_114_1710 ();
 FILLCELL_X16 FILLER_114_1742 ();
 FILLCELL_X4 FILLER_114_1758 ();
 FILLCELL_X32 FILLER_115_1 ();
 FILLCELL_X32 FILLER_115_33 ();
 FILLCELL_X32 FILLER_115_65 ();
 FILLCELL_X8 FILLER_115_97 ();
 FILLCELL_X4 FILLER_115_105 ();
 FILLCELL_X2 FILLER_115_109 ();
 FILLCELL_X1 FILLER_115_111 ();
 FILLCELL_X32 FILLER_115_129 ();
 FILLCELL_X32 FILLER_115_161 ();
 FILLCELL_X32 FILLER_115_193 ();
 FILLCELL_X32 FILLER_115_225 ();
 FILLCELL_X1 FILLER_115_257 ();
 FILLCELL_X4 FILLER_115_261 ();
 FILLCELL_X8 FILLER_115_270 ();
 FILLCELL_X1 FILLER_115_278 ();
 FILLCELL_X4 FILLER_115_284 ();
 FILLCELL_X2 FILLER_115_288 ();
 FILLCELL_X4 FILLER_115_294 ();
 FILLCELL_X4 FILLER_115_301 ();
 FILLCELL_X4 FILLER_115_309 ();
 FILLCELL_X4 FILLER_115_330 ();
 FILLCELL_X2 FILLER_115_334 ();
 FILLCELL_X1 FILLER_115_336 ();
 FILLCELL_X8 FILLER_115_354 ();
 FILLCELL_X2 FILLER_115_362 ();
 FILLCELL_X4 FILLER_115_367 ();
 FILLCELL_X4 FILLER_115_374 ();
 FILLCELL_X2 FILLER_115_378 ();
 FILLCELL_X32 FILLER_115_1518 ();
 FILLCELL_X32 FILLER_115_1550 ();
 FILLCELL_X32 FILLER_115_1582 ();
 FILLCELL_X32 FILLER_115_1614 ();
 FILLCELL_X32 FILLER_115_1646 ();
 FILLCELL_X32 FILLER_115_1678 ();
 FILLCELL_X32 FILLER_115_1710 ();
 FILLCELL_X16 FILLER_115_1742 ();
 FILLCELL_X4 FILLER_115_1758 ();
 FILLCELL_X32 FILLER_116_1 ();
 FILLCELL_X32 FILLER_116_33 ();
 FILLCELL_X32 FILLER_116_65 ();
 FILLCELL_X32 FILLER_116_97 ();
 FILLCELL_X32 FILLER_116_129 ();
 FILLCELL_X32 FILLER_116_161 ();
 FILLCELL_X32 FILLER_116_193 ();
 FILLCELL_X16 FILLER_116_225 ();
 FILLCELL_X8 FILLER_116_241 ();
 FILLCELL_X4 FILLER_116_249 ();
 FILLCELL_X2 FILLER_116_253 ();
 FILLCELL_X4 FILLER_116_272 ();
 FILLCELL_X4 FILLER_116_281 ();
 FILLCELL_X2 FILLER_116_285 ();
 FILLCELL_X1 FILLER_116_287 ();
 FILLCELL_X4 FILLER_116_293 ();
 FILLCELL_X4 FILLER_116_301 ();
 FILLCELL_X1 FILLER_116_305 ();
 FILLCELL_X4 FILLER_116_309 ();
 FILLCELL_X4 FILLER_116_316 ();
 FILLCELL_X8 FILLER_116_324 ();
 FILLCELL_X2 FILLER_116_332 ();
 FILLCELL_X4 FILLER_116_339 ();
 FILLCELL_X8 FILLER_116_347 ();
 FILLCELL_X4 FILLER_116_358 ();
 FILLCELL_X2 FILLER_116_362 ();
 FILLCELL_X4 FILLER_116_367 ();
 FILLCELL_X4 FILLER_116_374 ();
 FILLCELL_X2 FILLER_116_378 ();
 FILLCELL_X32 FILLER_116_1518 ();
 FILLCELL_X32 FILLER_116_1550 ();
 FILLCELL_X32 FILLER_116_1582 ();
 FILLCELL_X32 FILLER_116_1614 ();
 FILLCELL_X32 FILLER_116_1646 ();
 FILLCELL_X32 FILLER_116_1678 ();
 FILLCELL_X32 FILLER_116_1710 ();
 FILLCELL_X16 FILLER_116_1742 ();
 FILLCELL_X4 FILLER_116_1758 ();
 FILLCELL_X32 FILLER_117_1 ();
 FILLCELL_X32 FILLER_117_33 ();
 FILLCELL_X32 FILLER_117_65 ();
 FILLCELL_X32 FILLER_117_97 ();
 FILLCELL_X32 FILLER_117_129 ();
 FILLCELL_X32 FILLER_117_161 ();
 FILLCELL_X32 FILLER_117_193 ();
 FILLCELL_X16 FILLER_117_225 ();
 FILLCELL_X8 FILLER_117_241 ();
 FILLCELL_X1 FILLER_117_249 ();
 FILLCELL_X4 FILLER_117_253 ();
 FILLCELL_X4 FILLER_117_260 ();
 FILLCELL_X4 FILLER_117_267 ();
 FILLCELL_X2 FILLER_117_271 ();
 FILLCELL_X4 FILLER_117_276 ();
 FILLCELL_X1 FILLER_117_280 ();
 FILLCELL_X4 FILLER_117_285 ();
 FILLCELL_X2 FILLER_117_289 ();
 FILLCELL_X1 FILLER_117_291 ();
 FILLCELL_X4 FILLER_117_296 ();
 FILLCELL_X4 FILLER_117_302 ();
 FILLCELL_X4 FILLER_117_311 ();
 FILLCELL_X4 FILLER_117_320 ();
 FILLCELL_X2 FILLER_117_324 ();
 FILLCELL_X4 FILLER_117_331 ();
 FILLCELL_X4 FILLER_117_337 ();
 FILLCELL_X4 FILLER_117_345 ();
 FILLCELL_X2 FILLER_117_349 ();
 FILLCELL_X4 FILLER_117_354 ();
 FILLCELL_X4 FILLER_117_361 ();
 FILLCELL_X1 FILLER_117_365 ();
 FILLCELL_X4 FILLER_117_369 ();
 FILLCELL_X4 FILLER_117_376 ();
 FILLCELL_X32 FILLER_117_1518 ();
 FILLCELL_X32 FILLER_117_1550 ();
 FILLCELL_X32 FILLER_117_1582 ();
 FILLCELL_X32 FILLER_117_1614 ();
 FILLCELL_X32 FILLER_117_1646 ();
 FILLCELL_X32 FILLER_117_1678 ();
 FILLCELL_X32 FILLER_117_1710 ();
 FILLCELL_X8 FILLER_117_1742 ();
 FILLCELL_X4 FILLER_117_1750 ();
 FILLCELL_X1 FILLER_117_1754 ();
 FILLCELL_X4 FILLER_117_1758 ();
 FILLCELL_X32 FILLER_118_1 ();
 FILLCELL_X32 FILLER_118_33 ();
 FILLCELL_X32 FILLER_118_65 ();
 FILLCELL_X32 FILLER_118_97 ();
 FILLCELL_X32 FILLER_118_129 ();
 FILLCELL_X32 FILLER_118_161 ();
 FILLCELL_X32 FILLER_118_193 ();
 FILLCELL_X32 FILLER_118_225 ();
 FILLCELL_X1 FILLER_118_257 ();
 FILLCELL_X4 FILLER_118_261 ();
 FILLCELL_X4 FILLER_118_274 ();
 FILLCELL_X4 FILLER_118_281 ();
 FILLCELL_X4 FILLER_118_287 ();
 FILLCELL_X4 FILLER_118_296 ();
 FILLCELL_X4 FILLER_118_313 ();
 FILLCELL_X4 FILLER_118_320 ();
 FILLCELL_X1 FILLER_118_324 ();
 FILLCELL_X4 FILLER_118_334 ();
 FILLCELL_X1 FILLER_118_338 ();
 FILLCELL_X4 FILLER_118_343 ();
 FILLCELL_X8 FILLER_118_364 ();
 FILLCELL_X1 FILLER_118_372 ();
 FILLCELL_X4 FILLER_118_376 ();
 FILLCELL_X32 FILLER_118_1518 ();
 FILLCELL_X32 FILLER_118_1550 ();
 FILLCELL_X32 FILLER_118_1582 ();
 FILLCELL_X32 FILLER_118_1614 ();
 FILLCELL_X32 FILLER_118_1646 ();
 FILLCELL_X32 FILLER_118_1678 ();
 FILLCELL_X32 FILLER_118_1710 ();
 FILLCELL_X16 FILLER_118_1742 ();
 FILLCELL_X4 FILLER_118_1758 ();
 FILLCELL_X32 FILLER_119_1 ();
 FILLCELL_X32 FILLER_119_33 ();
 FILLCELL_X32 FILLER_119_65 ();
 FILLCELL_X32 FILLER_119_97 ();
 FILLCELL_X32 FILLER_119_129 ();
 FILLCELL_X32 FILLER_119_161 ();
 FILLCELL_X32 FILLER_119_193 ();
 FILLCELL_X16 FILLER_119_225 ();
 FILLCELL_X4 FILLER_119_241 ();
 FILLCELL_X4 FILLER_119_264 ();
 FILLCELL_X2 FILLER_119_268 ();
 FILLCELL_X1 FILLER_119_270 ();
 FILLCELL_X8 FILLER_119_282 ();
 FILLCELL_X4 FILLER_119_290 ();
 FILLCELL_X2 FILLER_119_294 ();
 FILLCELL_X4 FILLER_119_298 ();
 FILLCELL_X2 FILLER_119_302 ();
 FILLCELL_X4 FILLER_119_307 ();
 FILLCELL_X4 FILLER_119_314 ();
 FILLCELL_X4 FILLER_119_323 ();
 FILLCELL_X2 FILLER_119_327 ();
 FILLCELL_X1 FILLER_119_329 ();
 FILLCELL_X4 FILLER_119_333 ();
 FILLCELL_X4 FILLER_119_340 ();
 FILLCELL_X4 FILLER_119_349 ();
 FILLCELL_X4 FILLER_119_357 ();
 FILLCELL_X2 FILLER_119_361 ();
 FILLCELL_X4 FILLER_119_369 ();
 FILLCELL_X4 FILLER_119_376 ();
 FILLCELL_X32 FILLER_119_1518 ();
 FILLCELL_X32 FILLER_119_1550 ();
 FILLCELL_X32 FILLER_119_1582 ();
 FILLCELL_X32 FILLER_119_1614 ();
 FILLCELL_X32 FILLER_119_1646 ();
 FILLCELL_X32 FILLER_119_1678 ();
 FILLCELL_X32 FILLER_119_1710 ();
 FILLCELL_X16 FILLER_119_1742 ();
 FILLCELL_X4 FILLER_119_1758 ();
 FILLCELL_X32 FILLER_120_1 ();
 FILLCELL_X32 FILLER_120_33 ();
 FILLCELL_X32 FILLER_120_65 ();
 FILLCELL_X32 FILLER_120_97 ();
 FILLCELL_X32 FILLER_120_129 ();
 FILLCELL_X32 FILLER_120_161 ();
 FILLCELL_X32 FILLER_120_193 ();
 FILLCELL_X16 FILLER_120_225 ();
 FILLCELL_X4 FILLER_120_241 ();
 FILLCELL_X4 FILLER_120_248 ();
 FILLCELL_X4 FILLER_120_255 ();
 FILLCELL_X8 FILLER_120_264 ();
 FILLCELL_X1 FILLER_120_272 ();
 FILLCELL_X4 FILLER_120_278 ();
 FILLCELL_X4 FILLER_120_289 ();
 FILLCELL_X4 FILLER_120_297 ();
 FILLCELL_X4 FILLER_120_303 ();
 FILLCELL_X4 FILLER_120_311 ();
 FILLCELL_X4 FILLER_120_318 ();
 FILLCELL_X2 FILLER_120_322 ();
 FILLCELL_X1 FILLER_120_324 ();
 FILLCELL_X4 FILLER_120_330 ();
 FILLCELL_X4 FILLER_120_337 ();
 FILLCELL_X1 FILLER_120_341 ();
 FILLCELL_X4 FILLER_120_345 ();
 FILLCELL_X4 FILLER_120_355 ();
 FILLCELL_X8 FILLER_120_363 ();
 FILLCELL_X2 FILLER_120_371 ();
 FILLCELL_X4 FILLER_120_376 ();
 FILLCELL_X32 FILLER_120_1518 ();
 FILLCELL_X32 FILLER_120_1550 ();
 FILLCELL_X32 FILLER_120_1582 ();
 FILLCELL_X32 FILLER_120_1614 ();
 FILLCELL_X32 FILLER_120_1646 ();
 FILLCELL_X32 FILLER_120_1678 ();
 FILLCELL_X32 FILLER_120_1710 ();
 FILLCELL_X16 FILLER_120_1742 ();
 FILLCELL_X4 FILLER_120_1758 ();
 FILLCELL_X32 FILLER_121_1 ();
 FILLCELL_X32 FILLER_121_33 ();
 FILLCELL_X32 FILLER_121_65 ();
 FILLCELL_X32 FILLER_121_97 ();
 FILLCELL_X32 FILLER_121_129 ();
 FILLCELL_X32 FILLER_121_161 ();
 FILLCELL_X32 FILLER_121_193 ();
 FILLCELL_X16 FILLER_121_225 ();
 FILLCELL_X8 FILLER_121_241 ();
 FILLCELL_X2 FILLER_121_249 ();
 FILLCELL_X1 FILLER_121_251 ();
 FILLCELL_X4 FILLER_121_269 ();
 FILLCELL_X4 FILLER_121_278 ();
 FILLCELL_X8 FILLER_121_286 ();
 FILLCELL_X4 FILLER_121_298 ();
 FILLCELL_X4 FILLER_121_305 ();
 FILLCELL_X2 FILLER_121_309 ();
 FILLCELL_X1 FILLER_121_311 ();
 FILLCELL_X4 FILLER_121_315 ();
 FILLCELL_X4 FILLER_121_338 ();
 FILLCELL_X4 FILLER_121_345 ();
 FILLCELL_X2 FILLER_121_349 ();
 FILLCELL_X4 FILLER_121_368 ();
 FILLCELL_X1 FILLER_121_372 ();
 FILLCELL_X4 FILLER_121_376 ();
 FILLCELL_X32 FILLER_121_1518 ();
 FILLCELL_X32 FILLER_121_1550 ();
 FILLCELL_X32 FILLER_121_1582 ();
 FILLCELL_X32 FILLER_121_1614 ();
 FILLCELL_X32 FILLER_121_1646 ();
 FILLCELL_X32 FILLER_121_1678 ();
 FILLCELL_X32 FILLER_121_1710 ();
 FILLCELL_X16 FILLER_121_1742 ();
 FILLCELL_X4 FILLER_121_1758 ();
 FILLCELL_X4 FILLER_122_1 ();
 FILLCELL_X32 FILLER_122_8 ();
 FILLCELL_X32 FILLER_122_40 ();
 FILLCELL_X32 FILLER_122_72 ();
 FILLCELL_X32 FILLER_122_104 ();
 FILLCELL_X32 FILLER_122_136 ();
 FILLCELL_X32 FILLER_122_168 ();
 FILLCELL_X32 FILLER_122_200 ();
 FILLCELL_X16 FILLER_122_232 ();
 FILLCELL_X8 FILLER_122_248 ();
 FILLCELL_X1 FILLER_122_256 ();
 FILLCELL_X4 FILLER_122_260 ();
 FILLCELL_X4 FILLER_122_267 ();
 FILLCELL_X4 FILLER_122_274 ();
 FILLCELL_X4 FILLER_122_283 ();
 FILLCELL_X8 FILLER_122_292 ();
 FILLCELL_X1 FILLER_122_300 ();
 FILLCELL_X4 FILLER_122_306 ();
 FILLCELL_X4 FILLER_122_315 ();
 FILLCELL_X4 FILLER_122_323 ();
 FILLCELL_X1 FILLER_122_327 ();
 FILLCELL_X4 FILLER_122_332 ();
 FILLCELL_X8 FILLER_122_339 ();
 FILLCELL_X4 FILLER_122_350 ();
 FILLCELL_X2 FILLER_122_354 ();
 FILLCELL_X4 FILLER_122_359 ();
 FILLCELL_X1 FILLER_122_363 ();
 FILLCELL_X4 FILLER_122_367 ();
 FILLCELL_X4 FILLER_122_374 ();
 FILLCELL_X2 FILLER_122_378 ();
 FILLCELL_X32 FILLER_122_1518 ();
 FILLCELL_X32 FILLER_122_1550 ();
 FILLCELL_X32 FILLER_122_1582 ();
 FILLCELL_X32 FILLER_122_1614 ();
 FILLCELL_X32 FILLER_122_1646 ();
 FILLCELL_X32 FILLER_122_1678 ();
 FILLCELL_X32 FILLER_122_1710 ();
 FILLCELL_X16 FILLER_122_1742 ();
 FILLCELL_X4 FILLER_122_1758 ();
 FILLCELL_X32 FILLER_123_1 ();
 FILLCELL_X32 FILLER_123_33 ();
 FILLCELL_X32 FILLER_123_65 ();
 FILLCELL_X32 FILLER_123_97 ();
 FILLCELL_X32 FILLER_123_129 ();
 FILLCELL_X32 FILLER_123_161 ();
 FILLCELL_X32 FILLER_123_193 ();
 FILLCELL_X16 FILLER_123_225 ();
 FILLCELL_X8 FILLER_123_241 ();
 FILLCELL_X4 FILLER_123_249 ();
 FILLCELL_X2 FILLER_123_253 ();
 FILLCELL_X1 FILLER_123_255 ();
 FILLCELL_X4 FILLER_123_261 ();
 FILLCELL_X4 FILLER_123_268 ();
 FILLCELL_X4 FILLER_123_289 ();
 FILLCELL_X4 FILLER_123_310 ();
 FILLCELL_X4 FILLER_123_333 ();
 FILLCELL_X4 FILLER_123_344 ();
 FILLCELL_X4 FILLER_123_350 ();
 FILLCELL_X4 FILLER_123_357 ();
 FILLCELL_X8 FILLER_123_365 ();
 FILLCELL_X4 FILLER_123_376 ();
 FILLCELL_X32 FILLER_123_1518 ();
 FILLCELL_X32 FILLER_123_1550 ();
 FILLCELL_X32 FILLER_123_1582 ();
 FILLCELL_X32 FILLER_123_1614 ();
 FILLCELL_X32 FILLER_123_1646 ();
 FILLCELL_X32 FILLER_123_1678 ();
 FILLCELL_X32 FILLER_123_1710 ();
 FILLCELL_X16 FILLER_123_1742 ();
 FILLCELL_X4 FILLER_123_1758 ();
 FILLCELL_X32 FILLER_124_1 ();
 FILLCELL_X32 FILLER_124_33 ();
 FILLCELL_X32 FILLER_124_65 ();
 FILLCELL_X32 FILLER_124_97 ();
 FILLCELL_X32 FILLER_124_129 ();
 FILLCELL_X32 FILLER_124_161 ();
 FILLCELL_X32 FILLER_124_193 ();
 FILLCELL_X32 FILLER_124_225 ();
 FILLCELL_X8 FILLER_124_257 ();
 FILLCELL_X1 FILLER_124_265 ();
 FILLCELL_X8 FILLER_124_269 ();
 FILLCELL_X4 FILLER_124_277 ();
 FILLCELL_X1 FILLER_124_281 ();
 FILLCELL_X4 FILLER_124_285 ();
 FILLCELL_X4 FILLER_124_292 ();
 FILLCELL_X1 FILLER_124_296 ();
 FILLCELL_X4 FILLER_124_300 ();
 FILLCELL_X4 FILLER_124_307 ();
 FILLCELL_X8 FILLER_124_314 ();
 FILLCELL_X4 FILLER_124_322 ();
 FILLCELL_X2 FILLER_124_326 ();
 FILLCELL_X4 FILLER_124_333 ();
 FILLCELL_X4 FILLER_124_354 ();
 FILLCELL_X8 FILLER_124_364 ();
 FILLCELL_X1 FILLER_124_372 ();
 FILLCELL_X4 FILLER_124_376 ();
 FILLCELL_X32 FILLER_124_1518 ();
 FILLCELL_X32 FILLER_124_1550 ();
 FILLCELL_X32 FILLER_124_1582 ();
 FILLCELL_X32 FILLER_124_1614 ();
 FILLCELL_X32 FILLER_124_1646 ();
 FILLCELL_X32 FILLER_124_1678 ();
 FILLCELL_X32 FILLER_124_1710 ();
 FILLCELL_X16 FILLER_124_1742 ();
 FILLCELL_X4 FILLER_124_1758 ();
 FILLCELL_X32 FILLER_125_1 ();
 FILLCELL_X32 FILLER_125_33 ();
 FILLCELL_X32 FILLER_125_65 ();
 FILLCELL_X32 FILLER_125_97 ();
 FILLCELL_X32 FILLER_125_129 ();
 FILLCELL_X32 FILLER_125_161 ();
 FILLCELL_X32 FILLER_125_193 ();
 FILLCELL_X32 FILLER_125_225 ();
 FILLCELL_X16 FILLER_125_257 ();
 FILLCELL_X8 FILLER_125_273 ();
 FILLCELL_X4 FILLER_125_281 ();
 FILLCELL_X2 FILLER_125_285 ();
 FILLCELL_X16 FILLER_125_290 ();
 FILLCELL_X2 FILLER_125_306 ();
 FILLCELL_X32 FILLER_125_311 ();
 FILLCELL_X1 FILLER_125_343 ();
 FILLCELL_X4 FILLER_125_349 ();
 FILLCELL_X4 FILLER_125_359 ();
 FILLCELL_X4 FILLER_125_367 ();
 FILLCELL_X4 FILLER_125_374 ();
 FILLCELL_X2 FILLER_125_378 ();
 FILLCELL_X32 FILLER_125_1518 ();
 FILLCELL_X32 FILLER_125_1550 ();
 FILLCELL_X32 FILLER_125_1582 ();
 FILLCELL_X32 FILLER_125_1614 ();
 FILLCELL_X32 FILLER_125_1646 ();
 FILLCELL_X32 FILLER_125_1678 ();
 FILLCELL_X32 FILLER_125_1710 ();
 FILLCELL_X16 FILLER_125_1742 ();
 FILLCELL_X4 FILLER_125_1758 ();
 FILLCELL_X32 FILLER_126_1 ();
 FILLCELL_X32 FILLER_126_33 ();
 FILLCELL_X32 FILLER_126_65 ();
 FILLCELL_X32 FILLER_126_97 ();
 FILLCELL_X32 FILLER_126_129 ();
 FILLCELL_X32 FILLER_126_161 ();
 FILLCELL_X32 FILLER_126_193 ();
 FILLCELL_X32 FILLER_126_225 ();
 FILLCELL_X32 FILLER_126_257 ();
 FILLCELL_X32 FILLER_126_289 ();
 FILLCELL_X16 FILLER_126_321 ();
 FILLCELL_X2 FILLER_126_337 ();
 FILLCELL_X1 FILLER_126_339 ();
 FILLCELL_X4 FILLER_126_343 ();
 FILLCELL_X4 FILLER_126_364 ();
 FILLCELL_X8 FILLER_126_371 ();
 FILLCELL_X1 FILLER_126_379 ();
 FILLCELL_X32 FILLER_126_1518 ();
 FILLCELL_X32 FILLER_126_1550 ();
 FILLCELL_X32 FILLER_126_1582 ();
 FILLCELL_X32 FILLER_126_1614 ();
 FILLCELL_X32 FILLER_126_1646 ();
 FILLCELL_X32 FILLER_126_1678 ();
 FILLCELL_X32 FILLER_126_1710 ();
 FILLCELL_X8 FILLER_126_1742 ();
 FILLCELL_X2 FILLER_126_1750 ();
 FILLCELL_X1 FILLER_126_1752 ();
 FILLCELL_X4 FILLER_126_1758 ();
 FILLCELL_X32 FILLER_127_1 ();
 FILLCELL_X32 FILLER_127_33 ();
 FILLCELL_X32 FILLER_127_65 ();
 FILLCELL_X32 FILLER_127_97 ();
 FILLCELL_X32 FILLER_127_129 ();
 FILLCELL_X32 FILLER_127_161 ();
 FILLCELL_X32 FILLER_127_193 ();
 FILLCELL_X32 FILLER_127_225 ();
 FILLCELL_X32 FILLER_127_257 ();
 FILLCELL_X32 FILLER_127_289 ();
 FILLCELL_X16 FILLER_127_321 ();
 FILLCELL_X8 FILLER_127_337 ();
 FILLCELL_X2 FILLER_127_345 ();
 FILLCELL_X1 FILLER_127_347 ();
 FILLCELL_X4 FILLER_127_351 ();
 FILLCELL_X4 FILLER_127_360 ();
 FILLCELL_X2 FILLER_127_364 ();
 FILLCELL_X4 FILLER_127_369 ();
 FILLCELL_X4 FILLER_127_376 ();
 FILLCELL_X32 FILLER_127_1518 ();
 FILLCELL_X32 FILLER_127_1550 ();
 FILLCELL_X32 FILLER_127_1582 ();
 FILLCELL_X32 FILLER_127_1614 ();
 FILLCELL_X32 FILLER_127_1646 ();
 FILLCELL_X32 FILLER_127_1678 ();
 FILLCELL_X32 FILLER_127_1710 ();
 FILLCELL_X16 FILLER_127_1742 ();
 FILLCELL_X4 FILLER_127_1758 ();
 FILLCELL_X32 FILLER_128_1 ();
 FILLCELL_X32 FILLER_128_33 ();
 FILLCELL_X32 FILLER_128_65 ();
 FILLCELL_X32 FILLER_128_97 ();
 FILLCELL_X32 FILLER_128_129 ();
 FILLCELL_X32 FILLER_128_161 ();
 FILLCELL_X32 FILLER_128_193 ();
 FILLCELL_X32 FILLER_128_225 ();
 FILLCELL_X32 FILLER_128_257 ();
 FILLCELL_X32 FILLER_128_289 ();
 FILLCELL_X32 FILLER_128_321 ();
 FILLCELL_X16 FILLER_128_353 ();
 FILLCELL_X4 FILLER_128_369 ();
 FILLCELL_X4 FILLER_128_376 ();
 FILLCELL_X32 FILLER_128_1518 ();
 FILLCELL_X32 FILLER_128_1550 ();
 FILLCELL_X32 FILLER_128_1582 ();
 FILLCELL_X32 FILLER_128_1614 ();
 FILLCELL_X32 FILLER_128_1646 ();
 FILLCELL_X32 FILLER_128_1678 ();
 FILLCELL_X32 FILLER_128_1710 ();
 FILLCELL_X16 FILLER_128_1742 ();
 FILLCELL_X4 FILLER_128_1758 ();
 FILLCELL_X32 FILLER_129_1 ();
 FILLCELL_X32 FILLER_129_33 ();
 FILLCELL_X32 FILLER_129_65 ();
 FILLCELL_X32 FILLER_129_97 ();
 FILLCELL_X32 FILLER_129_129 ();
 FILLCELL_X32 FILLER_129_161 ();
 FILLCELL_X32 FILLER_129_193 ();
 FILLCELL_X32 FILLER_129_225 ();
 FILLCELL_X32 FILLER_129_257 ();
 FILLCELL_X32 FILLER_129_289 ();
 FILLCELL_X32 FILLER_129_321 ();
 FILLCELL_X16 FILLER_129_353 ();
 FILLCELL_X8 FILLER_129_369 ();
 FILLCELL_X2 FILLER_129_377 ();
 FILLCELL_X1 FILLER_129_379 ();
 FILLCELL_X32 FILLER_129_1518 ();
 FILLCELL_X32 FILLER_129_1550 ();
 FILLCELL_X32 FILLER_129_1582 ();
 FILLCELL_X32 FILLER_129_1614 ();
 FILLCELL_X32 FILLER_129_1646 ();
 FILLCELL_X32 FILLER_129_1678 ();
 FILLCELL_X32 FILLER_129_1710 ();
 FILLCELL_X16 FILLER_129_1742 ();
 FILLCELL_X4 FILLER_129_1758 ();
 FILLCELL_X32 FILLER_130_1 ();
 FILLCELL_X32 FILLER_130_33 ();
 FILLCELL_X32 FILLER_130_65 ();
 FILLCELL_X32 FILLER_130_97 ();
 FILLCELL_X32 FILLER_130_129 ();
 FILLCELL_X32 FILLER_130_161 ();
 FILLCELL_X32 FILLER_130_193 ();
 FILLCELL_X32 FILLER_130_225 ();
 FILLCELL_X32 FILLER_130_257 ();
 FILLCELL_X32 FILLER_130_289 ();
 FILLCELL_X32 FILLER_130_321 ();
 FILLCELL_X16 FILLER_130_353 ();
 FILLCELL_X8 FILLER_130_369 ();
 FILLCELL_X2 FILLER_130_377 ();
 FILLCELL_X1 FILLER_130_379 ();
 FILLCELL_X32 FILLER_130_1518 ();
 FILLCELL_X32 FILLER_130_1550 ();
 FILLCELL_X32 FILLER_130_1582 ();
 FILLCELL_X32 FILLER_130_1614 ();
 FILLCELL_X32 FILLER_130_1646 ();
 FILLCELL_X32 FILLER_130_1678 ();
 FILLCELL_X32 FILLER_130_1710 ();
 FILLCELL_X16 FILLER_130_1742 ();
 FILLCELL_X4 FILLER_130_1758 ();
 FILLCELL_X4 FILLER_131_1 ();
 FILLCELL_X32 FILLER_131_8 ();
 FILLCELL_X32 FILLER_131_40 ();
 FILLCELL_X32 FILLER_131_72 ();
 FILLCELL_X32 FILLER_131_104 ();
 FILLCELL_X32 FILLER_131_136 ();
 FILLCELL_X32 FILLER_131_168 ();
 FILLCELL_X32 FILLER_131_200 ();
 FILLCELL_X32 FILLER_131_232 ();
 FILLCELL_X32 FILLER_131_264 ();
 FILLCELL_X32 FILLER_131_296 ();
 FILLCELL_X32 FILLER_131_328 ();
 FILLCELL_X16 FILLER_131_360 ();
 FILLCELL_X4 FILLER_131_376 ();
 FILLCELL_X32 FILLER_131_1518 ();
 FILLCELL_X32 FILLER_131_1550 ();
 FILLCELL_X32 FILLER_131_1582 ();
 FILLCELL_X32 FILLER_131_1614 ();
 FILLCELL_X32 FILLER_131_1646 ();
 FILLCELL_X32 FILLER_131_1678 ();
 FILLCELL_X32 FILLER_131_1710 ();
 FILLCELL_X16 FILLER_131_1742 ();
 FILLCELL_X4 FILLER_131_1758 ();
 FILLCELL_X32 FILLER_132_1 ();
 FILLCELL_X32 FILLER_132_33 ();
 FILLCELL_X32 FILLER_132_65 ();
 FILLCELL_X32 FILLER_132_97 ();
 FILLCELL_X32 FILLER_132_129 ();
 FILLCELL_X32 FILLER_132_161 ();
 FILLCELL_X32 FILLER_132_193 ();
 FILLCELL_X32 FILLER_132_225 ();
 FILLCELL_X32 FILLER_132_257 ();
 FILLCELL_X32 FILLER_132_289 ();
 FILLCELL_X32 FILLER_132_321 ();
 FILLCELL_X16 FILLER_132_353 ();
 FILLCELL_X8 FILLER_132_369 ();
 FILLCELL_X2 FILLER_132_377 ();
 FILLCELL_X1 FILLER_132_379 ();
 FILLCELL_X32 FILLER_132_1518 ();
 FILLCELL_X32 FILLER_132_1550 ();
 FILLCELL_X32 FILLER_132_1582 ();
 FILLCELL_X32 FILLER_132_1614 ();
 FILLCELL_X32 FILLER_132_1646 ();
 FILLCELL_X32 FILLER_132_1678 ();
 FILLCELL_X32 FILLER_132_1710 ();
 FILLCELL_X16 FILLER_132_1742 ();
 FILLCELL_X4 FILLER_132_1758 ();
 FILLCELL_X32 FILLER_133_1 ();
 FILLCELL_X32 FILLER_133_33 ();
 FILLCELL_X32 FILLER_133_65 ();
 FILLCELL_X32 FILLER_133_97 ();
 FILLCELL_X32 FILLER_133_129 ();
 FILLCELL_X32 FILLER_133_161 ();
 FILLCELL_X32 FILLER_133_193 ();
 FILLCELL_X32 FILLER_133_225 ();
 FILLCELL_X32 FILLER_133_257 ();
 FILLCELL_X32 FILLER_133_289 ();
 FILLCELL_X32 FILLER_133_321 ();
 FILLCELL_X16 FILLER_133_353 ();
 FILLCELL_X8 FILLER_133_369 ();
 FILLCELL_X2 FILLER_133_377 ();
 FILLCELL_X1 FILLER_133_379 ();
 FILLCELL_X32 FILLER_133_1518 ();
 FILLCELL_X32 FILLER_133_1550 ();
 FILLCELL_X32 FILLER_133_1582 ();
 FILLCELL_X32 FILLER_133_1614 ();
 FILLCELL_X32 FILLER_133_1646 ();
 FILLCELL_X32 FILLER_133_1678 ();
 FILLCELL_X32 FILLER_133_1710 ();
 FILLCELL_X16 FILLER_133_1742 ();
 FILLCELL_X4 FILLER_133_1758 ();
 FILLCELL_X32 FILLER_134_1 ();
 FILLCELL_X32 FILLER_134_33 ();
 FILLCELL_X32 FILLER_134_65 ();
 FILLCELL_X32 FILLER_134_97 ();
 FILLCELL_X32 FILLER_134_129 ();
 FILLCELL_X32 FILLER_134_161 ();
 FILLCELL_X32 FILLER_134_193 ();
 FILLCELL_X32 FILLER_134_225 ();
 FILLCELL_X32 FILLER_134_257 ();
 FILLCELL_X32 FILLER_134_289 ();
 FILLCELL_X32 FILLER_134_321 ();
 FILLCELL_X16 FILLER_134_353 ();
 FILLCELL_X8 FILLER_134_369 ();
 FILLCELL_X2 FILLER_134_377 ();
 FILLCELL_X1 FILLER_134_379 ();
 FILLCELL_X32 FILLER_134_1518 ();
 FILLCELL_X32 FILLER_134_1550 ();
 FILLCELL_X32 FILLER_134_1582 ();
 FILLCELL_X32 FILLER_134_1614 ();
 FILLCELL_X32 FILLER_134_1646 ();
 FILLCELL_X32 FILLER_134_1678 ();
 FILLCELL_X32 FILLER_134_1710 ();
 FILLCELL_X16 FILLER_134_1742 ();
 FILLCELL_X4 FILLER_134_1758 ();
 FILLCELL_X32 FILLER_135_1 ();
 FILLCELL_X32 FILLER_135_33 ();
 FILLCELL_X32 FILLER_135_65 ();
 FILLCELL_X32 FILLER_135_97 ();
 FILLCELL_X32 FILLER_135_129 ();
 FILLCELL_X32 FILLER_135_161 ();
 FILLCELL_X32 FILLER_135_193 ();
 FILLCELL_X32 FILLER_135_225 ();
 FILLCELL_X32 FILLER_135_257 ();
 FILLCELL_X32 FILLER_135_289 ();
 FILLCELL_X32 FILLER_135_321 ();
 FILLCELL_X16 FILLER_135_353 ();
 FILLCELL_X8 FILLER_135_369 ();
 FILLCELL_X2 FILLER_135_377 ();
 FILLCELL_X1 FILLER_135_379 ();
 FILLCELL_X32 FILLER_135_1518 ();
 FILLCELL_X32 FILLER_135_1550 ();
 FILLCELL_X32 FILLER_135_1582 ();
 FILLCELL_X32 FILLER_135_1614 ();
 FILLCELL_X32 FILLER_135_1646 ();
 FILLCELL_X32 FILLER_135_1678 ();
 FILLCELL_X32 FILLER_135_1710 ();
 FILLCELL_X16 FILLER_135_1742 ();
 FILLCELL_X4 FILLER_135_1758 ();
 FILLCELL_X32 FILLER_136_1 ();
 FILLCELL_X32 FILLER_136_33 ();
 FILLCELL_X32 FILLER_136_65 ();
 FILLCELL_X32 FILLER_136_97 ();
 FILLCELL_X32 FILLER_136_129 ();
 FILLCELL_X32 FILLER_136_161 ();
 FILLCELL_X32 FILLER_136_193 ();
 FILLCELL_X32 FILLER_136_225 ();
 FILLCELL_X32 FILLER_136_257 ();
 FILLCELL_X32 FILLER_136_289 ();
 FILLCELL_X32 FILLER_136_321 ();
 FILLCELL_X16 FILLER_136_353 ();
 FILLCELL_X8 FILLER_136_369 ();
 FILLCELL_X2 FILLER_136_377 ();
 FILLCELL_X1 FILLER_136_379 ();
 FILLCELL_X32 FILLER_136_1518 ();
 FILLCELL_X32 FILLER_136_1550 ();
 FILLCELL_X32 FILLER_136_1582 ();
 FILLCELL_X32 FILLER_136_1614 ();
 FILLCELL_X32 FILLER_136_1646 ();
 FILLCELL_X32 FILLER_136_1678 ();
 FILLCELL_X32 FILLER_136_1710 ();
 FILLCELL_X8 FILLER_136_1742 ();
 FILLCELL_X4 FILLER_136_1750 ();
 FILLCELL_X1 FILLER_136_1754 ();
 FILLCELL_X4 FILLER_136_1758 ();
 FILLCELL_X32 FILLER_137_1 ();
 FILLCELL_X32 FILLER_137_33 ();
 FILLCELL_X32 FILLER_137_65 ();
 FILLCELL_X32 FILLER_137_97 ();
 FILLCELL_X32 FILLER_137_129 ();
 FILLCELL_X32 FILLER_137_161 ();
 FILLCELL_X32 FILLER_137_193 ();
 FILLCELL_X32 FILLER_137_225 ();
 FILLCELL_X32 FILLER_137_257 ();
 FILLCELL_X32 FILLER_137_289 ();
 FILLCELL_X32 FILLER_137_321 ();
 FILLCELL_X16 FILLER_137_353 ();
 FILLCELL_X8 FILLER_137_369 ();
 FILLCELL_X2 FILLER_137_377 ();
 FILLCELL_X1 FILLER_137_379 ();
 FILLCELL_X32 FILLER_137_1518 ();
 FILLCELL_X32 FILLER_137_1550 ();
 FILLCELL_X32 FILLER_137_1582 ();
 FILLCELL_X32 FILLER_137_1614 ();
 FILLCELL_X32 FILLER_137_1646 ();
 FILLCELL_X32 FILLER_137_1678 ();
 FILLCELL_X32 FILLER_137_1710 ();
 FILLCELL_X16 FILLER_137_1742 ();
 FILLCELL_X4 FILLER_137_1758 ();
 FILLCELL_X32 FILLER_138_1 ();
 FILLCELL_X32 FILLER_138_33 ();
 FILLCELL_X32 FILLER_138_65 ();
 FILLCELL_X32 FILLER_138_97 ();
 FILLCELL_X32 FILLER_138_129 ();
 FILLCELL_X32 FILLER_138_161 ();
 FILLCELL_X32 FILLER_138_193 ();
 FILLCELL_X32 FILLER_138_225 ();
 FILLCELL_X32 FILLER_138_257 ();
 FILLCELL_X32 FILLER_138_289 ();
 FILLCELL_X32 FILLER_138_321 ();
 FILLCELL_X16 FILLER_138_353 ();
 FILLCELL_X8 FILLER_138_369 ();
 FILLCELL_X2 FILLER_138_377 ();
 FILLCELL_X1 FILLER_138_379 ();
 FILLCELL_X32 FILLER_138_1518 ();
 FILLCELL_X32 FILLER_138_1550 ();
 FILLCELL_X32 FILLER_138_1582 ();
 FILLCELL_X32 FILLER_138_1614 ();
 FILLCELL_X32 FILLER_138_1646 ();
 FILLCELL_X32 FILLER_138_1678 ();
 FILLCELL_X32 FILLER_138_1710 ();
 FILLCELL_X16 FILLER_138_1742 ();
 FILLCELL_X4 FILLER_138_1758 ();
 FILLCELL_X32 FILLER_139_1 ();
 FILLCELL_X32 FILLER_139_33 ();
 FILLCELL_X32 FILLER_139_65 ();
 FILLCELL_X32 FILLER_139_97 ();
 FILLCELL_X32 FILLER_139_129 ();
 FILLCELL_X32 FILLER_139_161 ();
 FILLCELL_X32 FILLER_139_193 ();
 FILLCELL_X32 FILLER_139_225 ();
 FILLCELL_X32 FILLER_139_257 ();
 FILLCELL_X32 FILLER_139_289 ();
 FILLCELL_X32 FILLER_139_321 ();
 FILLCELL_X16 FILLER_139_353 ();
 FILLCELL_X8 FILLER_139_369 ();
 FILLCELL_X2 FILLER_139_377 ();
 FILLCELL_X1 FILLER_139_379 ();
 FILLCELL_X32 FILLER_139_1518 ();
 FILLCELL_X32 FILLER_139_1550 ();
 FILLCELL_X32 FILLER_139_1582 ();
 FILLCELL_X32 FILLER_139_1614 ();
 FILLCELL_X32 FILLER_139_1646 ();
 FILLCELL_X32 FILLER_139_1678 ();
 FILLCELL_X32 FILLER_139_1710 ();
 FILLCELL_X16 FILLER_139_1742 ();
 FILLCELL_X4 FILLER_139_1758 ();
 FILLCELL_X32 FILLER_140_1 ();
 FILLCELL_X32 FILLER_140_33 ();
 FILLCELL_X32 FILLER_140_65 ();
 FILLCELL_X32 FILLER_140_97 ();
 FILLCELL_X32 FILLER_140_129 ();
 FILLCELL_X32 FILLER_140_161 ();
 FILLCELL_X32 FILLER_140_193 ();
 FILLCELL_X32 FILLER_140_225 ();
 FILLCELL_X32 FILLER_140_257 ();
 FILLCELL_X32 FILLER_140_289 ();
 FILLCELL_X32 FILLER_140_321 ();
 FILLCELL_X16 FILLER_140_353 ();
 FILLCELL_X8 FILLER_140_369 ();
 FILLCELL_X2 FILLER_140_377 ();
 FILLCELL_X1 FILLER_140_379 ();
 FILLCELL_X32 FILLER_140_1518 ();
 FILLCELL_X32 FILLER_140_1550 ();
 FILLCELL_X32 FILLER_140_1582 ();
 FILLCELL_X32 FILLER_140_1614 ();
 FILLCELL_X32 FILLER_140_1646 ();
 FILLCELL_X32 FILLER_140_1678 ();
 FILLCELL_X32 FILLER_140_1710 ();
 FILLCELL_X16 FILLER_140_1742 ();
 FILLCELL_X4 FILLER_140_1758 ();
 FILLCELL_X4 FILLER_141_1 ();
 FILLCELL_X32 FILLER_141_8 ();
 FILLCELL_X32 FILLER_141_40 ();
 FILLCELL_X32 FILLER_141_72 ();
 FILLCELL_X32 FILLER_141_104 ();
 FILLCELL_X32 FILLER_141_136 ();
 FILLCELL_X32 FILLER_141_168 ();
 FILLCELL_X32 FILLER_141_200 ();
 FILLCELL_X32 FILLER_141_232 ();
 FILLCELL_X32 FILLER_141_264 ();
 FILLCELL_X32 FILLER_141_296 ();
 FILLCELL_X32 FILLER_141_328 ();
 FILLCELL_X16 FILLER_141_360 ();
 FILLCELL_X4 FILLER_141_376 ();
 FILLCELL_X32 FILLER_141_1518 ();
 FILLCELL_X32 FILLER_141_1550 ();
 FILLCELL_X32 FILLER_141_1582 ();
 FILLCELL_X32 FILLER_141_1614 ();
 FILLCELL_X32 FILLER_141_1646 ();
 FILLCELL_X32 FILLER_141_1678 ();
 FILLCELL_X32 FILLER_141_1710 ();
 FILLCELL_X16 FILLER_141_1742 ();
 FILLCELL_X4 FILLER_141_1758 ();
 FILLCELL_X32 FILLER_142_1 ();
 FILLCELL_X32 FILLER_142_33 ();
 FILLCELL_X32 FILLER_142_65 ();
 FILLCELL_X32 FILLER_142_97 ();
 FILLCELL_X32 FILLER_142_129 ();
 FILLCELL_X32 FILLER_142_161 ();
 FILLCELL_X32 FILLER_142_193 ();
 FILLCELL_X32 FILLER_142_225 ();
 FILLCELL_X32 FILLER_142_257 ();
 FILLCELL_X32 FILLER_142_289 ();
 FILLCELL_X32 FILLER_142_321 ();
 FILLCELL_X16 FILLER_142_353 ();
 FILLCELL_X8 FILLER_142_369 ();
 FILLCELL_X2 FILLER_142_377 ();
 FILLCELL_X1 FILLER_142_379 ();
 FILLCELL_X32 FILLER_142_1518 ();
 FILLCELL_X32 FILLER_142_1550 ();
 FILLCELL_X32 FILLER_142_1582 ();
 FILLCELL_X32 FILLER_142_1614 ();
 FILLCELL_X32 FILLER_142_1646 ();
 FILLCELL_X32 FILLER_142_1678 ();
 FILLCELL_X32 FILLER_142_1710 ();
 FILLCELL_X16 FILLER_142_1742 ();
 FILLCELL_X4 FILLER_142_1758 ();
 FILLCELL_X32 FILLER_143_1 ();
 FILLCELL_X32 FILLER_143_33 ();
 FILLCELL_X32 FILLER_143_65 ();
 FILLCELL_X32 FILLER_143_97 ();
 FILLCELL_X32 FILLER_143_129 ();
 FILLCELL_X32 FILLER_143_161 ();
 FILLCELL_X32 FILLER_143_193 ();
 FILLCELL_X32 FILLER_143_225 ();
 FILLCELL_X32 FILLER_143_257 ();
 FILLCELL_X32 FILLER_143_289 ();
 FILLCELL_X32 FILLER_143_321 ();
 FILLCELL_X16 FILLER_143_353 ();
 FILLCELL_X8 FILLER_143_369 ();
 FILLCELL_X2 FILLER_143_377 ();
 FILLCELL_X1 FILLER_143_379 ();
 FILLCELL_X32 FILLER_143_1518 ();
 FILLCELL_X32 FILLER_143_1550 ();
 FILLCELL_X32 FILLER_143_1582 ();
 FILLCELL_X32 FILLER_143_1614 ();
 FILLCELL_X32 FILLER_143_1646 ();
 FILLCELL_X32 FILLER_143_1678 ();
 FILLCELL_X32 FILLER_143_1710 ();
 FILLCELL_X16 FILLER_143_1742 ();
 FILLCELL_X4 FILLER_143_1758 ();
 FILLCELL_X32 FILLER_144_1 ();
 FILLCELL_X32 FILLER_144_33 ();
 FILLCELL_X32 FILLER_144_65 ();
 FILLCELL_X32 FILLER_144_97 ();
 FILLCELL_X32 FILLER_144_129 ();
 FILLCELL_X32 FILLER_144_161 ();
 FILLCELL_X32 FILLER_144_193 ();
 FILLCELL_X32 FILLER_144_225 ();
 FILLCELL_X32 FILLER_144_257 ();
 FILLCELL_X32 FILLER_144_289 ();
 FILLCELL_X32 FILLER_144_321 ();
 FILLCELL_X16 FILLER_144_353 ();
 FILLCELL_X8 FILLER_144_369 ();
 FILLCELL_X2 FILLER_144_377 ();
 FILLCELL_X1 FILLER_144_379 ();
 FILLCELL_X32 FILLER_144_1518 ();
 FILLCELL_X32 FILLER_144_1550 ();
 FILLCELL_X32 FILLER_144_1582 ();
 FILLCELL_X32 FILLER_144_1614 ();
 FILLCELL_X32 FILLER_144_1646 ();
 FILLCELL_X32 FILLER_144_1678 ();
 FILLCELL_X32 FILLER_144_1710 ();
 FILLCELL_X16 FILLER_144_1742 ();
 FILLCELL_X4 FILLER_144_1758 ();
 FILLCELL_X32 FILLER_145_1 ();
 FILLCELL_X32 FILLER_145_33 ();
 FILLCELL_X32 FILLER_145_65 ();
 FILLCELL_X32 FILLER_145_97 ();
 FILLCELL_X32 FILLER_145_129 ();
 FILLCELL_X32 FILLER_145_161 ();
 FILLCELL_X32 FILLER_145_193 ();
 FILLCELL_X32 FILLER_145_225 ();
 FILLCELL_X32 FILLER_145_257 ();
 FILLCELL_X32 FILLER_145_289 ();
 FILLCELL_X32 FILLER_145_321 ();
 FILLCELL_X16 FILLER_145_353 ();
 FILLCELL_X8 FILLER_145_369 ();
 FILLCELL_X2 FILLER_145_377 ();
 FILLCELL_X1 FILLER_145_379 ();
 FILLCELL_X32 FILLER_145_1518 ();
 FILLCELL_X32 FILLER_145_1550 ();
 FILLCELL_X32 FILLER_145_1582 ();
 FILLCELL_X32 FILLER_145_1614 ();
 FILLCELL_X32 FILLER_145_1646 ();
 FILLCELL_X32 FILLER_145_1678 ();
 FILLCELL_X32 FILLER_145_1710 ();
 FILLCELL_X16 FILLER_145_1742 ();
 FILLCELL_X4 FILLER_145_1758 ();
 FILLCELL_X32 FILLER_146_1 ();
 FILLCELL_X32 FILLER_146_33 ();
 FILLCELL_X32 FILLER_146_65 ();
 FILLCELL_X32 FILLER_146_97 ();
 FILLCELL_X32 FILLER_146_129 ();
 FILLCELL_X32 FILLER_146_161 ();
 FILLCELL_X32 FILLER_146_193 ();
 FILLCELL_X32 FILLER_146_225 ();
 FILLCELL_X32 FILLER_146_257 ();
 FILLCELL_X32 FILLER_146_289 ();
 FILLCELL_X32 FILLER_146_321 ();
 FILLCELL_X16 FILLER_146_353 ();
 FILLCELL_X8 FILLER_146_369 ();
 FILLCELL_X2 FILLER_146_377 ();
 FILLCELL_X1 FILLER_146_379 ();
 FILLCELL_X32 FILLER_146_1518 ();
 FILLCELL_X32 FILLER_146_1550 ();
 FILLCELL_X32 FILLER_146_1582 ();
 FILLCELL_X32 FILLER_146_1614 ();
 FILLCELL_X32 FILLER_146_1646 ();
 FILLCELL_X32 FILLER_146_1678 ();
 FILLCELL_X32 FILLER_146_1710 ();
 FILLCELL_X8 FILLER_146_1742 ();
 FILLCELL_X4 FILLER_146_1750 ();
 FILLCELL_X1 FILLER_146_1754 ();
 FILLCELL_X4 FILLER_146_1758 ();
 FILLCELL_X32 FILLER_147_1 ();
 FILLCELL_X32 FILLER_147_33 ();
 FILLCELL_X32 FILLER_147_65 ();
 FILLCELL_X32 FILLER_147_97 ();
 FILLCELL_X32 FILLER_147_129 ();
 FILLCELL_X32 FILLER_147_161 ();
 FILLCELL_X32 FILLER_147_193 ();
 FILLCELL_X32 FILLER_147_225 ();
 FILLCELL_X32 FILLER_147_257 ();
 FILLCELL_X32 FILLER_147_289 ();
 FILLCELL_X32 FILLER_147_321 ();
 FILLCELL_X16 FILLER_147_353 ();
 FILLCELL_X8 FILLER_147_369 ();
 FILLCELL_X2 FILLER_147_377 ();
 FILLCELL_X1 FILLER_147_379 ();
 FILLCELL_X32 FILLER_147_1518 ();
 FILLCELL_X32 FILLER_147_1550 ();
 FILLCELL_X32 FILLER_147_1582 ();
 FILLCELL_X32 FILLER_147_1614 ();
 FILLCELL_X32 FILLER_147_1646 ();
 FILLCELL_X32 FILLER_147_1678 ();
 FILLCELL_X32 FILLER_147_1710 ();
 FILLCELL_X16 FILLER_147_1742 ();
 FILLCELL_X4 FILLER_147_1758 ();
 FILLCELL_X32 FILLER_148_1 ();
 FILLCELL_X32 FILLER_148_33 ();
 FILLCELL_X32 FILLER_148_65 ();
 FILLCELL_X32 FILLER_148_97 ();
 FILLCELL_X32 FILLER_148_129 ();
 FILLCELL_X32 FILLER_148_161 ();
 FILLCELL_X32 FILLER_148_193 ();
 FILLCELL_X32 FILLER_148_225 ();
 FILLCELL_X32 FILLER_148_257 ();
 FILLCELL_X32 FILLER_148_289 ();
 FILLCELL_X32 FILLER_148_321 ();
 FILLCELL_X16 FILLER_148_353 ();
 FILLCELL_X8 FILLER_148_369 ();
 FILLCELL_X2 FILLER_148_377 ();
 FILLCELL_X1 FILLER_148_379 ();
 FILLCELL_X32 FILLER_148_1518 ();
 FILLCELL_X32 FILLER_148_1550 ();
 FILLCELL_X32 FILLER_148_1582 ();
 FILLCELL_X32 FILLER_148_1614 ();
 FILLCELL_X32 FILLER_148_1646 ();
 FILLCELL_X32 FILLER_148_1678 ();
 FILLCELL_X32 FILLER_148_1710 ();
 FILLCELL_X16 FILLER_148_1742 ();
 FILLCELL_X4 FILLER_148_1758 ();
 FILLCELL_X32 FILLER_149_1 ();
 FILLCELL_X32 FILLER_149_33 ();
 FILLCELL_X32 FILLER_149_65 ();
 FILLCELL_X32 FILLER_149_97 ();
 FILLCELL_X32 FILLER_149_129 ();
 FILLCELL_X32 FILLER_149_161 ();
 FILLCELL_X32 FILLER_149_193 ();
 FILLCELL_X32 FILLER_149_225 ();
 FILLCELL_X32 FILLER_149_257 ();
 FILLCELL_X32 FILLER_149_289 ();
 FILLCELL_X32 FILLER_149_321 ();
 FILLCELL_X16 FILLER_149_353 ();
 FILLCELL_X8 FILLER_149_369 ();
 FILLCELL_X2 FILLER_149_377 ();
 FILLCELL_X1 FILLER_149_379 ();
 FILLCELL_X32 FILLER_149_1518 ();
 FILLCELL_X32 FILLER_149_1550 ();
 FILLCELL_X32 FILLER_149_1582 ();
 FILLCELL_X32 FILLER_149_1614 ();
 FILLCELL_X32 FILLER_149_1646 ();
 FILLCELL_X32 FILLER_149_1678 ();
 FILLCELL_X32 FILLER_149_1710 ();
 FILLCELL_X16 FILLER_149_1742 ();
 FILLCELL_X4 FILLER_149_1758 ();
 FILLCELL_X4 FILLER_150_1 ();
 FILLCELL_X32 FILLER_150_9 ();
 FILLCELL_X32 FILLER_150_41 ();
 FILLCELL_X32 FILLER_150_73 ();
 FILLCELL_X32 FILLER_150_105 ();
 FILLCELL_X32 FILLER_150_137 ();
 FILLCELL_X32 FILLER_150_169 ();
 FILLCELL_X32 FILLER_150_201 ();
 FILLCELL_X32 FILLER_150_233 ();
 FILLCELL_X32 FILLER_150_265 ();
 FILLCELL_X32 FILLER_150_297 ();
 FILLCELL_X32 FILLER_150_329 ();
 FILLCELL_X16 FILLER_150_361 ();
 FILLCELL_X2 FILLER_150_377 ();
 FILLCELL_X1 FILLER_150_379 ();
 FILLCELL_X32 FILLER_150_1518 ();
 FILLCELL_X32 FILLER_150_1550 ();
 FILLCELL_X32 FILLER_150_1582 ();
 FILLCELL_X32 FILLER_150_1614 ();
 FILLCELL_X32 FILLER_150_1646 ();
 FILLCELL_X32 FILLER_150_1678 ();
 FILLCELL_X32 FILLER_150_1710 ();
 FILLCELL_X16 FILLER_150_1742 ();
 FILLCELL_X4 FILLER_150_1758 ();
 FILLCELL_X32 FILLER_151_1 ();
 FILLCELL_X32 FILLER_151_33 ();
 FILLCELL_X32 FILLER_151_65 ();
 FILLCELL_X32 FILLER_151_97 ();
 FILLCELL_X32 FILLER_151_129 ();
 FILLCELL_X32 FILLER_151_161 ();
 FILLCELL_X32 FILLER_151_193 ();
 FILLCELL_X32 FILLER_151_225 ();
 FILLCELL_X32 FILLER_151_257 ();
 FILLCELL_X32 FILLER_151_289 ();
 FILLCELL_X32 FILLER_151_321 ();
 FILLCELL_X16 FILLER_151_353 ();
 FILLCELL_X8 FILLER_151_369 ();
 FILLCELL_X2 FILLER_151_377 ();
 FILLCELL_X1 FILLER_151_379 ();
 FILLCELL_X32 FILLER_151_1518 ();
 FILLCELL_X32 FILLER_151_1550 ();
 FILLCELL_X32 FILLER_151_1582 ();
 FILLCELL_X32 FILLER_151_1614 ();
 FILLCELL_X32 FILLER_151_1646 ();
 FILLCELL_X32 FILLER_151_1678 ();
 FILLCELL_X32 FILLER_151_1710 ();
 FILLCELL_X16 FILLER_151_1742 ();
 FILLCELL_X4 FILLER_151_1758 ();
 FILLCELL_X32 FILLER_152_1 ();
 FILLCELL_X32 FILLER_152_33 ();
 FILLCELL_X32 FILLER_152_65 ();
 FILLCELL_X32 FILLER_152_97 ();
 FILLCELL_X32 FILLER_152_129 ();
 FILLCELL_X32 FILLER_152_161 ();
 FILLCELL_X32 FILLER_152_193 ();
 FILLCELL_X32 FILLER_152_225 ();
 FILLCELL_X32 FILLER_152_257 ();
 FILLCELL_X32 FILLER_152_289 ();
 FILLCELL_X32 FILLER_152_321 ();
 FILLCELL_X16 FILLER_152_353 ();
 FILLCELL_X8 FILLER_152_369 ();
 FILLCELL_X2 FILLER_152_377 ();
 FILLCELL_X1 FILLER_152_379 ();
 FILLCELL_X32 FILLER_152_1518 ();
 FILLCELL_X32 FILLER_152_1550 ();
 FILLCELL_X32 FILLER_152_1582 ();
 FILLCELL_X32 FILLER_152_1614 ();
 FILLCELL_X32 FILLER_152_1646 ();
 FILLCELL_X32 FILLER_152_1678 ();
 FILLCELL_X32 FILLER_152_1710 ();
 FILLCELL_X16 FILLER_152_1742 ();
 FILLCELL_X4 FILLER_152_1758 ();
 FILLCELL_X32 FILLER_153_1 ();
 FILLCELL_X32 FILLER_153_33 ();
 FILLCELL_X32 FILLER_153_65 ();
 FILLCELL_X32 FILLER_153_97 ();
 FILLCELL_X32 FILLER_153_129 ();
 FILLCELL_X32 FILLER_153_161 ();
 FILLCELL_X32 FILLER_153_193 ();
 FILLCELL_X32 FILLER_153_225 ();
 FILLCELL_X32 FILLER_153_257 ();
 FILLCELL_X32 FILLER_153_289 ();
 FILLCELL_X32 FILLER_153_321 ();
 FILLCELL_X16 FILLER_153_353 ();
 FILLCELL_X8 FILLER_153_369 ();
 FILLCELL_X2 FILLER_153_377 ();
 FILLCELL_X1 FILLER_153_379 ();
 FILLCELL_X32 FILLER_153_1518 ();
 FILLCELL_X32 FILLER_153_1550 ();
 FILLCELL_X32 FILLER_153_1582 ();
 FILLCELL_X32 FILLER_153_1614 ();
 FILLCELL_X32 FILLER_153_1646 ();
 FILLCELL_X32 FILLER_153_1678 ();
 FILLCELL_X32 FILLER_153_1710 ();
 FILLCELL_X16 FILLER_153_1742 ();
 FILLCELL_X4 FILLER_153_1758 ();
 FILLCELL_X32 FILLER_154_1 ();
 FILLCELL_X32 FILLER_154_33 ();
 FILLCELL_X32 FILLER_154_65 ();
 FILLCELL_X32 FILLER_154_97 ();
 FILLCELL_X32 FILLER_154_129 ();
 FILLCELL_X32 FILLER_154_161 ();
 FILLCELL_X32 FILLER_154_193 ();
 FILLCELL_X32 FILLER_154_225 ();
 FILLCELL_X32 FILLER_154_257 ();
 FILLCELL_X32 FILLER_154_289 ();
 FILLCELL_X32 FILLER_154_321 ();
 FILLCELL_X16 FILLER_154_353 ();
 FILLCELL_X8 FILLER_154_369 ();
 FILLCELL_X2 FILLER_154_377 ();
 FILLCELL_X1 FILLER_154_379 ();
 FILLCELL_X32 FILLER_154_1518 ();
 FILLCELL_X32 FILLER_154_1550 ();
 FILLCELL_X32 FILLER_154_1582 ();
 FILLCELL_X32 FILLER_154_1614 ();
 FILLCELL_X32 FILLER_154_1646 ();
 FILLCELL_X32 FILLER_154_1678 ();
 FILLCELL_X32 FILLER_154_1710 ();
 FILLCELL_X16 FILLER_154_1742 ();
 FILLCELL_X4 FILLER_154_1758 ();
 FILLCELL_X32 FILLER_155_1 ();
 FILLCELL_X32 FILLER_155_33 ();
 FILLCELL_X32 FILLER_155_65 ();
 FILLCELL_X32 FILLER_155_97 ();
 FILLCELL_X32 FILLER_155_129 ();
 FILLCELL_X32 FILLER_155_161 ();
 FILLCELL_X32 FILLER_155_193 ();
 FILLCELL_X32 FILLER_155_225 ();
 FILLCELL_X32 FILLER_155_257 ();
 FILLCELL_X32 FILLER_155_289 ();
 FILLCELL_X32 FILLER_155_321 ();
 FILLCELL_X16 FILLER_155_353 ();
 FILLCELL_X8 FILLER_155_369 ();
 FILLCELL_X2 FILLER_155_377 ();
 FILLCELL_X1 FILLER_155_379 ();
 FILLCELL_X32 FILLER_155_1518 ();
 FILLCELL_X32 FILLER_155_1550 ();
 FILLCELL_X32 FILLER_155_1582 ();
 FILLCELL_X32 FILLER_155_1614 ();
 FILLCELL_X32 FILLER_155_1646 ();
 FILLCELL_X32 FILLER_155_1678 ();
 FILLCELL_X32 FILLER_155_1710 ();
 FILLCELL_X8 FILLER_155_1742 ();
 FILLCELL_X4 FILLER_155_1750 ();
 FILLCELL_X1 FILLER_155_1754 ();
 FILLCELL_X4 FILLER_155_1758 ();
 FILLCELL_X32 FILLER_156_1 ();
 FILLCELL_X32 FILLER_156_33 ();
 FILLCELL_X32 FILLER_156_65 ();
 FILLCELL_X32 FILLER_156_97 ();
 FILLCELL_X32 FILLER_156_129 ();
 FILLCELL_X32 FILLER_156_161 ();
 FILLCELL_X32 FILLER_156_193 ();
 FILLCELL_X32 FILLER_156_225 ();
 FILLCELL_X32 FILLER_156_257 ();
 FILLCELL_X32 FILLER_156_289 ();
 FILLCELL_X32 FILLER_156_321 ();
 FILLCELL_X16 FILLER_156_353 ();
 FILLCELL_X8 FILLER_156_369 ();
 FILLCELL_X2 FILLER_156_377 ();
 FILLCELL_X1 FILLER_156_379 ();
 FILLCELL_X32 FILLER_156_1518 ();
 FILLCELL_X32 FILLER_156_1550 ();
 FILLCELL_X32 FILLER_156_1582 ();
 FILLCELL_X32 FILLER_156_1614 ();
 FILLCELL_X32 FILLER_156_1646 ();
 FILLCELL_X32 FILLER_156_1678 ();
 FILLCELL_X32 FILLER_156_1710 ();
 FILLCELL_X16 FILLER_156_1742 ();
 FILLCELL_X4 FILLER_156_1758 ();
 FILLCELL_X32 FILLER_157_1 ();
 FILLCELL_X32 FILLER_157_33 ();
 FILLCELL_X32 FILLER_157_65 ();
 FILLCELL_X32 FILLER_157_97 ();
 FILLCELL_X32 FILLER_157_129 ();
 FILLCELL_X32 FILLER_157_161 ();
 FILLCELL_X32 FILLER_157_193 ();
 FILLCELL_X32 FILLER_157_225 ();
 FILLCELL_X32 FILLER_157_257 ();
 FILLCELL_X32 FILLER_157_289 ();
 FILLCELL_X32 FILLER_157_321 ();
 FILLCELL_X16 FILLER_157_353 ();
 FILLCELL_X8 FILLER_157_369 ();
 FILLCELL_X2 FILLER_157_377 ();
 FILLCELL_X1 FILLER_157_379 ();
 FILLCELL_X32 FILLER_157_1518 ();
 FILLCELL_X32 FILLER_157_1550 ();
 FILLCELL_X32 FILLER_157_1582 ();
 FILLCELL_X32 FILLER_157_1614 ();
 FILLCELL_X32 FILLER_157_1646 ();
 FILLCELL_X32 FILLER_157_1678 ();
 FILLCELL_X32 FILLER_157_1710 ();
 FILLCELL_X16 FILLER_157_1742 ();
 FILLCELL_X4 FILLER_157_1758 ();
 FILLCELL_X32 FILLER_158_1 ();
 FILLCELL_X32 FILLER_158_33 ();
 FILLCELL_X32 FILLER_158_65 ();
 FILLCELL_X32 FILLER_158_97 ();
 FILLCELL_X32 FILLER_158_129 ();
 FILLCELL_X32 FILLER_158_161 ();
 FILLCELL_X32 FILLER_158_193 ();
 FILLCELL_X32 FILLER_158_225 ();
 FILLCELL_X32 FILLER_158_257 ();
 FILLCELL_X32 FILLER_158_289 ();
 FILLCELL_X32 FILLER_158_321 ();
 FILLCELL_X16 FILLER_158_353 ();
 FILLCELL_X8 FILLER_158_369 ();
 FILLCELL_X2 FILLER_158_377 ();
 FILLCELL_X1 FILLER_158_379 ();
 FILLCELL_X32 FILLER_158_1518 ();
 FILLCELL_X32 FILLER_158_1550 ();
 FILLCELL_X32 FILLER_158_1582 ();
 FILLCELL_X32 FILLER_158_1614 ();
 FILLCELL_X32 FILLER_158_1646 ();
 FILLCELL_X32 FILLER_158_1678 ();
 FILLCELL_X32 FILLER_158_1710 ();
 FILLCELL_X16 FILLER_158_1742 ();
 FILLCELL_X4 FILLER_158_1758 ();
 FILLCELL_X32 FILLER_159_1 ();
 FILLCELL_X32 FILLER_159_33 ();
 FILLCELL_X32 FILLER_159_65 ();
 FILLCELL_X32 FILLER_159_97 ();
 FILLCELL_X32 FILLER_159_129 ();
 FILLCELL_X32 FILLER_159_161 ();
 FILLCELL_X32 FILLER_159_193 ();
 FILLCELL_X32 FILLER_159_225 ();
 FILLCELL_X32 FILLER_159_257 ();
 FILLCELL_X32 FILLER_159_289 ();
 FILLCELL_X32 FILLER_159_321 ();
 FILLCELL_X16 FILLER_159_353 ();
 FILLCELL_X8 FILLER_159_369 ();
 FILLCELL_X2 FILLER_159_377 ();
 FILLCELL_X1 FILLER_159_379 ();
 FILLCELL_X32 FILLER_159_1518 ();
 FILLCELL_X32 FILLER_159_1550 ();
 FILLCELL_X32 FILLER_159_1582 ();
 FILLCELL_X32 FILLER_159_1614 ();
 FILLCELL_X32 FILLER_159_1646 ();
 FILLCELL_X32 FILLER_159_1678 ();
 FILLCELL_X32 FILLER_159_1710 ();
 FILLCELL_X16 FILLER_159_1742 ();
 FILLCELL_X4 FILLER_159_1758 ();
 FILLCELL_X4 FILLER_160_1 ();
 FILLCELL_X32 FILLER_160_10 ();
 FILLCELL_X32 FILLER_160_42 ();
 FILLCELL_X32 FILLER_160_74 ();
 FILLCELL_X32 FILLER_160_106 ();
 FILLCELL_X32 FILLER_160_138 ();
 FILLCELL_X32 FILLER_160_170 ();
 FILLCELL_X32 FILLER_160_202 ();
 FILLCELL_X32 FILLER_160_234 ();
 FILLCELL_X32 FILLER_160_266 ();
 FILLCELL_X32 FILLER_160_298 ();
 FILLCELL_X32 FILLER_160_330 ();
 FILLCELL_X16 FILLER_160_362 ();
 FILLCELL_X2 FILLER_160_378 ();
 FILLCELL_X32 FILLER_160_1518 ();
 FILLCELL_X32 FILLER_160_1550 ();
 FILLCELL_X32 FILLER_160_1582 ();
 FILLCELL_X32 FILLER_160_1614 ();
 FILLCELL_X32 FILLER_160_1646 ();
 FILLCELL_X32 FILLER_160_1678 ();
 FILLCELL_X32 FILLER_160_1710 ();
 FILLCELL_X16 FILLER_160_1742 ();
 FILLCELL_X4 FILLER_160_1758 ();
 FILLCELL_X32 FILLER_161_1 ();
 FILLCELL_X32 FILLER_161_33 ();
 FILLCELL_X32 FILLER_161_65 ();
 FILLCELL_X32 FILLER_161_97 ();
 FILLCELL_X32 FILLER_161_129 ();
 FILLCELL_X32 FILLER_161_161 ();
 FILLCELL_X32 FILLER_161_193 ();
 FILLCELL_X32 FILLER_161_225 ();
 FILLCELL_X32 FILLER_161_257 ();
 FILLCELL_X32 FILLER_161_289 ();
 FILLCELL_X32 FILLER_161_321 ();
 FILLCELL_X16 FILLER_161_353 ();
 FILLCELL_X8 FILLER_161_369 ();
 FILLCELL_X2 FILLER_161_377 ();
 FILLCELL_X1 FILLER_161_379 ();
 FILLCELL_X32 FILLER_161_1518 ();
 FILLCELL_X32 FILLER_161_1550 ();
 FILLCELL_X32 FILLER_161_1582 ();
 FILLCELL_X32 FILLER_161_1614 ();
 FILLCELL_X32 FILLER_161_1646 ();
 FILLCELL_X32 FILLER_161_1678 ();
 FILLCELL_X32 FILLER_161_1710 ();
 FILLCELL_X16 FILLER_161_1742 ();
 FILLCELL_X4 FILLER_161_1758 ();
 FILLCELL_X32 FILLER_162_1 ();
 FILLCELL_X32 FILLER_162_33 ();
 FILLCELL_X32 FILLER_162_65 ();
 FILLCELL_X32 FILLER_162_97 ();
 FILLCELL_X32 FILLER_162_129 ();
 FILLCELL_X32 FILLER_162_161 ();
 FILLCELL_X32 FILLER_162_193 ();
 FILLCELL_X32 FILLER_162_225 ();
 FILLCELL_X32 FILLER_162_257 ();
 FILLCELL_X32 FILLER_162_289 ();
 FILLCELL_X32 FILLER_162_321 ();
 FILLCELL_X16 FILLER_162_353 ();
 FILLCELL_X8 FILLER_162_369 ();
 FILLCELL_X2 FILLER_162_377 ();
 FILLCELL_X1 FILLER_162_379 ();
 FILLCELL_X32 FILLER_162_1518 ();
 FILLCELL_X32 FILLER_162_1550 ();
 FILLCELL_X32 FILLER_162_1582 ();
 FILLCELL_X32 FILLER_162_1614 ();
 FILLCELL_X32 FILLER_162_1646 ();
 FILLCELL_X32 FILLER_162_1678 ();
 FILLCELL_X32 FILLER_162_1710 ();
 FILLCELL_X16 FILLER_162_1742 ();
 FILLCELL_X4 FILLER_162_1758 ();
 FILLCELL_X32 FILLER_163_1 ();
 FILLCELL_X32 FILLER_163_33 ();
 FILLCELL_X32 FILLER_163_65 ();
 FILLCELL_X32 FILLER_163_97 ();
 FILLCELL_X32 FILLER_163_129 ();
 FILLCELL_X32 FILLER_163_161 ();
 FILLCELL_X32 FILLER_163_193 ();
 FILLCELL_X32 FILLER_163_225 ();
 FILLCELL_X32 FILLER_163_257 ();
 FILLCELL_X32 FILLER_163_289 ();
 FILLCELL_X32 FILLER_163_321 ();
 FILLCELL_X16 FILLER_163_353 ();
 FILLCELL_X8 FILLER_163_369 ();
 FILLCELL_X2 FILLER_163_377 ();
 FILLCELL_X1 FILLER_163_379 ();
 FILLCELL_X32 FILLER_163_1518 ();
 FILLCELL_X32 FILLER_163_1550 ();
 FILLCELL_X32 FILLER_163_1582 ();
 FILLCELL_X32 FILLER_163_1614 ();
 FILLCELL_X32 FILLER_163_1646 ();
 FILLCELL_X32 FILLER_163_1678 ();
 FILLCELL_X32 FILLER_163_1710 ();
 FILLCELL_X16 FILLER_163_1742 ();
 FILLCELL_X4 FILLER_163_1758 ();
 FILLCELL_X32 FILLER_164_1 ();
 FILLCELL_X32 FILLER_164_33 ();
 FILLCELL_X32 FILLER_164_65 ();
 FILLCELL_X32 FILLER_164_97 ();
 FILLCELL_X32 FILLER_164_129 ();
 FILLCELL_X32 FILLER_164_161 ();
 FILLCELL_X32 FILLER_164_193 ();
 FILLCELL_X32 FILLER_164_225 ();
 FILLCELL_X32 FILLER_164_257 ();
 FILLCELL_X32 FILLER_164_289 ();
 FILLCELL_X32 FILLER_164_321 ();
 FILLCELL_X16 FILLER_164_353 ();
 FILLCELL_X8 FILLER_164_369 ();
 FILLCELL_X2 FILLER_164_377 ();
 FILLCELL_X1 FILLER_164_379 ();
 FILLCELL_X32 FILLER_164_1518 ();
 FILLCELL_X32 FILLER_164_1550 ();
 FILLCELL_X32 FILLER_164_1582 ();
 FILLCELL_X32 FILLER_164_1614 ();
 FILLCELL_X32 FILLER_164_1646 ();
 FILLCELL_X32 FILLER_164_1678 ();
 FILLCELL_X32 FILLER_164_1710 ();
 FILLCELL_X16 FILLER_164_1742 ();
 FILLCELL_X4 FILLER_164_1758 ();
 FILLCELL_X32 FILLER_165_1 ();
 FILLCELL_X32 FILLER_165_33 ();
 FILLCELL_X32 FILLER_165_65 ();
 FILLCELL_X32 FILLER_165_97 ();
 FILLCELL_X32 FILLER_165_129 ();
 FILLCELL_X32 FILLER_165_161 ();
 FILLCELL_X32 FILLER_165_193 ();
 FILLCELL_X32 FILLER_165_225 ();
 FILLCELL_X32 FILLER_165_257 ();
 FILLCELL_X32 FILLER_165_289 ();
 FILLCELL_X32 FILLER_165_321 ();
 FILLCELL_X16 FILLER_165_353 ();
 FILLCELL_X8 FILLER_165_369 ();
 FILLCELL_X2 FILLER_165_377 ();
 FILLCELL_X1 FILLER_165_379 ();
 FILLCELL_X32 FILLER_165_1518 ();
 FILLCELL_X32 FILLER_165_1550 ();
 FILLCELL_X32 FILLER_165_1582 ();
 FILLCELL_X32 FILLER_165_1614 ();
 FILLCELL_X32 FILLER_165_1646 ();
 FILLCELL_X32 FILLER_165_1678 ();
 FILLCELL_X32 FILLER_165_1710 ();
 FILLCELL_X8 FILLER_165_1742 ();
 FILLCELL_X4 FILLER_165_1750 ();
 FILLCELL_X1 FILLER_165_1754 ();
 FILLCELL_X4 FILLER_165_1758 ();
 FILLCELL_X32 FILLER_166_1 ();
 FILLCELL_X32 FILLER_166_33 ();
 FILLCELL_X32 FILLER_166_65 ();
 FILLCELL_X32 FILLER_166_97 ();
 FILLCELL_X32 FILLER_166_129 ();
 FILLCELL_X32 FILLER_166_161 ();
 FILLCELL_X32 FILLER_166_193 ();
 FILLCELL_X32 FILLER_166_225 ();
 FILLCELL_X32 FILLER_166_257 ();
 FILLCELL_X32 FILLER_166_289 ();
 FILLCELL_X32 FILLER_166_321 ();
 FILLCELL_X16 FILLER_166_353 ();
 FILLCELL_X8 FILLER_166_369 ();
 FILLCELL_X2 FILLER_166_377 ();
 FILLCELL_X1 FILLER_166_379 ();
 FILLCELL_X32 FILLER_166_1518 ();
 FILLCELL_X32 FILLER_166_1550 ();
 FILLCELL_X32 FILLER_166_1582 ();
 FILLCELL_X32 FILLER_166_1614 ();
 FILLCELL_X32 FILLER_166_1646 ();
 FILLCELL_X32 FILLER_166_1678 ();
 FILLCELL_X32 FILLER_166_1710 ();
 FILLCELL_X16 FILLER_166_1742 ();
 FILLCELL_X4 FILLER_166_1758 ();
 FILLCELL_X32 FILLER_167_1 ();
 FILLCELL_X32 FILLER_167_33 ();
 FILLCELL_X32 FILLER_167_65 ();
 FILLCELL_X32 FILLER_167_97 ();
 FILLCELL_X32 FILLER_167_129 ();
 FILLCELL_X32 FILLER_167_161 ();
 FILLCELL_X32 FILLER_167_193 ();
 FILLCELL_X32 FILLER_167_225 ();
 FILLCELL_X32 FILLER_167_257 ();
 FILLCELL_X32 FILLER_167_289 ();
 FILLCELL_X32 FILLER_167_321 ();
 FILLCELL_X16 FILLER_167_353 ();
 FILLCELL_X8 FILLER_167_369 ();
 FILLCELL_X2 FILLER_167_377 ();
 FILLCELL_X1 FILLER_167_379 ();
 FILLCELL_X32 FILLER_167_1518 ();
 FILLCELL_X32 FILLER_167_1550 ();
 FILLCELL_X32 FILLER_167_1582 ();
 FILLCELL_X32 FILLER_167_1614 ();
 FILLCELL_X32 FILLER_167_1646 ();
 FILLCELL_X32 FILLER_167_1678 ();
 FILLCELL_X32 FILLER_167_1710 ();
 FILLCELL_X16 FILLER_167_1742 ();
 FILLCELL_X4 FILLER_167_1758 ();
 FILLCELL_X32 FILLER_168_1 ();
 FILLCELL_X32 FILLER_168_33 ();
 FILLCELL_X32 FILLER_168_65 ();
 FILLCELL_X32 FILLER_168_97 ();
 FILLCELL_X32 FILLER_168_129 ();
 FILLCELL_X32 FILLER_168_161 ();
 FILLCELL_X32 FILLER_168_193 ();
 FILLCELL_X32 FILLER_168_225 ();
 FILLCELL_X32 FILLER_168_257 ();
 FILLCELL_X32 FILLER_168_289 ();
 FILLCELL_X32 FILLER_168_321 ();
 FILLCELL_X16 FILLER_168_353 ();
 FILLCELL_X8 FILLER_168_369 ();
 FILLCELL_X2 FILLER_168_377 ();
 FILLCELL_X1 FILLER_168_379 ();
 FILLCELL_X32 FILLER_168_1518 ();
 FILLCELL_X32 FILLER_168_1550 ();
 FILLCELL_X32 FILLER_168_1582 ();
 FILLCELL_X32 FILLER_168_1614 ();
 FILLCELL_X32 FILLER_168_1646 ();
 FILLCELL_X32 FILLER_168_1678 ();
 FILLCELL_X32 FILLER_168_1710 ();
 FILLCELL_X16 FILLER_168_1742 ();
 FILLCELL_X4 FILLER_168_1758 ();
 FILLCELL_X32 FILLER_169_1 ();
 FILLCELL_X32 FILLER_169_33 ();
 FILLCELL_X32 FILLER_169_65 ();
 FILLCELL_X32 FILLER_169_97 ();
 FILLCELL_X32 FILLER_169_129 ();
 FILLCELL_X32 FILLER_169_161 ();
 FILLCELL_X32 FILLER_169_193 ();
 FILLCELL_X32 FILLER_169_225 ();
 FILLCELL_X32 FILLER_169_257 ();
 FILLCELL_X32 FILLER_169_289 ();
 FILLCELL_X32 FILLER_169_321 ();
 FILLCELL_X16 FILLER_169_353 ();
 FILLCELL_X8 FILLER_169_369 ();
 FILLCELL_X2 FILLER_169_377 ();
 FILLCELL_X1 FILLER_169_379 ();
 FILLCELL_X32 FILLER_169_1518 ();
 FILLCELL_X32 FILLER_169_1550 ();
 FILLCELL_X32 FILLER_169_1582 ();
 FILLCELL_X32 FILLER_169_1614 ();
 FILLCELL_X32 FILLER_169_1646 ();
 FILLCELL_X32 FILLER_169_1678 ();
 FILLCELL_X32 FILLER_169_1710 ();
 FILLCELL_X16 FILLER_169_1742 ();
 FILLCELL_X4 FILLER_169_1758 ();
 FILLCELL_X4 FILLER_170_1 ();
 FILLCELL_X32 FILLER_170_8 ();
 FILLCELL_X32 FILLER_170_40 ();
 FILLCELL_X32 FILLER_170_72 ();
 FILLCELL_X32 FILLER_170_104 ();
 FILLCELL_X32 FILLER_170_136 ();
 FILLCELL_X32 FILLER_170_168 ();
 FILLCELL_X32 FILLER_170_200 ();
 FILLCELL_X32 FILLER_170_232 ();
 FILLCELL_X32 FILLER_170_264 ();
 FILLCELL_X32 FILLER_170_296 ();
 FILLCELL_X32 FILLER_170_328 ();
 FILLCELL_X16 FILLER_170_360 ();
 FILLCELL_X4 FILLER_170_376 ();
 FILLCELL_X32 FILLER_170_1518 ();
 FILLCELL_X32 FILLER_170_1550 ();
 FILLCELL_X32 FILLER_170_1582 ();
 FILLCELL_X32 FILLER_170_1614 ();
 FILLCELL_X32 FILLER_170_1646 ();
 FILLCELL_X32 FILLER_170_1678 ();
 FILLCELL_X32 FILLER_170_1710 ();
 FILLCELL_X16 FILLER_170_1742 ();
 FILLCELL_X4 FILLER_170_1758 ();
 FILLCELL_X32 FILLER_171_1 ();
 FILLCELL_X32 FILLER_171_33 ();
 FILLCELL_X32 FILLER_171_65 ();
 FILLCELL_X32 FILLER_171_97 ();
 FILLCELL_X32 FILLER_171_129 ();
 FILLCELL_X32 FILLER_171_161 ();
 FILLCELL_X32 FILLER_171_193 ();
 FILLCELL_X32 FILLER_171_225 ();
 FILLCELL_X32 FILLER_171_257 ();
 FILLCELL_X32 FILLER_171_289 ();
 FILLCELL_X32 FILLER_171_321 ();
 FILLCELL_X16 FILLER_171_353 ();
 FILLCELL_X8 FILLER_171_369 ();
 FILLCELL_X2 FILLER_171_377 ();
 FILLCELL_X1 FILLER_171_379 ();
 FILLCELL_X32 FILLER_171_1518 ();
 FILLCELL_X32 FILLER_171_1550 ();
 FILLCELL_X32 FILLER_171_1582 ();
 FILLCELL_X32 FILLER_171_1614 ();
 FILLCELL_X32 FILLER_171_1646 ();
 FILLCELL_X32 FILLER_171_1678 ();
 FILLCELL_X32 FILLER_171_1710 ();
 FILLCELL_X16 FILLER_171_1742 ();
 FILLCELL_X4 FILLER_171_1758 ();
 FILLCELL_X32 FILLER_172_1 ();
 FILLCELL_X32 FILLER_172_33 ();
 FILLCELL_X32 FILLER_172_65 ();
 FILLCELL_X32 FILLER_172_97 ();
 FILLCELL_X32 FILLER_172_129 ();
 FILLCELL_X32 FILLER_172_161 ();
 FILLCELL_X32 FILLER_172_193 ();
 FILLCELL_X32 FILLER_172_225 ();
 FILLCELL_X32 FILLER_172_257 ();
 FILLCELL_X32 FILLER_172_289 ();
 FILLCELL_X32 FILLER_172_321 ();
 FILLCELL_X16 FILLER_172_353 ();
 FILLCELL_X8 FILLER_172_369 ();
 FILLCELL_X2 FILLER_172_377 ();
 FILLCELL_X1 FILLER_172_379 ();
 FILLCELL_X32 FILLER_172_1518 ();
 FILLCELL_X32 FILLER_172_1550 ();
 FILLCELL_X32 FILLER_172_1582 ();
 FILLCELL_X32 FILLER_172_1614 ();
 FILLCELL_X32 FILLER_172_1646 ();
 FILLCELL_X32 FILLER_172_1678 ();
 FILLCELL_X32 FILLER_172_1710 ();
 FILLCELL_X16 FILLER_172_1742 ();
 FILLCELL_X4 FILLER_172_1758 ();
 FILLCELL_X32 FILLER_173_1 ();
 FILLCELL_X32 FILLER_173_33 ();
 FILLCELL_X32 FILLER_173_65 ();
 FILLCELL_X32 FILLER_173_97 ();
 FILLCELL_X32 FILLER_173_129 ();
 FILLCELL_X32 FILLER_173_161 ();
 FILLCELL_X32 FILLER_173_193 ();
 FILLCELL_X32 FILLER_173_225 ();
 FILLCELL_X32 FILLER_173_257 ();
 FILLCELL_X32 FILLER_173_289 ();
 FILLCELL_X32 FILLER_173_321 ();
 FILLCELL_X16 FILLER_173_353 ();
 FILLCELL_X8 FILLER_173_369 ();
 FILLCELL_X2 FILLER_173_377 ();
 FILLCELL_X1 FILLER_173_379 ();
 FILLCELL_X32 FILLER_173_1518 ();
 FILLCELL_X32 FILLER_173_1550 ();
 FILLCELL_X32 FILLER_173_1582 ();
 FILLCELL_X32 FILLER_173_1614 ();
 FILLCELL_X32 FILLER_173_1646 ();
 FILLCELL_X32 FILLER_173_1678 ();
 FILLCELL_X32 FILLER_173_1710 ();
 FILLCELL_X16 FILLER_173_1742 ();
 FILLCELL_X4 FILLER_173_1758 ();
 FILLCELL_X32 FILLER_174_1 ();
 FILLCELL_X32 FILLER_174_33 ();
 FILLCELL_X32 FILLER_174_65 ();
 FILLCELL_X32 FILLER_174_97 ();
 FILLCELL_X32 FILLER_174_129 ();
 FILLCELL_X32 FILLER_174_161 ();
 FILLCELL_X32 FILLER_174_193 ();
 FILLCELL_X32 FILLER_174_225 ();
 FILLCELL_X32 FILLER_174_257 ();
 FILLCELL_X32 FILLER_174_289 ();
 FILLCELL_X32 FILLER_174_321 ();
 FILLCELL_X16 FILLER_174_353 ();
 FILLCELL_X8 FILLER_174_369 ();
 FILLCELL_X2 FILLER_174_377 ();
 FILLCELL_X1 FILLER_174_379 ();
 FILLCELL_X32 FILLER_174_1518 ();
 FILLCELL_X32 FILLER_174_1550 ();
 FILLCELL_X32 FILLER_174_1582 ();
 FILLCELL_X32 FILLER_174_1614 ();
 FILLCELL_X32 FILLER_174_1646 ();
 FILLCELL_X32 FILLER_174_1678 ();
 FILLCELL_X32 FILLER_174_1710 ();
 FILLCELL_X8 FILLER_174_1742 ();
 FILLCELL_X1 FILLER_174_1750 ();
 FILLCELL_X4 FILLER_174_1758 ();
 FILLCELL_X32 FILLER_175_1 ();
 FILLCELL_X32 FILLER_175_33 ();
 FILLCELL_X32 FILLER_175_65 ();
 FILLCELL_X32 FILLER_175_97 ();
 FILLCELL_X32 FILLER_175_129 ();
 FILLCELL_X32 FILLER_175_161 ();
 FILLCELL_X32 FILLER_175_193 ();
 FILLCELL_X32 FILLER_175_225 ();
 FILLCELL_X32 FILLER_175_257 ();
 FILLCELL_X32 FILLER_175_289 ();
 FILLCELL_X32 FILLER_175_321 ();
 FILLCELL_X16 FILLER_175_353 ();
 FILLCELL_X8 FILLER_175_369 ();
 FILLCELL_X2 FILLER_175_377 ();
 FILLCELL_X1 FILLER_175_379 ();
 FILLCELL_X32 FILLER_175_1518 ();
 FILLCELL_X32 FILLER_175_1550 ();
 FILLCELL_X32 FILLER_175_1582 ();
 FILLCELL_X32 FILLER_175_1614 ();
 FILLCELL_X32 FILLER_175_1646 ();
 FILLCELL_X32 FILLER_175_1678 ();
 FILLCELL_X32 FILLER_175_1710 ();
 FILLCELL_X16 FILLER_175_1742 ();
 FILLCELL_X4 FILLER_175_1758 ();
 FILLCELL_X32 FILLER_176_1 ();
 FILLCELL_X32 FILLER_176_33 ();
 FILLCELL_X32 FILLER_176_65 ();
 FILLCELL_X32 FILLER_176_97 ();
 FILLCELL_X32 FILLER_176_129 ();
 FILLCELL_X32 FILLER_176_161 ();
 FILLCELL_X32 FILLER_176_193 ();
 FILLCELL_X32 FILLER_176_225 ();
 FILLCELL_X32 FILLER_176_257 ();
 FILLCELL_X32 FILLER_176_289 ();
 FILLCELL_X32 FILLER_176_321 ();
 FILLCELL_X16 FILLER_176_353 ();
 FILLCELL_X8 FILLER_176_369 ();
 FILLCELL_X2 FILLER_176_377 ();
 FILLCELL_X1 FILLER_176_379 ();
 FILLCELL_X32 FILLER_176_1518 ();
 FILLCELL_X32 FILLER_176_1550 ();
 FILLCELL_X32 FILLER_176_1582 ();
 FILLCELL_X32 FILLER_176_1614 ();
 FILLCELL_X32 FILLER_176_1646 ();
 FILLCELL_X32 FILLER_176_1678 ();
 FILLCELL_X32 FILLER_176_1710 ();
 FILLCELL_X16 FILLER_176_1742 ();
 FILLCELL_X4 FILLER_176_1758 ();
 FILLCELL_X32 FILLER_177_1 ();
 FILLCELL_X32 FILLER_177_33 ();
 FILLCELL_X32 FILLER_177_65 ();
 FILLCELL_X32 FILLER_177_97 ();
 FILLCELL_X32 FILLER_177_129 ();
 FILLCELL_X32 FILLER_177_161 ();
 FILLCELL_X32 FILLER_177_193 ();
 FILLCELL_X32 FILLER_177_225 ();
 FILLCELL_X32 FILLER_177_257 ();
 FILLCELL_X32 FILLER_177_289 ();
 FILLCELL_X32 FILLER_177_321 ();
 FILLCELL_X16 FILLER_177_353 ();
 FILLCELL_X8 FILLER_177_369 ();
 FILLCELL_X2 FILLER_177_377 ();
 FILLCELL_X1 FILLER_177_379 ();
 FILLCELL_X32 FILLER_177_1518 ();
 FILLCELL_X32 FILLER_177_1550 ();
 FILLCELL_X32 FILLER_177_1582 ();
 FILLCELL_X32 FILLER_177_1614 ();
 FILLCELL_X32 FILLER_177_1646 ();
 FILLCELL_X32 FILLER_177_1678 ();
 FILLCELL_X32 FILLER_177_1710 ();
 FILLCELL_X16 FILLER_177_1742 ();
 FILLCELL_X4 FILLER_177_1758 ();
 FILLCELL_X32 FILLER_178_1 ();
 FILLCELL_X32 FILLER_178_33 ();
 FILLCELL_X32 FILLER_178_65 ();
 FILLCELL_X32 FILLER_178_97 ();
 FILLCELL_X32 FILLER_178_129 ();
 FILLCELL_X32 FILLER_178_161 ();
 FILLCELL_X32 FILLER_178_193 ();
 FILLCELL_X32 FILLER_178_225 ();
 FILLCELL_X32 FILLER_178_257 ();
 FILLCELL_X32 FILLER_178_289 ();
 FILLCELL_X32 FILLER_178_321 ();
 FILLCELL_X16 FILLER_178_353 ();
 FILLCELL_X8 FILLER_178_369 ();
 FILLCELL_X2 FILLER_178_377 ();
 FILLCELL_X1 FILLER_178_379 ();
 FILLCELL_X32 FILLER_178_1518 ();
 FILLCELL_X32 FILLER_178_1550 ();
 FILLCELL_X32 FILLER_178_1582 ();
 FILLCELL_X32 FILLER_178_1614 ();
 FILLCELL_X32 FILLER_178_1646 ();
 FILLCELL_X32 FILLER_178_1678 ();
 FILLCELL_X32 FILLER_178_1710 ();
 FILLCELL_X16 FILLER_178_1742 ();
 FILLCELL_X4 FILLER_178_1758 ();
 FILLCELL_X4 FILLER_179_1 ();
 FILLCELL_X32 FILLER_179_10 ();
 FILLCELL_X32 FILLER_179_42 ();
 FILLCELL_X32 FILLER_179_74 ();
 FILLCELL_X32 FILLER_179_106 ();
 FILLCELL_X32 FILLER_179_138 ();
 FILLCELL_X32 FILLER_179_170 ();
 FILLCELL_X32 FILLER_179_202 ();
 FILLCELL_X32 FILLER_179_234 ();
 FILLCELL_X32 FILLER_179_266 ();
 FILLCELL_X32 FILLER_179_298 ();
 FILLCELL_X32 FILLER_179_330 ();
 FILLCELL_X16 FILLER_179_362 ();
 FILLCELL_X2 FILLER_179_378 ();
 FILLCELL_X32 FILLER_179_1518 ();
 FILLCELL_X32 FILLER_179_1550 ();
 FILLCELL_X32 FILLER_179_1582 ();
 FILLCELL_X32 FILLER_179_1614 ();
 FILLCELL_X32 FILLER_179_1646 ();
 FILLCELL_X32 FILLER_179_1678 ();
 FILLCELL_X32 FILLER_179_1710 ();
 FILLCELL_X16 FILLER_179_1742 ();
 FILLCELL_X4 FILLER_179_1758 ();
 FILLCELL_X32 FILLER_180_1 ();
 FILLCELL_X32 FILLER_180_33 ();
 FILLCELL_X32 FILLER_180_65 ();
 FILLCELL_X32 FILLER_180_97 ();
 FILLCELL_X32 FILLER_180_129 ();
 FILLCELL_X32 FILLER_180_161 ();
 FILLCELL_X32 FILLER_180_193 ();
 FILLCELL_X32 FILLER_180_225 ();
 FILLCELL_X32 FILLER_180_257 ();
 FILLCELL_X32 FILLER_180_289 ();
 FILLCELL_X32 FILLER_180_321 ();
 FILLCELL_X16 FILLER_180_353 ();
 FILLCELL_X8 FILLER_180_369 ();
 FILLCELL_X2 FILLER_180_377 ();
 FILLCELL_X1 FILLER_180_379 ();
 FILLCELL_X32 FILLER_180_1518 ();
 FILLCELL_X32 FILLER_180_1550 ();
 FILLCELL_X32 FILLER_180_1582 ();
 FILLCELL_X32 FILLER_180_1614 ();
 FILLCELL_X32 FILLER_180_1646 ();
 FILLCELL_X32 FILLER_180_1678 ();
 FILLCELL_X32 FILLER_180_1710 ();
 FILLCELL_X16 FILLER_180_1742 ();
 FILLCELL_X4 FILLER_180_1758 ();
 FILLCELL_X32 FILLER_181_1 ();
 FILLCELL_X32 FILLER_181_33 ();
 FILLCELL_X32 FILLER_181_65 ();
 FILLCELL_X32 FILLER_181_97 ();
 FILLCELL_X32 FILLER_181_129 ();
 FILLCELL_X32 FILLER_181_161 ();
 FILLCELL_X32 FILLER_181_193 ();
 FILLCELL_X32 FILLER_181_225 ();
 FILLCELL_X32 FILLER_181_257 ();
 FILLCELL_X32 FILLER_181_289 ();
 FILLCELL_X32 FILLER_181_321 ();
 FILLCELL_X16 FILLER_181_353 ();
 FILLCELL_X8 FILLER_181_369 ();
 FILLCELL_X2 FILLER_181_377 ();
 FILLCELL_X1 FILLER_181_379 ();
 FILLCELL_X32 FILLER_181_1518 ();
 FILLCELL_X32 FILLER_181_1550 ();
 FILLCELL_X32 FILLER_181_1582 ();
 FILLCELL_X32 FILLER_181_1614 ();
 FILLCELL_X32 FILLER_181_1646 ();
 FILLCELL_X32 FILLER_181_1678 ();
 FILLCELL_X32 FILLER_181_1710 ();
 FILLCELL_X16 FILLER_181_1742 ();
 FILLCELL_X4 FILLER_181_1758 ();
 FILLCELL_X32 FILLER_182_1 ();
 FILLCELL_X32 FILLER_182_33 ();
 FILLCELL_X32 FILLER_182_65 ();
 FILLCELL_X32 FILLER_182_97 ();
 FILLCELL_X32 FILLER_182_129 ();
 FILLCELL_X32 FILLER_182_161 ();
 FILLCELL_X32 FILLER_182_193 ();
 FILLCELL_X32 FILLER_182_225 ();
 FILLCELL_X32 FILLER_182_257 ();
 FILLCELL_X32 FILLER_182_289 ();
 FILLCELL_X32 FILLER_182_321 ();
 FILLCELL_X16 FILLER_182_353 ();
 FILLCELL_X8 FILLER_182_369 ();
 FILLCELL_X2 FILLER_182_377 ();
 FILLCELL_X1 FILLER_182_379 ();
 FILLCELL_X32 FILLER_182_1518 ();
 FILLCELL_X32 FILLER_182_1550 ();
 FILLCELL_X32 FILLER_182_1582 ();
 FILLCELL_X32 FILLER_182_1614 ();
 FILLCELL_X32 FILLER_182_1646 ();
 FILLCELL_X32 FILLER_182_1678 ();
 FILLCELL_X32 FILLER_182_1710 ();
 FILLCELL_X16 FILLER_182_1742 ();
 FILLCELL_X4 FILLER_182_1758 ();
 FILLCELL_X32 FILLER_183_1 ();
 FILLCELL_X32 FILLER_183_33 ();
 FILLCELL_X32 FILLER_183_65 ();
 FILLCELL_X32 FILLER_183_97 ();
 FILLCELL_X32 FILLER_183_129 ();
 FILLCELL_X32 FILLER_183_161 ();
 FILLCELL_X32 FILLER_183_193 ();
 FILLCELL_X32 FILLER_183_225 ();
 FILLCELL_X32 FILLER_183_257 ();
 FILLCELL_X32 FILLER_183_289 ();
 FILLCELL_X32 FILLER_183_321 ();
 FILLCELL_X16 FILLER_183_353 ();
 FILLCELL_X8 FILLER_183_369 ();
 FILLCELL_X2 FILLER_183_377 ();
 FILLCELL_X1 FILLER_183_379 ();
 FILLCELL_X32 FILLER_183_1518 ();
 FILLCELL_X32 FILLER_183_1550 ();
 FILLCELL_X32 FILLER_183_1582 ();
 FILLCELL_X32 FILLER_183_1614 ();
 FILLCELL_X32 FILLER_183_1646 ();
 FILLCELL_X32 FILLER_183_1678 ();
 FILLCELL_X32 FILLER_183_1710 ();
 FILLCELL_X16 FILLER_183_1742 ();
 FILLCELL_X4 FILLER_183_1758 ();
 FILLCELL_X32 FILLER_184_1 ();
 FILLCELL_X32 FILLER_184_33 ();
 FILLCELL_X32 FILLER_184_65 ();
 FILLCELL_X32 FILLER_184_97 ();
 FILLCELL_X32 FILLER_184_129 ();
 FILLCELL_X32 FILLER_184_161 ();
 FILLCELL_X32 FILLER_184_193 ();
 FILLCELL_X32 FILLER_184_225 ();
 FILLCELL_X32 FILLER_184_257 ();
 FILLCELL_X32 FILLER_184_289 ();
 FILLCELL_X32 FILLER_184_321 ();
 FILLCELL_X16 FILLER_184_353 ();
 FILLCELL_X8 FILLER_184_369 ();
 FILLCELL_X2 FILLER_184_377 ();
 FILLCELL_X1 FILLER_184_379 ();
 FILLCELL_X32 FILLER_184_1518 ();
 FILLCELL_X32 FILLER_184_1550 ();
 FILLCELL_X32 FILLER_184_1582 ();
 FILLCELL_X32 FILLER_184_1614 ();
 FILLCELL_X32 FILLER_184_1646 ();
 FILLCELL_X32 FILLER_184_1678 ();
 FILLCELL_X32 FILLER_184_1710 ();
 FILLCELL_X8 FILLER_184_1742 ();
 FILLCELL_X4 FILLER_184_1750 ();
 FILLCELL_X1 FILLER_184_1754 ();
 FILLCELL_X4 FILLER_184_1758 ();
 FILLCELL_X32 FILLER_185_1 ();
 FILLCELL_X32 FILLER_185_33 ();
 FILLCELL_X32 FILLER_185_65 ();
 FILLCELL_X32 FILLER_185_97 ();
 FILLCELL_X32 FILLER_185_129 ();
 FILLCELL_X32 FILLER_185_161 ();
 FILLCELL_X32 FILLER_185_193 ();
 FILLCELL_X32 FILLER_185_225 ();
 FILLCELL_X32 FILLER_185_257 ();
 FILLCELL_X32 FILLER_185_289 ();
 FILLCELL_X32 FILLER_185_321 ();
 FILLCELL_X16 FILLER_185_353 ();
 FILLCELL_X8 FILLER_185_369 ();
 FILLCELL_X2 FILLER_185_377 ();
 FILLCELL_X1 FILLER_185_379 ();
 FILLCELL_X32 FILLER_185_1518 ();
 FILLCELL_X32 FILLER_185_1550 ();
 FILLCELL_X32 FILLER_185_1582 ();
 FILLCELL_X32 FILLER_185_1614 ();
 FILLCELL_X32 FILLER_185_1646 ();
 FILLCELL_X32 FILLER_185_1678 ();
 FILLCELL_X32 FILLER_185_1710 ();
 FILLCELL_X16 FILLER_185_1742 ();
 FILLCELL_X4 FILLER_185_1758 ();
 FILLCELL_X32 FILLER_186_1 ();
 FILLCELL_X32 FILLER_186_33 ();
 FILLCELL_X32 FILLER_186_65 ();
 FILLCELL_X32 FILLER_186_97 ();
 FILLCELL_X32 FILLER_186_129 ();
 FILLCELL_X32 FILLER_186_161 ();
 FILLCELL_X32 FILLER_186_193 ();
 FILLCELL_X32 FILLER_186_225 ();
 FILLCELL_X32 FILLER_186_257 ();
 FILLCELL_X32 FILLER_186_289 ();
 FILLCELL_X32 FILLER_186_321 ();
 FILLCELL_X16 FILLER_186_353 ();
 FILLCELL_X8 FILLER_186_369 ();
 FILLCELL_X2 FILLER_186_377 ();
 FILLCELL_X1 FILLER_186_379 ();
 FILLCELL_X32 FILLER_186_1518 ();
 FILLCELL_X32 FILLER_186_1550 ();
 FILLCELL_X32 FILLER_186_1582 ();
 FILLCELL_X32 FILLER_186_1614 ();
 FILLCELL_X32 FILLER_186_1646 ();
 FILLCELL_X32 FILLER_186_1678 ();
 FILLCELL_X32 FILLER_186_1710 ();
 FILLCELL_X16 FILLER_186_1742 ();
 FILLCELL_X4 FILLER_186_1758 ();
 FILLCELL_X32 FILLER_187_1 ();
 FILLCELL_X32 FILLER_187_33 ();
 FILLCELL_X32 FILLER_187_65 ();
 FILLCELL_X32 FILLER_187_97 ();
 FILLCELL_X32 FILLER_187_129 ();
 FILLCELL_X32 FILLER_187_161 ();
 FILLCELL_X32 FILLER_187_193 ();
 FILLCELL_X32 FILLER_187_225 ();
 FILLCELL_X32 FILLER_187_257 ();
 FILLCELL_X32 FILLER_187_289 ();
 FILLCELL_X32 FILLER_187_321 ();
 FILLCELL_X16 FILLER_187_353 ();
 FILLCELL_X8 FILLER_187_369 ();
 FILLCELL_X2 FILLER_187_377 ();
 FILLCELL_X1 FILLER_187_379 ();
 FILLCELL_X32 FILLER_187_1518 ();
 FILLCELL_X32 FILLER_187_1550 ();
 FILLCELL_X32 FILLER_187_1582 ();
 FILLCELL_X32 FILLER_187_1614 ();
 FILLCELL_X32 FILLER_187_1646 ();
 FILLCELL_X32 FILLER_187_1678 ();
 FILLCELL_X32 FILLER_187_1710 ();
 FILLCELL_X16 FILLER_187_1742 ();
 FILLCELL_X4 FILLER_187_1758 ();
 FILLCELL_X32 FILLER_188_1 ();
 FILLCELL_X32 FILLER_188_33 ();
 FILLCELL_X32 FILLER_188_65 ();
 FILLCELL_X32 FILLER_188_97 ();
 FILLCELL_X32 FILLER_188_129 ();
 FILLCELL_X32 FILLER_188_161 ();
 FILLCELL_X32 FILLER_188_193 ();
 FILLCELL_X32 FILLER_188_225 ();
 FILLCELL_X32 FILLER_188_257 ();
 FILLCELL_X32 FILLER_188_289 ();
 FILLCELL_X32 FILLER_188_321 ();
 FILLCELL_X16 FILLER_188_353 ();
 FILLCELL_X8 FILLER_188_369 ();
 FILLCELL_X2 FILLER_188_377 ();
 FILLCELL_X1 FILLER_188_379 ();
 FILLCELL_X32 FILLER_188_1518 ();
 FILLCELL_X32 FILLER_188_1550 ();
 FILLCELL_X32 FILLER_188_1582 ();
 FILLCELL_X32 FILLER_188_1614 ();
 FILLCELL_X32 FILLER_188_1646 ();
 FILLCELL_X32 FILLER_188_1678 ();
 FILLCELL_X32 FILLER_188_1710 ();
 FILLCELL_X16 FILLER_188_1742 ();
 FILLCELL_X4 FILLER_188_1758 ();
 FILLCELL_X4 FILLER_189_1 ();
 FILLCELL_X32 FILLER_189_10 ();
 FILLCELL_X32 FILLER_189_42 ();
 FILLCELL_X32 FILLER_189_74 ();
 FILLCELL_X32 FILLER_189_106 ();
 FILLCELL_X32 FILLER_189_138 ();
 FILLCELL_X32 FILLER_189_170 ();
 FILLCELL_X32 FILLER_189_202 ();
 FILLCELL_X32 FILLER_189_234 ();
 FILLCELL_X32 FILLER_189_266 ();
 FILLCELL_X32 FILLER_189_298 ();
 FILLCELL_X32 FILLER_189_330 ();
 FILLCELL_X16 FILLER_189_362 ();
 FILLCELL_X2 FILLER_189_378 ();
 FILLCELL_X32 FILLER_189_1518 ();
 FILLCELL_X32 FILLER_189_1550 ();
 FILLCELL_X32 FILLER_189_1582 ();
 FILLCELL_X32 FILLER_189_1614 ();
 FILLCELL_X32 FILLER_189_1646 ();
 FILLCELL_X32 FILLER_189_1678 ();
 FILLCELL_X32 FILLER_189_1710 ();
 FILLCELL_X16 FILLER_189_1742 ();
 FILLCELL_X4 FILLER_189_1758 ();
 FILLCELL_X32 FILLER_190_1 ();
 FILLCELL_X32 FILLER_190_33 ();
 FILLCELL_X32 FILLER_190_65 ();
 FILLCELL_X32 FILLER_190_97 ();
 FILLCELL_X32 FILLER_190_129 ();
 FILLCELL_X32 FILLER_190_161 ();
 FILLCELL_X32 FILLER_190_193 ();
 FILLCELL_X32 FILLER_190_225 ();
 FILLCELL_X32 FILLER_190_257 ();
 FILLCELL_X32 FILLER_190_289 ();
 FILLCELL_X32 FILLER_190_321 ();
 FILLCELL_X16 FILLER_190_353 ();
 FILLCELL_X8 FILLER_190_369 ();
 FILLCELL_X2 FILLER_190_377 ();
 FILLCELL_X1 FILLER_190_379 ();
 FILLCELL_X32 FILLER_190_1518 ();
 FILLCELL_X32 FILLER_190_1550 ();
 FILLCELL_X32 FILLER_190_1582 ();
 FILLCELL_X32 FILLER_190_1614 ();
 FILLCELL_X32 FILLER_190_1646 ();
 FILLCELL_X32 FILLER_190_1678 ();
 FILLCELL_X32 FILLER_190_1710 ();
 FILLCELL_X16 FILLER_190_1742 ();
 FILLCELL_X4 FILLER_190_1758 ();
 FILLCELL_X32 FILLER_191_1 ();
 FILLCELL_X32 FILLER_191_33 ();
 FILLCELL_X32 FILLER_191_65 ();
 FILLCELL_X32 FILLER_191_97 ();
 FILLCELL_X32 FILLER_191_129 ();
 FILLCELL_X32 FILLER_191_161 ();
 FILLCELL_X32 FILLER_191_193 ();
 FILLCELL_X32 FILLER_191_225 ();
 FILLCELL_X32 FILLER_191_257 ();
 FILLCELL_X32 FILLER_191_289 ();
 FILLCELL_X32 FILLER_191_321 ();
 FILLCELL_X16 FILLER_191_353 ();
 FILLCELL_X8 FILLER_191_369 ();
 FILLCELL_X2 FILLER_191_377 ();
 FILLCELL_X1 FILLER_191_379 ();
 FILLCELL_X32 FILLER_191_1518 ();
 FILLCELL_X32 FILLER_191_1550 ();
 FILLCELL_X32 FILLER_191_1582 ();
 FILLCELL_X32 FILLER_191_1614 ();
 FILLCELL_X32 FILLER_191_1646 ();
 FILLCELL_X32 FILLER_191_1678 ();
 FILLCELL_X32 FILLER_191_1710 ();
 FILLCELL_X16 FILLER_191_1742 ();
 FILLCELL_X4 FILLER_191_1758 ();
 FILLCELL_X32 FILLER_192_1 ();
 FILLCELL_X32 FILLER_192_33 ();
 FILLCELL_X32 FILLER_192_65 ();
 FILLCELL_X32 FILLER_192_97 ();
 FILLCELL_X32 FILLER_192_129 ();
 FILLCELL_X32 FILLER_192_161 ();
 FILLCELL_X32 FILLER_192_193 ();
 FILLCELL_X32 FILLER_192_225 ();
 FILLCELL_X32 FILLER_192_257 ();
 FILLCELL_X32 FILLER_192_289 ();
 FILLCELL_X32 FILLER_192_321 ();
 FILLCELL_X16 FILLER_192_353 ();
 FILLCELL_X8 FILLER_192_369 ();
 FILLCELL_X2 FILLER_192_377 ();
 FILLCELL_X1 FILLER_192_379 ();
 FILLCELL_X32 FILLER_192_1518 ();
 FILLCELL_X32 FILLER_192_1550 ();
 FILLCELL_X32 FILLER_192_1582 ();
 FILLCELL_X32 FILLER_192_1614 ();
 FILLCELL_X32 FILLER_192_1646 ();
 FILLCELL_X32 FILLER_192_1678 ();
 FILLCELL_X32 FILLER_192_1710 ();
 FILLCELL_X16 FILLER_192_1742 ();
 FILLCELL_X4 FILLER_192_1758 ();
 FILLCELL_X32 FILLER_193_1 ();
 FILLCELL_X32 FILLER_193_33 ();
 FILLCELL_X32 FILLER_193_65 ();
 FILLCELL_X32 FILLER_193_97 ();
 FILLCELL_X32 FILLER_193_129 ();
 FILLCELL_X32 FILLER_193_161 ();
 FILLCELL_X32 FILLER_193_193 ();
 FILLCELL_X32 FILLER_193_225 ();
 FILLCELL_X32 FILLER_193_257 ();
 FILLCELL_X32 FILLER_193_289 ();
 FILLCELL_X32 FILLER_193_321 ();
 FILLCELL_X16 FILLER_193_353 ();
 FILLCELL_X8 FILLER_193_369 ();
 FILLCELL_X2 FILLER_193_377 ();
 FILLCELL_X1 FILLER_193_379 ();
 FILLCELL_X32 FILLER_193_1518 ();
 FILLCELL_X32 FILLER_193_1550 ();
 FILLCELL_X32 FILLER_193_1582 ();
 FILLCELL_X32 FILLER_193_1614 ();
 FILLCELL_X32 FILLER_193_1646 ();
 FILLCELL_X32 FILLER_193_1678 ();
 FILLCELL_X32 FILLER_193_1710 ();
 FILLCELL_X16 FILLER_193_1742 ();
 FILLCELL_X4 FILLER_193_1758 ();
 FILLCELL_X32 FILLER_194_1 ();
 FILLCELL_X32 FILLER_194_33 ();
 FILLCELL_X32 FILLER_194_65 ();
 FILLCELL_X32 FILLER_194_97 ();
 FILLCELL_X32 FILLER_194_129 ();
 FILLCELL_X32 FILLER_194_161 ();
 FILLCELL_X32 FILLER_194_193 ();
 FILLCELL_X32 FILLER_194_225 ();
 FILLCELL_X32 FILLER_194_257 ();
 FILLCELL_X32 FILLER_194_289 ();
 FILLCELL_X32 FILLER_194_321 ();
 FILLCELL_X16 FILLER_194_353 ();
 FILLCELL_X8 FILLER_194_369 ();
 FILLCELL_X2 FILLER_194_377 ();
 FILLCELL_X1 FILLER_194_379 ();
 FILLCELL_X32 FILLER_194_1518 ();
 FILLCELL_X32 FILLER_194_1550 ();
 FILLCELL_X32 FILLER_194_1582 ();
 FILLCELL_X32 FILLER_194_1614 ();
 FILLCELL_X32 FILLER_194_1646 ();
 FILLCELL_X32 FILLER_194_1678 ();
 FILLCELL_X32 FILLER_194_1710 ();
 FILLCELL_X8 FILLER_194_1742 ();
 FILLCELL_X4 FILLER_194_1750 ();
 FILLCELL_X1 FILLER_194_1754 ();
 FILLCELL_X4 FILLER_194_1758 ();
 FILLCELL_X32 FILLER_195_1 ();
 FILLCELL_X32 FILLER_195_33 ();
 FILLCELL_X32 FILLER_195_65 ();
 FILLCELL_X32 FILLER_195_97 ();
 FILLCELL_X32 FILLER_195_129 ();
 FILLCELL_X32 FILLER_195_161 ();
 FILLCELL_X32 FILLER_195_193 ();
 FILLCELL_X32 FILLER_195_225 ();
 FILLCELL_X32 FILLER_195_257 ();
 FILLCELL_X32 FILLER_195_289 ();
 FILLCELL_X32 FILLER_195_321 ();
 FILLCELL_X16 FILLER_195_353 ();
 FILLCELL_X8 FILLER_195_369 ();
 FILLCELL_X2 FILLER_195_377 ();
 FILLCELL_X1 FILLER_195_379 ();
 FILLCELL_X32 FILLER_195_1518 ();
 FILLCELL_X32 FILLER_195_1550 ();
 FILLCELL_X32 FILLER_195_1582 ();
 FILLCELL_X32 FILLER_195_1614 ();
 FILLCELL_X32 FILLER_195_1646 ();
 FILLCELL_X32 FILLER_195_1678 ();
 FILLCELL_X32 FILLER_195_1710 ();
 FILLCELL_X16 FILLER_195_1742 ();
 FILLCELL_X4 FILLER_195_1758 ();
 FILLCELL_X32 FILLER_196_1 ();
 FILLCELL_X32 FILLER_196_33 ();
 FILLCELL_X32 FILLER_196_65 ();
 FILLCELL_X32 FILLER_196_97 ();
 FILLCELL_X32 FILLER_196_129 ();
 FILLCELL_X32 FILLER_196_161 ();
 FILLCELL_X32 FILLER_196_193 ();
 FILLCELL_X32 FILLER_196_225 ();
 FILLCELL_X32 FILLER_196_257 ();
 FILLCELL_X32 FILLER_196_289 ();
 FILLCELL_X32 FILLER_196_321 ();
 FILLCELL_X16 FILLER_196_353 ();
 FILLCELL_X8 FILLER_196_369 ();
 FILLCELL_X2 FILLER_196_377 ();
 FILLCELL_X1 FILLER_196_379 ();
 FILLCELL_X32 FILLER_196_1518 ();
 FILLCELL_X32 FILLER_196_1550 ();
 FILLCELL_X32 FILLER_196_1582 ();
 FILLCELL_X32 FILLER_196_1614 ();
 FILLCELL_X32 FILLER_196_1646 ();
 FILLCELL_X32 FILLER_196_1678 ();
 FILLCELL_X32 FILLER_196_1710 ();
 FILLCELL_X16 FILLER_196_1742 ();
 FILLCELL_X4 FILLER_196_1758 ();
 FILLCELL_X32 FILLER_197_1 ();
 FILLCELL_X32 FILLER_197_33 ();
 FILLCELL_X32 FILLER_197_65 ();
 FILLCELL_X32 FILLER_197_97 ();
 FILLCELL_X32 FILLER_197_129 ();
 FILLCELL_X32 FILLER_197_161 ();
 FILLCELL_X32 FILLER_197_193 ();
 FILLCELL_X32 FILLER_197_225 ();
 FILLCELL_X32 FILLER_197_257 ();
 FILLCELL_X32 FILLER_197_289 ();
 FILLCELL_X32 FILLER_197_321 ();
 FILLCELL_X16 FILLER_197_353 ();
 FILLCELL_X8 FILLER_197_369 ();
 FILLCELL_X2 FILLER_197_377 ();
 FILLCELL_X1 FILLER_197_379 ();
 FILLCELL_X32 FILLER_197_1518 ();
 FILLCELL_X32 FILLER_197_1550 ();
 FILLCELL_X32 FILLER_197_1582 ();
 FILLCELL_X32 FILLER_197_1614 ();
 FILLCELL_X32 FILLER_197_1646 ();
 FILLCELL_X32 FILLER_197_1678 ();
 FILLCELL_X32 FILLER_197_1710 ();
 FILLCELL_X16 FILLER_197_1742 ();
 FILLCELL_X4 FILLER_197_1758 ();
 FILLCELL_X4 FILLER_198_1 ();
 FILLCELL_X32 FILLER_198_8 ();
 FILLCELL_X32 FILLER_198_40 ();
 FILLCELL_X32 FILLER_198_72 ();
 FILLCELL_X32 FILLER_198_104 ();
 FILLCELL_X32 FILLER_198_136 ();
 FILLCELL_X32 FILLER_198_168 ();
 FILLCELL_X32 FILLER_198_200 ();
 FILLCELL_X32 FILLER_198_232 ();
 FILLCELL_X32 FILLER_198_264 ();
 FILLCELL_X32 FILLER_198_296 ();
 FILLCELL_X32 FILLER_198_328 ();
 FILLCELL_X16 FILLER_198_360 ();
 FILLCELL_X4 FILLER_198_376 ();
 FILLCELL_X32 FILLER_198_1518 ();
 FILLCELL_X32 FILLER_198_1550 ();
 FILLCELL_X32 FILLER_198_1582 ();
 FILLCELL_X32 FILLER_198_1614 ();
 FILLCELL_X32 FILLER_198_1646 ();
 FILLCELL_X32 FILLER_198_1678 ();
 FILLCELL_X32 FILLER_198_1710 ();
 FILLCELL_X16 FILLER_198_1742 ();
 FILLCELL_X4 FILLER_198_1758 ();
 FILLCELL_X32 FILLER_199_1 ();
 FILLCELL_X32 FILLER_199_33 ();
 FILLCELL_X32 FILLER_199_65 ();
 FILLCELL_X32 FILLER_199_97 ();
 FILLCELL_X32 FILLER_199_129 ();
 FILLCELL_X32 FILLER_199_161 ();
 FILLCELL_X32 FILLER_199_193 ();
 FILLCELL_X32 FILLER_199_225 ();
 FILLCELL_X32 FILLER_199_257 ();
 FILLCELL_X32 FILLER_199_289 ();
 FILLCELL_X32 FILLER_199_321 ();
 FILLCELL_X16 FILLER_199_353 ();
 FILLCELL_X8 FILLER_199_369 ();
 FILLCELL_X2 FILLER_199_377 ();
 FILLCELL_X1 FILLER_199_379 ();
 FILLCELL_X32 FILLER_199_1518 ();
 FILLCELL_X32 FILLER_199_1550 ();
 FILLCELL_X32 FILLER_199_1582 ();
 FILLCELL_X32 FILLER_199_1614 ();
 FILLCELL_X32 FILLER_199_1646 ();
 FILLCELL_X32 FILLER_199_1678 ();
 FILLCELL_X32 FILLER_199_1710 ();
 FILLCELL_X16 FILLER_199_1742 ();
 FILLCELL_X4 FILLER_199_1758 ();
 FILLCELL_X32 FILLER_200_1 ();
 FILLCELL_X32 FILLER_200_33 ();
 FILLCELL_X32 FILLER_200_65 ();
 FILLCELL_X32 FILLER_200_97 ();
 FILLCELL_X32 FILLER_200_129 ();
 FILLCELL_X32 FILLER_200_161 ();
 FILLCELL_X32 FILLER_200_193 ();
 FILLCELL_X32 FILLER_200_225 ();
 FILLCELL_X32 FILLER_200_257 ();
 FILLCELL_X32 FILLER_200_289 ();
 FILLCELL_X32 FILLER_200_321 ();
 FILLCELL_X16 FILLER_200_353 ();
 FILLCELL_X8 FILLER_200_369 ();
 FILLCELL_X2 FILLER_200_377 ();
 FILLCELL_X1 FILLER_200_379 ();
 FILLCELL_X32 FILLER_200_1518 ();
 FILLCELL_X32 FILLER_200_1550 ();
 FILLCELL_X32 FILLER_200_1582 ();
 FILLCELL_X32 FILLER_200_1614 ();
 FILLCELL_X32 FILLER_200_1646 ();
 FILLCELL_X32 FILLER_200_1678 ();
 FILLCELL_X32 FILLER_200_1710 ();
 FILLCELL_X16 FILLER_200_1742 ();
 FILLCELL_X4 FILLER_200_1758 ();
 FILLCELL_X32 FILLER_201_1 ();
 FILLCELL_X32 FILLER_201_33 ();
 FILLCELL_X32 FILLER_201_65 ();
 FILLCELL_X32 FILLER_201_97 ();
 FILLCELL_X32 FILLER_201_129 ();
 FILLCELL_X32 FILLER_201_161 ();
 FILLCELL_X32 FILLER_201_193 ();
 FILLCELL_X32 FILLER_201_225 ();
 FILLCELL_X32 FILLER_201_257 ();
 FILLCELL_X32 FILLER_201_289 ();
 FILLCELL_X32 FILLER_201_321 ();
 FILLCELL_X16 FILLER_201_353 ();
 FILLCELL_X8 FILLER_201_369 ();
 FILLCELL_X2 FILLER_201_377 ();
 FILLCELL_X1 FILLER_201_379 ();
 FILLCELL_X32 FILLER_201_1518 ();
 FILLCELL_X32 FILLER_201_1550 ();
 FILLCELL_X32 FILLER_201_1582 ();
 FILLCELL_X32 FILLER_201_1614 ();
 FILLCELL_X32 FILLER_201_1646 ();
 FILLCELL_X32 FILLER_201_1678 ();
 FILLCELL_X32 FILLER_201_1710 ();
 FILLCELL_X16 FILLER_201_1742 ();
 FILLCELL_X4 FILLER_201_1758 ();
 FILLCELL_X32 FILLER_202_1 ();
 FILLCELL_X32 FILLER_202_33 ();
 FILLCELL_X32 FILLER_202_65 ();
 FILLCELL_X32 FILLER_202_97 ();
 FILLCELL_X32 FILLER_202_129 ();
 FILLCELL_X32 FILLER_202_161 ();
 FILLCELL_X32 FILLER_202_193 ();
 FILLCELL_X32 FILLER_202_225 ();
 FILLCELL_X32 FILLER_202_257 ();
 FILLCELL_X32 FILLER_202_289 ();
 FILLCELL_X32 FILLER_202_321 ();
 FILLCELL_X16 FILLER_202_353 ();
 FILLCELL_X8 FILLER_202_369 ();
 FILLCELL_X2 FILLER_202_377 ();
 FILLCELL_X1 FILLER_202_379 ();
 FILLCELL_X32 FILLER_202_1518 ();
 FILLCELL_X32 FILLER_202_1550 ();
 FILLCELL_X32 FILLER_202_1582 ();
 FILLCELL_X32 FILLER_202_1614 ();
 FILLCELL_X32 FILLER_202_1646 ();
 FILLCELL_X32 FILLER_202_1678 ();
 FILLCELL_X32 FILLER_202_1710 ();
 FILLCELL_X16 FILLER_202_1742 ();
 FILLCELL_X4 FILLER_202_1758 ();
 FILLCELL_X32 FILLER_203_1 ();
 FILLCELL_X32 FILLER_203_33 ();
 FILLCELL_X32 FILLER_203_65 ();
 FILLCELL_X32 FILLER_203_97 ();
 FILLCELL_X32 FILLER_203_129 ();
 FILLCELL_X32 FILLER_203_161 ();
 FILLCELL_X32 FILLER_203_193 ();
 FILLCELL_X32 FILLER_203_225 ();
 FILLCELL_X32 FILLER_203_257 ();
 FILLCELL_X32 FILLER_203_289 ();
 FILLCELL_X32 FILLER_203_321 ();
 FILLCELL_X16 FILLER_203_353 ();
 FILLCELL_X8 FILLER_203_369 ();
 FILLCELL_X2 FILLER_203_377 ();
 FILLCELL_X1 FILLER_203_379 ();
 FILLCELL_X32 FILLER_203_1518 ();
 FILLCELL_X32 FILLER_203_1550 ();
 FILLCELL_X32 FILLER_203_1582 ();
 FILLCELL_X32 FILLER_203_1614 ();
 FILLCELL_X32 FILLER_203_1646 ();
 FILLCELL_X32 FILLER_203_1678 ();
 FILLCELL_X32 FILLER_203_1710 ();
 FILLCELL_X8 FILLER_203_1742 ();
 FILLCELL_X4 FILLER_203_1750 ();
 FILLCELL_X1 FILLER_203_1754 ();
 FILLCELL_X4 FILLER_203_1758 ();
 FILLCELL_X32 FILLER_204_1 ();
 FILLCELL_X32 FILLER_204_33 ();
 FILLCELL_X32 FILLER_204_65 ();
 FILLCELL_X32 FILLER_204_97 ();
 FILLCELL_X32 FILLER_204_129 ();
 FILLCELL_X32 FILLER_204_161 ();
 FILLCELL_X32 FILLER_204_193 ();
 FILLCELL_X32 FILLER_204_225 ();
 FILLCELL_X32 FILLER_204_257 ();
 FILLCELL_X32 FILLER_204_289 ();
 FILLCELL_X32 FILLER_204_321 ();
 FILLCELL_X16 FILLER_204_353 ();
 FILLCELL_X8 FILLER_204_369 ();
 FILLCELL_X2 FILLER_204_377 ();
 FILLCELL_X1 FILLER_204_379 ();
 FILLCELL_X32 FILLER_204_1518 ();
 FILLCELL_X32 FILLER_204_1550 ();
 FILLCELL_X32 FILLER_204_1582 ();
 FILLCELL_X32 FILLER_204_1614 ();
 FILLCELL_X32 FILLER_204_1646 ();
 FILLCELL_X32 FILLER_204_1678 ();
 FILLCELL_X32 FILLER_204_1710 ();
 FILLCELL_X16 FILLER_204_1742 ();
 FILLCELL_X4 FILLER_204_1758 ();
 FILLCELL_X32 FILLER_205_1 ();
 FILLCELL_X32 FILLER_205_33 ();
 FILLCELL_X32 FILLER_205_65 ();
 FILLCELL_X32 FILLER_205_97 ();
 FILLCELL_X32 FILLER_205_129 ();
 FILLCELL_X32 FILLER_205_161 ();
 FILLCELL_X32 FILLER_205_193 ();
 FILLCELL_X32 FILLER_205_225 ();
 FILLCELL_X32 FILLER_205_257 ();
 FILLCELL_X32 FILLER_205_289 ();
 FILLCELL_X32 FILLER_205_321 ();
 FILLCELL_X16 FILLER_205_353 ();
 FILLCELL_X8 FILLER_205_369 ();
 FILLCELL_X2 FILLER_205_377 ();
 FILLCELL_X1 FILLER_205_379 ();
 FILLCELL_X32 FILLER_205_1518 ();
 FILLCELL_X32 FILLER_205_1550 ();
 FILLCELL_X32 FILLER_205_1582 ();
 FILLCELL_X32 FILLER_205_1614 ();
 FILLCELL_X32 FILLER_205_1646 ();
 FILLCELL_X32 FILLER_205_1678 ();
 FILLCELL_X32 FILLER_205_1710 ();
 FILLCELL_X16 FILLER_205_1742 ();
 FILLCELL_X4 FILLER_205_1758 ();
 FILLCELL_X32 FILLER_206_1 ();
 FILLCELL_X32 FILLER_206_33 ();
 FILLCELL_X32 FILLER_206_65 ();
 FILLCELL_X32 FILLER_206_97 ();
 FILLCELL_X32 FILLER_206_129 ();
 FILLCELL_X32 FILLER_206_161 ();
 FILLCELL_X32 FILLER_206_193 ();
 FILLCELL_X32 FILLER_206_225 ();
 FILLCELL_X32 FILLER_206_257 ();
 FILLCELL_X32 FILLER_206_289 ();
 FILLCELL_X32 FILLER_206_321 ();
 FILLCELL_X16 FILLER_206_353 ();
 FILLCELL_X8 FILLER_206_369 ();
 FILLCELL_X2 FILLER_206_377 ();
 FILLCELL_X1 FILLER_206_379 ();
 FILLCELL_X32 FILLER_206_1518 ();
 FILLCELL_X32 FILLER_206_1550 ();
 FILLCELL_X32 FILLER_206_1582 ();
 FILLCELL_X32 FILLER_206_1614 ();
 FILLCELL_X32 FILLER_206_1646 ();
 FILLCELL_X32 FILLER_206_1678 ();
 FILLCELL_X32 FILLER_206_1710 ();
 FILLCELL_X16 FILLER_206_1742 ();
 FILLCELL_X4 FILLER_206_1758 ();
 FILLCELL_X32 FILLER_207_1 ();
 FILLCELL_X32 FILLER_207_33 ();
 FILLCELL_X32 FILLER_207_65 ();
 FILLCELL_X32 FILLER_207_97 ();
 FILLCELL_X32 FILLER_207_129 ();
 FILLCELL_X32 FILLER_207_161 ();
 FILLCELL_X32 FILLER_207_193 ();
 FILLCELL_X32 FILLER_207_225 ();
 FILLCELL_X32 FILLER_207_257 ();
 FILLCELL_X32 FILLER_207_289 ();
 FILLCELL_X32 FILLER_207_321 ();
 FILLCELL_X16 FILLER_207_353 ();
 FILLCELL_X8 FILLER_207_369 ();
 FILLCELL_X2 FILLER_207_377 ();
 FILLCELL_X1 FILLER_207_379 ();
 FILLCELL_X32 FILLER_207_1518 ();
 FILLCELL_X32 FILLER_207_1550 ();
 FILLCELL_X32 FILLER_207_1582 ();
 FILLCELL_X32 FILLER_207_1614 ();
 FILLCELL_X32 FILLER_207_1646 ();
 FILLCELL_X32 FILLER_207_1678 ();
 FILLCELL_X32 FILLER_207_1710 ();
 FILLCELL_X16 FILLER_207_1742 ();
 FILLCELL_X4 FILLER_207_1758 ();
 FILLCELL_X4 FILLER_208_1 ();
 FILLCELL_X32 FILLER_208_12 ();
 FILLCELL_X32 FILLER_208_44 ();
 FILLCELL_X32 FILLER_208_76 ();
 FILLCELL_X32 FILLER_208_108 ();
 FILLCELL_X32 FILLER_208_140 ();
 FILLCELL_X32 FILLER_208_172 ();
 FILLCELL_X32 FILLER_208_204 ();
 FILLCELL_X32 FILLER_208_236 ();
 FILLCELL_X32 FILLER_208_268 ();
 FILLCELL_X32 FILLER_208_300 ();
 FILLCELL_X32 FILLER_208_332 ();
 FILLCELL_X32 FILLER_208_364 ();
 FILLCELL_X32 FILLER_208_396 ();
 FILLCELL_X32 FILLER_208_428 ();
 FILLCELL_X32 FILLER_208_460 ();
 FILLCELL_X32 FILLER_208_492 ();
 FILLCELL_X32 FILLER_208_524 ();
 FILLCELL_X32 FILLER_208_556 ();
 FILLCELL_X32 FILLER_208_588 ();
 FILLCELL_X8 FILLER_208_620 ();
 FILLCELL_X2 FILLER_208_628 ();
 FILLCELL_X1 FILLER_208_630 ();
 FILLCELL_X32 FILLER_208_632 ();
 FILLCELL_X32 FILLER_208_664 ();
 FILLCELL_X32 FILLER_208_696 ();
 FILLCELL_X32 FILLER_208_728 ();
 FILLCELL_X32 FILLER_208_760 ();
 FILLCELL_X32 FILLER_208_792 ();
 FILLCELL_X32 FILLER_208_824 ();
 FILLCELL_X32 FILLER_208_856 ();
 FILLCELL_X32 FILLER_208_888 ();
 FILLCELL_X32 FILLER_208_920 ();
 FILLCELL_X32 FILLER_208_952 ();
 FILLCELL_X32 FILLER_208_984 ();
 FILLCELL_X32 FILLER_208_1016 ();
 FILLCELL_X32 FILLER_208_1048 ();
 FILLCELL_X32 FILLER_208_1080 ();
 FILLCELL_X32 FILLER_208_1112 ();
 FILLCELL_X32 FILLER_208_1144 ();
 FILLCELL_X32 FILLER_208_1176 ();
 FILLCELL_X32 FILLER_208_1208 ();
 FILLCELL_X16 FILLER_208_1240 ();
 FILLCELL_X4 FILLER_208_1256 ();
 FILLCELL_X2 FILLER_208_1260 ();
 FILLCELL_X32 FILLER_208_1263 ();
 FILLCELL_X32 FILLER_208_1295 ();
 FILLCELL_X32 FILLER_208_1327 ();
 FILLCELL_X32 FILLER_208_1359 ();
 FILLCELL_X32 FILLER_208_1391 ();
 FILLCELL_X32 FILLER_208_1423 ();
 FILLCELL_X32 FILLER_208_1455 ();
 FILLCELL_X32 FILLER_208_1487 ();
 FILLCELL_X32 FILLER_208_1519 ();
 FILLCELL_X32 FILLER_208_1551 ();
 FILLCELL_X32 FILLER_208_1583 ();
 FILLCELL_X32 FILLER_208_1615 ();
 FILLCELL_X32 FILLER_208_1647 ();
 FILLCELL_X32 FILLER_208_1679 ();
 FILLCELL_X32 FILLER_208_1711 ();
 FILLCELL_X16 FILLER_208_1743 ();
 FILLCELL_X2 FILLER_208_1759 ();
 FILLCELL_X1 FILLER_208_1761 ();
 FILLCELL_X32 FILLER_209_1 ();
 FILLCELL_X32 FILLER_209_33 ();
 FILLCELL_X32 FILLER_209_65 ();
 FILLCELL_X32 FILLER_209_97 ();
 FILLCELL_X32 FILLER_209_129 ();
 FILLCELL_X32 FILLER_209_161 ();
 FILLCELL_X32 FILLER_209_193 ();
 FILLCELL_X32 FILLER_209_225 ();
 FILLCELL_X32 FILLER_209_257 ();
 FILLCELL_X32 FILLER_209_289 ();
 FILLCELL_X32 FILLER_209_321 ();
 FILLCELL_X32 FILLER_209_353 ();
 FILLCELL_X32 FILLER_209_385 ();
 FILLCELL_X32 FILLER_209_417 ();
 FILLCELL_X32 FILLER_209_449 ();
 FILLCELL_X32 FILLER_209_481 ();
 FILLCELL_X32 FILLER_209_513 ();
 FILLCELL_X32 FILLER_209_545 ();
 FILLCELL_X32 FILLER_209_577 ();
 FILLCELL_X32 FILLER_209_609 ();
 FILLCELL_X32 FILLER_209_641 ();
 FILLCELL_X32 FILLER_209_673 ();
 FILLCELL_X32 FILLER_209_705 ();
 FILLCELL_X32 FILLER_209_737 ();
 FILLCELL_X32 FILLER_209_769 ();
 FILLCELL_X32 FILLER_209_801 ();
 FILLCELL_X32 FILLER_209_833 ();
 FILLCELL_X32 FILLER_209_865 ();
 FILLCELL_X32 FILLER_209_897 ();
 FILLCELL_X32 FILLER_209_929 ();
 FILLCELL_X32 FILLER_209_961 ();
 FILLCELL_X32 FILLER_209_993 ();
 FILLCELL_X32 FILLER_209_1025 ();
 FILLCELL_X32 FILLER_209_1057 ();
 FILLCELL_X32 FILLER_209_1089 ();
 FILLCELL_X32 FILLER_209_1121 ();
 FILLCELL_X32 FILLER_209_1153 ();
 FILLCELL_X32 FILLER_209_1185 ();
 FILLCELL_X32 FILLER_209_1217 ();
 FILLCELL_X8 FILLER_209_1249 ();
 FILLCELL_X4 FILLER_209_1257 ();
 FILLCELL_X2 FILLER_209_1261 ();
 FILLCELL_X32 FILLER_209_1264 ();
 FILLCELL_X32 FILLER_209_1296 ();
 FILLCELL_X32 FILLER_209_1328 ();
 FILLCELL_X32 FILLER_209_1360 ();
 FILLCELL_X32 FILLER_209_1392 ();
 FILLCELL_X32 FILLER_209_1424 ();
 FILLCELL_X32 FILLER_209_1456 ();
 FILLCELL_X32 FILLER_209_1488 ();
 FILLCELL_X32 FILLER_209_1520 ();
 FILLCELL_X32 FILLER_209_1552 ();
 FILLCELL_X32 FILLER_209_1584 ();
 FILLCELL_X32 FILLER_209_1616 ();
 FILLCELL_X32 FILLER_209_1648 ();
 FILLCELL_X32 FILLER_209_1680 ();
 FILLCELL_X32 FILLER_209_1712 ();
 FILLCELL_X16 FILLER_209_1744 ();
 FILLCELL_X2 FILLER_209_1760 ();
 FILLCELL_X32 FILLER_210_1 ();
 FILLCELL_X32 FILLER_210_33 ();
 FILLCELL_X32 FILLER_210_65 ();
 FILLCELL_X32 FILLER_210_97 ();
 FILLCELL_X32 FILLER_210_129 ();
 FILLCELL_X32 FILLER_210_161 ();
 FILLCELL_X32 FILLER_210_193 ();
 FILLCELL_X32 FILLER_210_225 ();
 FILLCELL_X32 FILLER_210_257 ();
 FILLCELL_X32 FILLER_210_289 ();
 FILLCELL_X32 FILLER_210_321 ();
 FILLCELL_X32 FILLER_210_353 ();
 FILLCELL_X32 FILLER_210_385 ();
 FILLCELL_X32 FILLER_210_417 ();
 FILLCELL_X32 FILLER_210_449 ();
 FILLCELL_X32 FILLER_210_481 ();
 FILLCELL_X32 FILLER_210_513 ();
 FILLCELL_X32 FILLER_210_545 ();
 FILLCELL_X32 FILLER_210_577 ();
 FILLCELL_X16 FILLER_210_609 ();
 FILLCELL_X4 FILLER_210_625 ();
 FILLCELL_X2 FILLER_210_629 ();
 FILLCELL_X32 FILLER_210_632 ();
 FILLCELL_X32 FILLER_210_664 ();
 FILLCELL_X32 FILLER_210_696 ();
 FILLCELL_X32 FILLER_210_728 ();
 FILLCELL_X32 FILLER_210_760 ();
 FILLCELL_X32 FILLER_210_792 ();
 FILLCELL_X32 FILLER_210_824 ();
 FILLCELL_X32 FILLER_210_856 ();
 FILLCELL_X32 FILLER_210_888 ();
 FILLCELL_X32 FILLER_210_920 ();
 FILLCELL_X32 FILLER_210_952 ();
 FILLCELL_X32 FILLER_210_984 ();
 FILLCELL_X32 FILLER_210_1016 ();
 FILLCELL_X32 FILLER_210_1048 ();
 FILLCELL_X32 FILLER_210_1080 ();
 FILLCELL_X32 FILLER_210_1112 ();
 FILLCELL_X32 FILLER_210_1144 ();
 FILLCELL_X32 FILLER_210_1176 ();
 FILLCELL_X32 FILLER_210_1208 ();
 FILLCELL_X32 FILLER_210_1240 ();
 FILLCELL_X32 FILLER_210_1272 ();
 FILLCELL_X32 FILLER_210_1304 ();
 FILLCELL_X32 FILLER_210_1336 ();
 FILLCELL_X32 FILLER_210_1368 ();
 FILLCELL_X32 FILLER_210_1400 ();
 FILLCELL_X32 FILLER_210_1432 ();
 FILLCELL_X32 FILLER_210_1464 ();
 FILLCELL_X32 FILLER_210_1496 ();
 FILLCELL_X32 FILLER_210_1528 ();
 FILLCELL_X32 FILLER_210_1560 ();
 FILLCELL_X32 FILLER_210_1592 ();
 FILLCELL_X32 FILLER_210_1624 ();
 FILLCELL_X32 FILLER_210_1656 ();
 FILLCELL_X32 FILLER_210_1688 ();
 FILLCELL_X32 FILLER_210_1720 ();
 FILLCELL_X8 FILLER_210_1752 ();
 FILLCELL_X2 FILLER_210_1760 ();
 FILLCELL_X32 FILLER_211_1 ();
 FILLCELL_X32 FILLER_211_33 ();
 FILLCELL_X32 FILLER_211_65 ();
 FILLCELL_X32 FILLER_211_97 ();
 FILLCELL_X32 FILLER_211_129 ();
 FILLCELL_X32 FILLER_211_161 ();
 FILLCELL_X32 FILLER_211_193 ();
 FILLCELL_X32 FILLER_211_225 ();
 FILLCELL_X32 FILLER_211_257 ();
 FILLCELL_X32 FILLER_211_289 ();
 FILLCELL_X32 FILLER_211_321 ();
 FILLCELL_X32 FILLER_211_353 ();
 FILLCELL_X32 FILLER_211_385 ();
 FILLCELL_X32 FILLER_211_417 ();
 FILLCELL_X32 FILLER_211_449 ();
 FILLCELL_X32 FILLER_211_481 ();
 FILLCELL_X32 FILLER_211_513 ();
 FILLCELL_X32 FILLER_211_545 ();
 FILLCELL_X32 FILLER_211_577 ();
 FILLCELL_X32 FILLER_211_609 ();
 FILLCELL_X32 FILLER_211_641 ();
 FILLCELL_X32 FILLER_211_673 ();
 FILLCELL_X32 FILLER_211_705 ();
 FILLCELL_X32 FILLER_211_737 ();
 FILLCELL_X32 FILLER_211_769 ();
 FILLCELL_X32 FILLER_211_801 ();
 FILLCELL_X32 FILLER_211_833 ();
 FILLCELL_X32 FILLER_211_865 ();
 FILLCELL_X32 FILLER_211_897 ();
 FILLCELL_X32 FILLER_211_929 ();
 FILLCELL_X32 FILLER_211_961 ();
 FILLCELL_X32 FILLER_211_993 ();
 FILLCELL_X32 FILLER_211_1025 ();
 FILLCELL_X32 FILLER_211_1057 ();
 FILLCELL_X32 FILLER_211_1089 ();
 FILLCELL_X32 FILLER_211_1121 ();
 FILLCELL_X32 FILLER_211_1153 ();
 FILLCELL_X32 FILLER_211_1185 ();
 FILLCELL_X32 FILLER_211_1217 ();
 FILLCELL_X8 FILLER_211_1249 ();
 FILLCELL_X4 FILLER_211_1257 ();
 FILLCELL_X2 FILLER_211_1261 ();
 FILLCELL_X32 FILLER_211_1264 ();
 FILLCELL_X32 FILLER_211_1296 ();
 FILLCELL_X32 FILLER_211_1328 ();
 FILLCELL_X32 FILLER_211_1360 ();
 FILLCELL_X32 FILLER_211_1392 ();
 FILLCELL_X32 FILLER_211_1424 ();
 FILLCELL_X32 FILLER_211_1456 ();
 FILLCELL_X32 FILLER_211_1488 ();
 FILLCELL_X32 FILLER_211_1520 ();
 FILLCELL_X32 FILLER_211_1552 ();
 FILLCELL_X32 FILLER_211_1584 ();
 FILLCELL_X32 FILLER_211_1616 ();
 FILLCELL_X32 FILLER_211_1648 ();
 FILLCELL_X32 FILLER_211_1680 ();
 FILLCELL_X32 FILLER_211_1712 ();
 FILLCELL_X16 FILLER_211_1744 ();
 FILLCELL_X2 FILLER_211_1760 ();
 FILLCELL_X32 FILLER_212_1 ();
 FILLCELL_X32 FILLER_212_33 ();
 FILLCELL_X32 FILLER_212_65 ();
 FILLCELL_X32 FILLER_212_97 ();
 FILLCELL_X32 FILLER_212_129 ();
 FILLCELL_X32 FILLER_212_161 ();
 FILLCELL_X32 FILLER_212_193 ();
 FILLCELL_X32 FILLER_212_225 ();
 FILLCELL_X32 FILLER_212_257 ();
 FILLCELL_X32 FILLER_212_289 ();
 FILLCELL_X32 FILLER_212_321 ();
 FILLCELL_X32 FILLER_212_353 ();
 FILLCELL_X32 FILLER_212_385 ();
 FILLCELL_X32 FILLER_212_417 ();
 FILLCELL_X32 FILLER_212_449 ();
 FILLCELL_X32 FILLER_212_481 ();
 FILLCELL_X32 FILLER_212_513 ();
 FILLCELL_X32 FILLER_212_545 ();
 FILLCELL_X32 FILLER_212_577 ();
 FILLCELL_X16 FILLER_212_609 ();
 FILLCELL_X4 FILLER_212_625 ();
 FILLCELL_X2 FILLER_212_629 ();
 FILLCELL_X32 FILLER_212_632 ();
 FILLCELL_X32 FILLER_212_664 ();
 FILLCELL_X32 FILLER_212_696 ();
 FILLCELL_X32 FILLER_212_728 ();
 FILLCELL_X32 FILLER_212_760 ();
 FILLCELL_X32 FILLER_212_792 ();
 FILLCELL_X32 FILLER_212_824 ();
 FILLCELL_X32 FILLER_212_856 ();
 FILLCELL_X32 FILLER_212_888 ();
 FILLCELL_X32 FILLER_212_920 ();
 FILLCELL_X32 FILLER_212_952 ();
 FILLCELL_X32 FILLER_212_984 ();
 FILLCELL_X32 FILLER_212_1016 ();
 FILLCELL_X32 FILLER_212_1048 ();
 FILLCELL_X32 FILLER_212_1080 ();
 FILLCELL_X32 FILLER_212_1112 ();
 FILLCELL_X32 FILLER_212_1144 ();
 FILLCELL_X32 FILLER_212_1176 ();
 FILLCELL_X32 FILLER_212_1208 ();
 FILLCELL_X32 FILLER_212_1240 ();
 FILLCELL_X32 FILLER_212_1272 ();
 FILLCELL_X32 FILLER_212_1304 ();
 FILLCELL_X32 FILLER_212_1336 ();
 FILLCELL_X32 FILLER_212_1368 ();
 FILLCELL_X32 FILLER_212_1400 ();
 FILLCELL_X32 FILLER_212_1432 ();
 FILLCELL_X32 FILLER_212_1464 ();
 FILLCELL_X32 FILLER_212_1496 ();
 FILLCELL_X32 FILLER_212_1528 ();
 FILLCELL_X32 FILLER_212_1560 ();
 FILLCELL_X32 FILLER_212_1592 ();
 FILLCELL_X32 FILLER_212_1624 ();
 FILLCELL_X32 FILLER_212_1656 ();
 FILLCELL_X32 FILLER_212_1688 ();
 FILLCELL_X32 FILLER_212_1720 ();
 FILLCELL_X8 FILLER_212_1752 ();
 FILLCELL_X2 FILLER_212_1760 ();
 FILLCELL_X32 FILLER_213_1 ();
 FILLCELL_X32 FILLER_213_33 ();
 FILLCELL_X32 FILLER_213_65 ();
 FILLCELL_X32 FILLER_213_97 ();
 FILLCELL_X32 FILLER_213_129 ();
 FILLCELL_X32 FILLER_213_161 ();
 FILLCELL_X32 FILLER_213_193 ();
 FILLCELL_X32 FILLER_213_225 ();
 FILLCELL_X32 FILLER_213_257 ();
 FILLCELL_X32 FILLER_213_289 ();
 FILLCELL_X32 FILLER_213_321 ();
 FILLCELL_X32 FILLER_213_353 ();
 FILLCELL_X32 FILLER_213_385 ();
 FILLCELL_X32 FILLER_213_417 ();
 FILLCELL_X32 FILLER_213_449 ();
 FILLCELL_X32 FILLER_213_481 ();
 FILLCELL_X32 FILLER_213_513 ();
 FILLCELL_X32 FILLER_213_545 ();
 FILLCELL_X32 FILLER_213_577 ();
 FILLCELL_X32 FILLER_213_609 ();
 FILLCELL_X32 FILLER_213_641 ();
 FILLCELL_X32 FILLER_213_673 ();
 FILLCELL_X32 FILLER_213_705 ();
 FILLCELL_X32 FILLER_213_737 ();
 FILLCELL_X32 FILLER_213_769 ();
 FILLCELL_X32 FILLER_213_801 ();
 FILLCELL_X32 FILLER_213_833 ();
 FILLCELL_X32 FILLER_213_865 ();
 FILLCELL_X32 FILLER_213_897 ();
 FILLCELL_X32 FILLER_213_929 ();
 FILLCELL_X32 FILLER_213_961 ();
 FILLCELL_X32 FILLER_213_993 ();
 FILLCELL_X32 FILLER_213_1025 ();
 FILLCELL_X32 FILLER_213_1057 ();
 FILLCELL_X32 FILLER_213_1089 ();
 FILLCELL_X32 FILLER_213_1121 ();
 FILLCELL_X32 FILLER_213_1153 ();
 FILLCELL_X32 FILLER_213_1185 ();
 FILLCELL_X32 FILLER_213_1217 ();
 FILLCELL_X8 FILLER_213_1249 ();
 FILLCELL_X4 FILLER_213_1257 ();
 FILLCELL_X2 FILLER_213_1261 ();
 FILLCELL_X32 FILLER_213_1264 ();
 FILLCELL_X32 FILLER_213_1296 ();
 FILLCELL_X32 FILLER_213_1328 ();
 FILLCELL_X32 FILLER_213_1360 ();
 FILLCELL_X32 FILLER_213_1392 ();
 FILLCELL_X32 FILLER_213_1424 ();
 FILLCELL_X32 FILLER_213_1456 ();
 FILLCELL_X32 FILLER_213_1488 ();
 FILLCELL_X32 FILLER_213_1520 ();
 FILLCELL_X32 FILLER_213_1552 ();
 FILLCELL_X32 FILLER_213_1584 ();
 FILLCELL_X32 FILLER_213_1616 ();
 FILLCELL_X32 FILLER_213_1648 ();
 FILLCELL_X32 FILLER_213_1680 ();
 FILLCELL_X32 FILLER_213_1712 ();
 FILLCELL_X4 FILLER_213_1744 ();
 FILLCELL_X2 FILLER_213_1748 ();
 FILLCELL_X1 FILLER_213_1750 ();
 FILLCELL_X4 FILLER_213_1758 ();
 FILLCELL_X32 FILLER_214_1 ();
 FILLCELL_X32 FILLER_214_33 ();
 FILLCELL_X32 FILLER_214_65 ();
 FILLCELL_X32 FILLER_214_97 ();
 FILLCELL_X32 FILLER_214_129 ();
 FILLCELL_X32 FILLER_214_161 ();
 FILLCELL_X32 FILLER_214_193 ();
 FILLCELL_X32 FILLER_214_225 ();
 FILLCELL_X32 FILLER_214_257 ();
 FILLCELL_X32 FILLER_214_289 ();
 FILLCELL_X32 FILLER_214_321 ();
 FILLCELL_X32 FILLER_214_353 ();
 FILLCELL_X32 FILLER_214_385 ();
 FILLCELL_X32 FILLER_214_417 ();
 FILLCELL_X32 FILLER_214_449 ();
 FILLCELL_X32 FILLER_214_481 ();
 FILLCELL_X32 FILLER_214_513 ();
 FILLCELL_X32 FILLER_214_545 ();
 FILLCELL_X32 FILLER_214_577 ();
 FILLCELL_X16 FILLER_214_609 ();
 FILLCELL_X4 FILLER_214_625 ();
 FILLCELL_X2 FILLER_214_629 ();
 FILLCELL_X32 FILLER_214_632 ();
 FILLCELL_X32 FILLER_214_664 ();
 FILLCELL_X32 FILLER_214_696 ();
 FILLCELL_X32 FILLER_214_728 ();
 FILLCELL_X32 FILLER_214_760 ();
 FILLCELL_X32 FILLER_214_792 ();
 FILLCELL_X32 FILLER_214_824 ();
 FILLCELL_X32 FILLER_214_856 ();
 FILLCELL_X32 FILLER_214_888 ();
 FILLCELL_X32 FILLER_214_920 ();
 FILLCELL_X32 FILLER_214_952 ();
 FILLCELL_X32 FILLER_214_984 ();
 FILLCELL_X32 FILLER_214_1016 ();
 FILLCELL_X32 FILLER_214_1048 ();
 FILLCELL_X32 FILLER_214_1080 ();
 FILLCELL_X32 FILLER_214_1112 ();
 FILLCELL_X32 FILLER_214_1144 ();
 FILLCELL_X32 FILLER_214_1176 ();
 FILLCELL_X32 FILLER_214_1208 ();
 FILLCELL_X32 FILLER_214_1240 ();
 FILLCELL_X32 FILLER_214_1272 ();
 FILLCELL_X32 FILLER_214_1304 ();
 FILLCELL_X32 FILLER_214_1336 ();
 FILLCELL_X32 FILLER_214_1368 ();
 FILLCELL_X32 FILLER_214_1400 ();
 FILLCELL_X32 FILLER_214_1432 ();
 FILLCELL_X32 FILLER_214_1464 ();
 FILLCELL_X32 FILLER_214_1496 ();
 FILLCELL_X32 FILLER_214_1528 ();
 FILLCELL_X32 FILLER_214_1560 ();
 FILLCELL_X32 FILLER_214_1592 ();
 FILLCELL_X32 FILLER_214_1624 ();
 FILLCELL_X32 FILLER_214_1656 ();
 FILLCELL_X32 FILLER_214_1688 ();
 FILLCELL_X32 FILLER_214_1720 ();
 FILLCELL_X8 FILLER_214_1752 ();
 FILLCELL_X2 FILLER_214_1760 ();
 FILLCELL_X32 FILLER_215_1 ();
 FILLCELL_X32 FILLER_215_33 ();
 FILLCELL_X32 FILLER_215_65 ();
 FILLCELL_X32 FILLER_215_97 ();
 FILLCELL_X32 FILLER_215_129 ();
 FILLCELL_X32 FILLER_215_161 ();
 FILLCELL_X32 FILLER_215_193 ();
 FILLCELL_X32 FILLER_215_225 ();
 FILLCELL_X32 FILLER_215_257 ();
 FILLCELL_X32 FILLER_215_289 ();
 FILLCELL_X32 FILLER_215_321 ();
 FILLCELL_X32 FILLER_215_353 ();
 FILLCELL_X32 FILLER_215_385 ();
 FILLCELL_X32 FILLER_215_417 ();
 FILLCELL_X32 FILLER_215_449 ();
 FILLCELL_X32 FILLER_215_481 ();
 FILLCELL_X32 FILLER_215_513 ();
 FILLCELL_X32 FILLER_215_545 ();
 FILLCELL_X32 FILLER_215_577 ();
 FILLCELL_X32 FILLER_215_609 ();
 FILLCELL_X32 FILLER_215_641 ();
 FILLCELL_X32 FILLER_215_673 ();
 FILLCELL_X32 FILLER_215_705 ();
 FILLCELL_X32 FILLER_215_737 ();
 FILLCELL_X32 FILLER_215_769 ();
 FILLCELL_X32 FILLER_215_801 ();
 FILLCELL_X32 FILLER_215_833 ();
 FILLCELL_X32 FILLER_215_865 ();
 FILLCELL_X32 FILLER_215_897 ();
 FILLCELL_X32 FILLER_215_929 ();
 FILLCELL_X32 FILLER_215_961 ();
 FILLCELL_X32 FILLER_215_993 ();
 FILLCELL_X32 FILLER_215_1025 ();
 FILLCELL_X32 FILLER_215_1057 ();
 FILLCELL_X32 FILLER_215_1089 ();
 FILLCELL_X32 FILLER_215_1121 ();
 FILLCELL_X32 FILLER_215_1153 ();
 FILLCELL_X32 FILLER_215_1185 ();
 FILLCELL_X32 FILLER_215_1217 ();
 FILLCELL_X8 FILLER_215_1249 ();
 FILLCELL_X4 FILLER_215_1257 ();
 FILLCELL_X2 FILLER_215_1261 ();
 FILLCELL_X32 FILLER_215_1264 ();
 FILLCELL_X32 FILLER_215_1296 ();
 FILLCELL_X32 FILLER_215_1328 ();
 FILLCELL_X32 FILLER_215_1360 ();
 FILLCELL_X32 FILLER_215_1392 ();
 FILLCELL_X32 FILLER_215_1424 ();
 FILLCELL_X32 FILLER_215_1456 ();
 FILLCELL_X32 FILLER_215_1488 ();
 FILLCELL_X32 FILLER_215_1520 ();
 FILLCELL_X32 FILLER_215_1552 ();
 FILLCELL_X32 FILLER_215_1584 ();
 FILLCELL_X32 FILLER_215_1616 ();
 FILLCELL_X32 FILLER_215_1648 ();
 FILLCELL_X32 FILLER_215_1680 ();
 FILLCELL_X32 FILLER_215_1712 ();
 FILLCELL_X16 FILLER_215_1744 ();
 FILLCELL_X2 FILLER_215_1760 ();
 FILLCELL_X32 FILLER_216_1 ();
 FILLCELL_X32 FILLER_216_33 ();
 FILLCELL_X32 FILLER_216_65 ();
 FILLCELL_X32 FILLER_216_97 ();
 FILLCELL_X32 FILLER_216_129 ();
 FILLCELL_X32 FILLER_216_161 ();
 FILLCELL_X32 FILLER_216_193 ();
 FILLCELL_X32 FILLER_216_225 ();
 FILLCELL_X32 FILLER_216_257 ();
 FILLCELL_X32 FILLER_216_289 ();
 FILLCELL_X32 FILLER_216_321 ();
 FILLCELL_X32 FILLER_216_353 ();
 FILLCELL_X32 FILLER_216_385 ();
 FILLCELL_X32 FILLER_216_417 ();
 FILLCELL_X32 FILLER_216_449 ();
 FILLCELL_X32 FILLER_216_481 ();
 FILLCELL_X32 FILLER_216_513 ();
 FILLCELL_X32 FILLER_216_545 ();
 FILLCELL_X32 FILLER_216_577 ();
 FILLCELL_X16 FILLER_216_609 ();
 FILLCELL_X4 FILLER_216_625 ();
 FILLCELL_X2 FILLER_216_629 ();
 FILLCELL_X32 FILLER_216_632 ();
 FILLCELL_X32 FILLER_216_664 ();
 FILLCELL_X32 FILLER_216_696 ();
 FILLCELL_X32 FILLER_216_728 ();
 FILLCELL_X32 FILLER_216_760 ();
 FILLCELL_X32 FILLER_216_792 ();
 FILLCELL_X32 FILLER_216_824 ();
 FILLCELL_X32 FILLER_216_856 ();
 FILLCELL_X32 FILLER_216_888 ();
 FILLCELL_X32 FILLER_216_920 ();
 FILLCELL_X32 FILLER_216_952 ();
 FILLCELL_X32 FILLER_216_984 ();
 FILLCELL_X32 FILLER_216_1016 ();
 FILLCELL_X32 FILLER_216_1048 ();
 FILLCELL_X32 FILLER_216_1080 ();
 FILLCELL_X32 FILLER_216_1112 ();
 FILLCELL_X32 FILLER_216_1144 ();
 FILLCELL_X32 FILLER_216_1176 ();
 FILLCELL_X32 FILLER_216_1208 ();
 FILLCELL_X32 FILLER_216_1240 ();
 FILLCELL_X32 FILLER_216_1272 ();
 FILLCELL_X32 FILLER_216_1304 ();
 FILLCELL_X32 FILLER_216_1336 ();
 FILLCELL_X32 FILLER_216_1368 ();
 FILLCELL_X32 FILLER_216_1400 ();
 FILLCELL_X32 FILLER_216_1432 ();
 FILLCELL_X32 FILLER_216_1464 ();
 FILLCELL_X32 FILLER_216_1496 ();
 FILLCELL_X32 FILLER_216_1528 ();
 FILLCELL_X32 FILLER_216_1560 ();
 FILLCELL_X32 FILLER_216_1592 ();
 FILLCELL_X32 FILLER_216_1624 ();
 FILLCELL_X32 FILLER_216_1656 ();
 FILLCELL_X32 FILLER_216_1688 ();
 FILLCELL_X32 FILLER_216_1720 ();
 FILLCELL_X8 FILLER_216_1752 ();
 FILLCELL_X2 FILLER_216_1760 ();
 FILLCELL_X32 FILLER_217_1 ();
 FILLCELL_X32 FILLER_217_33 ();
 FILLCELL_X32 FILLER_217_65 ();
 FILLCELL_X32 FILLER_217_97 ();
 FILLCELL_X32 FILLER_217_129 ();
 FILLCELL_X32 FILLER_217_161 ();
 FILLCELL_X32 FILLER_217_193 ();
 FILLCELL_X32 FILLER_217_225 ();
 FILLCELL_X32 FILLER_217_257 ();
 FILLCELL_X32 FILLER_217_289 ();
 FILLCELL_X32 FILLER_217_321 ();
 FILLCELL_X32 FILLER_217_353 ();
 FILLCELL_X32 FILLER_217_385 ();
 FILLCELL_X32 FILLER_217_417 ();
 FILLCELL_X32 FILLER_217_449 ();
 FILLCELL_X32 FILLER_217_481 ();
 FILLCELL_X32 FILLER_217_513 ();
 FILLCELL_X32 FILLER_217_545 ();
 FILLCELL_X32 FILLER_217_577 ();
 FILLCELL_X32 FILLER_217_609 ();
 FILLCELL_X32 FILLER_217_641 ();
 FILLCELL_X32 FILLER_217_673 ();
 FILLCELL_X32 FILLER_217_705 ();
 FILLCELL_X32 FILLER_217_737 ();
 FILLCELL_X32 FILLER_217_769 ();
 FILLCELL_X32 FILLER_217_801 ();
 FILLCELL_X32 FILLER_217_833 ();
 FILLCELL_X32 FILLER_217_865 ();
 FILLCELL_X32 FILLER_217_897 ();
 FILLCELL_X32 FILLER_217_929 ();
 FILLCELL_X32 FILLER_217_961 ();
 FILLCELL_X32 FILLER_217_993 ();
 FILLCELL_X32 FILLER_217_1025 ();
 FILLCELL_X32 FILLER_217_1057 ();
 FILLCELL_X32 FILLER_217_1089 ();
 FILLCELL_X32 FILLER_217_1121 ();
 FILLCELL_X32 FILLER_217_1153 ();
 FILLCELL_X32 FILLER_217_1185 ();
 FILLCELL_X32 FILLER_217_1217 ();
 FILLCELL_X8 FILLER_217_1249 ();
 FILLCELL_X4 FILLER_217_1257 ();
 FILLCELL_X2 FILLER_217_1261 ();
 FILLCELL_X32 FILLER_217_1264 ();
 FILLCELL_X32 FILLER_217_1296 ();
 FILLCELL_X32 FILLER_217_1328 ();
 FILLCELL_X32 FILLER_217_1360 ();
 FILLCELL_X32 FILLER_217_1392 ();
 FILLCELL_X32 FILLER_217_1424 ();
 FILLCELL_X32 FILLER_217_1456 ();
 FILLCELL_X32 FILLER_217_1488 ();
 FILLCELL_X32 FILLER_217_1520 ();
 FILLCELL_X32 FILLER_217_1552 ();
 FILLCELL_X32 FILLER_217_1584 ();
 FILLCELL_X32 FILLER_217_1616 ();
 FILLCELL_X32 FILLER_217_1648 ();
 FILLCELL_X32 FILLER_217_1680 ();
 FILLCELL_X32 FILLER_217_1712 ();
 FILLCELL_X16 FILLER_217_1744 ();
 FILLCELL_X2 FILLER_217_1760 ();
 FILLCELL_X4 FILLER_218_1 ();
 FILLCELL_X32 FILLER_218_12 ();
 FILLCELL_X32 FILLER_218_44 ();
 FILLCELL_X32 FILLER_218_76 ();
 FILLCELL_X32 FILLER_218_108 ();
 FILLCELL_X32 FILLER_218_140 ();
 FILLCELL_X32 FILLER_218_172 ();
 FILLCELL_X32 FILLER_218_204 ();
 FILLCELL_X32 FILLER_218_236 ();
 FILLCELL_X32 FILLER_218_268 ();
 FILLCELL_X32 FILLER_218_300 ();
 FILLCELL_X32 FILLER_218_332 ();
 FILLCELL_X32 FILLER_218_364 ();
 FILLCELL_X32 FILLER_218_396 ();
 FILLCELL_X32 FILLER_218_428 ();
 FILLCELL_X32 FILLER_218_460 ();
 FILLCELL_X32 FILLER_218_492 ();
 FILLCELL_X32 FILLER_218_524 ();
 FILLCELL_X32 FILLER_218_556 ();
 FILLCELL_X32 FILLER_218_588 ();
 FILLCELL_X8 FILLER_218_620 ();
 FILLCELL_X2 FILLER_218_628 ();
 FILLCELL_X1 FILLER_218_630 ();
 FILLCELL_X32 FILLER_218_632 ();
 FILLCELL_X32 FILLER_218_664 ();
 FILLCELL_X32 FILLER_218_696 ();
 FILLCELL_X32 FILLER_218_728 ();
 FILLCELL_X32 FILLER_218_760 ();
 FILLCELL_X32 FILLER_218_792 ();
 FILLCELL_X32 FILLER_218_824 ();
 FILLCELL_X32 FILLER_218_856 ();
 FILLCELL_X32 FILLER_218_888 ();
 FILLCELL_X32 FILLER_218_920 ();
 FILLCELL_X32 FILLER_218_952 ();
 FILLCELL_X32 FILLER_218_984 ();
 FILLCELL_X32 FILLER_218_1016 ();
 FILLCELL_X32 FILLER_218_1048 ();
 FILLCELL_X32 FILLER_218_1080 ();
 FILLCELL_X32 FILLER_218_1112 ();
 FILLCELL_X32 FILLER_218_1144 ();
 FILLCELL_X32 FILLER_218_1176 ();
 FILLCELL_X32 FILLER_218_1208 ();
 FILLCELL_X32 FILLER_218_1240 ();
 FILLCELL_X32 FILLER_218_1272 ();
 FILLCELL_X32 FILLER_218_1304 ();
 FILLCELL_X32 FILLER_218_1336 ();
 FILLCELL_X32 FILLER_218_1368 ();
 FILLCELL_X32 FILLER_218_1400 ();
 FILLCELL_X32 FILLER_218_1432 ();
 FILLCELL_X32 FILLER_218_1464 ();
 FILLCELL_X32 FILLER_218_1496 ();
 FILLCELL_X32 FILLER_218_1528 ();
 FILLCELL_X32 FILLER_218_1560 ();
 FILLCELL_X32 FILLER_218_1592 ();
 FILLCELL_X32 FILLER_218_1624 ();
 FILLCELL_X32 FILLER_218_1656 ();
 FILLCELL_X32 FILLER_218_1688 ();
 FILLCELL_X32 FILLER_218_1720 ();
 FILLCELL_X8 FILLER_218_1752 ();
 FILLCELL_X2 FILLER_218_1760 ();
 FILLCELL_X32 FILLER_219_1 ();
 FILLCELL_X32 FILLER_219_33 ();
 FILLCELL_X32 FILLER_219_65 ();
 FILLCELL_X32 FILLER_219_97 ();
 FILLCELL_X32 FILLER_219_129 ();
 FILLCELL_X32 FILLER_219_161 ();
 FILLCELL_X32 FILLER_219_193 ();
 FILLCELL_X32 FILLER_219_225 ();
 FILLCELL_X32 FILLER_219_257 ();
 FILLCELL_X32 FILLER_219_289 ();
 FILLCELL_X32 FILLER_219_321 ();
 FILLCELL_X32 FILLER_219_353 ();
 FILLCELL_X32 FILLER_219_385 ();
 FILLCELL_X32 FILLER_219_417 ();
 FILLCELL_X32 FILLER_219_449 ();
 FILLCELL_X32 FILLER_219_481 ();
 FILLCELL_X32 FILLER_219_513 ();
 FILLCELL_X32 FILLER_219_545 ();
 FILLCELL_X32 FILLER_219_577 ();
 FILLCELL_X32 FILLER_219_609 ();
 FILLCELL_X32 FILLER_219_641 ();
 FILLCELL_X32 FILLER_219_673 ();
 FILLCELL_X32 FILLER_219_705 ();
 FILLCELL_X32 FILLER_219_737 ();
 FILLCELL_X32 FILLER_219_769 ();
 FILLCELL_X32 FILLER_219_801 ();
 FILLCELL_X32 FILLER_219_833 ();
 FILLCELL_X32 FILLER_219_865 ();
 FILLCELL_X32 FILLER_219_897 ();
 FILLCELL_X32 FILLER_219_929 ();
 FILLCELL_X32 FILLER_219_961 ();
 FILLCELL_X32 FILLER_219_993 ();
 FILLCELL_X32 FILLER_219_1025 ();
 FILLCELL_X32 FILLER_219_1057 ();
 FILLCELL_X32 FILLER_219_1089 ();
 FILLCELL_X32 FILLER_219_1121 ();
 FILLCELL_X32 FILLER_219_1153 ();
 FILLCELL_X32 FILLER_219_1185 ();
 FILLCELL_X32 FILLER_219_1217 ();
 FILLCELL_X8 FILLER_219_1249 ();
 FILLCELL_X4 FILLER_219_1257 ();
 FILLCELL_X2 FILLER_219_1261 ();
 FILLCELL_X32 FILLER_219_1264 ();
 FILLCELL_X32 FILLER_219_1296 ();
 FILLCELL_X32 FILLER_219_1328 ();
 FILLCELL_X32 FILLER_219_1360 ();
 FILLCELL_X32 FILLER_219_1392 ();
 FILLCELL_X32 FILLER_219_1424 ();
 FILLCELL_X32 FILLER_219_1456 ();
 FILLCELL_X32 FILLER_219_1488 ();
 FILLCELL_X32 FILLER_219_1520 ();
 FILLCELL_X32 FILLER_219_1552 ();
 FILLCELL_X32 FILLER_219_1584 ();
 FILLCELL_X32 FILLER_219_1616 ();
 FILLCELL_X32 FILLER_219_1648 ();
 FILLCELL_X32 FILLER_219_1680 ();
 FILLCELL_X32 FILLER_219_1712 ();
 FILLCELL_X16 FILLER_219_1744 ();
 FILLCELL_X2 FILLER_219_1760 ();
 FILLCELL_X32 FILLER_220_1 ();
 FILLCELL_X32 FILLER_220_33 ();
 FILLCELL_X32 FILLER_220_65 ();
 FILLCELL_X32 FILLER_220_97 ();
 FILLCELL_X32 FILLER_220_129 ();
 FILLCELL_X32 FILLER_220_161 ();
 FILLCELL_X32 FILLER_220_193 ();
 FILLCELL_X32 FILLER_220_225 ();
 FILLCELL_X32 FILLER_220_257 ();
 FILLCELL_X32 FILLER_220_289 ();
 FILLCELL_X32 FILLER_220_321 ();
 FILLCELL_X32 FILLER_220_353 ();
 FILLCELL_X32 FILLER_220_385 ();
 FILLCELL_X32 FILLER_220_417 ();
 FILLCELL_X32 FILLER_220_449 ();
 FILLCELL_X32 FILLER_220_481 ();
 FILLCELL_X32 FILLER_220_513 ();
 FILLCELL_X32 FILLER_220_545 ();
 FILLCELL_X32 FILLER_220_577 ();
 FILLCELL_X16 FILLER_220_609 ();
 FILLCELL_X4 FILLER_220_625 ();
 FILLCELL_X2 FILLER_220_629 ();
 FILLCELL_X32 FILLER_220_632 ();
 FILLCELL_X32 FILLER_220_664 ();
 FILLCELL_X32 FILLER_220_696 ();
 FILLCELL_X32 FILLER_220_728 ();
 FILLCELL_X32 FILLER_220_760 ();
 FILLCELL_X32 FILLER_220_792 ();
 FILLCELL_X32 FILLER_220_824 ();
 FILLCELL_X32 FILLER_220_856 ();
 FILLCELL_X32 FILLER_220_888 ();
 FILLCELL_X32 FILLER_220_920 ();
 FILLCELL_X32 FILLER_220_952 ();
 FILLCELL_X32 FILLER_220_984 ();
 FILLCELL_X32 FILLER_220_1016 ();
 FILLCELL_X32 FILLER_220_1048 ();
 FILLCELL_X32 FILLER_220_1080 ();
 FILLCELL_X32 FILLER_220_1112 ();
 FILLCELL_X32 FILLER_220_1144 ();
 FILLCELL_X32 FILLER_220_1176 ();
 FILLCELL_X32 FILLER_220_1208 ();
 FILLCELL_X32 FILLER_220_1240 ();
 FILLCELL_X32 FILLER_220_1272 ();
 FILLCELL_X32 FILLER_220_1304 ();
 FILLCELL_X32 FILLER_220_1336 ();
 FILLCELL_X32 FILLER_220_1368 ();
 FILLCELL_X32 FILLER_220_1400 ();
 FILLCELL_X32 FILLER_220_1432 ();
 FILLCELL_X32 FILLER_220_1464 ();
 FILLCELL_X32 FILLER_220_1496 ();
 FILLCELL_X32 FILLER_220_1528 ();
 FILLCELL_X32 FILLER_220_1560 ();
 FILLCELL_X32 FILLER_220_1592 ();
 FILLCELL_X32 FILLER_220_1624 ();
 FILLCELL_X32 FILLER_220_1656 ();
 FILLCELL_X32 FILLER_220_1688 ();
 FILLCELL_X32 FILLER_220_1720 ();
 FILLCELL_X8 FILLER_220_1752 ();
 FILLCELL_X2 FILLER_220_1760 ();
 FILLCELL_X32 FILLER_221_1 ();
 FILLCELL_X32 FILLER_221_33 ();
 FILLCELL_X32 FILLER_221_65 ();
 FILLCELL_X32 FILLER_221_97 ();
 FILLCELL_X32 FILLER_221_129 ();
 FILLCELL_X32 FILLER_221_161 ();
 FILLCELL_X32 FILLER_221_193 ();
 FILLCELL_X32 FILLER_221_225 ();
 FILLCELL_X32 FILLER_221_257 ();
 FILLCELL_X32 FILLER_221_289 ();
 FILLCELL_X32 FILLER_221_321 ();
 FILLCELL_X32 FILLER_221_353 ();
 FILLCELL_X32 FILLER_221_385 ();
 FILLCELL_X32 FILLER_221_417 ();
 FILLCELL_X32 FILLER_221_449 ();
 FILLCELL_X32 FILLER_221_481 ();
 FILLCELL_X32 FILLER_221_513 ();
 FILLCELL_X32 FILLER_221_545 ();
 FILLCELL_X32 FILLER_221_577 ();
 FILLCELL_X32 FILLER_221_609 ();
 FILLCELL_X32 FILLER_221_641 ();
 FILLCELL_X32 FILLER_221_673 ();
 FILLCELL_X32 FILLER_221_705 ();
 FILLCELL_X32 FILLER_221_737 ();
 FILLCELL_X32 FILLER_221_769 ();
 FILLCELL_X32 FILLER_221_801 ();
 FILLCELL_X32 FILLER_221_833 ();
 FILLCELL_X32 FILLER_221_865 ();
 FILLCELL_X32 FILLER_221_897 ();
 FILLCELL_X32 FILLER_221_929 ();
 FILLCELL_X32 FILLER_221_961 ();
 FILLCELL_X32 FILLER_221_993 ();
 FILLCELL_X32 FILLER_221_1025 ();
 FILLCELL_X32 FILLER_221_1057 ();
 FILLCELL_X32 FILLER_221_1089 ();
 FILLCELL_X32 FILLER_221_1121 ();
 FILLCELL_X32 FILLER_221_1153 ();
 FILLCELL_X32 FILLER_221_1185 ();
 FILLCELL_X32 FILLER_221_1217 ();
 FILLCELL_X8 FILLER_221_1249 ();
 FILLCELL_X4 FILLER_221_1257 ();
 FILLCELL_X2 FILLER_221_1261 ();
 FILLCELL_X32 FILLER_221_1264 ();
 FILLCELL_X32 FILLER_221_1296 ();
 FILLCELL_X32 FILLER_221_1328 ();
 FILLCELL_X32 FILLER_221_1360 ();
 FILLCELL_X32 FILLER_221_1392 ();
 FILLCELL_X32 FILLER_221_1424 ();
 FILLCELL_X32 FILLER_221_1456 ();
 FILLCELL_X32 FILLER_221_1488 ();
 FILLCELL_X32 FILLER_221_1520 ();
 FILLCELL_X32 FILLER_221_1552 ();
 FILLCELL_X32 FILLER_221_1584 ();
 FILLCELL_X32 FILLER_221_1616 ();
 FILLCELL_X32 FILLER_221_1648 ();
 FILLCELL_X32 FILLER_221_1680 ();
 FILLCELL_X32 FILLER_221_1712 ();
 FILLCELL_X16 FILLER_221_1744 ();
 FILLCELL_X2 FILLER_221_1760 ();
 FILLCELL_X32 FILLER_222_1 ();
 FILLCELL_X32 FILLER_222_33 ();
 FILLCELL_X32 FILLER_222_65 ();
 FILLCELL_X32 FILLER_222_97 ();
 FILLCELL_X32 FILLER_222_129 ();
 FILLCELL_X32 FILLER_222_161 ();
 FILLCELL_X32 FILLER_222_193 ();
 FILLCELL_X32 FILLER_222_225 ();
 FILLCELL_X32 FILLER_222_257 ();
 FILLCELL_X32 FILLER_222_289 ();
 FILLCELL_X32 FILLER_222_321 ();
 FILLCELL_X32 FILLER_222_353 ();
 FILLCELL_X32 FILLER_222_385 ();
 FILLCELL_X32 FILLER_222_417 ();
 FILLCELL_X32 FILLER_222_449 ();
 FILLCELL_X32 FILLER_222_481 ();
 FILLCELL_X32 FILLER_222_513 ();
 FILLCELL_X32 FILLER_222_545 ();
 FILLCELL_X32 FILLER_222_577 ();
 FILLCELL_X16 FILLER_222_609 ();
 FILLCELL_X4 FILLER_222_625 ();
 FILLCELL_X2 FILLER_222_629 ();
 FILLCELL_X32 FILLER_222_632 ();
 FILLCELL_X32 FILLER_222_664 ();
 FILLCELL_X32 FILLER_222_696 ();
 FILLCELL_X32 FILLER_222_728 ();
 FILLCELL_X32 FILLER_222_760 ();
 FILLCELL_X32 FILLER_222_792 ();
 FILLCELL_X32 FILLER_222_824 ();
 FILLCELL_X32 FILLER_222_856 ();
 FILLCELL_X32 FILLER_222_888 ();
 FILLCELL_X32 FILLER_222_920 ();
 FILLCELL_X32 FILLER_222_952 ();
 FILLCELL_X32 FILLER_222_984 ();
 FILLCELL_X32 FILLER_222_1016 ();
 FILLCELL_X32 FILLER_222_1048 ();
 FILLCELL_X32 FILLER_222_1080 ();
 FILLCELL_X32 FILLER_222_1112 ();
 FILLCELL_X32 FILLER_222_1144 ();
 FILLCELL_X32 FILLER_222_1176 ();
 FILLCELL_X32 FILLER_222_1208 ();
 FILLCELL_X32 FILLER_222_1240 ();
 FILLCELL_X32 FILLER_222_1272 ();
 FILLCELL_X32 FILLER_222_1304 ();
 FILLCELL_X32 FILLER_222_1336 ();
 FILLCELL_X32 FILLER_222_1368 ();
 FILLCELL_X32 FILLER_222_1400 ();
 FILLCELL_X32 FILLER_222_1432 ();
 FILLCELL_X32 FILLER_222_1464 ();
 FILLCELL_X32 FILLER_222_1496 ();
 FILLCELL_X32 FILLER_222_1528 ();
 FILLCELL_X32 FILLER_222_1560 ();
 FILLCELL_X32 FILLER_222_1592 ();
 FILLCELL_X32 FILLER_222_1624 ();
 FILLCELL_X32 FILLER_222_1656 ();
 FILLCELL_X32 FILLER_222_1688 ();
 FILLCELL_X16 FILLER_222_1720 ();
 FILLCELL_X8 FILLER_222_1736 ();
 FILLCELL_X4 FILLER_222_1744 ();
 FILLCELL_X2 FILLER_222_1748 ();
 FILLCELL_X1 FILLER_222_1750 ();
 FILLCELL_X4 FILLER_222_1758 ();
 FILLCELL_X32 FILLER_223_1 ();
 FILLCELL_X32 FILLER_223_33 ();
 FILLCELL_X32 FILLER_223_65 ();
 FILLCELL_X32 FILLER_223_97 ();
 FILLCELL_X32 FILLER_223_129 ();
 FILLCELL_X32 FILLER_223_161 ();
 FILLCELL_X32 FILLER_223_193 ();
 FILLCELL_X32 FILLER_223_225 ();
 FILLCELL_X32 FILLER_223_257 ();
 FILLCELL_X32 FILLER_223_289 ();
 FILLCELL_X32 FILLER_223_321 ();
 FILLCELL_X32 FILLER_223_353 ();
 FILLCELL_X32 FILLER_223_385 ();
 FILLCELL_X32 FILLER_223_417 ();
 FILLCELL_X32 FILLER_223_449 ();
 FILLCELL_X32 FILLER_223_481 ();
 FILLCELL_X32 FILLER_223_513 ();
 FILLCELL_X32 FILLER_223_545 ();
 FILLCELL_X32 FILLER_223_577 ();
 FILLCELL_X32 FILLER_223_609 ();
 FILLCELL_X32 FILLER_223_641 ();
 FILLCELL_X32 FILLER_223_673 ();
 FILLCELL_X32 FILLER_223_705 ();
 FILLCELL_X32 FILLER_223_737 ();
 FILLCELL_X32 FILLER_223_769 ();
 FILLCELL_X32 FILLER_223_801 ();
 FILLCELL_X32 FILLER_223_833 ();
 FILLCELL_X32 FILLER_223_865 ();
 FILLCELL_X32 FILLER_223_897 ();
 FILLCELL_X32 FILLER_223_929 ();
 FILLCELL_X32 FILLER_223_961 ();
 FILLCELL_X32 FILLER_223_993 ();
 FILLCELL_X32 FILLER_223_1025 ();
 FILLCELL_X32 FILLER_223_1057 ();
 FILLCELL_X32 FILLER_223_1089 ();
 FILLCELL_X32 FILLER_223_1121 ();
 FILLCELL_X32 FILLER_223_1153 ();
 FILLCELL_X32 FILLER_223_1185 ();
 FILLCELL_X32 FILLER_223_1217 ();
 FILLCELL_X8 FILLER_223_1249 ();
 FILLCELL_X4 FILLER_223_1257 ();
 FILLCELL_X2 FILLER_223_1261 ();
 FILLCELL_X32 FILLER_223_1264 ();
 FILLCELL_X32 FILLER_223_1296 ();
 FILLCELL_X32 FILLER_223_1328 ();
 FILLCELL_X32 FILLER_223_1360 ();
 FILLCELL_X32 FILLER_223_1392 ();
 FILLCELL_X32 FILLER_223_1424 ();
 FILLCELL_X32 FILLER_223_1456 ();
 FILLCELL_X32 FILLER_223_1488 ();
 FILLCELL_X32 FILLER_223_1520 ();
 FILLCELL_X32 FILLER_223_1552 ();
 FILLCELL_X32 FILLER_223_1584 ();
 FILLCELL_X32 FILLER_223_1616 ();
 FILLCELL_X32 FILLER_223_1648 ();
 FILLCELL_X32 FILLER_223_1680 ();
 FILLCELL_X32 FILLER_223_1712 ();
 FILLCELL_X16 FILLER_223_1744 ();
 FILLCELL_X2 FILLER_223_1760 ();
 FILLCELL_X32 FILLER_224_1 ();
 FILLCELL_X32 FILLER_224_33 ();
 FILLCELL_X32 FILLER_224_65 ();
 FILLCELL_X32 FILLER_224_97 ();
 FILLCELL_X32 FILLER_224_129 ();
 FILLCELL_X32 FILLER_224_161 ();
 FILLCELL_X32 FILLER_224_193 ();
 FILLCELL_X32 FILLER_224_225 ();
 FILLCELL_X32 FILLER_224_257 ();
 FILLCELL_X32 FILLER_224_289 ();
 FILLCELL_X32 FILLER_224_321 ();
 FILLCELL_X32 FILLER_224_353 ();
 FILLCELL_X32 FILLER_224_385 ();
 FILLCELL_X32 FILLER_224_417 ();
 FILLCELL_X32 FILLER_224_449 ();
 FILLCELL_X32 FILLER_224_481 ();
 FILLCELL_X32 FILLER_224_513 ();
 FILLCELL_X32 FILLER_224_545 ();
 FILLCELL_X32 FILLER_224_577 ();
 FILLCELL_X16 FILLER_224_609 ();
 FILLCELL_X4 FILLER_224_625 ();
 FILLCELL_X2 FILLER_224_629 ();
 FILLCELL_X32 FILLER_224_632 ();
 FILLCELL_X32 FILLER_224_664 ();
 FILLCELL_X32 FILLER_224_696 ();
 FILLCELL_X32 FILLER_224_728 ();
 FILLCELL_X32 FILLER_224_760 ();
 FILLCELL_X32 FILLER_224_792 ();
 FILLCELL_X32 FILLER_224_824 ();
 FILLCELL_X32 FILLER_224_856 ();
 FILLCELL_X32 FILLER_224_888 ();
 FILLCELL_X32 FILLER_224_920 ();
 FILLCELL_X32 FILLER_224_952 ();
 FILLCELL_X32 FILLER_224_984 ();
 FILLCELL_X32 FILLER_224_1016 ();
 FILLCELL_X32 FILLER_224_1048 ();
 FILLCELL_X32 FILLER_224_1080 ();
 FILLCELL_X32 FILLER_224_1112 ();
 FILLCELL_X32 FILLER_224_1144 ();
 FILLCELL_X32 FILLER_224_1176 ();
 FILLCELL_X32 FILLER_224_1208 ();
 FILLCELL_X32 FILLER_224_1240 ();
 FILLCELL_X32 FILLER_224_1272 ();
 FILLCELL_X32 FILLER_224_1304 ();
 FILLCELL_X32 FILLER_224_1336 ();
 FILLCELL_X32 FILLER_224_1368 ();
 FILLCELL_X32 FILLER_224_1400 ();
 FILLCELL_X32 FILLER_224_1432 ();
 FILLCELL_X32 FILLER_224_1464 ();
 FILLCELL_X32 FILLER_224_1496 ();
 FILLCELL_X32 FILLER_224_1528 ();
 FILLCELL_X32 FILLER_224_1560 ();
 FILLCELL_X32 FILLER_224_1592 ();
 FILLCELL_X32 FILLER_224_1624 ();
 FILLCELL_X32 FILLER_224_1656 ();
 FILLCELL_X32 FILLER_224_1688 ();
 FILLCELL_X32 FILLER_224_1720 ();
 FILLCELL_X8 FILLER_224_1752 ();
 FILLCELL_X2 FILLER_224_1760 ();
 FILLCELL_X32 FILLER_225_1 ();
 FILLCELL_X32 FILLER_225_33 ();
 FILLCELL_X32 FILLER_225_65 ();
 FILLCELL_X32 FILLER_225_97 ();
 FILLCELL_X32 FILLER_225_129 ();
 FILLCELL_X32 FILLER_225_161 ();
 FILLCELL_X32 FILLER_225_193 ();
 FILLCELL_X32 FILLER_225_225 ();
 FILLCELL_X32 FILLER_225_257 ();
 FILLCELL_X32 FILLER_225_289 ();
 FILLCELL_X32 FILLER_225_321 ();
 FILLCELL_X32 FILLER_225_353 ();
 FILLCELL_X32 FILLER_225_385 ();
 FILLCELL_X32 FILLER_225_417 ();
 FILLCELL_X32 FILLER_225_449 ();
 FILLCELL_X32 FILLER_225_481 ();
 FILLCELL_X32 FILLER_225_513 ();
 FILLCELL_X32 FILLER_225_545 ();
 FILLCELL_X32 FILLER_225_577 ();
 FILLCELL_X32 FILLER_225_609 ();
 FILLCELL_X32 FILLER_225_641 ();
 FILLCELL_X32 FILLER_225_673 ();
 FILLCELL_X32 FILLER_225_705 ();
 FILLCELL_X32 FILLER_225_737 ();
 FILLCELL_X32 FILLER_225_769 ();
 FILLCELL_X32 FILLER_225_801 ();
 FILLCELL_X32 FILLER_225_833 ();
 FILLCELL_X32 FILLER_225_865 ();
 FILLCELL_X32 FILLER_225_897 ();
 FILLCELL_X32 FILLER_225_929 ();
 FILLCELL_X32 FILLER_225_961 ();
 FILLCELL_X32 FILLER_225_993 ();
 FILLCELL_X32 FILLER_225_1025 ();
 FILLCELL_X32 FILLER_225_1057 ();
 FILLCELL_X32 FILLER_225_1089 ();
 FILLCELL_X32 FILLER_225_1121 ();
 FILLCELL_X32 FILLER_225_1153 ();
 FILLCELL_X32 FILLER_225_1185 ();
 FILLCELL_X32 FILLER_225_1217 ();
 FILLCELL_X8 FILLER_225_1249 ();
 FILLCELL_X4 FILLER_225_1257 ();
 FILLCELL_X2 FILLER_225_1261 ();
 FILLCELL_X32 FILLER_225_1264 ();
 FILLCELL_X32 FILLER_225_1296 ();
 FILLCELL_X32 FILLER_225_1328 ();
 FILLCELL_X32 FILLER_225_1360 ();
 FILLCELL_X32 FILLER_225_1392 ();
 FILLCELL_X32 FILLER_225_1424 ();
 FILLCELL_X32 FILLER_225_1456 ();
 FILLCELL_X32 FILLER_225_1488 ();
 FILLCELL_X32 FILLER_225_1520 ();
 FILLCELL_X32 FILLER_225_1552 ();
 FILLCELL_X32 FILLER_225_1584 ();
 FILLCELL_X32 FILLER_225_1616 ();
 FILLCELL_X32 FILLER_225_1648 ();
 FILLCELL_X32 FILLER_225_1680 ();
 FILLCELL_X32 FILLER_225_1712 ();
 FILLCELL_X16 FILLER_225_1744 ();
 FILLCELL_X2 FILLER_225_1760 ();
 FILLCELL_X32 FILLER_226_1 ();
 FILLCELL_X32 FILLER_226_33 ();
 FILLCELL_X32 FILLER_226_65 ();
 FILLCELL_X32 FILLER_226_97 ();
 FILLCELL_X32 FILLER_226_129 ();
 FILLCELL_X32 FILLER_226_161 ();
 FILLCELL_X32 FILLER_226_193 ();
 FILLCELL_X32 FILLER_226_225 ();
 FILLCELL_X32 FILLER_226_257 ();
 FILLCELL_X32 FILLER_226_289 ();
 FILLCELL_X32 FILLER_226_321 ();
 FILLCELL_X32 FILLER_226_353 ();
 FILLCELL_X32 FILLER_226_385 ();
 FILLCELL_X32 FILLER_226_417 ();
 FILLCELL_X32 FILLER_226_449 ();
 FILLCELL_X32 FILLER_226_481 ();
 FILLCELL_X32 FILLER_226_513 ();
 FILLCELL_X32 FILLER_226_545 ();
 FILLCELL_X32 FILLER_226_577 ();
 FILLCELL_X16 FILLER_226_609 ();
 FILLCELL_X4 FILLER_226_625 ();
 FILLCELL_X2 FILLER_226_629 ();
 FILLCELL_X32 FILLER_226_632 ();
 FILLCELL_X32 FILLER_226_664 ();
 FILLCELL_X32 FILLER_226_696 ();
 FILLCELL_X32 FILLER_226_728 ();
 FILLCELL_X32 FILLER_226_760 ();
 FILLCELL_X32 FILLER_226_792 ();
 FILLCELL_X32 FILLER_226_824 ();
 FILLCELL_X32 FILLER_226_856 ();
 FILLCELL_X32 FILLER_226_888 ();
 FILLCELL_X32 FILLER_226_920 ();
 FILLCELL_X32 FILLER_226_952 ();
 FILLCELL_X32 FILLER_226_984 ();
 FILLCELL_X32 FILLER_226_1016 ();
 FILLCELL_X32 FILLER_226_1048 ();
 FILLCELL_X32 FILLER_226_1080 ();
 FILLCELL_X32 FILLER_226_1112 ();
 FILLCELL_X32 FILLER_226_1144 ();
 FILLCELL_X32 FILLER_226_1176 ();
 FILLCELL_X32 FILLER_226_1208 ();
 FILLCELL_X32 FILLER_226_1240 ();
 FILLCELL_X32 FILLER_226_1272 ();
 FILLCELL_X32 FILLER_226_1304 ();
 FILLCELL_X32 FILLER_226_1336 ();
 FILLCELL_X32 FILLER_226_1368 ();
 FILLCELL_X32 FILLER_226_1400 ();
 FILLCELL_X32 FILLER_226_1432 ();
 FILLCELL_X32 FILLER_226_1464 ();
 FILLCELL_X32 FILLER_226_1496 ();
 FILLCELL_X32 FILLER_226_1528 ();
 FILLCELL_X32 FILLER_226_1560 ();
 FILLCELL_X32 FILLER_226_1592 ();
 FILLCELL_X32 FILLER_226_1624 ();
 FILLCELL_X32 FILLER_226_1656 ();
 FILLCELL_X32 FILLER_226_1688 ();
 FILLCELL_X32 FILLER_226_1720 ();
 FILLCELL_X8 FILLER_226_1752 ();
 FILLCELL_X2 FILLER_226_1760 ();
 FILLCELL_X4 FILLER_227_1 ();
 FILLCELL_X32 FILLER_227_9 ();
 FILLCELL_X32 FILLER_227_41 ();
 FILLCELL_X32 FILLER_227_73 ();
 FILLCELL_X32 FILLER_227_105 ();
 FILLCELL_X32 FILLER_227_137 ();
 FILLCELL_X32 FILLER_227_169 ();
 FILLCELL_X32 FILLER_227_201 ();
 FILLCELL_X32 FILLER_227_233 ();
 FILLCELL_X32 FILLER_227_265 ();
 FILLCELL_X32 FILLER_227_297 ();
 FILLCELL_X32 FILLER_227_329 ();
 FILLCELL_X32 FILLER_227_361 ();
 FILLCELL_X32 FILLER_227_393 ();
 FILLCELL_X32 FILLER_227_425 ();
 FILLCELL_X32 FILLER_227_457 ();
 FILLCELL_X32 FILLER_227_489 ();
 FILLCELL_X32 FILLER_227_521 ();
 FILLCELL_X32 FILLER_227_553 ();
 FILLCELL_X32 FILLER_227_585 ();
 FILLCELL_X32 FILLER_227_617 ();
 FILLCELL_X32 FILLER_227_649 ();
 FILLCELL_X32 FILLER_227_681 ();
 FILLCELL_X32 FILLER_227_713 ();
 FILLCELL_X32 FILLER_227_745 ();
 FILLCELL_X32 FILLER_227_777 ();
 FILLCELL_X32 FILLER_227_809 ();
 FILLCELL_X32 FILLER_227_841 ();
 FILLCELL_X32 FILLER_227_873 ();
 FILLCELL_X32 FILLER_227_905 ();
 FILLCELL_X32 FILLER_227_937 ();
 FILLCELL_X32 FILLER_227_969 ();
 FILLCELL_X32 FILLER_227_1001 ();
 FILLCELL_X32 FILLER_227_1033 ();
 FILLCELL_X32 FILLER_227_1065 ();
 FILLCELL_X32 FILLER_227_1097 ();
 FILLCELL_X32 FILLER_227_1129 ();
 FILLCELL_X32 FILLER_227_1161 ();
 FILLCELL_X32 FILLER_227_1193 ();
 FILLCELL_X32 FILLER_227_1225 ();
 FILLCELL_X4 FILLER_227_1257 ();
 FILLCELL_X2 FILLER_227_1261 ();
 FILLCELL_X32 FILLER_227_1264 ();
 FILLCELL_X32 FILLER_227_1296 ();
 FILLCELL_X32 FILLER_227_1328 ();
 FILLCELL_X32 FILLER_227_1360 ();
 FILLCELL_X32 FILLER_227_1392 ();
 FILLCELL_X32 FILLER_227_1424 ();
 FILLCELL_X32 FILLER_227_1456 ();
 FILLCELL_X32 FILLER_227_1488 ();
 FILLCELL_X32 FILLER_227_1520 ();
 FILLCELL_X32 FILLER_227_1552 ();
 FILLCELL_X32 FILLER_227_1584 ();
 FILLCELL_X32 FILLER_227_1616 ();
 FILLCELL_X32 FILLER_227_1648 ();
 FILLCELL_X32 FILLER_227_1680 ();
 FILLCELL_X32 FILLER_227_1712 ();
 FILLCELL_X16 FILLER_227_1744 ();
 FILLCELL_X2 FILLER_227_1760 ();
 FILLCELL_X32 FILLER_228_1 ();
 FILLCELL_X32 FILLER_228_33 ();
 FILLCELL_X32 FILLER_228_65 ();
 FILLCELL_X32 FILLER_228_97 ();
 FILLCELL_X32 FILLER_228_129 ();
 FILLCELL_X32 FILLER_228_161 ();
 FILLCELL_X32 FILLER_228_193 ();
 FILLCELL_X32 FILLER_228_225 ();
 FILLCELL_X32 FILLER_228_257 ();
 FILLCELL_X32 FILLER_228_289 ();
 FILLCELL_X32 FILLER_228_321 ();
 FILLCELL_X32 FILLER_228_353 ();
 FILLCELL_X32 FILLER_228_385 ();
 FILLCELL_X32 FILLER_228_417 ();
 FILLCELL_X32 FILLER_228_449 ();
 FILLCELL_X32 FILLER_228_481 ();
 FILLCELL_X32 FILLER_228_513 ();
 FILLCELL_X32 FILLER_228_545 ();
 FILLCELL_X32 FILLER_228_577 ();
 FILLCELL_X16 FILLER_228_609 ();
 FILLCELL_X4 FILLER_228_625 ();
 FILLCELL_X2 FILLER_228_629 ();
 FILLCELL_X32 FILLER_228_632 ();
 FILLCELL_X32 FILLER_228_664 ();
 FILLCELL_X32 FILLER_228_696 ();
 FILLCELL_X32 FILLER_228_728 ();
 FILLCELL_X32 FILLER_228_760 ();
 FILLCELL_X32 FILLER_228_792 ();
 FILLCELL_X32 FILLER_228_824 ();
 FILLCELL_X32 FILLER_228_856 ();
 FILLCELL_X32 FILLER_228_888 ();
 FILLCELL_X32 FILLER_228_920 ();
 FILLCELL_X32 FILLER_228_952 ();
 FILLCELL_X32 FILLER_228_984 ();
 FILLCELL_X32 FILLER_228_1016 ();
 FILLCELL_X32 FILLER_228_1048 ();
 FILLCELL_X32 FILLER_228_1080 ();
 FILLCELL_X32 FILLER_228_1112 ();
 FILLCELL_X32 FILLER_228_1144 ();
 FILLCELL_X32 FILLER_228_1176 ();
 FILLCELL_X32 FILLER_228_1208 ();
 FILLCELL_X32 FILLER_228_1240 ();
 FILLCELL_X32 FILLER_228_1272 ();
 FILLCELL_X32 FILLER_228_1304 ();
 FILLCELL_X32 FILLER_228_1336 ();
 FILLCELL_X32 FILLER_228_1368 ();
 FILLCELL_X32 FILLER_228_1400 ();
 FILLCELL_X32 FILLER_228_1432 ();
 FILLCELL_X32 FILLER_228_1464 ();
 FILLCELL_X32 FILLER_228_1496 ();
 FILLCELL_X32 FILLER_228_1528 ();
 FILLCELL_X32 FILLER_228_1560 ();
 FILLCELL_X32 FILLER_228_1592 ();
 FILLCELL_X32 FILLER_228_1624 ();
 FILLCELL_X32 FILLER_228_1656 ();
 FILLCELL_X32 FILLER_228_1688 ();
 FILLCELL_X32 FILLER_228_1720 ();
 FILLCELL_X8 FILLER_228_1752 ();
 FILLCELL_X2 FILLER_228_1760 ();
 FILLCELL_X32 FILLER_229_1 ();
 FILLCELL_X32 FILLER_229_33 ();
 FILLCELL_X32 FILLER_229_65 ();
 FILLCELL_X32 FILLER_229_97 ();
 FILLCELL_X32 FILLER_229_129 ();
 FILLCELL_X32 FILLER_229_161 ();
 FILLCELL_X32 FILLER_229_193 ();
 FILLCELL_X32 FILLER_229_225 ();
 FILLCELL_X32 FILLER_229_257 ();
 FILLCELL_X32 FILLER_229_289 ();
 FILLCELL_X32 FILLER_229_321 ();
 FILLCELL_X32 FILLER_229_353 ();
 FILLCELL_X32 FILLER_229_385 ();
 FILLCELL_X32 FILLER_229_417 ();
 FILLCELL_X32 FILLER_229_449 ();
 FILLCELL_X32 FILLER_229_481 ();
 FILLCELL_X32 FILLER_229_513 ();
 FILLCELL_X32 FILLER_229_545 ();
 FILLCELL_X32 FILLER_229_577 ();
 FILLCELL_X32 FILLER_229_609 ();
 FILLCELL_X32 FILLER_229_641 ();
 FILLCELL_X32 FILLER_229_673 ();
 FILLCELL_X32 FILLER_229_705 ();
 FILLCELL_X32 FILLER_229_737 ();
 FILLCELL_X32 FILLER_229_769 ();
 FILLCELL_X32 FILLER_229_801 ();
 FILLCELL_X32 FILLER_229_833 ();
 FILLCELL_X32 FILLER_229_865 ();
 FILLCELL_X32 FILLER_229_897 ();
 FILLCELL_X32 FILLER_229_929 ();
 FILLCELL_X32 FILLER_229_961 ();
 FILLCELL_X32 FILLER_229_993 ();
 FILLCELL_X32 FILLER_229_1025 ();
 FILLCELL_X32 FILLER_229_1057 ();
 FILLCELL_X32 FILLER_229_1089 ();
 FILLCELL_X32 FILLER_229_1121 ();
 FILLCELL_X32 FILLER_229_1153 ();
 FILLCELL_X32 FILLER_229_1185 ();
 FILLCELL_X32 FILLER_229_1217 ();
 FILLCELL_X8 FILLER_229_1249 ();
 FILLCELL_X4 FILLER_229_1257 ();
 FILLCELL_X2 FILLER_229_1261 ();
 FILLCELL_X32 FILLER_229_1264 ();
 FILLCELL_X32 FILLER_229_1296 ();
 FILLCELL_X32 FILLER_229_1328 ();
 FILLCELL_X32 FILLER_229_1360 ();
 FILLCELL_X32 FILLER_229_1392 ();
 FILLCELL_X32 FILLER_229_1424 ();
 FILLCELL_X32 FILLER_229_1456 ();
 FILLCELL_X32 FILLER_229_1488 ();
 FILLCELL_X32 FILLER_229_1520 ();
 FILLCELL_X32 FILLER_229_1552 ();
 FILLCELL_X32 FILLER_229_1584 ();
 FILLCELL_X32 FILLER_229_1616 ();
 FILLCELL_X32 FILLER_229_1648 ();
 FILLCELL_X32 FILLER_229_1680 ();
 FILLCELL_X32 FILLER_229_1712 ();
 FILLCELL_X16 FILLER_229_1744 ();
 FILLCELL_X2 FILLER_229_1760 ();
 FILLCELL_X32 FILLER_230_1 ();
 FILLCELL_X32 FILLER_230_33 ();
 FILLCELL_X32 FILLER_230_65 ();
 FILLCELL_X32 FILLER_230_97 ();
 FILLCELL_X32 FILLER_230_129 ();
 FILLCELL_X32 FILLER_230_161 ();
 FILLCELL_X32 FILLER_230_193 ();
 FILLCELL_X32 FILLER_230_225 ();
 FILLCELL_X32 FILLER_230_257 ();
 FILLCELL_X32 FILLER_230_289 ();
 FILLCELL_X32 FILLER_230_321 ();
 FILLCELL_X32 FILLER_230_353 ();
 FILLCELL_X32 FILLER_230_385 ();
 FILLCELL_X32 FILLER_230_417 ();
 FILLCELL_X32 FILLER_230_449 ();
 FILLCELL_X32 FILLER_230_481 ();
 FILLCELL_X32 FILLER_230_513 ();
 FILLCELL_X32 FILLER_230_545 ();
 FILLCELL_X32 FILLER_230_577 ();
 FILLCELL_X16 FILLER_230_609 ();
 FILLCELL_X4 FILLER_230_625 ();
 FILLCELL_X2 FILLER_230_629 ();
 FILLCELL_X32 FILLER_230_632 ();
 FILLCELL_X32 FILLER_230_664 ();
 FILLCELL_X32 FILLER_230_696 ();
 FILLCELL_X32 FILLER_230_728 ();
 FILLCELL_X32 FILLER_230_760 ();
 FILLCELL_X32 FILLER_230_792 ();
 FILLCELL_X32 FILLER_230_824 ();
 FILLCELL_X32 FILLER_230_856 ();
 FILLCELL_X32 FILLER_230_888 ();
 FILLCELL_X32 FILLER_230_920 ();
 FILLCELL_X32 FILLER_230_952 ();
 FILLCELL_X32 FILLER_230_984 ();
 FILLCELL_X32 FILLER_230_1016 ();
 FILLCELL_X32 FILLER_230_1048 ();
 FILLCELL_X32 FILLER_230_1080 ();
 FILLCELL_X32 FILLER_230_1112 ();
 FILLCELL_X32 FILLER_230_1144 ();
 FILLCELL_X32 FILLER_230_1176 ();
 FILLCELL_X32 FILLER_230_1208 ();
 FILLCELL_X32 FILLER_230_1240 ();
 FILLCELL_X32 FILLER_230_1272 ();
 FILLCELL_X32 FILLER_230_1304 ();
 FILLCELL_X32 FILLER_230_1336 ();
 FILLCELL_X32 FILLER_230_1368 ();
 FILLCELL_X32 FILLER_230_1400 ();
 FILLCELL_X32 FILLER_230_1432 ();
 FILLCELL_X32 FILLER_230_1464 ();
 FILLCELL_X32 FILLER_230_1496 ();
 FILLCELL_X32 FILLER_230_1528 ();
 FILLCELL_X32 FILLER_230_1560 ();
 FILLCELL_X32 FILLER_230_1592 ();
 FILLCELL_X32 FILLER_230_1624 ();
 FILLCELL_X32 FILLER_230_1656 ();
 FILLCELL_X32 FILLER_230_1688 ();
 FILLCELL_X32 FILLER_230_1720 ();
 FILLCELL_X8 FILLER_230_1752 ();
 FILLCELL_X2 FILLER_230_1760 ();
 FILLCELL_X32 FILLER_231_1 ();
 FILLCELL_X32 FILLER_231_33 ();
 FILLCELL_X32 FILLER_231_65 ();
 FILLCELL_X32 FILLER_231_97 ();
 FILLCELL_X32 FILLER_231_129 ();
 FILLCELL_X32 FILLER_231_161 ();
 FILLCELL_X32 FILLER_231_193 ();
 FILLCELL_X32 FILLER_231_225 ();
 FILLCELL_X32 FILLER_231_257 ();
 FILLCELL_X32 FILLER_231_289 ();
 FILLCELL_X32 FILLER_231_321 ();
 FILLCELL_X32 FILLER_231_353 ();
 FILLCELL_X32 FILLER_231_385 ();
 FILLCELL_X32 FILLER_231_417 ();
 FILLCELL_X32 FILLER_231_449 ();
 FILLCELL_X32 FILLER_231_481 ();
 FILLCELL_X32 FILLER_231_513 ();
 FILLCELL_X32 FILLER_231_545 ();
 FILLCELL_X32 FILLER_231_577 ();
 FILLCELL_X32 FILLER_231_609 ();
 FILLCELL_X32 FILLER_231_641 ();
 FILLCELL_X32 FILLER_231_673 ();
 FILLCELL_X32 FILLER_231_705 ();
 FILLCELL_X32 FILLER_231_737 ();
 FILLCELL_X32 FILLER_231_769 ();
 FILLCELL_X32 FILLER_231_801 ();
 FILLCELL_X32 FILLER_231_833 ();
 FILLCELL_X32 FILLER_231_865 ();
 FILLCELL_X32 FILLER_231_897 ();
 FILLCELL_X32 FILLER_231_929 ();
 FILLCELL_X32 FILLER_231_961 ();
 FILLCELL_X32 FILLER_231_993 ();
 FILLCELL_X32 FILLER_231_1025 ();
 FILLCELL_X32 FILLER_231_1057 ();
 FILLCELL_X32 FILLER_231_1089 ();
 FILLCELL_X32 FILLER_231_1121 ();
 FILLCELL_X32 FILLER_231_1153 ();
 FILLCELL_X32 FILLER_231_1185 ();
 FILLCELL_X32 FILLER_231_1217 ();
 FILLCELL_X8 FILLER_231_1249 ();
 FILLCELL_X4 FILLER_231_1257 ();
 FILLCELL_X2 FILLER_231_1261 ();
 FILLCELL_X32 FILLER_231_1264 ();
 FILLCELL_X32 FILLER_231_1296 ();
 FILLCELL_X32 FILLER_231_1328 ();
 FILLCELL_X32 FILLER_231_1360 ();
 FILLCELL_X32 FILLER_231_1392 ();
 FILLCELL_X32 FILLER_231_1424 ();
 FILLCELL_X32 FILLER_231_1456 ();
 FILLCELL_X32 FILLER_231_1488 ();
 FILLCELL_X32 FILLER_231_1520 ();
 FILLCELL_X32 FILLER_231_1552 ();
 FILLCELL_X32 FILLER_231_1584 ();
 FILLCELL_X32 FILLER_231_1616 ();
 FILLCELL_X32 FILLER_231_1648 ();
 FILLCELL_X32 FILLER_231_1680 ();
 FILLCELL_X32 FILLER_231_1712 ();
 FILLCELL_X16 FILLER_231_1744 ();
 FILLCELL_X2 FILLER_231_1760 ();
 FILLCELL_X32 FILLER_232_1 ();
 FILLCELL_X32 FILLER_232_33 ();
 FILLCELL_X32 FILLER_232_65 ();
 FILLCELL_X32 FILLER_232_97 ();
 FILLCELL_X32 FILLER_232_129 ();
 FILLCELL_X32 FILLER_232_161 ();
 FILLCELL_X32 FILLER_232_193 ();
 FILLCELL_X32 FILLER_232_225 ();
 FILLCELL_X32 FILLER_232_257 ();
 FILLCELL_X32 FILLER_232_289 ();
 FILLCELL_X32 FILLER_232_321 ();
 FILLCELL_X32 FILLER_232_353 ();
 FILLCELL_X32 FILLER_232_385 ();
 FILLCELL_X32 FILLER_232_417 ();
 FILLCELL_X32 FILLER_232_449 ();
 FILLCELL_X32 FILLER_232_481 ();
 FILLCELL_X32 FILLER_232_513 ();
 FILLCELL_X32 FILLER_232_545 ();
 FILLCELL_X32 FILLER_232_577 ();
 FILLCELL_X16 FILLER_232_609 ();
 FILLCELL_X4 FILLER_232_625 ();
 FILLCELL_X2 FILLER_232_629 ();
 FILLCELL_X32 FILLER_232_632 ();
 FILLCELL_X32 FILLER_232_664 ();
 FILLCELL_X32 FILLER_232_696 ();
 FILLCELL_X32 FILLER_232_728 ();
 FILLCELL_X32 FILLER_232_760 ();
 FILLCELL_X32 FILLER_232_792 ();
 FILLCELL_X32 FILLER_232_824 ();
 FILLCELL_X32 FILLER_232_856 ();
 FILLCELL_X32 FILLER_232_888 ();
 FILLCELL_X32 FILLER_232_920 ();
 FILLCELL_X32 FILLER_232_952 ();
 FILLCELL_X32 FILLER_232_984 ();
 FILLCELL_X32 FILLER_232_1016 ();
 FILLCELL_X32 FILLER_232_1048 ();
 FILLCELL_X32 FILLER_232_1080 ();
 FILLCELL_X32 FILLER_232_1112 ();
 FILLCELL_X32 FILLER_232_1144 ();
 FILLCELL_X32 FILLER_232_1176 ();
 FILLCELL_X32 FILLER_232_1208 ();
 FILLCELL_X32 FILLER_232_1240 ();
 FILLCELL_X32 FILLER_232_1272 ();
 FILLCELL_X32 FILLER_232_1304 ();
 FILLCELL_X32 FILLER_232_1336 ();
 FILLCELL_X32 FILLER_232_1368 ();
 FILLCELL_X32 FILLER_232_1400 ();
 FILLCELL_X32 FILLER_232_1432 ();
 FILLCELL_X32 FILLER_232_1464 ();
 FILLCELL_X32 FILLER_232_1496 ();
 FILLCELL_X32 FILLER_232_1528 ();
 FILLCELL_X32 FILLER_232_1560 ();
 FILLCELL_X32 FILLER_232_1592 ();
 FILLCELL_X32 FILLER_232_1624 ();
 FILLCELL_X32 FILLER_232_1656 ();
 FILLCELL_X32 FILLER_232_1688 ();
 FILLCELL_X16 FILLER_232_1720 ();
 FILLCELL_X8 FILLER_232_1736 ();
 FILLCELL_X4 FILLER_232_1744 ();
 FILLCELL_X2 FILLER_232_1748 ();
 FILLCELL_X1 FILLER_232_1750 ();
 FILLCELL_X4 FILLER_232_1758 ();
 FILLCELL_X32 FILLER_233_1 ();
 FILLCELL_X32 FILLER_233_33 ();
 FILLCELL_X32 FILLER_233_65 ();
 FILLCELL_X32 FILLER_233_97 ();
 FILLCELL_X32 FILLER_233_129 ();
 FILLCELL_X32 FILLER_233_161 ();
 FILLCELL_X32 FILLER_233_193 ();
 FILLCELL_X32 FILLER_233_225 ();
 FILLCELL_X32 FILLER_233_257 ();
 FILLCELL_X32 FILLER_233_289 ();
 FILLCELL_X32 FILLER_233_321 ();
 FILLCELL_X32 FILLER_233_353 ();
 FILLCELL_X32 FILLER_233_385 ();
 FILLCELL_X32 FILLER_233_417 ();
 FILLCELL_X32 FILLER_233_449 ();
 FILLCELL_X32 FILLER_233_481 ();
 FILLCELL_X32 FILLER_233_513 ();
 FILLCELL_X32 FILLER_233_545 ();
 FILLCELL_X32 FILLER_233_577 ();
 FILLCELL_X32 FILLER_233_609 ();
 FILLCELL_X32 FILLER_233_641 ();
 FILLCELL_X32 FILLER_233_673 ();
 FILLCELL_X32 FILLER_233_705 ();
 FILLCELL_X32 FILLER_233_737 ();
 FILLCELL_X32 FILLER_233_769 ();
 FILLCELL_X32 FILLER_233_801 ();
 FILLCELL_X32 FILLER_233_833 ();
 FILLCELL_X32 FILLER_233_865 ();
 FILLCELL_X32 FILLER_233_897 ();
 FILLCELL_X32 FILLER_233_929 ();
 FILLCELL_X32 FILLER_233_961 ();
 FILLCELL_X32 FILLER_233_993 ();
 FILLCELL_X32 FILLER_233_1025 ();
 FILLCELL_X32 FILLER_233_1057 ();
 FILLCELL_X32 FILLER_233_1089 ();
 FILLCELL_X32 FILLER_233_1121 ();
 FILLCELL_X32 FILLER_233_1153 ();
 FILLCELL_X32 FILLER_233_1185 ();
 FILLCELL_X32 FILLER_233_1217 ();
 FILLCELL_X8 FILLER_233_1249 ();
 FILLCELL_X4 FILLER_233_1257 ();
 FILLCELL_X2 FILLER_233_1261 ();
 FILLCELL_X32 FILLER_233_1264 ();
 FILLCELL_X32 FILLER_233_1296 ();
 FILLCELL_X32 FILLER_233_1328 ();
 FILLCELL_X32 FILLER_233_1360 ();
 FILLCELL_X32 FILLER_233_1392 ();
 FILLCELL_X32 FILLER_233_1424 ();
 FILLCELL_X32 FILLER_233_1456 ();
 FILLCELL_X32 FILLER_233_1488 ();
 FILLCELL_X32 FILLER_233_1520 ();
 FILLCELL_X32 FILLER_233_1552 ();
 FILLCELL_X32 FILLER_233_1584 ();
 FILLCELL_X32 FILLER_233_1616 ();
 FILLCELL_X32 FILLER_233_1648 ();
 FILLCELL_X32 FILLER_233_1680 ();
 FILLCELL_X32 FILLER_233_1712 ();
 FILLCELL_X16 FILLER_233_1744 ();
 FILLCELL_X2 FILLER_233_1760 ();
 FILLCELL_X32 FILLER_234_1 ();
 FILLCELL_X32 FILLER_234_33 ();
 FILLCELL_X32 FILLER_234_65 ();
 FILLCELL_X32 FILLER_234_97 ();
 FILLCELL_X32 FILLER_234_129 ();
 FILLCELL_X32 FILLER_234_161 ();
 FILLCELL_X32 FILLER_234_193 ();
 FILLCELL_X32 FILLER_234_225 ();
 FILLCELL_X32 FILLER_234_257 ();
 FILLCELL_X32 FILLER_234_289 ();
 FILLCELL_X32 FILLER_234_321 ();
 FILLCELL_X32 FILLER_234_353 ();
 FILLCELL_X32 FILLER_234_385 ();
 FILLCELL_X32 FILLER_234_417 ();
 FILLCELL_X32 FILLER_234_449 ();
 FILLCELL_X32 FILLER_234_481 ();
 FILLCELL_X32 FILLER_234_513 ();
 FILLCELL_X32 FILLER_234_545 ();
 FILLCELL_X32 FILLER_234_577 ();
 FILLCELL_X16 FILLER_234_609 ();
 FILLCELL_X4 FILLER_234_625 ();
 FILLCELL_X2 FILLER_234_629 ();
 FILLCELL_X32 FILLER_234_632 ();
 FILLCELL_X32 FILLER_234_664 ();
 FILLCELL_X32 FILLER_234_696 ();
 FILLCELL_X32 FILLER_234_728 ();
 FILLCELL_X32 FILLER_234_760 ();
 FILLCELL_X32 FILLER_234_792 ();
 FILLCELL_X32 FILLER_234_824 ();
 FILLCELL_X32 FILLER_234_856 ();
 FILLCELL_X32 FILLER_234_888 ();
 FILLCELL_X32 FILLER_234_920 ();
 FILLCELL_X32 FILLER_234_952 ();
 FILLCELL_X32 FILLER_234_984 ();
 FILLCELL_X32 FILLER_234_1016 ();
 FILLCELL_X32 FILLER_234_1048 ();
 FILLCELL_X32 FILLER_234_1080 ();
 FILLCELL_X32 FILLER_234_1112 ();
 FILLCELL_X32 FILLER_234_1144 ();
 FILLCELL_X32 FILLER_234_1176 ();
 FILLCELL_X32 FILLER_234_1208 ();
 FILLCELL_X32 FILLER_234_1240 ();
 FILLCELL_X32 FILLER_234_1272 ();
 FILLCELL_X32 FILLER_234_1304 ();
 FILLCELL_X32 FILLER_234_1336 ();
 FILLCELL_X32 FILLER_234_1368 ();
 FILLCELL_X32 FILLER_234_1400 ();
 FILLCELL_X32 FILLER_234_1432 ();
 FILLCELL_X32 FILLER_234_1464 ();
 FILLCELL_X32 FILLER_234_1496 ();
 FILLCELL_X32 FILLER_234_1528 ();
 FILLCELL_X32 FILLER_234_1560 ();
 FILLCELL_X32 FILLER_234_1592 ();
 FILLCELL_X32 FILLER_234_1624 ();
 FILLCELL_X32 FILLER_234_1656 ();
 FILLCELL_X32 FILLER_234_1688 ();
 FILLCELL_X32 FILLER_234_1720 ();
 FILLCELL_X8 FILLER_234_1752 ();
 FILLCELL_X2 FILLER_234_1760 ();
 FILLCELL_X32 FILLER_235_1 ();
 FILLCELL_X32 FILLER_235_33 ();
 FILLCELL_X32 FILLER_235_65 ();
 FILLCELL_X32 FILLER_235_97 ();
 FILLCELL_X32 FILLER_235_129 ();
 FILLCELL_X32 FILLER_235_161 ();
 FILLCELL_X32 FILLER_235_193 ();
 FILLCELL_X32 FILLER_235_225 ();
 FILLCELL_X32 FILLER_235_257 ();
 FILLCELL_X32 FILLER_235_289 ();
 FILLCELL_X32 FILLER_235_321 ();
 FILLCELL_X32 FILLER_235_353 ();
 FILLCELL_X32 FILLER_235_385 ();
 FILLCELL_X32 FILLER_235_417 ();
 FILLCELL_X32 FILLER_235_449 ();
 FILLCELL_X32 FILLER_235_481 ();
 FILLCELL_X32 FILLER_235_513 ();
 FILLCELL_X32 FILLER_235_545 ();
 FILLCELL_X32 FILLER_235_577 ();
 FILLCELL_X32 FILLER_235_609 ();
 FILLCELL_X32 FILLER_235_641 ();
 FILLCELL_X32 FILLER_235_673 ();
 FILLCELL_X32 FILLER_235_705 ();
 FILLCELL_X32 FILLER_235_737 ();
 FILLCELL_X32 FILLER_235_769 ();
 FILLCELL_X32 FILLER_235_801 ();
 FILLCELL_X32 FILLER_235_833 ();
 FILLCELL_X32 FILLER_235_865 ();
 FILLCELL_X32 FILLER_235_897 ();
 FILLCELL_X32 FILLER_235_929 ();
 FILLCELL_X32 FILLER_235_961 ();
 FILLCELL_X32 FILLER_235_993 ();
 FILLCELL_X32 FILLER_235_1025 ();
 FILLCELL_X32 FILLER_235_1057 ();
 FILLCELL_X32 FILLER_235_1089 ();
 FILLCELL_X32 FILLER_235_1121 ();
 FILLCELL_X32 FILLER_235_1153 ();
 FILLCELL_X32 FILLER_235_1185 ();
 FILLCELL_X32 FILLER_235_1217 ();
 FILLCELL_X8 FILLER_235_1249 ();
 FILLCELL_X4 FILLER_235_1257 ();
 FILLCELL_X2 FILLER_235_1261 ();
 FILLCELL_X32 FILLER_235_1264 ();
 FILLCELL_X32 FILLER_235_1296 ();
 FILLCELL_X32 FILLER_235_1328 ();
 FILLCELL_X32 FILLER_235_1360 ();
 FILLCELL_X32 FILLER_235_1392 ();
 FILLCELL_X32 FILLER_235_1424 ();
 FILLCELL_X32 FILLER_235_1456 ();
 FILLCELL_X32 FILLER_235_1488 ();
 FILLCELL_X32 FILLER_235_1520 ();
 FILLCELL_X32 FILLER_235_1552 ();
 FILLCELL_X32 FILLER_235_1584 ();
 FILLCELL_X32 FILLER_235_1616 ();
 FILLCELL_X32 FILLER_235_1648 ();
 FILLCELL_X32 FILLER_235_1680 ();
 FILLCELL_X32 FILLER_235_1712 ();
 FILLCELL_X16 FILLER_235_1744 ();
 FILLCELL_X2 FILLER_235_1760 ();
 FILLCELL_X4 FILLER_236_1 ();
 FILLCELL_X32 FILLER_236_8 ();
 FILLCELL_X32 FILLER_236_40 ();
 FILLCELL_X32 FILLER_236_72 ();
 FILLCELL_X32 FILLER_236_104 ();
 FILLCELL_X32 FILLER_236_136 ();
 FILLCELL_X32 FILLER_236_168 ();
 FILLCELL_X32 FILLER_236_200 ();
 FILLCELL_X32 FILLER_236_232 ();
 FILLCELL_X32 FILLER_236_264 ();
 FILLCELL_X32 FILLER_236_296 ();
 FILLCELL_X32 FILLER_236_328 ();
 FILLCELL_X32 FILLER_236_360 ();
 FILLCELL_X32 FILLER_236_392 ();
 FILLCELL_X32 FILLER_236_424 ();
 FILLCELL_X32 FILLER_236_456 ();
 FILLCELL_X32 FILLER_236_488 ();
 FILLCELL_X32 FILLER_236_520 ();
 FILLCELL_X32 FILLER_236_552 ();
 FILLCELL_X32 FILLER_236_584 ();
 FILLCELL_X8 FILLER_236_616 ();
 FILLCELL_X4 FILLER_236_624 ();
 FILLCELL_X2 FILLER_236_628 ();
 FILLCELL_X1 FILLER_236_630 ();
 FILLCELL_X32 FILLER_236_632 ();
 FILLCELL_X32 FILLER_236_664 ();
 FILLCELL_X32 FILLER_236_696 ();
 FILLCELL_X32 FILLER_236_728 ();
 FILLCELL_X32 FILLER_236_760 ();
 FILLCELL_X32 FILLER_236_792 ();
 FILLCELL_X32 FILLER_236_824 ();
 FILLCELL_X32 FILLER_236_856 ();
 FILLCELL_X32 FILLER_236_888 ();
 FILLCELL_X32 FILLER_236_920 ();
 FILLCELL_X32 FILLER_236_952 ();
 FILLCELL_X32 FILLER_236_984 ();
 FILLCELL_X32 FILLER_236_1016 ();
 FILLCELL_X32 FILLER_236_1048 ();
 FILLCELL_X32 FILLER_236_1080 ();
 FILLCELL_X32 FILLER_236_1112 ();
 FILLCELL_X32 FILLER_236_1144 ();
 FILLCELL_X32 FILLER_236_1176 ();
 FILLCELL_X32 FILLER_236_1208 ();
 FILLCELL_X32 FILLER_236_1240 ();
 FILLCELL_X32 FILLER_236_1272 ();
 FILLCELL_X32 FILLER_236_1304 ();
 FILLCELL_X32 FILLER_236_1336 ();
 FILLCELL_X32 FILLER_236_1368 ();
 FILLCELL_X32 FILLER_236_1400 ();
 FILLCELL_X32 FILLER_236_1432 ();
 FILLCELL_X32 FILLER_236_1464 ();
 FILLCELL_X32 FILLER_236_1496 ();
 FILLCELL_X32 FILLER_236_1528 ();
 FILLCELL_X32 FILLER_236_1560 ();
 FILLCELL_X32 FILLER_236_1592 ();
 FILLCELL_X32 FILLER_236_1624 ();
 FILLCELL_X32 FILLER_236_1656 ();
 FILLCELL_X32 FILLER_236_1688 ();
 FILLCELL_X32 FILLER_236_1720 ();
 FILLCELL_X8 FILLER_236_1752 ();
 FILLCELL_X2 FILLER_236_1760 ();
 FILLCELL_X8 FILLER_237_1 ();
 FILLCELL_X32 FILLER_237_12 ();
 FILLCELL_X32 FILLER_237_44 ();
 FILLCELL_X4 FILLER_237_76 ();
 FILLCELL_X32 FILLER_237_83 ();
 FILLCELL_X32 FILLER_237_115 ();
 FILLCELL_X2 FILLER_237_147 ();
 FILLCELL_X1 FILLER_237_149 ();
 FILLCELL_X32 FILLER_237_153 ();
 FILLCELL_X32 FILLER_237_185 ();
 FILLCELL_X4 FILLER_237_217 ();
 FILLCELL_X32 FILLER_237_224 ();
 FILLCELL_X32 FILLER_237_256 ();
 FILLCELL_X4 FILLER_237_288 ();
 FILLCELL_X32 FILLER_237_295 ();
 FILLCELL_X32 FILLER_237_327 ();
 FILLCELL_X4 FILLER_237_359 ();
 FILLCELL_X32 FILLER_237_366 ();
 FILLCELL_X32 FILLER_237_398 ();
 FILLCELL_X2 FILLER_237_430 ();
 FILLCELL_X1 FILLER_237_432 ();
 FILLCELL_X32 FILLER_237_436 ();
 FILLCELL_X32 FILLER_237_468 ();
 FILLCELL_X4 FILLER_237_500 ();
 FILLCELL_X32 FILLER_237_507 ();
 FILLCELL_X32 FILLER_237_539 ();
 FILLCELL_X4 FILLER_237_571 ();
 FILLCELL_X32 FILLER_237_582 ();
 FILLCELL_X16 FILLER_237_614 ();
 FILLCELL_X1 FILLER_237_630 ();
 FILLCELL_X8 FILLER_237_632 ();
 FILLCELL_X4 FILLER_237_640 ();
 FILLCELL_X2 FILLER_237_644 ();
 FILLCELL_X32 FILLER_237_653 ();
 FILLCELL_X16 FILLER_237_685 ();
 FILLCELL_X8 FILLER_237_701 ();
 FILLCELL_X4 FILLER_237_709 ();
 FILLCELL_X2 FILLER_237_713 ();
 FILLCELL_X1 FILLER_237_715 ();
 FILLCELL_X32 FILLER_237_719 ();
 FILLCELL_X32 FILLER_237_751 ();
 FILLCELL_X4 FILLER_237_783 ();
 FILLCELL_X32 FILLER_237_794 ();
 FILLCELL_X32 FILLER_237_826 ();
 FILLCELL_X32 FILLER_237_861 ();
 FILLCELL_X32 FILLER_237_893 ();
 FILLCELL_X2 FILLER_237_925 ();
 FILLCELL_X1 FILLER_237_927 ();
 FILLCELL_X32 FILLER_237_931 ();
 FILLCELL_X32 FILLER_237_963 ();
 FILLCELL_X4 FILLER_237_995 ();
 FILLCELL_X32 FILLER_237_1006 ();
 FILLCELL_X32 FILLER_237_1038 ();
 FILLCELL_X32 FILLER_237_1077 ();
 FILLCELL_X32 FILLER_237_1109 ();
 FILLCELL_X32 FILLER_237_1144 ();
 FILLCELL_X32 FILLER_237_1176 ();
 FILLCELL_X2 FILLER_237_1208 ();
 FILLCELL_X1 FILLER_237_1210 ();
 FILLCELL_X32 FILLER_237_1214 ();
 FILLCELL_X16 FILLER_237_1246 ();
 FILLCELL_X16 FILLER_237_1263 ();
 FILLCELL_X2 FILLER_237_1279 ();
 FILLCELL_X1 FILLER_237_1281 ();
 FILLCELL_X32 FILLER_237_1285 ();
 FILLCELL_X32 FILLER_237_1317 ();
 FILLCELL_X4 FILLER_237_1349 ();
 FILLCELL_X32 FILLER_237_1356 ();
 FILLCELL_X32 FILLER_237_1388 ();
 FILLCELL_X4 FILLER_237_1420 ();
 FILLCELL_X32 FILLER_237_1427 ();
 FILLCELL_X32 FILLER_237_1459 ();
 FILLCELL_X2 FILLER_237_1491 ();
 FILLCELL_X1 FILLER_237_1493 ();
 FILLCELL_X32 FILLER_237_1497 ();
 FILLCELL_X32 FILLER_237_1529 ();
 FILLCELL_X4 FILLER_237_1561 ();
 FILLCELL_X32 FILLER_237_1568 ();
 FILLCELL_X32 FILLER_237_1600 ();
 FILLCELL_X4 FILLER_237_1632 ();
 FILLCELL_X32 FILLER_237_1639 ();
 FILLCELL_X32 FILLER_237_1671 ();
 FILLCELL_X4 FILLER_237_1703 ();
 FILLCELL_X32 FILLER_237_1714 ();
 FILLCELL_X8 FILLER_237_1746 ();
 FILLCELL_X1 FILLER_237_1754 ();
 FILLCELL_X4 FILLER_237_1758 ();
 assign init_done = curr_state[1];
 assign valid_out = valid_reg_out;
endmodule
