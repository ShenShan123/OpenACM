module sram_multiplier_system (clk,
    init_done,
    init_enable,
    pe_ce,
    rst_n,
    valid_out,
    data_in,
    data_out);
 input clk;
 output init_done;
 input init_enable;
 input pe_ce;
 input rst_n;
 output valid_out;
 input [15:0] data_in;
 output [31:0] data_out;

 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire \u_multiplier/_0827_ ;
 wire \u_multiplier/_0828_ ;
 wire \u_multiplier/_0829_ ;
 wire \u_multiplier/_0830_ ;
 wire \u_multiplier/_0831_ ;
 wire \u_multiplier/_0832_ ;
 wire \u_multiplier/_0833_ ;
 wire \u_multiplier/_0834_ ;
 wire \u_multiplier/_0835_ ;
 wire \u_multiplier/_0836_ ;
 wire \u_multiplier/_0837_ ;
 wire \u_multiplier/_0838_ ;
 wire \u_multiplier/_0839_ ;
 wire \u_multiplier/_0840_ ;
 wire \u_multiplier/_0841_ ;
 wire \u_multiplier/_0842_ ;
 wire \u_multiplier/_0843_ ;
 wire \u_multiplier/_0844_ ;
 wire \u_multiplier/_0845_ ;
 wire \u_multiplier/_0846_ ;
 wire \u_multiplier/_0917_ ;
 wire \u_multiplier/_0918_ ;
 wire \u_multiplier/_0919_ ;
 wire \u_multiplier/_0920_ ;
 wire \u_multiplier/_0921_ ;
 wire \u_multiplier/_0922_ ;
 wire \u_multiplier/_0923_ ;
 wire \u_multiplier/_0924_ ;
 wire \u_multiplier/_0925_ ;
 wire \u_multiplier/_0926_ ;
 wire \u_multiplier/_0927_ ;
 wire \u_multiplier/_0928_ ;
 wire \u_multiplier/_0929_ ;
 wire \u_multiplier/_0930_ ;
 wire \u_multiplier/_0931_ ;
 wire \u_multiplier/_0932_ ;
 wire \u_multiplier/_0933_ ;
 wire \u_multiplier/_0934_ ;
 wire \u_multiplier/_0935_ ;
 wire \u_multiplier/_0936_ ;
 wire \u_multiplier/_0937_ ;
 wire \u_multiplier/_0938_ ;
 wire \u_multiplier/_0939_ ;
 wire \u_multiplier/_0940_ ;
 wire \u_multiplier/_0941_ ;
 wire \u_multiplier/_0942_ ;
 wire \u_multiplier/_0943_ ;
 wire \u_multiplier/_0944_ ;
 wire \u_multiplier/_0945_ ;
 wire \u_multiplier/_0946_ ;
 wire \u_multiplier/_0947_ ;
 wire \u_multiplier/_0948_ ;
 wire \u_multiplier/_0949_ ;
 wire \u_multiplier/_0950_ ;
 wire \u_multiplier/_0951_ ;
 wire \u_multiplier/_0952_ ;
 wire \u_multiplier/_0953_ ;
 wire \u_multiplier/_0954_ ;
 wire \u_multiplier/_0955_ ;
 wire \u_multiplier/_0956_ ;
 wire \u_multiplier/_0957_ ;
 wire \u_multiplier/_0958_ ;
 wire \u_multiplier/_0959_ ;
 wire \u_multiplier/_0960_ ;
 wire \u_multiplier/_0961_ ;
 wire \u_multiplier/_0962_ ;
 wire \u_multiplier/_0963_ ;
 wire \u_multiplier/_0964_ ;
 wire \u_multiplier/_0965_ ;
 wire \u_multiplier/_0966_ ;
 wire \u_multiplier/_0967_ ;
 wire \u_multiplier/_0968_ ;
 wire \u_multiplier/_0969_ ;
 wire \u_multiplier/_0970_ ;
 wire \u_multiplier/_0971_ ;
 wire \u_multiplier/_0972_ ;
 wire \u_multiplier/_0973_ ;
 wire \u_multiplier/_0974_ ;
 wire \u_multiplier/_0975_ ;
 wire \u_multiplier/_0976_ ;
 wire \u_multiplier/_0977_ ;
 wire \u_multiplier/_0978_ ;
 wire \u_multiplier/_0979_ ;
 wire \u_multiplier/_0980_ ;
 wire \u_multiplier/_0981_ ;
 wire \u_multiplier/_0982_ ;
 wire \u_multiplier/_0983_ ;
 wire \u_multiplier/_0984_ ;
 wire \u_multiplier/_0985_ ;
 wire \u_multiplier/_0986_ ;
 wire \u_multiplier/_0987_ ;
 wire \u_multiplier/_0988_ ;
 wire \u_multiplier/_0989_ ;
 wire \u_multiplier/_0990_ ;
 wire \u_multiplier/_0991_ ;
 wire \u_multiplier/_0992_ ;
 wire \u_multiplier/_0993_ ;
 wire \u_multiplier/_0994_ ;
 wire \u_multiplier/_0995_ ;
 wire \u_multiplier/_0996_ ;
 wire \u_multiplier/_0997_ ;
 wire \u_multiplier/_0998_ ;
 wire \u_multiplier/_0999_ ;
 wire \u_multiplier/_1000_ ;
 wire \u_multiplier/_1001_ ;
 wire \u_multiplier/_1002_ ;
 wire \u_multiplier/_1003_ ;
 wire \u_multiplier/_1004_ ;
 wire \u_multiplier/_1005_ ;
 wire \u_multiplier/_1006_ ;
 wire \u_multiplier/_1007_ ;
 wire \u_multiplier/_1008_ ;
 wire \u_multiplier/_1009_ ;
 wire \u_multiplier/_1010_ ;
 wire \u_multiplier/_1011_ ;
 wire \u_multiplier/_1012_ ;
 wire \u_multiplier/_1013_ ;
 wire \u_multiplier/_1014_ ;
 wire \u_multiplier/_1015_ ;
 wire \u_multiplier/_1016_ ;
 wire \u_multiplier/_1017_ ;
 wire \u_multiplier/_1018_ ;
 wire \u_multiplier/_1019_ ;
 wire \u_multiplier/_1020_ ;
 wire \u_multiplier/_1021_ ;
 wire \u_multiplier/_1022_ ;
 wire \u_multiplier/_1023_ ;
 wire \u_multiplier/_1024_ ;
 wire \u_multiplier/_1025_ ;
 wire \u_multiplier/_1026_ ;
 wire \u_multiplier/_1027_ ;
 wire \u_multiplier/_1028_ ;
 wire \u_multiplier/_1029_ ;
 wire \u_multiplier/_1030_ ;
 wire \u_multiplier/_1031_ ;
 wire \u_multiplier/_1032_ ;
 wire \u_multiplier/_1033_ ;
 wire \u_multiplier/_1034_ ;
 wire \u_multiplier/_1035_ ;
 wire \u_multiplier/_1036_ ;
 wire \u_multiplier/_1037_ ;
 wire \u_multiplier/_1038_ ;
 wire \u_multiplier/_1039_ ;
 wire \u_multiplier/_1040_ ;
 wire \u_multiplier/_1041_ ;
 wire \u_multiplier/_1042_ ;
 wire \u_multiplier/_1043_ ;
 wire \u_multiplier/_1044_ ;
 wire \u_multiplier/_1045_ ;
 wire \u_multiplier/_1046_ ;
 wire \u_multiplier/_1047_ ;
 wire \u_multiplier/_1048_ ;
 wire \u_multiplier/_1049_ ;
 wire \u_multiplier/_1050_ ;
 wire \u_multiplier/_1051_ ;
 wire \u_multiplier/_1052_ ;
 wire \u_multiplier/_1053_ ;
 wire \u_multiplier/_1054_ ;
 wire \u_multiplier/_1055_ ;
 wire \u_multiplier/_1056_ ;
 wire \u_multiplier/_1057_ ;
 wire \u_multiplier/_1058_ ;
 wire \u_multiplier/_1059_ ;
 wire \u_multiplier/_1060_ ;
 wire \u_multiplier/_1061_ ;
 wire \u_multiplier/_1062_ ;
 wire \u_multiplier/_1063_ ;
 wire \u_multiplier/_1064_ ;
 wire \u_multiplier/_1065_ ;
 wire \u_multiplier/_1066_ ;
 wire \u_multiplier/_1067_ ;
 wire \u_multiplier/_1068_ ;
 wire \u_multiplier/_1069_ ;
 wire \u_multiplier/_1070_ ;
 wire \u_multiplier/_1071_ ;
 wire \u_multiplier/_1072_ ;
 wire \u_multiplier/_1073_ ;
 wire \u_multiplier/_1074_ ;
 wire \u_multiplier/_1075_ ;
 wire \u_multiplier/_1076_ ;
 wire \u_multiplier/_1077_ ;
 wire \u_multiplier/_1078_ ;
 wire \u_multiplier/_1079_ ;
 wire \u_multiplier/_1080_ ;
 wire \u_multiplier/_1081_ ;
 wire \u_multiplier/_1082_ ;
 wire \u_multiplier/_1083_ ;
 wire \u_multiplier/_1084_ ;
 wire \u_multiplier/_1085_ ;
 wire \u_multiplier/_1086_ ;
 wire \u_multiplier/_1087_ ;
 wire \u_multiplier/_1088_ ;
 wire \u_multiplier/_1089_ ;
 wire \u_multiplier/_1090_ ;
 wire \u_multiplier/_1091_ ;
 wire \u_multiplier/_1092_ ;
 wire \u_multiplier/_1093_ ;
 wire \u_multiplier/_1094_ ;
 wire \u_multiplier/_1095_ ;
 wire \u_multiplier/_1096_ ;
 wire \u_multiplier/_1097_ ;
 wire \u_multiplier/_1098_ ;
 wire \u_multiplier/_1099_ ;
 wire \u_multiplier/_1100_ ;
 wire \u_multiplier/_1101_ ;
 wire \u_multiplier/_1102_ ;
 wire \u_multiplier/_1103_ ;
 wire \u_multiplier/_1104_ ;
 wire \u_multiplier/_1105_ ;
 wire \u_multiplier/_1106_ ;
 wire \u_multiplier/_1107_ ;
 wire \u_multiplier/_1108_ ;
 wire \u_multiplier/_1109_ ;
 wire \u_multiplier/_1110_ ;
 wire \u_multiplier/_1111_ ;
 wire \u_multiplier/_1112_ ;
 wire \u_multiplier/_1113_ ;
 wire \u_multiplier/_1114_ ;
 wire \u_multiplier/_1115_ ;
 wire \u_multiplier/_1116_ ;
 wire \u_multiplier/_1117_ ;
 wire \u_multiplier/_1118_ ;
 wire \u_multiplier/_1119_ ;
 wire \u_multiplier/_1120_ ;
 wire \u_multiplier/_1121_ ;
 wire \u_multiplier/_1122_ ;
 wire \u_multiplier/_1123_ ;
 wire \u_multiplier/_1124_ ;
 wire \u_multiplier/_1125_ ;
 wire \u_multiplier/_1126_ ;
 wire \u_multiplier/_1127_ ;
 wire \u_multiplier/_1128_ ;
 wire \u_multiplier/_1129_ ;
 wire \u_multiplier/_1130_ ;
 wire \u_multiplier/_1131_ ;
 wire \u_multiplier/_1132_ ;
 wire \u_multiplier/_1133_ ;
 wire \u_multiplier/_1134_ ;
 wire \u_multiplier/_1135_ ;
 wire \u_multiplier/_1136_ ;
 wire \u_multiplier/_1137_ ;
 wire \u_multiplier/_1138_ ;
 wire \u_multiplier/_1139_ ;
 wire \u_multiplier/_1140_ ;
 wire \u_multiplier/_1141_ ;
 wire \u_multiplier/_1142_ ;
 wire \u_multiplier/_1143_ ;
 wire \u_multiplier/_1144_ ;
 wire \u_multiplier/_1145_ ;
 wire \u_multiplier/_1146_ ;
 wire \u_multiplier/_1147_ ;
 wire \u_multiplier/_1148_ ;
 wire \u_multiplier/_1149_ ;
 wire \u_multiplier/_1150_ ;
 wire \u_multiplier/_1151_ ;
 wire \u_multiplier/_1152_ ;
 wire \u_multiplier/_1153_ ;
 wire \u_multiplier/_1154_ ;
 wire \u_multiplier/_1155_ ;
 wire \u_multiplier/_1156_ ;
 wire \u_multiplier/_1157_ ;
 wire \u_multiplier/_1158_ ;
 wire \u_multiplier/_1159_ ;
 wire \u_multiplier/_1160_ ;
 wire \u_multiplier/_1161_ ;
 wire \u_multiplier/_1162_ ;
 wire \u_multiplier/_1163_ ;
 wire \u_multiplier/_1164_ ;
 wire \u_multiplier/_1165_ ;
 wire \u_multiplier/_1166_ ;
 wire \u_multiplier/_1167_ ;
 wire \u_multiplier/_1168_ ;
 wire \u_multiplier/_1169_ ;
 wire \u_multiplier/_1170_ ;
 wire \u_multiplier/_1171_ ;
 wire \u_multiplier/_1172_ ;
 wire \u_multiplier/_1173_ ;
 wire \u_multiplier/_1174_ ;
 wire \u_multiplier/_1175_ ;
 wire \u_multiplier/_1176_ ;
 wire \u_multiplier/_1177_ ;
 wire \u_multiplier/_1178_ ;
 wire \u_multiplier/_1179_ ;
 wire \u_multiplier/_1180_ ;
 wire \u_multiplier/_1181_ ;
 wire \u_multiplier/_1182_ ;
 wire \u_multiplier/_1183_ ;
 wire \u_multiplier/_1184_ ;
 wire \u_multiplier/_1185_ ;
 wire \u_multiplier/_1186_ ;
 wire \u_multiplier/_1187_ ;
 wire \u_multiplier/_1188_ ;
 wire \u_multiplier/_1189_ ;
 wire \u_multiplier/_1190_ ;
 wire \u_multiplier/_1191_ ;
 wire \u_multiplier/_1192_ ;
 wire \u_multiplier/_1193_ ;
 wire \u_multiplier/_1194_ ;
 wire \u_multiplier/_1195_ ;
 wire \u_multiplier/_1196_ ;
 wire \u_multiplier/_1197_ ;
 wire \u_multiplier/_1198_ ;
 wire \u_multiplier/_1199_ ;
 wire \u_multiplier/_1200_ ;
 wire \u_multiplier/_1201_ ;
 wire \u_multiplier/_1202_ ;
 wire \u_multiplier/_1203_ ;
 wire \u_multiplier/_1204_ ;
 wire \u_multiplier/_1205_ ;
 wire \u_multiplier/_1206_ ;
 wire \u_multiplier/_1207_ ;
 wire \u_multiplier/_1208_ ;
 wire \u_multiplier/_1209_ ;
 wire \u_multiplier/_1210_ ;
 wire \u_multiplier/_1211_ ;
 wire \u_multiplier/_1212_ ;
 wire \u_multiplier/_1213_ ;
 wire \u_multiplier/_1214_ ;
 wire \u_multiplier/_1215_ ;
 wire \u_multiplier/_1216_ ;
 wire \u_multiplier/_1217_ ;
 wire \u_multiplier/_1218_ ;
 wire \u_multiplier/_1219_ ;
 wire \u_multiplier/_1220_ ;
 wire \u_multiplier/_1221_ ;
 wire \u_multiplier/_1222_ ;
 wire \u_multiplier/_1223_ ;
 wire \u_multiplier/_1224_ ;
 wire \u_multiplier/_1225_ ;
 wire \u_multiplier/_1226_ ;
 wire \u_multiplier/_1227_ ;
 wire \u_multiplier/_1228_ ;
 wire \u_multiplier/_1229_ ;
 wire \u_multiplier/_1230_ ;
 wire \u_multiplier/_1231_ ;
 wire \u_multiplier/_1232_ ;
 wire \u_multiplier/_1233_ ;
 wire \u_multiplier/_1234_ ;
 wire \u_multiplier/_1235_ ;
 wire \u_multiplier/_1236_ ;
 wire \u_multiplier/_1237_ ;
 wire \u_multiplier/_1238_ ;
 wire \u_multiplier/_1239_ ;
 wire \u_multiplier/_1240_ ;
 wire \u_multiplier/_1241_ ;
 wire \u_multiplier/_1242_ ;
 wire \u_multiplier/_1243_ ;
 wire \u_multiplier/_1244_ ;
 wire \u_multiplier/_1245_ ;
 wire \u_multiplier/_1246_ ;
 wire \u_multiplier/_1247_ ;
 wire \u_multiplier/_1248_ ;
 wire \u_multiplier/_1249_ ;
 wire \u_multiplier/_1250_ ;
 wire \u_multiplier/_1251_ ;
 wire \u_multiplier/_1252_ ;
 wire \u_multiplier/_1253_ ;
 wire \u_multiplier/_1254_ ;
 wire \u_multiplier/_1255_ ;
 wire \u_multiplier/_1256_ ;
 wire \u_multiplier/_1257_ ;
 wire \u_multiplier/_1258_ ;
 wire \u_multiplier/_1259_ ;
 wire \u_multiplier/_1260_ ;
 wire \u_multiplier/_1261_ ;
 wire \u_multiplier/_1262_ ;
 wire \u_multiplier/_1263_ ;
 wire \u_multiplier/_1264_ ;
 wire \u_multiplier/_1265_ ;
 wire \u_multiplier/_1266_ ;
 wire \u_multiplier/_1267_ ;
 wire \u_multiplier/_1268_ ;
 wire \u_multiplier/_1269_ ;
 wire \u_multiplier/_1270_ ;
 wire \u_multiplier/_1271_ ;
 wire \u_multiplier/_1272_ ;
 wire \u_multiplier/_1273_ ;
 wire \u_multiplier/_1274_ ;
 wire \u_multiplier/_1275_ ;
 wire \u_multiplier/_1276_ ;
 wire \u_multiplier/_1277_ ;
 wire \u_multiplier/_1278_ ;
 wire \u_multiplier/_1279_ ;
 wire \u_multiplier/_1280_ ;
 wire \u_multiplier/_1281_ ;
 wire \u_multiplier/_1282_ ;
 wire \u_multiplier/_1283_ ;
 wire \u_multiplier/_1284_ ;
 wire \u_multiplier/_1285_ ;
 wire \u_multiplier/_1286_ ;
 wire \u_multiplier/_1287_ ;
 wire \u_multiplier/_1288_ ;
 wire \u_multiplier/_1289_ ;
 wire \u_multiplier/_1290_ ;
 wire \u_multiplier/_1291_ ;
 wire \u_multiplier/_1292_ ;
 wire \u_multiplier/_1293_ ;
 wire \u_multiplier/_1294_ ;
 wire \u_multiplier/_1295_ ;
 wire \u_multiplier/_1296_ ;
 wire \u_multiplier/_1297_ ;
 wire \u_multiplier/_1298_ ;
 wire \u_multiplier/_1299_ ;
 wire \u_multiplier/_1300_ ;
 wire \u_multiplier/_1301_ ;
 wire \u_multiplier/_1302_ ;
 wire \u_multiplier/_1303_ ;
 wire \u_multiplier/_1304_ ;
 wire \u_multiplier/_1305_ ;
 wire \u_multiplier/_1306_ ;
 wire \u_multiplier/_1307_ ;
 wire \u_multiplier/_1308_ ;
 wire \u_multiplier/_1309_ ;
 wire \u_multiplier/_1310_ ;
 wire \u_multiplier/_1311_ ;
 wire \u_multiplier/_1312_ ;
 wire \u_multiplier/_1313_ ;
 wire \u_multiplier/_1314_ ;
 wire \u_multiplier/_1315_ ;
 wire \u_multiplier/_1316_ ;
 wire \u_multiplier/_1317_ ;
 wire \u_multiplier/_1318_ ;
 wire \u_multiplier/_1319_ ;
 wire \u_multiplier/_1320_ ;
 wire \u_multiplier/_1321_ ;
 wire \u_multiplier/_1322_ ;
 wire \u_multiplier/_1323_ ;
 wire \u_multiplier/_1324_ ;
 wire \u_multiplier/_1325_ ;
 wire \u_multiplier/_1326_ ;
 wire \u_multiplier/_1327_ ;
 wire \u_multiplier/_1328_ ;
 wire \u_multiplier/_1329_ ;
 wire \u_multiplier/_1330_ ;
 wire \u_multiplier/_1331_ ;
 wire \u_multiplier/_1332_ ;
 wire \u_multiplier/_1333_ ;
 wire \u_multiplier/_1334_ ;
 wire \u_multiplier/_1335_ ;
 wire \u_multiplier/_1336_ ;
 wire \u_multiplier/_1337_ ;
 wire \u_multiplier/_1338_ ;
 wire \u_multiplier/_1339_ ;
 wire \u_multiplier/_1340_ ;
 wire \u_multiplier/_1341_ ;
 wire \u_multiplier/_1342_ ;
 wire \u_multiplier/_1343_ ;
 wire \u_multiplier/_1344_ ;
 wire \u_multiplier/_1345_ ;
 wire \u_multiplier/_1346_ ;
 wire \u_multiplier/_1347_ ;
 wire \u_multiplier/_1348_ ;
 wire \u_multiplier/_1349_ ;
 wire \u_multiplier/_1350_ ;
 wire \u_multiplier/_1351_ ;
 wire \u_multiplier/_1352_ ;
 wire \u_multiplier/_1353_ ;
 wire \u_multiplier/_1354_ ;
 wire \u_multiplier/_1355_ ;
 wire \u_multiplier/_1356_ ;
 wire \u_multiplier/_1357_ ;
 wire \u_multiplier/_1358_ ;
 wire \u_multiplier/_1359_ ;
 wire \u_multiplier/_1360_ ;
 wire \u_multiplier/_1361_ ;
 wire \u_multiplier/_1362_ ;
 wire \u_multiplier/_1363_ ;
 wire \u_multiplier/_1364_ ;
 wire \u_multiplier/_1365_ ;
 wire \u_multiplier/_1366_ ;
 wire \u_multiplier/_1367_ ;
 wire \u_multiplier/_1368_ ;
 wire \u_multiplier/_1369_ ;
 wire \u_multiplier/_1370_ ;
 wire \u_multiplier/_1371_ ;
 wire \u_multiplier/_1372_ ;
 wire \u_multiplier/_1373_ ;
 wire \u_multiplier/_1374_ ;
 wire \u_multiplier/_1375_ ;
 wire \u_multiplier/_1376_ ;
 wire \u_multiplier/_1377_ ;
 wire \u_multiplier/_1378_ ;
 wire \u_multiplier/_1379_ ;
 wire \u_multiplier/_1380_ ;
 wire \u_multiplier/_1381_ ;
 wire \u_multiplier/_1382_ ;
 wire \u_multiplier/_1383_ ;
 wire \u_multiplier/_1384_ ;
 wire \u_multiplier/_1385_ ;
 wire \u_multiplier/_1386_ ;
 wire \u_multiplier/_1387_ ;
 wire \u_multiplier/_1388_ ;
 wire \u_multiplier/_1389_ ;
 wire \u_multiplier/_1390_ ;
 wire \u_multiplier/_1391_ ;
 wire \u_multiplier/_1392_ ;
 wire \u_multiplier/_1393_ ;
 wire \u_multiplier/_1394_ ;
 wire \u_multiplier/_1395_ ;
 wire \u_multiplier/_1396_ ;
 wire \u_multiplier/_1397_ ;
 wire \u_multiplier/_1398_ ;
 wire \u_multiplier/_1399_ ;
 wire \u_multiplier/_1400_ ;
 wire \u_multiplier/_1401_ ;
 wire \u_multiplier/_1402_ ;
 wire \u_multiplier/_1403_ ;
 wire \u_multiplier/_1404_ ;
 wire \u_multiplier/_1405_ ;
 wire \u_multiplier/_1406_ ;
 wire \u_multiplier/_1407_ ;
 wire \u_multiplier/_1408_ ;
 wire \u_multiplier/_1409_ ;
 wire \u_multiplier/_1410_ ;
 wire \u_multiplier/_1411_ ;
 wire \u_multiplier/_1412_ ;
 wire \u_multiplier/_1413_ ;
 wire \u_multiplier/_1414_ ;
 wire \u_multiplier/_1415_ ;
 wire \u_multiplier/_1416_ ;
 wire \u_multiplier/_1417_ ;
 wire \u_multiplier/_1418_ ;
 wire \u_multiplier/_1419_ ;
 wire \u_multiplier/_1420_ ;
 wire \u_multiplier/_1421_ ;
 wire \u_multiplier/_1422_ ;
 wire \u_multiplier/_1423_ ;
 wire \u_multiplier/_1424_ ;
 wire \u_multiplier/_1425_ ;
 wire \u_multiplier/_1426_ ;
 wire \u_multiplier/_1427_ ;
 wire \u_multiplier/_1428_ ;
 wire \u_multiplier/_1429_ ;
 wire \u_multiplier/_1430_ ;
 wire \u_multiplier/_1431_ ;
 wire \u_multiplier/_1432_ ;
 wire \u_multiplier/_1433_ ;
 wire \u_multiplier/_1434_ ;
 wire \u_multiplier/_1435_ ;
 wire \u_multiplier/_1436_ ;
 wire \u_multiplier/_1437_ ;
 wire \u_multiplier/_1438_ ;
 wire \u_multiplier/_1439_ ;
 wire \u_multiplier/_1440_ ;
 wire \u_multiplier/_1441_ ;
 wire \u_multiplier/_1442_ ;
 wire \u_multiplier/_1443_ ;
 wire \u_multiplier/_1444_ ;
 wire \u_multiplier/_1445_ ;
 wire \u_multiplier/_1446_ ;
 wire \u_multiplier/_1447_ ;
 wire \u_multiplier/_1448_ ;
 wire \u_multiplier/_1449_ ;
 wire \u_multiplier/_1450_ ;
 wire \u_multiplier/_1451_ ;
 wire \u_multiplier/_1452_ ;
 wire \u_multiplier/_1453_ ;
 wire \u_multiplier/_1454_ ;
 wire \u_multiplier/_1455_ ;
 wire \u_multiplier/_1456_ ;
 wire \u_multiplier/_1457_ ;
 wire \u_multiplier/_1458_ ;
 wire \u_multiplier/_1459_ ;
 wire \u_multiplier/_1460_ ;
 wire \u_multiplier/_1461_ ;
 wire \u_multiplier/_1462_ ;
 wire \u_multiplier/_1463_ ;
 wire \u_multiplier/_1464_ ;
 wire \u_multiplier/_1465_ ;
 wire \u_multiplier/_1466_ ;
 wire \u_multiplier/_1467_ ;
 wire \u_multiplier/_1468_ ;
 wire \u_multiplier/_1469_ ;
 wire \u_multiplier/_1470_ ;
 wire \u_multiplier/_1471_ ;
 wire \u_multiplier/_1472_ ;
 wire \u_multiplier/_1473_ ;
 wire \u_multiplier/_1474_ ;
 wire \u_multiplier/_1475_ ;
 wire \u_multiplier/_1476_ ;
 wire \u_multiplier/_1477_ ;
 wire \u_multiplier/_1478_ ;
 wire \u_multiplier/_1479_ ;
 wire \u_multiplier/_1480_ ;
 wire \u_multiplier/_1481_ ;
 wire \u_multiplier/_1482_ ;
 wire \u_multiplier/_1483_ ;
 wire \u_multiplier/_1484_ ;
 wire \u_multiplier/_1485_ ;
 wire \u_multiplier/_1486_ ;
 wire \u_multiplier/_1487_ ;
 wire \u_multiplier/_1488_ ;
 wire \u_multiplier/_1489_ ;
 wire \u_multiplier/_1490_ ;
 wire \u_multiplier/_1491_ ;
 wire \u_multiplier/_1492_ ;
 wire \u_multiplier/_1493_ ;
 wire \u_multiplier/_1494_ ;
 wire \u_multiplier/_1495_ ;
 wire \u_multiplier/_1496_ ;
 wire \u_multiplier/_1497_ ;
 wire \u_multiplier/_1498_ ;
 wire \u_multiplier/_1499_ ;
 wire \u_multiplier/_1500_ ;
 wire \u_multiplier/_1501_ ;
 wire \u_multiplier/_1502_ ;
 wire \u_multiplier/_1503_ ;
 wire \u_multiplier/_1504_ ;
 wire \u_multiplier/_1505_ ;
 wire \u_multiplier/_1506_ ;
 wire \u_multiplier/_1507_ ;
 wire \u_multiplier/_1508_ ;
 wire \u_multiplier/_1509_ ;
 wire \u_multiplier/_1510_ ;
 wire \u_multiplier/_1511_ ;
 wire \u_multiplier/_1512_ ;
 wire \u_multiplier/_1513_ ;
 wire \u_multiplier/_1514_ ;
 wire \u_multiplier/_1515_ ;
 wire \u_multiplier/_1516_ ;
 wire \u_multiplier/_1517_ ;
 wire \u_multiplier/_1518_ ;
 wire \u_multiplier/_1519_ ;
 wire \u_multiplier/_1520_ ;
 wire \u_multiplier/_1521_ ;
 wire \u_multiplier/_1522_ ;
 wire \u_multiplier/_1523_ ;
 wire \u_multiplier/_1524_ ;
 wire \u_multiplier/_1525_ ;
 wire \u_multiplier/_1526_ ;
 wire \u_multiplier/_1527_ ;
 wire \u_multiplier/_1528_ ;
 wire \u_multiplier/_1529_ ;
 wire \u_multiplier/_1530_ ;
 wire \u_multiplier/_1531_ ;
 wire \u_multiplier/_1532_ ;
 wire \u_multiplier/_1533_ ;
 wire \u_multiplier/_1534_ ;
 wire \u_multiplier/_1535_ ;
 wire \u_multiplier/_1536_ ;
 wire \u_multiplier/_1537_ ;
 wire \u_multiplier/_1538_ ;
 wire \u_multiplier/_1539_ ;
 wire \u_multiplier/_1540_ ;
 wire \u_multiplier/_1541_ ;
 wire \u_multiplier/_1542_ ;
 wire \u_multiplier/_1543_ ;
 wire \u_multiplier/_1544_ ;
 wire \u_multiplier/_1545_ ;
 wire \u_multiplier/_1546_ ;
 wire \u_multiplier/_1547_ ;
 wire \u_multiplier/_1548_ ;
 wire \u_multiplier/_1549_ ;
 wire \u_multiplier/_1550_ ;
 wire \u_multiplier/_1551_ ;
 wire \u_multiplier/_1552_ ;
 wire \u_multiplier/_1553_ ;
 wire \u_multiplier/_1554_ ;
 wire \u_multiplier/_1555_ ;
 wire \u_multiplier/_1556_ ;
 wire \u_multiplier/_1557_ ;
 wire \u_multiplier/_1558_ ;
 wire \u_multiplier/_1559_ ;
 wire \u_multiplier/_1560_ ;
 wire \u_multiplier/_1561_ ;
 wire \u_multiplier/_1562_ ;
 wire \u_multiplier/_1563_ ;
 wire \u_multiplier/_1564_ ;
 wire \u_multiplier/_1565_ ;
 wire \u_multiplier/_1566_ ;
 wire \u_multiplier/_1567_ ;
 wire \u_multiplier/_1568_ ;
 wire \u_multiplier/_1569_ ;
 wire \u_multiplier/_1570_ ;
 wire \u_multiplier/_1571_ ;
 wire \u_multiplier/_1572_ ;
 wire \u_multiplier/_1573_ ;
 wire \u_multiplier/_1574_ ;
 wire \u_multiplier/_1575_ ;
 wire \u_multiplier/_1576_ ;
 wire \u_multiplier/_1577_ ;
 wire \u_multiplier/_1578_ ;
 wire \u_multiplier/_1579_ ;
 wire \u_multiplier/_1580_ ;
 wire \u_multiplier/_1581_ ;
 wire \u_multiplier/_1582_ ;
 wire \u_multiplier/_1583_ ;
 wire \u_multiplier/_1584_ ;
 wire \u_multiplier/_1585_ ;
 wire \u_multiplier/_1586_ ;
 wire \u_multiplier/_1587_ ;
 wire \u_multiplier/_1588_ ;
 wire \u_multiplier/_1589_ ;
 wire \u_multiplier/_1590_ ;
 wire \u_multiplier/_1591_ ;
 wire \u_multiplier/_1592_ ;
 wire \u_multiplier/_1593_ ;
 wire \u_multiplier/_1594_ ;
 wire \u_multiplier/_1595_ ;
 wire \u_multiplier/_1596_ ;
 wire \u_multiplier/_1597_ ;
 wire \u_multiplier/_1598_ ;
 wire \u_multiplier/_1599_ ;
 wire \u_multiplier/_1600_ ;
 wire \u_multiplier/_1601_ ;
 wire \u_multiplier/_1602_ ;
 wire \u_multiplier/_1603_ ;
 wire \u_multiplier/_1604_ ;
 wire \u_multiplier/_1605_ ;
 wire \u_multiplier/_1606_ ;
 wire \u_multiplier/_1607_ ;
 wire \u_multiplier/_1608_ ;
 wire \u_multiplier/_1609_ ;
 wire \u_multiplier/_1610_ ;
 wire \u_multiplier/_1611_ ;
 wire \u_multiplier/_1612_ ;
 wire \u_multiplier/_1613_ ;
 wire \u_multiplier/_1614_ ;
 wire \u_multiplier/_1615_ ;
 wire \u_multiplier/_1616_ ;
 wire \u_multiplier/_1617_ ;
 wire \u_multiplier/_1618_ ;
 wire \u_multiplier/_1619_ ;
 wire \u_multiplier/_1620_ ;
 wire \u_multiplier/_1621_ ;
 wire \u_multiplier/_1622_ ;
 wire \u_multiplier/_1623_ ;
 wire \u_multiplier/_1624_ ;
 wire \u_multiplier/_1625_ ;
 wire \u_multiplier/_1626_ ;
 wire \u_multiplier/_1627_ ;
 wire \u_multiplier/_1628_ ;
 wire \u_multiplier/_1629_ ;
 wire \u_multiplier/_1630_ ;
 wire \u_multiplier/_1631_ ;
 wire \u_multiplier/_1632_ ;
 wire \u_multiplier/_1633_ ;
 wire \u_multiplier/_1634_ ;
 wire \u_multiplier/_1635_ ;
 wire \u_multiplier/_1636_ ;
 wire \u_multiplier/_1637_ ;
 wire \u_multiplier/_1638_ ;
 wire \u_multiplier/_1639_ ;
 wire \u_multiplier/_1640_ ;
 wire \u_multiplier/_1641_ ;
 wire \u_multiplier/_1642_ ;
 wire \u_multiplier/_1643_ ;
 wire \u_multiplier/_1644_ ;
 wire \u_multiplier/_1645_ ;
 wire \u_multiplier/_1646_ ;
 wire \u_multiplier/_1647_ ;
 wire \u_multiplier/_1648_ ;
 wire \u_multiplier/_1649_ ;
 wire \u_multiplier/_1650_ ;
 wire \u_multiplier/_1651_ ;
 wire \u_multiplier/_1652_ ;
 wire \u_multiplier/_1653_ ;
 wire \u_multiplier/_1654_ ;
 wire \u_multiplier/_1655_ ;
 wire \u_multiplier/_1656_ ;
 wire \u_multiplier/_1657_ ;
 wire \u_multiplier/_1658_ ;
 wire \u_multiplier/_1659_ ;
 wire \u_multiplier/_1660_ ;
 wire \u_multiplier/_1661_ ;
 wire \u_multiplier/_1662_ ;
 wire \u_multiplier/_1663_ ;
 wire \u_multiplier/_1664_ ;
 wire \u_multiplier/_1665_ ;
 wire \u_multiplier/_1666_ ;
 wire \u_multiplier/_1667_ ;
 wire \u_multiplier/_1668_ ;
 wire \u_multiplier/_1669_ ;
 wire \u_multiplier/_1670_ ;
 wire \u_multiplier/_1671_ ;
 wire \u_multiplier/_1672_ ;
 wire \u_multiplier/_1673_ ;
 wire \u_multiplier/_1674_ ;
 wire \u_multiplier/_1675_ ;
 wire \u_multiplier/_1676_ ;
 wire \u_multiplier/_1677_ ;
 wire \u_multiplier/_1678_ ;
 wire \u_multiplier/_1679_ ;
 wire \u_multiplier/_1680_ ;
 wire \u_multiplier/_1681_ ;
 wire \u_multiplier/_1682_ ;
 wire \u_multiplier/_1683_ ;
 wire \u_multiplier/_1684_ ;
 wire \u_multiplier/_1685_ ;
 wire \u_multiplier/_1686_ ;
 wire \u_multiplier/_1687_ ;
 wire \u_multiplier/_1688_ ;
 wire \u_multiplier/_1689_ ;
 wire \u_multiplier/_1690_ ;
 wire \u_multiplier/_1691_ ;
 wire \u_multiplier/_1692_ ;
 wire \u_multiplier/_1693_ ;
 wire \u_multiplier/_1694_ ;
 wire \u_multiplier/_1695_ ;
 wire \u_multiplier/_1696_ ;
 wire \u_multiplier/_1697_ ;
 wire \u_multiplier/_1698_ ;
 wire \u_multiplier/_1699_ ;
 wire \u_multiplier/_1700_ ;
 wire \u_multiplier/_1701_ ;
 wire \u_multiplier/_1702_ ;
 wire \u_multiplier/_1703_ ;
 wire \u_multiplier/_1704_ ;
 wire \u_multiplier/_1705_ ;
 wire \u_multiplier/_1706_ ;
 wire \u_multiplier/_1707_ ;
 wire \u_multiplier/_1708_ ;
 wire \u_multiplier/_1709_ ;
 wire \u_multiplier/_1710_ ;
 wire \u_multiplier/_1711_ ;
 wire \u_multiplier/_1712_ ;
 wire \u_multiplier/_1713_ ;
 wire \u_multiplier/_1714_ ;
 wire \u_multiplier/_1715_ ;
 wire \u_multiplier/_1716_ ;
 wire \u_multiplier/_1717_ ;
 wire \u_multiplier/_1718_ ;
 wire \u_multiplier/_1719_ ;
 wire \u_multiplier/_1720_ ;
 wire \u_multiplier/_1721_ ;
 wire \u_multiplier/_1722_ ;
 wire \u_multiplier/_1723_ ;
 wire \u_multiplier/_1724_ ;
 wire \u_multiplier/_1725_ ;
 wire \u_multiplier/_1726_ ;
 wire \u_multiplier/_1727_ ;
 wire \u_multiplier/_1728_ ;
 wire \u_multiplier/_1729_ ;
 wire \u_multiplier/_1730_ ;
 wire \u_multiplier/_1731_ ;
 wire \u_multiplier/_1732_ ;
 wire \u_multiplier/_1733_ ;
 wire \u_multiplier/_1734_ ;
 wire \u_multiplier/_1735_ ;
 wire \u_multiplier/_1736_ ;
 wire \u_multiplier/_1737_ ;
 wire \u_multiplier/_1738_ ;
 wire \u_multiplier/_1739_ ;
 wire net55;
 wire \u_multiplier/zero_x ;
 wire \u_multiplier/zero_y ;
 wire \u_multiplier/LODx/_26_ ;
 wire \u_multiplier/LODx/_27_ ;
 wire \u_multiplier/LODx/_28_ ;
 wire \u_multiplier/LODx/_29_ ;
 wire \u_multiplier/LODx/lod4_0/_09_ ;
 wire \u_multiplier/LODx/lod4_0/_10_ ;
 wire \u_multiplier/LODx/lod4_0/_11_ ;
 wire \u_multiplier/LODx/lod4_1/_09_ ;
 wire \u_multiplier/LODx/lod4_1/_10_ ;
 wire \u_multiplier/LODx/lod4_1/_11_ ;
 wire \u_multiplier/LODx/lod4_2/_09_ ;
 wire \u_multiplier/LODx/lod4_2/_10_ ;
 wire \u_multiplier/LODx/lod4_2/_11_ ;
 wire \u_multiplier/LODx/lod4_3/_09_ ;
 wire \u_multiplier/LODx/lod4_3/_10_ ;
 wire \u_multiplier/LODx/lod4_3/_11_ ;
 wire \u_multiplier/LODx/lod4_middle/_09_ ;
 wire \u_multiplier/LODx/lod4_middle/_10_ ;
 wire \u_multiplier/LODx/lod4_middle/_11_ ;
 wire \u_multiplier/LODy/_26_ ;
 wire \u_multiplier/LODy/_27_ ;
 wire \u_multiplier/LODy/_28_ ;
 wire \u_multiplier/LODy/_29_ ;
 wire \u_multiplier/LODy/lod4_0/_09_ ;
 wire \u_multiplier/LODy/lod4_0/_10_ ;
 wire \u_multiplier/LODy/lod4_0/_11_ ;
 wire \u_multiplier/LODy/lod4_1/_09_ ;
 wire \u_multiplier/LODy/lod4_1/_10_ ;
 wire \u_multiplier/LODy/lod4_1/_11_ ;
 wire \u_multiplier/LODy/lod4_2/_09_ ;
 wire \u_multiplier/LODy/lod4_2/_10_ ;
 wire \u_multiplier/LODy/lod4_2/_11_ ;
 wire \u_multiplier/LODy/lod4_3/_09_ ;
 wire \u_multiplier/LODy/lod4_3/_10_ ;
 wire \u_multiplier/LODy/lod4_3/_11_ ;
 wire \u_multiplier/LODy/lod4_middle/_09_ ;
 wire \u_multiplier/LODy/lod4_middle/_10_ ;
 wire \u_multiplier/LODy/lod4_middle/_11_ ;
 wire \u_multiplier/NOD/_11_ ;
 wire \u_multiplier/NOD/_12_ ;
 wire \u_multiplier/NOD/_13_ ;
 wire net56;
 wire \u_multiplier/NOD/nod_basic_unit15/_5_ ;
 wire \u_multiplier/NOD/nod_cels[10].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[10].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[10].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[10].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[11].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[11].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[11].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[11].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[12].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[12].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[12].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[12].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[13].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[13].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[13].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[13].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[2].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[2].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[2].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[2].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[3].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[3].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[3].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[3].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[4].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[4].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[4].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[4].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[5].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[5].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[5].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[5].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[6].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[6].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[6].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[6].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[7].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[7].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[7].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[7].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[8].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[8].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[8].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[8].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[9].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[9].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[9].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[9].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/PE/code0/_15_ ;
 wire \u_multiplier/PE/code0/_16_ ;
 wire \u_multiplier/PE/code1/_15_ ;
 wire \u_multiplier/PE/code1/_16_ ;
 wire \u_multiplier/PE/code2/_15_ ;
 wire \u_multiplier/PE/code2/_16_ ;
 wire \u_multiplier/PE/code3/_15_ ;
 wire \u_multiplier/PE/code3/_16_ ;
 wire \u_multiplier/PEx/code0/_15_ ;
 wire \u_multiplier/PEx/code0/_16_ ;
 wire \u_multiplier/PEx/code1/_15_ ;
 wire \u_multiplier/PEx/code1/_16_ ;
 wire \u_multiplier/PEx/code2/_15_ ;
 wire \u_multiplier/PEx/code2/_16_ ;
 wire \u_multiplier/PEx/code3/_15_ ;
 wire \u_multiplier/PEx/code3/_16_ ;
 wire \u_multiplier/PEy/code0/_15_ ;
 wire \u_multiplier/PEy/code0/_16_ ;
 wire \u_multiplier/PEy/code1/_15_ ;
 wire \u_multiplier/PEy/code1/_16_ ;
 wire \u_multiplier/PEy/code2/_15_ ;
 wire \u_multiplier/PEy/code2/_16_ ;
 wire \u_multiplier/PEy/code3/_15_ ;
 wire \u_multiplier/PEy/code3/_16_ ;
 wire \u_multiplier/dec/_068_ ;
 wire \u_multiplier/dec/_069_ ;
 wire \u_multiplier/dec/_070_ ;
 wire \u_multiplier/dec/_071_ ;
 wire \u_multiplier/dec/_072_ ;
 wire \u_multiplier/dec/_073_ ;
 wire \u_multiplier/dec/_074_ ;
 wire \u_multiplier/dec/_075_ ;
 wire \u_multiplier/dec/_076_ ;
 wire \u_multiplier/dec/_077_ ;
 wire \u_multiplier/dec/_078_ ;
 wire \u_multiplier/dec/_079_ ;
 wire \u_multiplier/dec/_080_ ;
 wire \u_multiplier/dec/_081_ ;
 wire \u_multiplier/dec/_082_ ;
 wire \u_multiplier/dec/_083_ ;
 wire \u_multiplier/dec/_084_ ;
 wire \u_multiplier/dec/_085_ ;
 wire \u_multiplier/dec/_086_ ;
 wire \u_multiplier/dec/_087_ ;
 wire \u_multiplier/dec/_088_ ;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire valid_reg_out;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire clknet_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire net1;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire [4:0] addr_ptr;
 wire [2:0] curr_state;
 wire [15:0] data_in_reg;
 wire [4:0] init_count;
 wire [31:0] product;
 wire [15:0] sram_rdata;
 wire [15:0] sram_rdata_reg;
 wire [3:0] \u_multiplier/K ;
 wire [3:0] \u_multiplier/LODx/select ;
 wire [15:0] \u_multiplier/LODx/z ;
 wire [3:0] \u_multiplier/LODy/select ;
 wire [15:0] \u_multiplier/LODy/z ;
 wire [12:0] \u_multiplier/NOD/t_in ;
 wire [15:0] \u_multiplier/NOD_Q1 ;
 wire [3:0] \u_multiplier/code_x ;
 wire [3:0] \u_multiplier/code_y ;
 wire [31:0] \u_multiplier/dec_out ;
 wire [15:0] \u_multiplier/kx ;
 wire [15:0] \u_multiplier/ky ;

 INV_X1 _420_ (.A(net20),
    .ZN(_238_));
 INV_X2 _421_ (.A(net19),
    .ZN(_196_));
 INV_X1 _422_ (.A(curr_state[2]),
    .ZN(_239_));
 INV_X1 _423_ (.A(net93),
    .ZN(_240_));
 INV_X1 _424_ (.A(_409_),
    .ZN(_241_));
 INV_X1 _425_ (.A(addr_ptr[0]),
    .ZN(_242_));
 INV_X1 _426_ (.A(_402_),
    .ZN(_243_));
 AND2_X4 _427_ (.A1(net20),
    .A2(net21),
    .ZN(_192_));
 INV_X1 _428_ (.A(_192_),
    .ZN(_244_));
 NAND2_X2 _429_ (.A1(net20),
    .A2(net114),
    .ZN(_197_));
 NAND2_X1 _430_ (.A1(init_count[1]),
    .A2(init_count[0]),
    .ZN(_245_));
 AND3_X1 _431_ (.A1(init_count[1]),
    .A2(init_count[0]),
    .A3(init_count[2]),
    .ZN(_246_));
 AND4_X2 _432_ (.A1(init_count[1]),
    .A2(init_count[0]),
    .A3(init_count[3]),
    .A4(init_count[2]),
    .ZN(_247_));
 AND3_X1 _433_ (.A1(net19),
    .A2(init_count[4]),
    .A3(_247_),
    .ZN(_248_));
 NOR2_X1 _434_ (.A1(_192_),
    .A2(_248_),
    .ZN(_249_));
 AOI21_X1 _435_ (.A(_249_),
    .B1(_197_),
    .B2(_244_),
    .ZN(_194_));
 NOR2_X2 _436_ (.A1(_238_),
    .A2(_196_),
    .ZN(_250_));
 NAND2_X2 _437_ (.A1(net20),
    .A2(net19),
    .ZN(_251_));
 NAND3_X1 _438_ (.A1(net18),
    .A2(net93),
    .A3(_250_),
    .ZN(_252_));
 OAI21_X1 _439_ (.A(_252_),
    .B1(_248_),
    .B2(_197_),
    .ZN(_195_));
 AOI22_X1 _440_ (.A1(net20),
    .A2(net94),
    .B1(_250_),
    .B2(net18),
    .ZN(_193_));
 AND2_X1 _441_ (.A1(net20),
    .A2(sram_rdata[0]),
    .ZN(_176_));
 AND2_X1 _442_ (.A1(net20),
    .A2(sram_rdata[1]),
    .ZN(_183_));
 AND2_X1 _443_ (.A1(net20),
    .A2(sram_rdata[2]),
    .ZN(_184_));
 AND2_X1 _444_ (.A1(net20),
    .A2(sram_rdata[3]),
    .ZN(_185_));
 AND2_X1 _445_ (.A1(net20),
    .A2(sram_rdata[4]),
    .ZN(_186_));
 AND2_X1 _446_ (.A1(net20),
    .A2(sram_rdata[5]),
    .ZN(_187_));
 AND2_X1 _447_ (.A1(net20),
    .A2(sram_rdata[6]),
    .ZN(_188_));
 AND2_X1 _448_ (.A1(net20),
    .A2(sram_rdata[7]),
    .ZN(_189_));
 AND2_X1 _449_ (.A1(net20),
    .A2(sram_rdata[8]),
    .ZN(_190_));
 AND2_X1 _450_ (.A1(net20),
    .A2(sram_rdata[9]),
    .ZN(_191_));
 AND2_X1 _451_ (.A1(net20),
    .A2(sram_rdata[10]),
    .ZN(_177_));
 AND2_X1 _452_ (.A1(net20),
    .A2(sram_rdata[11]),
    .ZN(_178_));
 AND2_X1 _453_ (.A1(net20),
    .A2(sram_rdata[12]),
    .ZN(_179_));
 AND2_X1 _454_ (.A1(net20),
    .A2(sram_rdata[13]),
    .ZN(_180_));
 AND2_X1 _455_ (.A1(net20),
    .A2(sram_rdata[14]),
    .ZN(_181_));
 AND2_X1 _456_ (.A1(net20),
    .A2(sram_rdata[15]),
    .ZN(_182_));
 AND2_X1 _457_ (.A1(product[0]),
    .A2(_192_),
    .ZN(_139_));
 AND2_X1 _458_ (.A1(product[1]),
    .A2(_192_),
    .ZN(_150_));
 AND2_X1 _459_ (.A1(product[2]),
    .A2(_192_),
    .ZN(_161_));
 AND2_X1 _460_ (.A1(product[3]),
    .A2(_192_),
    .ZN(_164_));
 AND2_X1 _461_ (.A1(product[4]),
    .A2(_192_),
    .ZN(_165_));
 AND2_X1 _462_ (.A1(product[5]),
    .A2(_192_),
    .ZN(_166_));
 AND2_X2 _463_ (.A1(product[6]),
    .A2(_192_),
    .ZN(_167_));
 AND2_X1 _464_ (.A1(product[7]),
    .A2(_192_),
    .ZN(_168_));
 AND2_X2 _465_ (.A1(product[8]),
    .A2(_192_),
    .ZN(_169_));
 AND2_X1 _466_ (.A1(product[9]),
    .A2(_192_),
    .ZN(_170_));
 AND2_X1 _467_ (.A1(product[10]),
    .A2(_192_),
    .ZN(_140_));
 AND2_X1 _468_ (.A1(product[11]),
    .A2(_192_),
    .ZN(_141_));
 AND2_X2 _469_ (.A1(product[12]),
    .A2(_192_),
    .ZN(_142_));
 AND2_X1 _470_ (.A1(product[13]),
    .A2(_192_),
    .ZN(_143_));
 AND2_X1 _471_ (.A1(product[14]),
    .A2(_192_),
    .ZN(_144_));
 AND2_X1 _472_ (.A1(product[15]),
    .A2(_192_),
    .ZN(_145_));
 AND2_X2 _473_ (.A1(product[16]),
    .A2(_192_),
    .ZN(_146_));
 AND2_X1 _474_ (.A1(product[17]),
    .A2(_192_),
    .ZN(_147_));
 AND2_X2 _475_ (.A1(product[18]),
    .A2(_192_),
    .ZN(_148_));
 AND2_X1 _476_ (.A1(product[19]),
    .A2(_192_),
    .ZN(_149_));
 AND2_X1 _477_ (.A1(product[20]),
    .A2(_192_),
    .ZN(_151_));
 AND2_X1 _478_ (.A1(product[21]),
    .A2(_192_),
    .ZN(_152_));
 AND2_X1 _479_ (.A1(product[22]),
    .A2(_192_),
    .ZN(_153_));
 AND2_X1 _480_ (.A1(product[23]),
    .A2(_192_),
    .ZN(_154_));
 AND2_X1 _481_ (.A1(product[24]),
    .A2(_192_),
    .ZN(_155_));
 AND2_X1 _482_ (.A1(product[25]),
    .A2(_192_),
    .ZN(_156_));
 AND2_X1 _483_ (.A1(product[26]),
    .A2(_192_),
    .ZN(_157_));
 AND2_X1 _484_ (.A1(product[27]),
    .A2(_192_),
    .ZN(_158_));
 AND2_X1 _485_ (.A1(product[28]),
    .A2(_192_),
    .ZN(_159_));
 AND2_X1 _486_ (.A1(product[29]),
    .A2(_192_),
    .ZN(_160_));
 AND2_X1 _487_ (.A1(product[30]),
    .A2(_192_),
    .ZN(_162_));
 AND2_X1 _488_ (.A1(product[31]),
    .A2(_192_),
    .ZN(_163_));
 AND2_X1 _489_ (.A1(net20),
    .A2(net2),
    .ZN(_123_));
 AND2_X1 _490_ (.A1(net20),
    .A2(net9),
    .ZN(_130_));
 AND2_X1 _491_ (.A1(net20),
    .A2(net10),
    .ZN(_131_));
 AND2_X1 _492_ (.A1(net20),
    .A2(net11),
    .ZN(_132_));
 AND2_X1 _493_ (.A1(net20),
    .A2(net12),
    .ZN(_133_));
 AND2_X1 _494_ (.A1(net20),
    .A2(net13),
    .ZN(_134_));
 AND2_X1 _495_ (.A1(net20),
    .A2(net14),
    .ZN(_135_));
 AND2_X1 _496_ (.A1(net20),
    .A2(net15),
    .ZN(_136_));
 AND2_X1 _497_ (.A1(net20),
    .A2(net16),
    .ZN(_137_));
 AND2_X1 _498_ (.A1(net20),
    .A2(net17),
    .ZN(_138_));
 AND2_X1 _499_ (.A1(net20),
    .A2(net3),
    .ZN(_124_));
 AND2_X1 _500_ (.A1(net20),
    .A2(net4),
    .ZN(_125_));
 AND2_X1 _501_ (.A1(net20),
    .A2(net5),
    .ZN(_126_));
 AND2_X1 _502_ (.A1(net20),
    .A2(net6),
    .ZN(_127_));
 AND2_X1 _503_ (.A1(net20),
    .A2(net7),
    .ZN(_128_));
 AND2_X1 _504_ (.A1(net20),
    .A2(net8),
    .ZN(_129_));
 NAND2_X2 _505_ (.A1(net20),
    .A2(_196_),
    .ZN(_253_));
 NAND2_X2 _506_ (.A1(_241_),
    .A2(_247_),
    .ZN(_254_));
 XNOR2_X1 _507_ (.A(net116),
    .B(_254_),
    .ZN(_255_));
 AOI22_X1 _508_ (.A1(init_count[0]),
    .A2(net21),
    .B1(_255_),
    .B2(curr_state[2]),
    .ZN(_256_));
 OAI22_X1 _509_ (.A1(net117),
    .A2(_253_),
    .B1(_256_),
    .B2(_251_),
    .ZN(_171_));
 XNOR2_X1 _510_ (.A(init_count[1]),
    .B(init_count[0]),
    .ZN(_257_));
 AOI21_X1 _511_ (.A(_239_),
    .B1(_254_),
    .B2(_257_),
    .ZN(_258_));
 AOI21_X1 _512_ (.A(_258_),
    .B1(net21),
    .B2(init_count[1]),
    .ZN(_259_));
 OAI22_X1 _513_ (.A1(net106),
    .A2(_253_),
    .B1(_259_),
    .B2(_251_),
    .ZN(_172_));
 XNOR2_X1 _514_ (.A(_407_),
    .B(_245_),
    .ZN(_260_));
 AOI21_X1 _515_ (.A(_239_),
    .B1(_254_),
    .B2(_260_),
    .ZN(_261_));
 AOI21_X1 _516_ (.A(_261_),
    .B1(net21),
    .B2(init_count[2]),
    .ZN(_262_));
 OAI22_X1 _517_ (.A1(net103),
    .A2(_253_),
    .B1(_262_),
    .B2(_251_),
    .ZN(_173_));
 OAI21_X1 _518_ (.A(curr_state[2]),
    .B1(_246_),
    .B2(init_count[3]),
    .ZN(_263_));
 AOI21_X1 _519_ (.A(_263_),
    .B1(_247_),
    .B2(_409_),
    .ZN(_264_));
 AOI21_X1 _520_ (.A(_264_),
    .B1(net21),
    .B2(init_count[3]),
    .ZN(_265_));
 OAI22_X1 _521_ (.A1(net56),
    .A2(_253_),
    .B1(_265_),
    .B2(_251_),
    .ZN(_174_));
 AND2_X1 _522_ (.A1(init_count[4]),
    .A2(net21),
    .ZN(_266_));
 OAI221_X1 _523_ (.A(_250_),
    .B1(_266_),
    .B2(curr_state[2]),
    .C1(_247_),
    .C2(init_count[4]),
    .ZN(_267_));
 OAI21_X1 _524_ (.A(_267_),
    .B1(_253_),
    .B2(net125),
    .ZN(_175_));
 AND2_X1 _525_ (.A1(curr_state[2]),
    .A2(net83),
    .ZN(_268_));
 AOI22_X1 _526_ (.A1(net21),
    .A2(_242_),
    .B1(_254_),
    .B2(_268_),
    .ZN(_269_));
 OAI22_X1 _527_ (.A1(net84),
    .A2(_253_),
    .B1(_269_),
    .B2(_251_),
    .ZN(_118_));
 AOI21_X2 _528_ (.A(_239_),
    .B1(_247_),
    .B2(init_count[4]),
    .ZN(_270_));
 AND2_X1 _529_ (.A1(addr_ptr[0]),
    .A2(addr_ptr[1]),
    .ZN(_271_));
 NOR2_X1 _530_ (.A1(_251_),
    .A2(_271_),
    .ZN(_272_));
 OAI221_X1 _531_ (.A(_272_),
    .B1(addr_ptr[1]),
    .B2(addr_ptr[0]),
    .C1(net21),
    .C2(_270_),
    .ZN(_273_));
 OAI21_X1 _532_ (.A(_273_),
    .B1(_253_),
    .B2(net78),
    .ZN(_119_));
 NAND4_X1 _533_ (.A1(addr_ptr[3]),
    .A2(addr_ptr[2]),
    .A3(net80),
    .A4(_271_),
    .ZN(_274_));
 AOI21_X2 _534_ (.A(_270_),
    .B1(_274_),
    .B2(net21),
    .ZN(_275_));
 XNOR2_X1 _535_ (.A(net119),
    .B(_271_),
    .ZN(_276_));
 NAND2_X1 _536_ (.A1(_250_),
    .A2(_276_),
    .ZN(_277_));
 OAI22_X1 _537_ (.A1(net120),
    .A2(_253_),
    .B1(_275_),
    .B2(_277_),
    .ZN(_120_));
 NAND3_X1 _538_ (.A1(net19),
    .A2(_243_),
    .A3(_271_),
    .ZN(_278_));
 XNOR2_X1 _539_ (.A(net90),
    .B(_278_),
    .ZN(_279_));
 AOI211_X1 _540_ (.A(_238_),
    .B(net91),
    .C1(_275_),
    .C2(net19),
    .ZN(_121_));
 NAND4_X1 _541_ (.A1(net19),
    .A2(addr_ptr[3]),
    .A3(addr_ptr[2]),
    .A4(_271_),
    .ZN(_280_));
 XNOR2_X1 _542_ (.A(net97),
    .B(_280_),
    .ZN(_281_));
 AOI211_X1 _543_ (.A(_238_),
    .B(net98),
    .C1(_275_),
    .C2(net19),
    .ZN(_122_));
 DFF_X1 _544_ (.D(_193_),
    .CK(clknet_3_2_0_clk),
    .Q(curr_state[0]),
    .QN(_332_));
 DFF_X2 _545_ (.D(_194_),
    .CK(clknet_3_3_0_clk),
    .Q(net21),
    .QN(_333_));
 DFF_X2 _546_ (.D(net115),
    .CK(clknet_3_2_0_clk),
    .Q(curr_state[2]),
    .QN(_334_));
 DFF_X1 _547_ (.D(_139_),
    .CK(clknet_3_6_0_clk),
    .Q(net22),
    .QN(_335_));
 DFF_X1 _548_ (.D(_150_),
    .CK(clknet_3_7_0_clk),
    .Q(net33),
    .QN(_336_));
 DFF_X1 _549_ (.D(_161_),
    .CK(clknet_3_6_0_clk),
    .Q(net44),
    .QN(_337_));
 DFF_X2 _550_ (.D(_164_),
    .CK(clknet_3_5_0_clk),
    .Q(net47),
    .QN(_338_));
 DFF_X2 _551_ (.D(_165_),
    .CK(clknet_3_5_0_clk),
    .Q(net48),
    .QN(_339_));
 DFF_X2 _552_ (.D(_166_),
    .CK(clknet_3_6_0_clk),
    .Q(net49),
    .QN(_340_));
 DFF_X1 _553_ (.D(_167_),
    .CK(clknet_3_3_0_clk),
    .Q(net50),
    .QN(_341_));
 DFF_X2 _554_ (.D(_168_),
    .CK(clknet_3_7_0_clk),
    .Q(net51),
    .QN(_342_));
 DFF_X1 _555_ (.D(_169_),
    .CK(clknet_3_3_0_clk),
    .Q(net52),
    .QN(_343_));
 DFF_X2 _556_ (.D(_170_),
    .CK(clknet_3_7_0_clk),
    .Q(net53),
    .QN(_344_));
 DFF_X2 _557_ (.D(_140_),
    .CK(clknet_3_7_0_clk),
    .Q(net23),
    .QN(_345_));
 DFF_X1 _558_ (.D(_141_),
    .CK(clknet_3_4_0_clk),
    .Q(net24),
    .QN(_346_));
 DFF_X2 _559_ (.D(_142_),
    .CK(clknet_3_3_0_clk),
    .Q(net25),
    .QN(_347_));
 DFF_X2 _560_ (.D(_143_),
    .CK(clknet_3_5_0_clk),
    .Q(net26),
    .QN(_348_));
 DFF_X2 _561_ (.D(_144_),
    .CK(clknet_3_6_0_clk),
    .Q(net27),
    .QN(_349_));
 DFF_X1 _562_ (.D(_145_),
    .CK(clknet_3_7_0_clk),
    .Q(net28),
    .QN(_350_));
 DFF_X2 _563_ (.D(_146_),
    .CK(clknet_3_2_0_clk),
    .Q(net29),
    .QN(_351_));
 DFF_X2 _564_ (.D(_147_),
    .CK(clknet_3_7_0_clk),
    .Q(net30),
    .QN(_352_));
 DFF_X2 _565_ (.D(_148_),
    .CK(clknet_3_3_0_clk),
    .Q(net31),
    .QN(_353_));
 DFF_X1 _566_ (.D(_149_),
    .CK(clknet_3_7_0_clk),
    .Q(net32),
    .QN(_354_));
 DFF_X1 _567_ (.D(_151_),
    .CK(clknet_3_2_0_clk),
    .Q(net34),
    .QN(_355_));
 DFF_X2 _568_ (.D(_152_),
    .CK(clknet_3_6_0_clk),
    .Q(net35),
    .QN(_356_));
 DFF_X2 _569_ (.D(_153_),
    .CK(clknet_3_7_0_clk),
    .Q(net36),
    .QN(_357_));
 DFF_X2 _570_ (.D(_154_),
    .CK(clknet_3_6_0_clk),
    .Q(net37),
    .QN(_358_));
 DFF_X2 _571_ (.D(_155_),
    .CK(clknet_3_6_0_clk),
    .Q(net38),
    .QN(_359_));
 DFF_X1 _572_ (.D(_156_),
    .CK(clknet_3_6_0_clk),
    .Q(net39),
    .QN(_360_));
 DFF_X2 _573_ (.D(_157_),
    .CK(clknet_3_5_0_clk),
    .Q(net40),
    .QN(_361_));
 DFF_X1 _574_ (.D(_158_),
    .CK(clknet_3_7_0_clk),
    .Q(net41),
    .QN(_362_));
 DFF_X1 _575_ (.D(_159_),
    .CK(clknet_3_5_0_clk),
    .Q(net42),
    .QN(_363_));
 DFF_X2 _576_ (.D(_160_),
    .CK(clknet_3_7_0_clk),
    .Q(net43),
    .QN(_364_));
 DFF_X2 _577_ (.D(_162_),
    .CK(clknet_3_3_0_clk),
    .Q(net45),
    .QN(_365_));
 DFF_X2 _578_ (.D(_163_),
    .CK(clknet_3_3_0_clk),
    .Q(net46),
    .QN(_366_));
 DFF_X2 _579_ (.D(_123_),
    .CK(clknet_3_6_0_clk),
    .Q(data_in_reg[0]),
    .QN(_367_));
 DFF_X2 _580_ (.D(_130_),
    .CK(clknet_3_0_0_clk),
    .Q(data_in_reg[1]),
    .QN(_368_));
 DFF_X2 _581_ (.D(_131_),
    .CK(clknet_3_5_0_clk),
    .Q(data_in_reg[2]),
    .QN(_369_));
 DFF_X2 _582_ (.D(_132_),
    .CK(clknet_3_4_0_clk),
    .Q(\u_multiplier/LODx/z [3]),
    .QN(_370_));
 DFF_X2 _583_ (.D(_133_),
    .CK(clknet_3_0_0_clk),
    .Q(data_in_reg[4]),
    .QN(_371_));
 DFF_X2 _584_ (.D(_134_),
    .CK(clknet_3_4_0_clk),
    .Q(data_in_reg[5]),
    .QN(_372_));
 DFF_X2 _585_ (.D(_135_),
    .CK(clknet_3_5_0_clk),
    .Q(data_in_reg[6]),
    .QN(_373_));
 DFF_X2 _586_ (.D(_136_),
    .CK(clknet_3_7_0_clk),
    .Q(\u_multiplier/LODx/z [7]),
    .QN(_374_));
 DFF_X2 _587_ (.D(_137_),
    .CK(clknet_3_0_0_clk),
    .Q(data_in_reg[8]),
    .QN(_375_));
 DFF_X2 _588_ (.D(_138_),
    .CK(clknet_3_0_0_clk),
    .Q(data_in_reg[9]),
    .QN(_376_));
 DFF_X2 _589_ (.D(_124_),
    .CK(clknet_3_4_0_clk),
    .Q(data_in_reg[10]),
    .QN(_377_));
 DFF_X2 _590_ (.D(_125_),
    .CK(clknet_3_5_0_clk),
    .Q(\u_multiplier/LODx/z [11]),
    .QN(_378_));
 DFF_X2 _591_ (.D(_126_),
    .CK(clknet_3_5_0_clk),
    .Q(data_in_reg[12]),
    .QN(_379_));
 DFF_X2 _592_ (.D(_127_),
    .CK(clknet_3_4_0_clk),
    .Q(data_in_reg[13]),
    .QN(_380_));
 DFF_X2 _593_ (.D(_128_),
    .CK(clknet_3_4_0_clk),
    .Q(data_in_reg[14]),
    .QN(_381_));
 DFF_X2 _594_ (.D(_129_),
    .CK(clknet_3_4_0_clk),
    .Q(\u_multiplier/LODx/z [15]),
    .QN(_382_));
 DFF_X2 _595_ (.D(_176_),
    .CK(clknet_3_0_0_clk),
    .Q(sram_rdata_reg[0]),
    .QN(_383_));
 DFF_X2 _596_ (.D(_183_),
    .CK(clknet_3_0_0_clk),
    .Q(sram_rdata_reg[1]),
    .QN(_384_));
 DFF_X2 _597_ (.D(_184_),
    .CK(clknet_3_0_0_clk),
    .Q(sram_rdata_reg[2]),
    .QN(_385_));
 DFF_X2 _598_ (.D(_185_),
    .CK(clknet_3_0_0_clk),
    .Q(\u_multiplier/LODy/z [3]),
    .QN(_386_));
 DFF_X2 _599_ (.D(_186_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[4]),
    .QN(_387_));
 DFF_X2 _600_ (.D(_187_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[5]),
    .QN(_388_));
 DFF_X2 _601_ (.D(_188_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[6]),
    .QN(_389_));
 DFF_X2 _602_ (.D(_189_),
    .CK(clknet_3_1_0_clk),
    .Q(\u_multiplier/LODy/z [7]),
    .QN(_390_));
 DFF_X2 _603_ (.D(_190_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[8]),
    .QN(_391_));
 DFF_X2 _604_ (.D(_191_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[9]),
    .QN(_392_));
 DFF_X2 _605_ (.D(_177_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[10]),
    .QN(_393_));
 DFF_X2 _606_ (.D(_178_),
    .CK(clknet_3_1_0_clk),
    .Q(\u_multiplier/LODy/z [11]),
    .QN(_394_));
 DFF_X2 _607_ (.D(_179_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[12]),
    .QN(_395_));
 DFF_X2 _608_ (.D(_180_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[13]),
    .QN(_396_));
 DFF_X2 _609_ (.D(_181_),
    .CK(clknet_3_1_0_clk),
    .Q(sram_rdata_reg[14]),
    .QN(_397_));
 DFF_X2 _610_ (.D(_182_),
    .CK(clknet_3_1_0_clk),
    .Q(\u_multiplier/LODy/z [15]),
    .QN(_398_));
 DFF_X1 _611_ (.D(_192_),
    .CK(clknet_3_7_0_clk),
    .Q(net54),
    .QN(_399_));
 DFF_X1 _612_ (.D(net85),
    .CK(clknet_3_3_0_clk),
    .Q(addr_ptr[0]),
    .QN(_400_));
 DFF_X1 _613_ (.D(net79),
    .CK(clknet_3_3_0_clk),
    .Q(addr_ptr[1]),
    .QN(_401_));
 DFF_X1 _614_ (.D(net121),
    .CK(clknet_3_3_0_clk),
    .Q(addr_ptr[2]),
    .QN(_402_));
 DFF_X1 _615_ (.D(net92),
    .CK(clknet_3_3_0_clk),
    .Q(addr_ptr[3]),
    .QN(_403_));
 DFF_X1 _616_ (.D(_122_),
    .CK(clknet_3_2_0_clk),
    .Q(addr_ptr[4]),
    .QN(_404_));
 DFF_X2 _617_ (.D(net118),
    .CK(clknet_3_2_0_clk),
    .Q(init_count[0]),
    .QN(_405_));
 DFF_X2 _618_ (.D(net107),
    .CK(clknet_3_2_0_clk),
    .Q(init_count[1]),
    .QN(_406_));
 DFF_X1 _619_ (.D(net104),
    .CK(clknet_3_2_0_clk),
    .Q(init_count[2]),
    .QN(_407_));
 DFF_X1 _620_ (.D(net57),
    .CK(clknet_3_2_0_clk),
    .Q(init_count[3]),
    .QN(_408_));
 DFF_X1 _621_ (.D(net126),
    .CK(clknet_3_3_0_clk),
    .Q(init_count[4]),
    .QN(_409_));
 SRAM_6T_CORE_32x16_MC_TB sram_inst (.ce_in(_196_),
    .we_in(_197_),
    .clk(clknet_3_0_0_clk),
    .addr_in({net81,
    net101,
    net109,
    net88,
    net112}),
    .rd_out({sram_rdata[15],
    sram_rdata[14],
    sram_rdata[13],
    sram_rdata[12],
    sram_rdata[11],
    sram_rdata[10],
    sram_rdata[9],
    sram_rdata[8],
    sram_rdata[7],
    sram_rdata[6],
    sram_rdata[5],
    sram_rdata[4],
    sram_rdata[3],
    sram_rdata[2],
    sram_rdata[1],
    sram_rdata[0]}),
    .wd_in({net123,
    net1,
    net128,
    net73,
    net82,
    net74,
    net99,
    net95,
    net110,
    net89,
    net75,
    net72,
    net76,
    net96,
    net86,
    net113}));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_0/_09_  (.A1(\u_multiplier/LODx/z [1]),
    .A2(\u_multiplier/LODx/select [0]),
    .ZN(\u_multiplier/kx [1]));
 AND2_X1 \u_multiplier/LODx/Inst_MUX214_0/_10_  (.A1(\u_multiplier/LODx/select [0]),
    .A2(\u_multiplier/LODx/z [0]),
    .ZN(\u_multiplier/kx [0]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_0/_11_  (.A1(\u_multiplier/LODx/select [0]),
    .A2(\u_multiplier/LODx/z [3]),
    .ZN(\u_multiplier/kx [3]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_0/_12_  (.A1(\u_multiplier/LODx/select [0]),
    .A2(\u_multiplier/LODx/z [2]),
    .ZN(\u_multiplier/kx [2]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_1/_09_  (.A1(\u_multiplier/LODx/z [5]),
    .A2(\u_multiplier/LODx/select [1]),
    .ZN(\u_multiplier/kx [5]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_1/_10_  (.A1(\u_multiplier/LODx/select [1]),
    .A2(\u_multiplier/LODx/z [4]),
    .ZN(\u_multiplier/kx [4]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_1/_11_  (.A1(\u_multiplier/LODx/select [1]),
    .A2(\u_multiplier/LODx/z [7]),
    .ZN(\u_multiplier/kx [7]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_1/_12_  (.A1(\u_multiplier/LODx/select [1]),
    .A2(\u_multiplier/LODx/z [6]),
    .ZN(\u_multiplier/kx [6]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_2/_09_  (.A1(\u_multiplier/LODx/z [9]),
    .A2(\u_multiplier/LODx/select [2]),
    .ZN(\u_multiplier/kx [9]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_2/_10_  (.A1(\u_multiplier/LODx/select [2]),
    .A2(\u_multiplier/LODx/z [8]),
    .ZN(\u_multiplier/kx [8]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_2/_11_  (.A1(\u_multiplier/LODx/select [2]),
    .A2(\u_multiplier/LODx/z [11]),
    .ZN(\u_multiplier/kx [11]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_2/_12_  (.A1(\u_multiplier/LODx/select [2]),
    .A2(\u_multiplier/LODx/z [10]),
    .ZN(\u_multiplier/kx [10]));
 AND2_X4 \u_multiplier/LODx/Inst_MUX214_3/_09_  (.A1(\u_multiplier/LODx/z [13]),
    .A2(\u_multiplier/LODx/select [3]),
    .ZN(\u_multiplier/kx [13]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_3/_10_  (.A1(\u_multiplier/LODx/select [3]),
    .A2(\u_multiplier/LODx/z [12]),
    .ZN(\u_multiplier/kx [12]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_3/_11_  (.A1(\u_multiplier/LODx/select [3]),
    .A2(\u_multiplier/LODx/z [15]),
    .ZN(\u_multiplier/kx [15]));
 AND2_X4 \u_multiplier/LODx/Inst_MUX214_3/_12_  (.A1(\u_multiplier/LODx/select [3]),
    .A2(\u_multiplier/LODx/z [14]),
    .ZN(\u_multiplier/kx [14]));
 OR4_X4 \u_multiplier/LODx/_31_  (.A1(data_in_reg[14]),
    .A2(\u_multiplier/LODx/z [15]),
    .A3(data_in_reg[13]),
    .A4(data_in_reg[12]),
    .ZN(\u_multiplier/LODx/select [3]));
 OR4_X4 \u_multiplier/LODx/_32_  (.A1(data_in_reg[10]),
    .A2(\u_multiplier/LODx/z [11]),
    .A3(data_in_reg[9]),
    .A4(data_in_reg[8]),
    .ZN(\u_multiplier/LODx/_28_ ));
 OR4_X2 \u_multiplier/LODx/_33_  (.A1(data_in_reg[6]),
    .A2(\u_multiplier/LODx/z [7]),
    .A3(data_in_reg[5]),
    .A4(data_in_reg[4]),
    .ZN(\u_multiplier/LODx/_27_ ));
 OR4_X1 \u_multiplier/LODx/_34_  (.A1(data_in_reg[2]),
    .A2(\u_multiplier/LODx/z [3]),
    .A3(data_in_reg[1]),
    .A4(data_in_reg[0]),
    .ZN(\u_multiplier/LODx/_26_ ));
 NOR4_X2 \u_multiplier/LODx/_35_  (.A1(\u_multiplier/LODx/select [3]),
    .A2(\u_multiplier/LODx/_28_ ),
    .A3(\u_multiplier/LODx/_27_ ),
    .A4(\u_multiplier/LODx/_26_ ),
    .ZN(\u_multiplier/zero_x ));
 INV_X1 \u_multiplier/LODx/lod4_0/_12_  (.A(data_in_reg[2]),
    .ZN(\u_multiplier/LODx/lod4_0/_10_ ));
 INV_X1 \u_multiplier/LODx/lod4_0/_13_  (.A(data_in_reg[1]),
    .ZN(\u_multiplier/LODx/lod4_0/_11_ ));
 INV_X1 \u_multiplier/LODx/lod4_0/_14_  (.A(data_in_reg[0]),
    .ZN(\u_multiplier/LODx/lod4_0/_09_ ));
 NOR2_X1 \u_multiplier/LODx/lod4_0/_15_  (.A1(\u_multiplier/LODx/lod4_0/_10_ ),
    .A2(\u_multiplier/LODx/z [3]),
    .ZN(\u_multiplier/LODx/z [2]));
 NOR3_X1 \u_multiplier/LODx/lod4_0/_16_  (.A1(data_in_reg[2]),
    .A2(\u_multiplier/LODx/z [3]),
    .A3(\u_multiplier/LODx/lod4_0/_11_ ),
    .ZN(\u_multiplier/LODx/z [1]));
 NOR4_X1 \u_multiplier/LODx/lod4_0/_17_  (.A1(data_in_reg[2]),
    .A2(\u_multiplier/LODx/z [3]),
    .A3(data_in_reg[1]),
    .A4(\u_multiplier/LODx/lod4_0/_09_ ),
    .ZN(\u_multiplier/LODx/z [0]));
 INV_X1 \u_multiplier/LODx/lod4_1/_12_  (.A(data_in_reg[6]),
    .ZN(\u_multiplier/LODx/lod4_1/_10_ ));
 INV_X1 \u_multiplier/LODx/lod4_1/_13_  (.A(data_in_reg[5]),
    .ZN(\u_multiplier/LODx/lod4_1/_11_ ));
 INV_X1 \u_multiplier/LODx/lod4_1/_14_  (.A(data_in_reg[4]),
    .ZN(\u_multiplier/LODx/lod4_1/_09_ ));
 NOR2_X1 \u_multiplier/LODx/lod4_1/_15_  (.A1(\u_multiplier/LODx/lod4_1/_10_ ),
    .A2(\u_multiplier/LODx/z [7]),
    .ZN(\u_multiplier/LODx/z [6]));
 NOR3_X1 \u_multiplier/LODx/lod4_1/_16_  (.A1(data_in_reg[6]),
    .A2(\u_multiplier/LODx/z [7]),
    .A3(\u_multiplier/LODx/lod4_1/_11_ ),
    .ZN(\u_multiplier/LODx/z [5]));
 NOR4_X1 \u_multiplier/LODx/lod4_1/_17_  (.A1(data_in_reg[6]),
    .A2(\u_multiplier/LODx/z [7]),
    .A3(data_in_reg[5]),
    .A4(\u_multiplier/LODx/lod4_1/_09_ ),
    .ZN(\u_multiplier/LODx/z [4]));
 INV_X1 \u_multiplier/LODx/lod4_2/_12_  (.A(data_in_reg[10]),
    .ZN(\u_multiplier/LODx/lod4_2/_10_ ));
 INV_X1 \u_multiplier/LODx/lod4_2/_13_  (.A(data_in_reg[9]),
    .ZN(\u_multiplier/LODx/lod4_2/_11_ ));
 INV_X1 \u_multiplier/LODx/lod4_2/_14_  (.A(data_in_reg[8]),
    .ZN(\u_multiplier/LODx/lod4_2/_09_ ));
 NOR2_X1 \u_multiplier/LODx/lod4_2/_15_  (.A1(\u_multiplier/LODx/lod4_2/_10_ ),
    .A2(\u_multiplier/LODx/z [11]),
    .ZN(\u_multiplier/LODx/z [10]));
 NOR3_X1 \u_multiplier/LODx/lod4_2/_16_  (.A1(data_in_reg[10]),
    .A2(\u_multiplier/LODx/z [11]),
    .A3(\u_multiplier/LODx/lod4_2/_11_ ),
    .ZN(\u_multiplier/LODx/z [9]));
 NOR4_X1 \u_multiplier/LODx/lod4_2/_17_  (.A1(data_in_reg[10]),
    .A2(\u_multiplier/LODx/z [11]),
    .A3(data_in_reg[9]),
    .A4(\u_multiplier/LODx/lod4_2/_09_ ),
    .ZN(\u_multiplier/LODx/z [8]));
 INV_X1 \u_multiplier/LODx/lod4_3/_12_  (.A(data_in_reg[14]),
    .ZN(\u_multiplier/LODx/lod4_3/_10_ ));
 INV_X1 \u_multiplier/LODx/lod4_3/_13_  (.A(data_in_reg[13]),
    .ZN(\u_multiplier/LODx/lod4_3/_11_ ));
 INV_X1 \u_multiplier/LODx/lod4_3/_14_  (.A(data_in_reg[12]),
    .ZN(\u_multiplier/LODx/lod4_3/_09_ ));
 NOR2_X1 \u_multiplier/LODx/lod4_3/_15_  (.A1(\u_multiplier/LODx/lod4_3/_10_ ),
    .A2(\u_multiplier/LODx/z [15]),
    .ZN(\u_multiplier/LODx/z [14]));
 NOR3_X1 \u_multiplier/LODx/lod4_3/_16_  (.A1(data_in_reg[14]),
    .A2(\u_multiplier/LODx/z [15]),
    .A3(\u_multiplier/LODx/lod4_3/_11_ ),
    .ZN(\u_multiplier/LODx/z [13]));
 NOR4_X1 \u_multiplier/LODx/lod4_3/_17_  (.A1(data_in_reg[14]),
    .A2(\u_multiplier/LODx/z [15]),
    .A3(data_in_reg[13]),
    .A4(\u_multiplier/LODx/lod4_3/_09_ ),
    .ZN(\u_multiplier/LODx/z [12]));
 INV_X1 \u_multiplier/LODx/lod4_middle/_12_  (.A(\u_multiplier/LODx/_28_ ),
    .ZN(\u_multiplier/LODx/lod4_middle/_10_ ));
 INV_X1 \u_multiplier/LODx/lod4_middle/_13_  (.A(\u_multiplier/LODx/_27_ ),
    .ZN(\u_multiplier/LODx/lod4_middle/_11_ ));
 INV_X1 \u_multiplier/LODx/lod4_middle/_14_  (.A(\u_multiplier/LODx/_26_ ),
    .ZN(\u_multiplier/LODx/lod4_middle/_09_ ));
 NOR2_X2 \u_multiplier/LODx/lod4_middle/_15_  (.A1(\u_multiplier/LODx/lod4_middle/_10_ ),
    .A2(\u_multiplier/LODx/select [3]),
    .ZN(\u_multiplier/LODx/select [2]));
 NOR3_X2 \u_multiplier/LODx/lod4_middle/_16_  (.A1(\u_multiplier/LODx/_28_ ),
    .A2(\u_multiplier/LODx/select [3]),
    .A3(\u_multiplier/LODx/lod4_middle/_11_ ),
    .ZN(\u_multiplier/LODx/select [1]));
 NOR4_X4 \u_multiplier/LODx/lod4_middle/_17_  (.A1(\u_multiplier/LODx/_28_ ),
    .A2(\u_multiplier/LODx/select [3]),
    .A3(\u_multiplier/LODx/_27_ ),
    .A4(\u_multiplier/LODx/lod4_middle/_09_ ),
    .ZN(\u_multiplier/LODx/select [0]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_0/_09_  (.A1(\u_multiplier/LODy/z [1]),
    .A2(\u_multiplier/LODy/select [0]),
    .ZN(\u_multiplier/ky [1]));
 AND2_X1 \u_multiplier/LODy/Inst_MUX214_0/_10_  (.A1(\u_multiplier/LODy/select [0]),
    .A2(\u_multiplier/LODy/z [0]),
    .ZN(\u_multiplier/ky [0]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_0/_11_  (.A1(\u_multiplier/LODy/select [0]),
    .A2(\u_multiplier/LODy/z [3]),
    .ZN(\u_multiplier/ky [3]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_0/_12_  (.A1(\u_multiplier/LODy/select [0]),
    .A2(\u_multiplier/LODy/z [2]),
    .ZN(\u_multiplier/ky [2]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_1/_09_  (.A1(\u_multiplier/LODy/z [5]),
    .A2(\u_multiplier/LODy/select [1]),
    .ZN(\u_multiplier/ky [5]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_1/_10_  (.A1(\u_multiplier/LODy/select [1]),
    .A2(\u_multiplier/LODy/z [4]),
    .ZN(\u_multiplier/ky [4]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_1/_11_  (.A1(\u_multiplier/LODy/select [1]),
    .A2(\u_multiplier/LODy/z [7]),
    .ZN(\u_multiplier/ky [7]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_1/_12_  (.A1(\u_multiplier/LODy/select [1]),
    .A2(\u_multiplier/LODy/z [6]),
    .ZN(\u_multiplier/ky [6]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_2/_09_  (.A1(\u_multiplier/LODy/z [9]),
    .A2(\u_multiplier/LODy/select [2]),
    .ZN(\u_multiplier/ky [9]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_2/_10_  (.A1(\u_multiplier/LODy/select [2]),
    .A2(\u_multiplier/LODy/z [8]),
    .ZN(\u_multiplier/ky [8]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_2/_11_  (.A1(\u_multiplier/LODy/select [2]),
    .A2(\u_multiplier/LODy/z [11]),
    .ZN(\u_multiplier/ky [11]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_2/_12_  (.A1(\u_multiplier/LODy/select [2]),
    .A2(\u_multiplier/LODy/z [10]),
    .ZN(\u_multiplier/ky [10]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_3/_09_  (.A1(\u_multiplier/LODy/z [13]),
    .A2(\u_multiplier/LODy/select [3]),
    .ZN(\u_multiplier/ky [13]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_3/_10_  (.A1(\u_multiplier/LODy/select [3]),
    .A2(\u_multiplier/LODy/z [12]),
    .ZN(\u_multiplier/ky [12]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_3/_11_  (.A1(\u_multiplier/LODy/select [3]),
    .A2(\u_multiplier/LODy/z [15]),
    .ZN(\u_multiplier/ky [15]));
 AND2_X4 \u_multiplier/LODy/Inst_MUX214_3/_12_  (.A1(\u_multiplier/LODy/select [3]),
    .A2(\u_multiplier/LODy/z [14]),
    .ZN(\u_multiplier/ky [14]));
 OR4_X4 \u_multiplier/LODy/_31_  (.A1(sram_rdata_reg[14]),
    .A2(\u_multiplier/LODy/z [15]),
    .A3(sram_rdata_reg[13]),
    .A4(sram_rdata_reg[12]),
    .ZN(\u_multiplier/LODy/select [3]));
 OR4_X4 \u_multiplier/LODy/_32_  (.A1(sram_rdata_reg[10]),
    .A2(\u_multiplier/LODy/z [11]),
    .A3(sram_rdata_reg[9]),
    .A4(sram_rdata_reg[8]),
    .ZN(\u_multiplier/LODy/_28_ ));
 OR4_X2 \u_multiplier/LODy/_33_  (.A1(sram_rdata_reg[6]),
    .A2(\u_multiplier/LODy/z [7]),
    .A3(sram_rdata_reg[5]),
    .A4(sram_rdata_reg[4]),
    .ZN(\u_multiplier/LODy/_27_ ));
 OR4_X1 \u_multiplier/LODy/_34_  (.A1(sram_rdata_reg[2]),
    .A2(\u_multiplier/LODy/z [3]),
    .A3(sram_rdata_reg[1]),
    .A4(sram_rdata_reg[0]),
    .ZN(\u_multiplier/LODy/_26_ ));
 NOR4_X2 \u_multiplier/LODy/_35_  (.A1(\u_multiplier/LODy/select [3]),
    .A2(\u_multiplier/LODy/_28_ ),
    .A3(\u_multiplier/LODy/_27_ ),
    .A4(\u_multiplier/LODy/_26_ ),
    .ZN(\u_multiplier/zero_y ));
 INV_X1 \u_multiplier/LODy/lod4_0/_12_  (.A(sram_rdata_reg[2]),
    .ZN(\u_multiplier/LODy/lod4_0/_10_ ));
 INV_X1 \u_multiplier/LODy/lod4_0/_13_  (.A(sram_rdata_reg[1]),
    .ZN(\u_multiplier/LODy/lod4_0/_11_ ));
 INV_X1 \u_multiplier/LODy/lod4_0/_14_  (.A(sram_rdata_reg[0]),
    .ZN(\u_multiplier/LODy/lod4_0/_09_ ));
 NOR2_X1 \u_multiplier/LODy/lod4_0/_15_  (.A1(\u_multiplier/LODy/lod4_0/_10_ ),
    .A2(\u_multiplier/LODy/z [3]),
    .ZN(\u_multiplier/LODy/z [2]));
 NOR3_X1 \u_multiplier/LODy/lod4_0/_16_  (.A1(sram_rdata_reg[2]),
    .A2(\u_multiplier/LODy/z [3]),
    .A3(\u_multiplier/LODy/lod4_0/_11_ ),
    .ZN(\u_multiplier/LODy/z [1]));
 NOR4_X1 \u_multiplier/LODy/lod4_0/_17_  (.A1(sram_rdata_reg[2]),
    .A2(\u_multiplier/LODy/z [3]),
    .A3(sram_rdata_reg[1]),
    .A4(\u_multiplier/LODy/lod4_0/_09_ ),
    .ZN(\u_multiplier/LODy/z [0]));
 INV_X1 \u_multiplier/LODy/lod4_1/_12_  (.A(sram_rdata_reg[6]),
    .ZN(\u_multiplier/LODy/lod4_1/_10_ ));
 INV_X1 \u_multiplier/LODy/lod4_1/_13_  (.A(sram_rdata_reg[5]),
    .ZN(\u_multiplier/LODy/lod4_1/_11_ ));
 INV_X1 \u_multiplier/LODy/lod4_1/_14_  (.A(sram_rdata_reg[4]),
    .ZN(\u_multiplier/LODy/lod4_1/_09_ ));
 NOR2_X1 \u_multiplier/LODy/lod4_1/_15_  (.A1(\u_multiplier/LODy/lod4_1/_10_ ),
    .A2(\u_multiplier/LODy/z [7]),
    .ZN(\u_multiplier/LODy/z [6]));
 NOR3_X1 \u_multiplier/LODy/lod4_1/_16_  (.A1(sram_rdata_reg[6]),
    .A2(\u_multiplier/LODy/z [7]),
    .A3(\u_multiplier/LODy/lod4_1/_11_ ),
    .ZN(\u_multiplier/LODy/z [5]));
 NOR4_X1 \u_multiplier/LODy/lod4_1/_17_  (.A1(sram_rdata_reg[6]),
    .A2(\u_multiplier/LODy/z [7]),
    .A3(sram_rdata_reg[5]),
    .A4(\u_multiplier/LODy/lod4_1/_09_ ),
    .ZN(\u_multiplier/LODy/z [4]));
 INV_X1 \u_multiplier/LODy/lod4_2/_12_  (.A(sram_rdata_reg[10]),
    .ZN(\u_multiplier/LODy/lod4_2/_10_ ));
 INV_X1 \u_multiplier/LODy/lod4_2/_13_  (.A(sram_rdata_reg[9]),
    .ZN(\u_multiplier/LODy/lod4_2/_11_ ));
 INV_X1 \u_multiplier/LODy/lod4_2/_14_  (.A(sram_rdata_reg[8]),
    .ZN(\u_multiplier/LODy/lod4_2/_09_ ));
 NOR2_X1 \u_multiplier/LODy/lod4_2/_15_  (.A1(\u_multiplier/LODy/lod4_2/_10_ ),
    .A2(\u_multiplier/LODy/z [11]),
    .ZN(\u_multiplier/LODy/z [10]));
 NOR3_X1 \u_multiplier/LODy/lod4_2/_16_  (.A1(sram_rdata_reg[10]),
    .A2(\u_multiplier/LODy/z [11]),
    .A3(\u_multiplier/LODy/lod4_2/_11_ ),
    .ZN(\u_multiplier/LODy/z [9]));
 NOR4_X1 \u_multiplier/LODy/lod4_2/_17_  (.A1(sram_rdata_reg[10]),
    .A2(\u_multiplier/LODy/z [11]),
    .A3(sram_rdata_reg[9]),
    .A4(\u_multiplier/LODy/lod4_2/_09_ ),
    .ZN(\u_multiplier/LODy/z [8]));
 INV_X1 \u_multiplier/LODy/lod4_3/_12_  (.A(sram_rdata_reg[14]),
    .ZN(\u_multiplier/LODy/lod4_3/_10_ ));
 INV_X1 \u_multiplier/LODy/lod4_3/_13_  (.A(sram_rdata_reg[13]),
    .ZN(\u_multiplier/LODy/lod4_3/_11_ ));
 INV_X1 \u_multiplier/LODy/lod4_3/_14_  (.A(sram_rdata_reg[12]),
    .ZN(\u_multiplier/LODy/lod4_3/_09_ ));
 NOR2_X1 \u_multiplier/LODy/lod4_3/_15_  (.A1(\u_multiplier/LODy/lod4_3/_10_ ),
    .A2(\u_multiplier/LODy/z [15]),
    .ZN(\u_multiplier/LODy/z [14]));
 NOR3_X1 \u_multiplier/LODy/lod4_3/_16_  (.A1(sram_rdata_reg[14]),
    .A2(\u_multiplier/LODy/z [15]),
    .A3(\u_multiplier/LODy/lod4_3/_11_ ),
    .ZN(\u_multiplier/LODy/z [13]));
 NOR4_X1 \u_multiplier/LODy/lod4_3/_17_  (.A1(sram_rdata_reg[14]),
    .A2(\u_multiplier/LODy/z [15]),
    .A3(sram_rdata_reg[13]),
    .A4(\u_multiplier/LODy/lod4_3/_09_ ),
    .ZN(\u_multiplier/LODy/z [12]));
 INV_X1 \u_multiplier/LODy/lod4_middle/_12_  (.A(\u_multiplier/LODy/_28_ ),
    .ZN(\u_multiplier/LODy/lod4_middle/_10_ ));
 INV_X1 \u_multiplier/LODy/lod4_middle/_13_  (.A(\u_multiplier/LODy/_27_ ),
    .ZN(\u_multiplier/LODy/lod4_middle/_11_ ));
 INV_X1 \u_multiplier/LODy/lod4_middle/_14_  (.A(\u_multiplier/LODy/_26_ ),
    .ZN(\u_multiplier/LODy/lod4_middle/_09_ ));
 NOR2_X2 \u_multiplier/LODy/lod4_middle/_15_  (.A1(\u_multiplier/LODy/lod4_middle/_10_ ),
    .A2(\u_multiplier/LODy/select [3]),
    .ZN(\u_multiplier/LODy/select [2]));
 NOR3_X2 \u_multiplier/LODy/lod4_middle/_16_  (.A1(\u_multiplier/LODy/_28_ ),
    .A2(\u_multiplier/LODy/select [3]),
    .A3(\u_multiplier/LODy/lod4_middle/_11_ ),
    .ZN(\u_multiplier/LODy/select [1]));
 NOR4_X4 \u_multiplier/LODy/lod4_middle/_17_  (.A1(\u_multiplier/LODy/_28_ ),
    .A2(\u_multiplier/LODy/select [3]),
    .A3(\u_multiplier/LODy/_27_ ),
    .A4(\u_multiplier/LODy/lod4_middle/_09_ ),
    .ZN(\u_multiplier/LODy/select [0]));
 INV_X1 \u_multiplier/NOD/_15_  (.A(\u_multiplier/NOD/t_in [1]),
    .ZN(\u_multiplier/NOD/_11_ ));
 INV_X1 \u_multiplier/NOD/_16_  (.A(\u_multiplier/_0833_ ),
    .ZN(\u_multiplier/NOD/_12_ ));
 INV_X1 \u_multiplier/NOD/_17_  (.A(\u_multiplier/_0827_ ),
    .ZN(\u_multiplier/NOD/_13_ ));
 NOR4_X4 \u_multiplier/NOD/_18_  (.A1(\u_multiplier/_0834_ ),
    .A2(\u_multiplier/NOD/_11_ ),
    .A3(\u_multiplier/NOD/_12_ ),
    .A4(\u_multiplier/_0827_ ),
    .ZN(\u_multiplier/NOD_Q1 [1]));
 AND2_X2 \u_multiplier/NOD/_19_  (.A1(\u_multiplier/_0831_ ),
    .A2(\u_multiplier/_0832_ ),
    .ZN(\u_multiplier/NOD_Q1 [15]));
 NOR4_X1 \u_multiplier/NOD/_20_  (.A1(\u_multiplier/_0834_ ),
    .A2(\u_multiplier/NOD/_11_ ),
    .A3(\u_multiplier/_0833_ ),
    .A4(\u_multiplier/NOD/_13_ ),
    .ZN(\u_multiplier/NOD_Q1 [0]));
 AOI21_X2 \u_multiplier/NOD/nod_basic_unit15/_7_  (.A(\u_multiplier/_0832_ ),
    .B1(\u_multiplier/_0830_ ),
    .B2(\u_multiplier/_0831_ ),
    .ZN(\u_multiplier/NOD/nod_basic_unit15/_5_ ));
 AOI21_X4 \u_multiplier/NOD/nod_basic_unit15/_8_  (.A(\u_multiplier/NOD/nod_basic_unit15/_5_ ),
    .B1(\u_multiplier/_0832_ ),
    .B2(\u_multiplier/_0831_ ),
    .ZN(\u_multiplier/NOD_Q1 [14]));
 INV_X1 \u_multiplier/NOD/nod_cels[10].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [10]),
    .ZN(\u_multiplier/NOD/nod_cels[10].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[10].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[10].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[10].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[10].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[10].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0829_ ),
    .ZN(\u_multiplier/NOD/t_in [9]));
 NOR3_X4 \u_multiplier/NOD/nod_cels[10].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[10].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0829_ ),
    .A3(\u_multiplier/NOD/nod_cels[10].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [10]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[10].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_0828_ ),
    .B1(\u_multiplier/_0840_ ),
    .B2(\u_multiplier/_0841_ ),
    .ZN(\u_multiplier/NOD/nod_cels[10].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[10].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[10].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_0828_ ),
    .B2(\u_multiplier/_0841_ ),
    .ZN(\u_multiplier/NOD/nod_cels[10].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[11].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [11]),
    .ZN(\u_multiplier/NOD/nod_cels[11].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[11].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[11].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[11].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[11].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[11].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0830_ ),
    .ZN(\u_multiplier/NOD/t_in [10]));
 NOR3_X4 \u_multiplier/NOD/nod_cels[11].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[11].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0830_ ),
    .A3(\u_multiplier/NOD/nod_cels[11].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [11]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[11].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_0829_ ),
    .B1(\u_multiplier/_0841_ ),
    .B2(\u_multiplier/_0828_ ),
    .ZN(\u_multiplier/NOD/nod_cels[11].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[11].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[11].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_0829_ ),
    .B2(\u_multiplier/_0828_ ),
    .ZN(\u_multiplier/NOD/nod_cels[11].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[12].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [12]),
    .ZN(\u_multiplier/NOD/nod_cels[12].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[12].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[12].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[12].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[12].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[12].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0831_ ),
    .ZN(\u_multiplier/NOD/t_in [11]));
 NOR3_X4 \u_multiplier/NOD/nod_cels[12].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[12].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0831_ ),
    .A3(\u_multiplier/NOD/nod_cels[12].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [12]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[12].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_0830_ ),
    .B1(\u_multiplier/_0828_ ),
    .B2(\u_multiplier/_0829_ ),
    .ZN(\u_multiplier/NOD/nod_cels[12].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[12].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[12].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_0830_ ),
    .B2(\u_multiplier/_0829_ ),
    .ZN(\u_multiplier/NOD/nod_cels[12].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[13].Nod_bits/_07_  (.A(net55),
    .ZN(\u_multiplier/NOD/nod_cels[13].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[13].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[13].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[13].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[13].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[13].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0832_ ),
    .ZN(\u_multiplier/NOD/t_in [12]));
 NOR3_X4 \u_multiplier/NOD/nod_cels[13].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[13].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0832_ ),
    .A3(\u_multiplier/NOD/nod_cels[13].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [13]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[13].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_0831_ ),
    .B1(\u_multiplier/_0829_ ),
    .B2(\u_multiplier/_0830_ ),
    .ZN(\u_multiplier/NOD/nod_cels[13].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[13].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[13].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_0831_ ),
    .B2(\u_multiplier/_0830_ ),
    .ZN(\u_multiplier/NOD/nod_cels[13].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[2].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [2]),
    .ZN(\u_multiplier/NOD/nod_cels[2].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[2].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[2].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[2].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[2].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[2].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0835_ ),
    .ZN(\u_multiplier/NOD/t_in [1]));
 NOR3_X2 \u_multiplier/NOD/nod_cels[2].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[2].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0835_ ),
    .A3(\u_multiplier/NOD/nod_cels[2].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [2]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[2].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_0834_ ),
    .B1(\u_multiplier/_0827_ ),
    .B2(\u_multiplier/_0833_ ),
    .ZN(\u_multiplier/NOD/nod_cels[2].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[2].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[2].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_0834_ ),
    .B2(\u_multiplier/_0833_ ),
    .ZN(\u_multiplier/NOD/nod_cels[2].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[3].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [3]),
    .ZN(\u_multiplier/NOD/nod_cels[3].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[3].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[3].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[3].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[3].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[3].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0836_ ),
    .ZN(\u_multiplier/NOD/t_in [2]));
 NOR3_X2 \u_multiplier/NOD/nod_cels[3].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[3].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0836_ ),
    .A3(\u_multiplier/NOD/nod_cels[3].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [3]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[3].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_0835_ ),
    .B1(\u_multiplier/_0833_ ),
    .B2(\u_multiplier/_0834_ ),
    .ZN(\u_multiplier/NOD/nod_cels[3].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[3].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[3].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_0835_ ),
    .B2(\u_multiplier/_0834_ ),
    .ZN(\u_multiplier/NOD/nod_cels[3].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[4].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [4]),
    .ZN(\u_multiplier/NOD/nod_cels[4].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[4].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[4].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[4].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[4].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[4].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0837_ ),
    .ZN(\u_multiplier/NOD/t_in [3]));
 NOR3_X2 \u_multiplier/NOD/nod_cels[4].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[4].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0837_ ),
    .A3(\u_multiplier/NOD/nod_cels[4].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [4]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[4].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_0836_ ),
    .B1(\u_multiplier/_0834_ ),
    .B2(\u_multiplier/_0835_ ),
    .ZN(\u_multiplier/NOD/nod_cels[4].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[4].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[4].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_0836_ ),
    .B2(\u_multiplier/_0835_ ),
    .ZN(\u_multiplier/NOD/nod_cels[4].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[5].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [5]),
    .ZN(\u_multiplier/NOD/nod_cels[5].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[5].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[5].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[5].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[5].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[5].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0838_ ),
    .ZN(\u_multiplier/NOD/t_in [4]));
 NOR3_X4 \u_multiplier/NOD/nod_cels[5].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[5].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0838_ ),
    .A3(\u_multiplier/NOD/nod_cels[5].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [5]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[5].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_0837_ ),
    .B1(\u_multiplier/_0835_ ),
    .B2(\u_multiplier/_0836_ ),
    .ZN(\u_multiplier/NOD/nod_cels[5].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[5].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[5].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_0837_ ),
    .B2(\u_multiplier/_0836_ ),
    .ZN(\u_multiplier/NOD/nod_cels[5].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[6].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [6]),
    .ZN(\u_multiplier/NOD/nod_cels[6].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[6].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[6].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[6].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[6].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[6].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0839_ ),
    .ZN(\u_multiplier/NOD/t_in [5]));
 NOR3_X4 \u_multiplier/NOD/nod_cels[6].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[6].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0839_ ),
    .A3(\u_multiplier/NOD/nod_cels[6].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [6]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[6].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_0838_ ),
    .B1(\u_multiplier/_0836_ ),
    .B2(\u_multiplier/_0837_ ),
    .ZN(\u_multiplier/NOD/nod_cels[6].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[6].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[6].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_0838_ ),
    .B2(\u_multiplier/_0837_ ),
    .ZN(\u_multiplier/NOD/nod_cels[6].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[7].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [7]),
    .ZN(\u_multiplier/NOD/nod_cels[7].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[7].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[7].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[7].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[7].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[7].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0840_ ),
    .ZN(\u_multiplier/NOD/t_in [6]));
 NOR3_X4 \u_multiplier/NOD/nod_cels[7].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[7].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0840_ ),
    .A3(\u_multiplier/NOD/nod_cels[7].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [7]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[7].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_0839_ ),
    .B1(\u_multiplier/_0837_ ),
    .B2(\u_multiplier/_0838_ ),
    .ZN(\u_multiplier/NOD/nod_cels[7].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[7].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[7].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_0839_ ),
    .B2(\u_multiplier/_0838_ ),
    .ZN(\u_multiplier/NOD/nod_cels[7].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[8].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [8]),
    .ZN(\u_multiplier/NOD/nod_cels[8].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[8].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[8].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[8].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[8].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[8].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0841_ ),
    .ZN(\u_multiplier/NOD/t_in [7]));
 NOR3_X2 \u_multiplier/NOD/nod_cels[8].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[8].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0841_ ),
    .A3(\u_multiplier/NOD/nod_cels[8].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [8]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[8].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_0840_ ),
    .B1(\u_multiplier/_0838_ ),
    .B2(\u_multiplier/_0839_ ),
    .ZN(\u_multiplier/NOD/nod_cels[8].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[8].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[8].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_0840_ ),
    .B2(\u_multiplier/_0839_ ),
    .ZN(\u_multiplier/NOD/nod_cels[8].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[9].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [9]),
    .ZN(\u_multiplier/NOD/nod_cels[9].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[9].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[9].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[9].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[9].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[9].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0828_ ),
    .ZN(\u_multiplier/NOD/t_in [8]));
 NOR3_X4 \u_multiplier/NOD/nod_cels[9].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[9].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0828_ ),
    .A3(\u_multiplier/NOD/nod_cels[9].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [9]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[9].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_0841_ ),
    .B1(\u_multiplier/_0839_ ),
    .B2(\u_multiplier/_0840_ ),
    .ZN(\u_multiplier/NOD/nod_cels[9].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[9].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[9].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_0841_ ),
    .B2(\u_multiplier/_0840_ ),
    .ZN(\u_multiplier/NOD/nod_cels[9].Nod_bits/tmp1 ));
 NOR4_X2 \u_multiplier/PE/code0/_17_  (.A1(\u_multiplier/NOD_Q1 [11]),
    .A2(\u_multiplier/NOD_Q1 [3]),
    .A3(\u_multiplier/NOD_Q1 [15]),
    .A4(\u_multiplier/NOD_Q1 [7]),
    .ZN(\u_multiplier/PE/code0/_15_ ));
 NOR4_X4 \u_multiplier/PE/code0/_18_  (.A1(\u_multiplier/NOD_Q1 [9]),
    .A2(\u_multiplier/NOD_Q1 [1]),
    .A3(\u_multiplier/NOD_Q1 [13]),
    .A4(\u_multiplier/NOD_Q1 [5]),
    .ZN(\u_multiplier/PE/code0/_16_ ));
 NAND2_X4 \u_multiplier/PE/code0/_19_  (.A1(\u_multiplier/PE/code0/_15_ ),
    .A2(\u_multiplier/PE/code0/_16_ ),
    .ZN(\u_multiplier/K [0]));
 NOR4_X2 \u_multiplier/PE/code1/_17_  (.A1(\u_multiplier/NOD_Q1 [11]),
    .A2(\u_multiplier/NOD_Q1 [3]),
    .A3(\u_multiplier/NOD_Q1 [15]),
    .A4(\u_multiplier/NOD_Q1 [7]),
    .ZN(\u_multiplier/PE/code1/_15_ ));
 NOR4_X4 \u_multiplier/PE/code1/_18_  (.A1(\u_multiplier/NOD_Q1 [10]),
    .A2(\u_multiplier/NOD_Q1 [2]),
    .A3(\u_multiplier/NOD_Q1 [14]),
    .A4(\u_multiplier/NOD_Q1 [6]),
    .ZN(\u_multiplier/PE/code1/_16_ ));
 NAND2_X4 \u_multiplier/PE/code1/_19_  (.A1(\u_multiplier/PE/code1/_15_ ),
    .A2(\u_multiplier/PE/code1/_16_ ),
    .ZN(\u_multiplier/K [1]));
 NOR4_X2 \u_multiplier/PE/code2/_17_  (.A1(\u_multiplier/NOD_Q1 [13]),
    .A2(\u_multiplier/NOD_Q1 [5]),
    .A3(\u_multiplier/NOD_Q1 [15]),
    .A4(\u_multiplier/NOD_Q1 [7]),
    .ZN(\u_multiplier/PE/code2/_15_ ));
 NOR4_X4 \u_multiplier/PE/code2/_18_  (.A1(\u_multiplier/NOD_Q1 [12]),
    .A2(\u_multiplier/NOD_Q1 [4]),
    .A3(\u_multiplier/NOD_Q1 [14]),
    .A4(\u_multiplier/NOD_Q1 [6]),
    .ZN(\u_multiplier/PE/code2/_16_ ));
 NAND2_X4 \u_multiplier/PE/code2/_19_  (.A1(\u_multiplier/PE/code2/_15_ ),
    .A2(\u_multiplier/PE/code2/_16_ ),
    .ZN(\u_multiplier/K [2]));
 NOR4_X2 \u_multiplier/PE/code3/_17_  (.A1(\u_multiplier/NOD_Q1 [13]),
    .A2(\u_multiplier/NOD_Q1 [9]),
    .A3(\u_multiplier/NOD_Q1 [15]),
    .A4(\u_multiplier/NOD_Q1 [11]),
    .ZN(\u_multiplier/PE/code3/_15_ ));
 NOR4_X4 \u_multiplier/PE/code3/_18_  (.A1(\u_multiplier/NOD_Q1 [12]),
    .A2(\u_multiplier/NOD_Q1 [8]),
    .A3(\u_multiplier/NOD_Q1 [14]),
    .A4(\u_multiplier/NOD_Q1 [10]),
    .ZN(\u_multiplier/PE/code3/_16_ ));
 NAND2_X4 \u_multiplier/PE/code3/_19_  (.A1(\u_multiplier/PE/code3/_15_ ),
    .A2(\u_multiplier/PE/code3/_16_ ),
    .ZN(\u_multiplier/K [3]));
 NOR4_X2 \u_multiplier/PEx/code0/_17_  (.A1(\u_multiplier/kx [11]),
    .A2(\u_multiplier/kx [3]),
    .A3(\u_multiplier/kx [15]),
    .A4(\u_multiplier/kx [7]),
    .ZN(\u_multiplier/PEx/code0/_15_ ));
 NOR4_X4 \u_multiplier/PEx/code0/_18_  (.A1(\u_multiplier/kx [9]),
    .A2(\u_multiplier/kx [1]),
    .A3(\u_multiplier/kx [13]),
    .A4(\u_multiplier/kx [5]),
    .ZN(\u_multiplier/PEx/code0/_16_ ));
 NAND2_X4 \u_multiplier/PEx/code0/_19_  (.A1(\u_multiplier/PEx/code0/_15_ ),
    .A2(\u_multiplier/PEx/code0/_16_ ),
    .ZN(\u_multiplier/code_x [0]));
 NOR4_X4 \u_multiplier/PEx/code1/_17_  (.A1(\u_multiplier/kx [11]),
    .A2(\u_multiplier/kx [3]),
    .A3(\u_multiplier/kx [15]),
    .A4(\u_multiplier/kx [7]),
    .ZN(\u_multiplier/PEx/code1/_15_ ));
 NOR4_X2 \u_multiplier/PEx/code1/_18_  (.A1(\u_multiplier/kx [10]),
    .A2(\u_multiplier/kx [2]),
    .A3(\u_multiplier/kx [14]),
    .A4(\u_multiplier/kx [6]),
    .ZN(\u_multiplier/PEx/code1/_16_ ));
 NAND2_X4 \u_multiplier/PEx/code1/_19_  (.A1(\u_multiplier/PEx/code1/_15_ ),
    .A2(\u_multiplier/PEx/code1/_16_ ),
    .ZN(\u_multiplier/code_x [1]));
 NOR4_X4 \u_multiplier/PEx/code2/_17_  (.A1(\u_multiplier/kx [13]),
    .A2(\u_multiplier/kx [5]),
    .A3(\u_multiplier/kx [15]),
    .A4(\u_multiplier/kx [7]),
    .ZN(\u_multiplier/PEx/code2/_15_ ));
 NOR4_X4 \u_multiplier/PEx/code2/_18_  (.A1(\u_multiplier/kx [12]),
    .A2(\u_multiplier/kx [4]),
    .A3(\u_multiplier/kx [14]),
    .A4(\u_multiplier/kx [6]),
    .ZN(\u_multiplier/PEx/code2/_16_ ));
 NAND2_X4 \u_multiplier/PEx/code2/_19_  (.A1(\u_multiplier/PEx/code2/_15_ ),
    .A2(\u_multiplier/PEx/code2/_16_ ),
    .ZN(\u_multiplier/code_x [2]));
 NOR4_X4 \u_multiplier/PEx/code3/_17_  (.A1(\u_multiplier/kx [13]),
    .A2(\u_multiplier/kx [9]),
    .A3(\u_multiplier/kx [15]),
    .A4(\u_multiplier/kx [11]),
    .ZN(\u_multiplier/PEx/code3/_15_ ));
 NOR4_X4 \u_multiplier/PEx/code3/_18_  (.A1(\u_multiplier/kx [12]),
    .A2(\u_multiplier/kx [8]),
    .A3(\u_multiplier/kx [14]),
    .A4(\u_multiplier/kx [10]),
    .ZN(\u_multiplier/PEx/code3/_16_ ));
 NAND2_X4 \u_multiplier/PEx/code3/_19_  (.A1(\u_multiplier/PEx/code3/_15_ ),
    .A2(\u_multiplier/PEx/code3/_16_ ),
    .ZN(\u_multiplier/code_x [3]));
 NOR4_X2 \u_multiplier/PEy/code0/_17_  (.A1(\u_multiplier/ky [11]),
    .A2(\u_multiplier/ky [3]),
    .A3(\u_multiplier/ky [15]),
    .A4(\u_multiplier/ky [7]),
    .ZN(\u_multiplier/PEy/code0/_15_ ));
 NOR4_X2 \u_multiplier/PEy/code0/_18_  (.A1(\u_multiplier/ky [9]),
    .A2(\u_multiplier/ky [1]),
    .A3(\u_multiplier/ky [13]),
    .A4(\u_multiplier/ky [5]),
    .ZN(\u_multiplier/PEy/code0/_16_ ));
 NAND2_X4 \u_multiplier/PEy/code0/_19_  (.A1(\u_multiplier/PEy/code0/_15_ ),
    .A2(\u_multiplier/PEy/code0/_16_ ),
    .ZN(\u_multiplier/code_y [0]));
 NOR4_X2 \u_multiplier/PEy/code1/_17_  (.A1(\u_multiplier/ky [11]),
    .A2(\u_multiplier/ky [3]),
    .A3(\u_multiplier/ky [15]),
    .A4(\u_multiplier/ky [7]),
    .ZN(\u_multiplier/PEy/code1/_15_ ));
 NOR4_X4 \u_multiplier/PEy/code1/_18_  (.A1(\u_multiplier/ky [10]),
    .A2(\u_multiplier/ky [2]),
    .A3(\u_multiplier/ky [14]),
    .A4(\u_multiplier/ky [6]),
    .ZN(\u_multiplier/PEy/code1/_16_ ));
 NAND2_X4 \u_multiplier/PEy/code1/_19_  (.A1(\u_multiplier/PEy/code1/_15_ ),
    .A2(\u_multiplier/PEy/code1/_16_ ),
    .ZN(\u_multiplier/code_y [1]));
 NOR4_X2 \u_multiplier/PEy/code2/_17_  (.A1(\u_multiplier/ky [13]),
    .A2(\u_multiplier/ky [5]),
    .A3(\u_multiplier/ky [15]),
    .A4(\u_multiplier/ky [7]),
    .ZN(\u_multiplier/PEy/code2/_15_ ));
 NOR4_X4 \u_multiplier/PEy/code2/_18_  (.A1(\u_multiplier/ky [12]),
    .A2(\u_multiplier/ky [4]),
    .A3(\u_multiplier/ky [14]),
    .A4(\u_multiplier/ky [6]),
    .ZN(\u_multiplier/PEy/code2/_16_ ));
 NAND2_X4 \u_multiplier/PEy/code2/_19_  (.A1(\u_multiplier/PEy/code2/_15_ ),
    .A2(\u_multiplier/PEy/code2/_16_ ),
    .ZN(\u_multiplier/code_y [2]));
 NOR4_X2 \u_multiplier/PEy/code3/_17_  (.A1(\u_multiplier/ky [13]),
    .A2(\u_multiplier/ky [9]),
    .A3(\u_multiplier/ky [15]),
    .A4(\u_multiplier/ky [11]),
    .ZN(\u_multiplier/PEy/code3/_15_ ));
 NOR4_X2 \u_multiplier/PEy/code3/_18_  (.A1(\u_multiplier/ky [12]),
    .A2(\u_multiplier/ky [8]),
    .A3(\u_multiplier/ky [14]),
    .A4(\u_multiplier/ky [10]),
    .ZN(\u_multiplier/PEy/code3/_16_ ));
 NAND2_X4 \u_multiplier/PEy/code3/_19_  (.A1(\u_multiplier/PEy/code3/_15_ ),
    .A2(\u_multiplier/PEy/code3/_16_ ),
    .ZN(\u_multiplier/code_y [3]));
 INV_X2 \u_multiplier/_1804_  (.A(\u_multiplier/code_y [0]),
    .ZN(\u_multiplier/_0930_ ));
 INV_X4 \u_multiplier/_1805_  (.A(\u_multiplier/code_y [2]),
    .ZN(\u_multiplier/_0931_ ));
 INV_X4 \u_multiplier/_1806_  (.A(\u_multiplier/code_y [3]),
    .ZN(\u_multiplier/_0932_ ));
 INV_X4 \u_multiplier/_1807_  (.A(\u_multiplier/code_x [3]),
    .ZN(\u_multiplier/_0933_ ));
 INV_X2 \u_multiplier/_1808_  (.A(\u_multiplier/code_x [0]),
    .ZN(\u_multiplier/_0934_ ));
 INV_X4 \u_multiplier/_1809_  (.A(\u_multiplier/code_x [2]),
    .ZN(\u_multiplier/_0935_ ));
 INV_X4 \u_multiplier/_1810_  (.A(\u_multiplier/K [1]),
    .ZN(\u_multiplier/_0936_ ));
 INV_X4 \u_multiplier/_1811_  (.A(\u_multiplier/K [0]),
    .ZN(\u_multiplier/_0937_ ));
 INV_X4 \u_multiplier/_1812_  (.A(\u_multiplier/K [2]),
    .ZN(\u_multiplier/_0938_ ));
 INV_X8 \u_multiplier/_1813_  (.A(\u_multiplier/K [3]),
    .ZN(\u_multiplier/_0939_ ));
 INV_X1 \u_multiplier/_1814_  (.A(\u_multiplier/dec_out [2]),
    .ZN(\u_multiplier/_0940_ ));
 INV_X1 \u_multiplier/_1815_  (.A(\u_multiplier/dec_out [26]),
    .ZN(\u_multiplier/_0941_ ));
 INV_X1 \u_multiplier/_1816_  (.A(\u_multiplier/dec_out [31]),
    .ZN(\u_multiplier/_0942_ ));
 OR2_X4 \u_multiplier/_1817_  (.A1(\u_multiplier/zero_y ),
    .A2(\u_multiplier/zero_x ),
    .ZN(\u_multiplier/_0943_ ));
 INV_X4 \u_multiplier/_1818_  (.A(\u_multiplier/_0943_ ),
    .ZN(\u_multiplier/_1739_ ));
 XOR2_X2 \u_multiplier/_1819_  (.A(\u_multiplier/ky [0]),
    .B(sram_rdata_reg[0]),
    .Z(\u_multiplier/_0944_ ));
 XNOR2_X2 \u_multiplier/_1820_  (.A(\u_multiplier/ky [0]),
    .B(sram_rdata_reg[0]),
    .ZN(\u_multiplier/_0945_ ));
 XOR2_X2 \u_multiplier/_1821_  (.A(\u_multiplier/ky [9]),
    .B(sram_rdata_reg[9]),
    .Z(\u_multiplier/_0946_ ));
 XNOR2_X2 \u_multiplier/_1822_  (.A(\u_multiplier/ky [9]),
    .B(sram_rdata_reg[9]),
    .ZN(\u_multiplier/_0947_ ));
 XOR2_X2 \u_multiplier/_1823_  (.A(\u_multiplier/kx [9]),
    .B(data_in_reg[9]),
    .Z(\u_multiplier/_0948_ ));
 NOR2_X1 \u_multiplier/_1824_  (.A1(\u_multiplier/_0947_ ),
    .A2(\u_multiplier/_0948_ ),
    .ZN(\u_multiplier/_0949_ ));
 XOR2_X2 \u_multiplier/_1825_  (.A(\u_multiplier/ky [8]),
    .B(sram_rdata_reg[8]),
    .Z(\u_multiplier/_0950_ ));
 XNOR2_X2 \u_multiplier/_1826_  (.A(\u_multiplier/ky [8]),
    .B(sram_rdata_reg[8]),
    .ZN(\u_multiplier/_0951_ ));
 XOR2_X2 \u_multiplier/_1827_  (.A(\u_multiplier/kx [8]),
    .B(data_in_reg[8]),
    .Z(\u_multiplier/_0952_ ));
 AND2_X1 \u_multiplier/_1828_  (.A1(\u_multiplier/_0951_ ),
    .A2(\u_multiplier/_0952_ ),
    .ZN(\u_multiplier/_0953_ ));
 AOI21_X2 \u_multiplier/_1829_  (.A(\u_multiplier/_0953_ ),
    .B1(\u_multiplier/_0948_ ),
    .B2(\u_multiplier/_0947_ ),
    .ZN(\u_multiplier/_0954_ ));
 NOR2_X1 \u_multiplier/_1830_  (.A1(\u_multiplier/_0949_ ),
    .A2(\u_multiplier/_0954_ ),
    .ZN(\u_multiplier/_0955_ ));
 XOR2_X2 \u_multiplier/_1831_  (.A(\u_multiplier/ky [7]),
    .B(\u_multiplier/LODy/z [7]),
    .Z(\u_multiplier/_0956_ ));
 XNOR2_X2 \u_multiplier/_1832_  (.A(\u_multiplier/ky [7]),
    .B(\u_multiplier/LODy/z [7]),
    .ZN(\u_multiplier/_0957_ ));
 XOR2_X2 \u_multiplier/_1833_  (.A(\u_multiplier/kx [7]),
    .B(\u_multiplier/LODx/z [7]),
    .Z(\u_multiplier/_0958_ ));
 NAND2_X1 \u_multiplier/_1834_  (.A1(\u_multiplier/_0957_ ),
    .A2(\u_multiplier/_0958_ ),
    .ZN(\u_multiplier/_0959_ ));
 XOR2_X2 \u_multiplier/_1835_  (.A(\u_multiplier/ky [6]),
    .B(sram_rdata_reg[6]),
    .Z(\u_multiplier/_0960_ ));
 XOR2_X2 \u_multiplier/_1836_  (.A(\u_multiplier/kx [6]),
    .B(data_in_reg[6]),
    .Z(\u_multiplier/_0961_ ));
 XNOR2_X2 \u_multiplier/_1837_  (.A(\u_multiplier/kx [6]),
    .B(data_in_reg[6]),
    .ZN(\u_multiplier/_0962_ ));
 NAND2_X2 \u_multiplier/_1838_  (.A1(\u_multiplier/_0960_ ),
    .A2(\u_multiplier/_0962_ ),
    .ZN(\u_multiplier/_0963_ ));
 INV_X1 \u_multiplier/_1839_  (.A(\u_multiplier/_0963_ ),
    .ZN(\u_multiplier/_0964_ ));
 XOR2_X2 \u_multiplier/_1840_  (.A(\u_multiplier/kx [0]),
    .B(data_in_reg[0]),
    .Z(\u_multiplier/_0965_ ));
 XNOR2_X2 \u_multiplier/_1841_  (.A(\u_multiplier/kx [0]),
    .B(data_in_reg[0]),
    .ZN(\u_multiplier/_0966_ ));
 XOR2_X2 \u_multiplier/_1842_  (.A(\u_multiplier/ky [1]),
    .B(sram_rdata_reg[1]),
    .Z(\u_multiplier/_0967_ ));
 XNOR2_X2 \u_multiplier/_1843_  (.A(\u_multiplier/ky [1]),
    .B(sram_rdata_reg[1]),
    .ZN(\u_multiplier/_0968_ ));
 XOR2_X2 \u_multiplier/_1844_  (.A(\u_multiplier/kx [1]),
    .B(data_in_reg[1]),
    .Z(\u_multiplier/_0969_ ));
 XNOR2_X2 \u_multiplier/_1845_  (.A(\u_multiplier/kx [1]),
    .B(data_in_reg[1]),
    .ZN(\u_multiplier/_0970_ ));
 AOI211_X1 \u_multiplier/_1846_  (.A(\u_multiplier/_0945_ ),
    .B(\u_multiplier/_0965_ ),
    .C1(\u_multiplier/_0968_ ),
    .C2(\u_multiplier/_0969_ ),
    .ZN(\u_multiplier/_0971_ ));
 OAI211_X1 \u_multiplier/_1847_  (.A(\u_multiplier/_0944_ ),
    .B(\u_multiplier/_0966_ ),
    .C1(\u_multiplier/_0967_ ),
    .C2(\u_multiplier/_0970_ ),
    .ZN(\u_multiplier/_0972_ ));
 XOR2_X2 \u_multiplier/_1848_  (.A(\u_multiplier/ky [2]),
    .B(sram_rdata_reg[2]),
    .Z(\u_multiplier/_0973_ ));
 XNOR2_X2 \u_multiplier/_1849_  (.A(\u_multiplier/ky [2]),
    .B(sram_rdata_reg[2]),
    .ZN(\u_multiplier/_0974_ ));
 XOR2_X2 \u_multiplier/_1850_  (.A(\u_multiplier/kx [2]),
    .B(data_in_reg[2]),
    .Z(\u_multiplier/_0975_ ));
 XNOR2_X2 \u_multiplier/_1851_  (.A(\u_multiplier/kx [2]),
    .B(data_in_reg[2]),
    .ZN(\u_multiplier/_0976_ ));
 AOI22_X4 \u_multiplier/_1852_  (.A1(\u_multiplier/_0967_ ),
    .A2(\u_multiplier/_0970_ ),
    .B1(\u_multiplier/_0973_ ),
    .B2(\u_multiplier/_0976_ ),
    .ZN(\u_multiplier/_0977_ ));
 OAI22_X1 \u_multiplier/_1853_  (.A1(\u_multiplier/_0968_ ),
    .A2(\u_multiplier/_0969_ ),
    .B1(\u_multiplier/_0974_ ),
    .B2(\u_multiplier/_0975_ ),
    .ZN(\u_multiplier/_0978_ ));
 XOR2_X2 \u_multiplier/_1854_  (.A(\u_multiplier/ky [3]),
    .B(\u_multiplier/LODy/z [3]),
    .Z(\u_multiplier/_0979_ ));
 XNOR2_X2 \u_multiplier/_1855_  (.A(\u_multiplier/ky [3]),
    .B(\u_multiplier/LODy/z [3]),
    .ZN(\u_multiplier/_0980_ ));
 XOR2_X2 \u_multiplier/_1856_  (.A(\u_multiplier/kx [3]),
    .B(\u_multiplier/LODx/z [3]),
    .Z(\u_multiplier/_0981_ ));
 XNOR2_X1 \u_multiplier/_1857_  (.A(\u_multiplier/kx [3]),
    .B(\u_multiplier/LODx/z [3]),
    .ZN(\u_multiplier/_0982_ ));
 AOI22_X2 \u_multiplier/_1858_  (.A1(\u_multiplier/_0974_ ),
    .A2(\u_multiplier/_0975_ ),
    .B1(\u_multiplier/_0980_ ),
    .B2(\u_multiplier/_0981_ ),
    .ZN(\u_multiplier/_0983_ ));
 AOI222_X2 \u_multiplier/_1859_  (.A1(\u_multiplier/_0974_ ),
    .A2(\u_multiplier/_0975_ ),
    .B1(\u_multiplier/_0980_ ),
    .B2(\u_multiplier/_0981_ ),
    .C1(\u_multiplier/_0977_ ),
    .C2(\u_multiplier/_0972_ ),
    .ZN(\u_multiplier/_0984_ ));
 OAI21_X1 \u_multiplier/_1860_  (.A(\u_multiplier/_0983_ ),
    .B1(\u_multiplier/_0978_ ),
    .B2(\u_multiplier/_0971_ ),
    .ZN(\u_multiplier/_0985_ ));
 NOR2_X1 \u_multiplier/_1861_  (.A1(\u_multiplier/_0980_ ),
    .A2(\u_multiplier/_0981_ ),
    .ZN(\u_multiplier/_0986_ ));
 NAND2_X1 \u_multiplier/_1862_  (.A1(\u_multiplier/_0979_ ),
    .A2(\u_multiplier/_0982_ ),
    .ZN(\u_multiplier/_0987_ ));
 XOR2_X2 \u_multiplier/_1863_  (.A(\u_multiplier/ky [4]),
    .B(sram_rdata_reg[4]),
    .Z(\u_multiplier/_0988_ ));
 XNOR2_X1 \u_multiplier/_1864_  (.A(\u_multiplier/ky [4]),
    .B(sram_rdata_reg[4]),
    .ZN(\u_multiplier/_0989_ ));
 XOR2_X2 \u_multiplier/_1865_  (.A(\u_multiplier/kx [4]),
    .B(data_in_reg[4]),
    .Z(\u_multiplier/_0990_ ));
 XOR2_X2 \u_multiplier/_1866_  (.A(\u_multiplier/ky [5]),
    .B(sram_rdata_reg[5]),
    .Z(\u_multiplier/_0991_ ));
 XNOR2_X2 \u_multiplier/_1867_  (.A(\u_multiplier/ky [5]),
    .B(sram_rdata_reg[5]),
    .ZN(\u_multiplier/_0992_ ));
 XOR2_X2 \u_multiplier/_1868_  (.A(\u_multiplier/kx [5]),
    .B(data_in_reg[5]),
    .Z(\u_multiplier/_0993_ ));
 XNOR2_X1 \u_multiplier/_1869_  (.A(\u_multiplier/kx [5]),
    .B(data_in_reg[5]),
    .ZN(\u_multiplier/_0994_ ));
 XNOR2_X2 \u_multiplier/_1870_  (.A(\u_multiplier/_0991_ ),
    .B(\u_multiplier/_0993_ ),
    .ZN(\u_multiplier/_0995_ ));
 XNOR2_X2 \u_multiplier/_1871_  (.A(\u_multiplier/_0988_ ),
    .B(\u_multiplier/_0990_ ),
    .ZN(\u_multiplier/_0996_ ));
 AND3_X1 \u_multiplier/_1872_  (.A1(\u_multiplier/_0987_ ),
    .A2(\u_multiplier/_0995_ ),
    .A3(\u_multiplier/_0996_ ),
    .ZN(\u_multiplier/_0997_ ));
 NAND3_X1 \u_multiplier/_1873_  (.A1(\u_multiplier/_0987_ ),
    .A2(\u_multiplier/_0995_ ),
    .A3(\u_multiplier/_0996_ ),
    .ZN(\u_multiplier/_0998_ ));
 OAI211_X2 \u_multiplier/_1874_  (.A(\u_multiplier/_0989_ ),
    .B(\u_multiplier/_0990_ ),
    .C1(\u_multiplier/_0992_ ),
    .C2(\u_multiplier/_0993_ ),
    .ZN(\u_multiplier/_0999_ ));
 NOR2_X2 \u_multiplier/_1875_  (.A1(\u_multiplier/_0960_ ),
    .A2(\u_multiplier/_0962_ ),
    .ZN(\u_multiplier/_1000_ ));
 AOI21_X1 \u_multiplier/_1876_  (.A(\u_multiplier/_1000_ ),
    .B1(\u_multiplier/_0993_ ),
    .B2(\u_multiplier/_0992_ ),
    .ZN(\u_multiplier/_1001_ ));
 OAI21_X1 \u_multiplier/_1877_  (.A(\u_multiplier/_0999_ ),
    .B1(\u_multiplier/_0994_ ),
    .B2(\u_multiplier/_0991_ ),
    .ZN(\u_multiplier/_1002_ ));
 AOI211_X1 \u_multiplier/_1878_  (.A(\u_multiplier/_1000_ ),
    .B(\u_multiplier/_1002_ ),
    .C1(\u_multiplier/_0985_ ),
    .C2(\u_multiplier/_0997_ ),
    .ZN(\u_multiplier/_1003_ ));
 OAI211_X1 \u_multiplier/_1879_  (.A(\u_multiplier/_0999_ ),
    .B(\u_multiplier/_1001_ ),
    .C1(\u_multiplier/_0984_ ),
    .C2(\u_multiplier/_0998_ ),
    .ZN(\u_multiplier/_1004_ ));
 AOI22_X2 \u_multiplier/_1880_  (.A1(\u_multiplier/_0957_ ),
    .A2(\u_multiplier/_0958_ ),
    .B1(\u_multiplier/_0963_ ),
    .B2(\u_multiplier/_1004_ ),
    .ZN(\u_multiplier/_1005_ ));
 OAI21_X1 \u_multiplier/_1881_  (.A(\u_multiplier/_0959_ ),
    .B1(\u_multiplier/_0964_ ),
    .B2(\u_multiplier/_1003_ ),
    .ZN(\u_multiplier/_1006_ ));
 NOR2_X1 \u_multiplier/_1882_  (.A1(\u_multiplier/_0957_ ),
    .A2(\u_multiplier/_0958_ ),
    .ZN(\u_multiplier/_1007_ ));
 OAI22_X2 \u_multiplier/_1883_  (.A1(\u_multiplier/_0947_ ),
    .A2(\u_multiplier/_0948_ ),
    .B1(\u_multiplier/_0951_ ),
    .B2(\u_multiplier/_0952_ ),
    .ZN(\u_multiplier/_1008_ ));
 AOI211_X2 \u_multiplier/_1884_  (.A(\u_multiplier/_0953_ ),
    .B(\u_multiplier/_1008_ ),
    .C1(\u_multiplier/_0947_ ),
    .C2(\u_multiplier/_0948_ ),
    .ZN(\u_multiplier/_1009_ ));
 INV_X1 \u_multiplier/_1885_  (.A(\u_multiplier/_1009_ ),
    .ZN(\u_multiplier/_1010_ ));
 NOR2_X1 \u_multiplier/_1886_  (.A1(\u_multiplier/_1007_ ),
    .A2(\u_multiplier/_1010_ ),
    .ZN(\u_multiplier/_1011_ ));
 OAI21_X1 \u_multiplier/_1887_  (.A(\u_multiplier/_1009_ ),
    .B1(\u_multiplier/_0958_ ),
    .B2(\u_multiplier/_0957_ ),
    .ZN(\u_multiplier/_1012_ ));
 AOI21_X1 \u_multiplier/_1888_  (.A(\u_multiplier/_0955_ ),
    .B1(\u_multiplier/_1006_ ),
    .B2(\u_multiplier/_1011_ ),
    .ZN(\u_multiplier/_1013_ ));
 OAI22_X2 \u_multiplier/_1889_  (.A1(\u_multiplier/_0949_ ),
    .A2(\u_multiplier/_0954_ ),
    .B1(\u_multiplier/_1005_ ),
    .B2(\u_multiplier/_1012_ ),
    .ZN(\u_multiplier/_1014_ ));
 XOR2_X2 \u_multiplier/_1890_  (.A(\u_multiplier/ky [13]),
    .B(sram_rdata_reg[13]),
    .Z(\u_multiplier/_1015_ ));
 XOR2_X2 \u_multiplier/_1891_  (.A(\u_multiplier/kx [13]),
    .B(data_in_reg[13]),
    .Z(\u_multiplier/_1016_ ));
 INV_X1 \u_multiplier/_1892_  (.A(\u_multiplier/_1016_ ),
    .ZN(\u_multiplier/_1017_ ));
 NOR2_X1 \u_multiplier/_1893_  (.A1(\u_multiplier/_1015_ ),
    .A2(\u_multiplier/_1017_ ),
    .ZN(\u_multiplier/_1018_ ));
 XOR2_X2 \u_multiplier/_1894_  (.A(\u_multiplier/ky [12]),
    .B(sram_rdata_reg[12]),
    .Z(\u_multiplier/_1019_ ));
 INV_X1 \u_multiplier/_1895_  (.A(\u_multiplier/_1019_ ),
    .ZN(\u_multiplier/_1020_ ));
 XOR2_X2 \u_multiplier/_1896_  (.A(\u_multiplier/kx [12]),
    .B(data_in_reg[12]),
    .Z(\u_multiplier/_1021_ ));
 AND2_X1 \u_multiplier/_1897_  (.A1(\u_multiplier/_1015_ ),
    .A2(\u_multiplier/_1017_ ),
    .ZN(\u_multiplier/_1022_ ));
 XOR2_X1 \u_multiplier/_1898_  (.A(\u_multiplier/_1019_ ),
    .B(\u_multiplier/_1021_ ),
    .Z(\u_multiplier/_1023_ ));
 OR3_X1 \u_multiplier/_1899_  (.A1(\u_multiplier/_1018_ ),
    .A2(\u_multiplier/_1022_ ),
    .A3(\u_multiplier/_1023_ ),
    .ZN(\u_multiplier/_1024_ ));
 XOR2_X2 \u_multiplier/_1900_  (.A(\u_multiplier/ky [11]),
    .B(\u_multiplier/LODy/z [11]),
    .Z(\u_multiplier/_1025_ ));
 XNOR2_X1 \u_multiplier/_1901_  (.A(\u_multiplier/ky [11]),
    .B(\u_multiplier/LODy/z [11]),
    .ZN(\u_multiplier/_1026_ ));
 XOR2_X2 \u_multiplier/_1902_  (.A(\u_multiplier/kx [11]),
    .B(\u_multiplier/LODx/z [11]),
    .Z(\u_multiplier/_1027_ ));
 NAND2_X1 \u_multiplier/_1903_  (.A1(\u_multiplier/_1026_ ),
    .A2(\u_multiplier/_1027_ ),
    .ZN(\u_multiplier/_1028_ ));
 XOR2_X2 \u_multiplier/_1904_  (.A(\u_multiplier/ky [10]),
    .B(sram_rdata_reg[10]),
    .Z(\u_multiplier/_1029_ ));
 INV_X1 \u_multiplier/_1905_  (.A(\u_multiplier/_1029_ ),
    .ZN(\u_multiplier/_1030_ ));
 XOR2_X2 \u_multiplier/_1906_  (.A(\u_multiplier/kx [10]),
    .B(data_in_reg[10]),
    .Z(\u_multiplier/_1031_ ));
 OR2_X1 \u_multiplier/_1907_  (.A1(\u_multiplier/_1026_ ),
    .A2(\u_multiplier/_1027_ ),
    .ZN(\u_multiplier/_1032_ ));
 XNOR2_X1 \u_multiplier/_1908_  (.A(\u_multiplier/_1029_ ),
    .B(\u_multiplier/_1031_ ),
    .ZN(\u_multiplier/_1033_ ));
 NAND3_X1 \u_multiplier/_1909_  (.A1(\u_multiplier/_1028_ ),
    .A2(\u_multiplier/_1032_ ),
    .A3(\u_multiplier/_1033_ ),
    .ZN(\u_multiplier/_1034_ ));
 OR2_X2 \u_multiplier/_1910_  (.A1(\u_multiplier/_1024_ ),
    .A2(\u_multiplier/_1034_ ),
    .ZN(\u_multiplier/_1035_ ));
 INV_X1 \u_multiplier/_1911_  (.A(\u_multiplier/_1035_ ),
    .ZN(\u_multiplier/_1036_ ));
 NAND3_X1 \u_multiplier/_1912_  (.A1(\u_multiplier/_1030_ ),
    .A2(\u_multiplier/_1031_ ),
    .A3(\u_multiplier/_1032_ ),
    .ZN(\u_multiplier/_1037_ ));
 AOI21_X2 \u_multiplier/_1913_  (.A(\u_multiplier/_1024_ ),
    .B1(\u_multiplier/_1028_ ),
    .B2(\u_multiplier/_1037_ ),
    .ZN(\u_multiplier/_1038_ ));
 XOR2_X2 \u_multiplier/_1914_  (.A(\u_multiplier/ky [14]),
    .B(sram_rdata_reg[14]),
    .Z(\u_multiplier/_1039_ ));
 XNOR2_X2 \u_multiplier/_1915_  (.A(\u_multiplier/ky [14]),
    .B(sram_rdata_reg[14]),
    .ZN(\u_multiplier/_1040_ ));
 XOR2_X2 \u_multiplier/_1916_  (.A(\u_multiplier/kx [14]),
    .B(data_in_reg[14]),
    .Z(\u_multiplier/_1041_ ));
 XNOR2_X2 \u_multiplier/_1917_  (.A(\u_multiplier/kx [14]),
    .B(data_in_reg[14]),
    .ZN(\u_multiplier/_1042_ ));
 NOR2_X1 \u_multiplier/_1918_  (.A1(\u_multiplier/_1039_ ),
    .A2(\u_multiplier/_1042_ ),
    .ZN(\u_multiplier/_1043_ ));
 AOI21_X1 \u_multiplier/_1919_  (.A(\u_multiplier/_1018_ ),
    .B1(\u_multiplier/_1020_ ),
    .B2(\u_multiplier/_1021_ ),
    .ZN(\u_multiplier/_1044_ ));
 OAI22_X2 \u_multiplier/_1920_  (.A1(\u_multiplier/_1039_ ),
    .A2(\u_multiplier/_1042_ ),
    .B1(\u_multiplier/_1044_ ),
    .B2(\u_multiplier/_1022_ ),
    .ZN(\u_multiplier/_1045_ ));
 NOR2_X1 \u_multiplier/_1921_  (.A1(\u_multiplier/_1038_ ),
    .A2(\u_multiplier/_1045_ ),
    .ZN(\u_multiplier/_1046_ ));
 AOI211_X2 \u_multiplier/_1922_  (.A(\u_multiplier/_1038_ ),
    .B(\u_multiplier/_1045_ ),
    .C1(\u_multiplier/_1014_ ),
    .C2(\u_multiplier/_1036_ ),
    .ZN(\u_multiplier/_1047_ ));
 OAI21_X2 \u_multiplier/_1923_  (.A(\u_multiplier/_1046_ ),
    .B1(\u_multiplier/_1035_ ),
    .B2(\u_multiplier/_1013_ ),
    .ZN(\u_multiplier/_1048_ ));
 NOR2_X2 \u_multiplier/_1924_  (.A1(\u_multiplier/_1040_ ),
    .A2(\u_multiplier/_1041_ ),
    .ZN(\u_multiplier/_1049_ ));
 NOR2_X1 \u_multiplier/_1925_  (.A1(\u_multiplier/_0944_ ),
    .A2(\u_multiplier/_0966_ ),
    .ZN(\u_multiplier/_1050_ ));
 OR4_X1 \u_multiplier/_1926_  (.A1(\u_multiplier/_1007_ ),
    .A2(\u_multiplier/_1043_ ),
    .A3(\u_multiplier/_1049_ ),
    .A4(\u_multiplier/_1050_ ),
    .ZN(\u_multiplier/_1051_ ));
 OAI22_X2 \u_multiplier/_1927_  (.A1(\u_multiplier/_0945_ ),
    .A2(\u_multiplier/_0965_ ),
    .B1(\u_multiplier/_0967_ ),
    .B2(\u_multiplier/_0970_ ),
    .ZN(\u_multiplier/_1052_ ));
 NOR4_X2 \u_multiplier/_1928_  (.A1(\u_multiplier/_0986_ ),
    .A2(\u_multiplier/_1000_ ),
    .A3(\u_multiplier/_1051_ ),
    .A4(\u_multiplier/_1052_ ),
    .ZN(\u_multiplier/_1053_ ));
 NAND4_X2 \u_multiplier/_1929_  (.A1(\u_multiplier/_0995_ ),
    .A2(\u_multiplier/_0996_ ),
    .A3(\u_multiplier/_1009_ ),
    .A4(\u_multiplier/_1053_ ),
    .ZN(\u_multiplier/_1054_ ));
 NAND4_X2 \u_multiplier/_1930_  (.A1(\u_multiplier/_0959_ ),
    .A2(\u_multiplier/_0963_ ),
    .A3(\u_multiplier/_0977_ ),
    .A4(\u_multiplier/_0983_ ),
    .ZN(\u_multiplier/_1055_ ));
 NOR3_X4 \u_multiplier/_1931_  (.A1(\u_multiplier/_1035_ ),
    .A2(\u_multiplier/_1054_ ),
    .A3(\u_multiplier/_1055_ ),
    .ZN(\u_multiplier/_1056_ ));
 NOR2_X2 \u_multiplier/_1932_  (.A1(\u_multiplier/_1049_ ),
    .A2(\u_multiplier/_1056_ ),
    .ZN(\u_multiplier/_1057_ ));
 OR2_X2 \u_multiplier/_1933_  (.A1(\u_multiplier/_1049_ ),
    .A2(\u_multiplier/_1056_ ),
    .ZN(\u_multiplier/_1058_ ));
 NAND2_X4 \u_multiplier/_1934_  (.A1(\u_multiplier/_1048_ ),
    .A2(\u_multiplier/_1057_ ),
    .ZN(\u_multiplier/_1059_ ));
 NOR3_X4 \u_multiplier/_1935_  (.A1(\u_multiplier/_0945_ ),
    .A2(\u_multiplier/_1047_ ),
    .A3(\u_multiplier/_1058_ ),
    .ZN(\u_multiplier/_1060_ ));
 AOI21_X4 \u_multiplier/_1936_  (.A(\u_multiplier/_1060_ ),
    .B1(\u_multiplier/_1059_ ),
    .B2(\u_multiplier/_0965_ ),
    .ZN(\u_multiplier/_1061_ ));
 NOR3_X1 \u_multiplier/_1937_  (.A1(\u_multiplier/K [1]),
    .A2(\u_multiplier/K [0]),
    .A3(\u_multiplier/_1061_ ),
    .ZN(\u_multiplier/_1062_ ));
 NOR4_X4 \u_multiplier/_1938_  (.A1(\u_multiplier/K [1]),
    .A2(\u_multiplier/K [0]),
    .A3(\u_multiplier/K [2]),
    .A4(\u_multiplier/_1061_ ),
    .ZN(\u_multiplier/_1063_ ));
 AOI21_X2 \u_multiplier/_1939_  (.A(\u_multiplier/dec_out [0]),
    .B1(\u_multiplier/_1063_ ),
    .B2(\u_multiplier/_0939_ ),
    .ZN(\u_multiplier/_1064_ ));
 NOR2_X1 \u_multiplier/_1940_  (.A1(\u_multiplier/code_x [0]),
    .A2(\u_multiplier/_0945_ ),
    .ZN(\u_multiplier/_1065_ ));
 NOR4_X4 \u_multiplier/_1941_  (.A1(\u_multiplier/code_x [0]),
    .A2(\u_multiplier/code_x [1]),
    .A3(\u_multiplier/code_x [2]),
    .A4(\u_multiplier/_0945_ ),
    .ZN(\u_multiplier/_1066_ ));
 NAND2_X1 \u_multiplier/_1942_  (.A1(\u_multiplier/_0933_ ),
    .A2(\u_multiplier/_1066_ ),
    .ZN(\u_multiplier/_1067_ ));
 NOR3_X2 \u_multiplier/_1943_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/code_y [0]),
    .A3(\u_multiplier/_0966_ ),
    .ZN(\u_multiplier/_1068_ ));
 NAND2_X1 \u_multiplier/_1944_  (.A1(\u_multiplier/_0931_ ),
    .A2(\u_multiplier/_1068_ ),
    .ZN(\u_multiplier/_1069_ ));
 NOR2_X1 \u_multiplier/_1945_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_1069_ ),
    .ZN(\u_multiplier/_1070_ ));
 NAND3_X1 \u_multiplier/_1946_  (.A1(\u_multiplier/_0933_ ),
    .A2(\u_multiplier/_1066_ ),
    .A3(\u_multiplier/_1070_ ),
    .ZN(\u_multiplier/_1071_ ));
 XOR2_X2 \u_multiplier/_1947_  (.A(\u_multiplier/_1067_ ),
    .B(\u_multiplier/_1070_ ),
    .Z(\u_multiplier/_1072_ ));
 OAI21_X1 \u_multiplier/_1948_  (.A(\u_multiplier/_1739_ ),
    .B1(\u_multiplier/_1064_ ),
    .B2(\u_multiplier/_1072_ ),
    .ZN(\u_multiplier/_1073_ ));
 AOI21_X1 \u_multiplier/_1949_  (.A(\u_multiplier/_1073_ ),
    .B1(\u_multiplier/_1072_ ),
    .B2(\u_multiplier/_1064_ ),
    .ZN(product[0]));
 OAI21_X2 \u_multiplier/_1950_  (.A(\u_multiplier/_1071_ ),
    .B1(\u_multiplier/_1072_ ),
    .B2(\u_multiplier/_1064_ ),
    .ZN(\u_multiplier/_1074_ ));
 AOI21_X2 \u_multiplier/_1951_  (.A(\u_multiplier/_0970_ ),
    .B1(\u_multiplier/_1048_ ),
    .B2(\u_multiplier/_1057_ ),
    .ZN(\u_multiplier/_1075_ ));
 NOR3_X2 \u_multiplier/_1952_  (.A1(\u_multiplier/_0968_ ),
    .A2(\u_multiplier/_1047_ ),
    .A3(\u_multiplier/_1058_ ),
    .ZN(\u_multiplier/_1076_ ));
 NOR3_X2 \u_multiplier/_1953_  (.A1(\u_multiplier/K [0]),
    .A2(\u_multiplier/_1075_ ),
    .A3(\u_multiplier/_1076_ ),
    .ZN(\u_multiplier/_1077_ ));
 AOI211_X2 \u_multiplier/_1954_  (.A(\u_multiplier/_0937_ ),
    .B(\u_multiplier/_1060_ ),
    .C1(\u_multiplier/_1059_ ),
    .C2(\u_multiplier/_0965_ ),
    .ZN(\u_multiplier/_1078_ ));
 OR2_X1 \u_multiplier/_1955_  (.A1(\u_multiplier/_1077_ ),
    .A2(\u_multiplier/_1078_ ),
    .ZN(\u_multiplier/_1079_ ));
 NOR2_X1 \u_multiplier/_1956_  (.A1(\u_multiplier/K [1]),
    .A2(\u_multiplier/_1079_ ),
    .ZN(\u_multiplier/_1080_ ));
 NOR4_X4 \u_multiplier/_1957_  (.A1(\u_multiplier/K [1]),
    .A2(\u_multiplier/K [2]),
    .A3(\u_multiplier/_1077_ ),
    .A4(\u_multiplier/_1078_ ),
    .ZN(\u_multiplier/_1081_ ));
 AND2_X1 \u_multiplier/_1958_  (.A1(\u_multiplier/_0939_ ),
    .A2(\u_multiplier/_1081_ ),
    .ZN(\u_multiplier/_1082_ ));
 AOI21_X1 \u_multiplier/_1959_  (.A(\u_multiplier/dec_out [1]),
    .B1(\u_multiplier/_1081_ ),
    .B2(\u_multiplier/_0939_ ),
    .ZN(\u_multiplier/_1083_ ));
 MUX2_X1 \u_multiplier/_1960_  (.A(\u_multiplier/_0945_ ),
    .B(\u_multiplier/_0968_ ),
    .S(\u_multiplier/_0934_ ),
    .Z(\u_multiplier/_1084_ ));
 OR2_X1 \u_multiplier/_1961_  (.A1(\u_multiplier/code_x [1]),
    .A2(\u_multiplier/_1084_ ),
    .ZN(\u_multiplier/_1085_ ));
 OR2_X1 \u_multiplier/_1962_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_1085_ ),
    .ZN(\u_multiplier/_1086_ ));
 MUX2_X1 \u_multiplier/_1963_  (.A(\u_multiplier/_0966_ ),
    .B(\u_multiplier/_0970_ ),
    .S(\u_multiplier/_0930_ ),
    .Z(\u_multiplier/_1087_ ));
 OR2_X1 \u_multiplier/_1964_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_1087_ ),
    .ZN(\u_multiplier/_1088_ ));
 OR2_X1 \u_multiplier/_1965_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_1088_ ),
    .ZN(\u_multiplier/_1089_ ));
 OAI22_X1 \u_multiplier/_1966_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_1086_ ),
    .B1(\u_multiplier/_1089_ ),
    .B2(\u_multiplier/code_y [3]),
    .ZN(\u_multiplier/_1090_ ));
 OR4_X2 \u_multiplier/_1967_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/code_x [3]),
    .A3(\u_multiplier/_1086_ ),
    .A4(\u_multiplier/_1089_ ),
    .ZN(\u_multiplier/_1091_ ));
 AND2_X1 \u_multiplier/_1968_  (.A1(\u_multiplier/_1090_ ),
    .A2(\u_multiplier/_1091_ ),
    .ZN(\u_multiplier/_1092_ ));
 OAI21_X2 \u_multiplier/_1969_  (.A(\u_multiplier/_1092_ ),
    .B1(\u_multiplier/_1082_ ),
    .B2(\u_multiplier/dec_out [1]),
    .ZN(\u_multiplier/_1093_ ));
 XNOR2_X1 \u_multiplier/_1970_  (.A(\u_multiplier/_1083_ ),
    .B(\u_multiplier/_1092_ ),
    .ZN(\u_multiplier/_1094_ ));
 AND2_X1 \u_multiplier/_1971_  (.A1(\u_multiplier/_1074_ ),
    .A2(\u_multiplier/_1094_ ),
    .ZN(\u_multiplier/_1095_ ));
 NAND2_X1 \u_multiplier/_1972_  (.A1(\u_multiplier/_1074_ ),
    .A2(\u_multiplier/_1094_ ),
    .ZN(\u_multiplier/_1096_ ));
 OAI21_X1 \u_multiplier/_1973_  (.A(\u_multiplier/_1739_ ),
    .B1(\u_multiplier/_1074_ ),
    .B2(\u_multiplier/_1094_ ),
    .ZN(\u_multiplier/_1097_ ));
 NOR2_X1 \u_multiplier/_1974_  (.A1(\u_multiplier/_1095_ ),
    .A2(\u_multiplier/_1097_ ),
    .ZN(product[1]));
 NAND2_X1 \u_multiplier/_1975_  (.A1(\u_multiplier/_1091_ ),
    .A2(\u_multiplier/_1093_ ),
    .ZN(\u_multiplier/_1098_ ));
 NOR3_X1 \u_multiplier/_1976_  (.A1(\u_multiplier/_0974_ ),
    .A2(\u_multiplier/_1047_ ),
    .A3(\u_multiplier/_1058_ ),
    .ZN(\u_multiplier/_1099_ ));
 AOI21_X1 \u_multiplier/_1977_  (.A(\u_multiplier/_0975_ ),
    .B1(\u_multiplier/_1048_ ),
    .B2(\u_multiplier/_1057_ ),
    .ZN(\u_multiplier/_1100_ ));
 NOR3_X1 \u_multiplier/_1978_  (.A1(\u_multiplier/_0973_ ),
    .A2(\u_multiplier/_1047_ ),
    .A3(\u_multiplier/_1058_ ),
    .ZN(\u_multiplier/_1101_ ));
 NOR2_X1 \u_multiplier/_1979_  (.A1(\u_multiplier/_1100_ ),
    .A2(\u_multiplier/_1101_ ),
    .ZN(\u_multiplier/_1102_ ));
 NOR3_X2 \u_multiplier/_1980_  (.A1(\u_multiplier/_0937_ ),
    .A2(\u_multiplier/_1075_ ),
    .A3(\u_multiplier/_1076_ ),
    .ZN(\u_multiplier/_1103_ ));
 AOI211_X2 \u_multiplier/_1981_  (.A(\u_multiplier/K [0]),
    .B(\u_multiplier/_1099_ ),
    .C1(\u_multiplier/_1059_ ),
    .C2(\u_multiplier/_0975_ ),
    .ZN(\u_multiplier/_1104_ ));
 OAI21_X1 \u_multiplier/_1982_  (.A(\u_multiplier/K [1]),
    .B1(\u_multiplier/K [0]),
    .B2(\u_multiplier/_1061_ ),
    .ZN(\u_multiplier/_1105_ ));
 OAI21_X2 \u_multiplier/_1983_  (.A(\u_multiplier/_0936_ ),
    .B1(\u_multiplier/_1103_ ),
    .B2(\u_multiplier/_1104_ ),
    .ZN(\u_multiplier/_1106_ ));
 NAND2_X1 \u_multiplier/_1984_  (.A1(\u_multiplier/_1105_ ),
    .A2(\u_multiplier/_1106_ ),
    .ZN(\u_multiplier/_1107_ ));
 NAND4_X2 \u_multiplier/_1985_  (.A1(\u_multiplier/_0938_ ),
    .A2(\u_multiplier/_0939_ ),
    .A3(\u_multiplier/_1105_ ),
    .A4(\u_multiplier/_1106_ ),
    .ZN(\u_multiplier/_1108_ ));
 MUX2_X1 \u_multiplier/_1986_  (.A(\u_multiplier/_0967_ ),
    .B(\u_multiplier/_0973_ ),
    .S(\u_multiplier/_0934_ ),
    .Z(\u_multiplier/_1109_ ));
 MUX2_X1 \u_multiplier/_1987_  (.A(\u_multiplier/_1109_ ),
    .B(\u_multiplier/_1065_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_1110_ ));
 NAND2_X1 \u_multiplier/_1988_  (.A1(\u_multiplier/_0935_ ),
    .A2(\u_multiplier/_1110_ ),
    .ZN(\u_multiplier/_1111_ ));
 NOR2_X1 \u_multiplier/_1989_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_1111_ ),
    .ZN(\u_multiplier/_1112_ ));
 MUX2_X1 \u_multiplier/_1990_  (.A(\u_multiplier/_0969_ ),
    .B(\u_multiplier/_0975_ ),
    .S(\u_multiplier/_0930_ ),
    .Z(\u_multiplier/_1113_ ));
 INV_X1 \u_multiplier/_1991_  (.A(\u_multiplier/_1113_ ),
    .ZN(\u_multiplier/_1114_ ));
 NAND3_X1 \u_multiplier/_1992_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_0930_ ),
    .A3(\u_multiplier/_0965_ ),
    .ZN(\u_multiplier/_1115_ ));
 OAI21_X2 \u_multiplier/_1993_  (.A(\u_multiplier/_1115_ ),
    .B1(\u_multiplier/_1114_ ),
    .B2(\u_multiplier/code_y [1]),
    .ZN(\u_multiplier/_1116_ ));
 NAND2_X1 \u_multiplier/_1994_  (.A1(\u_multiplier/_0931_ ),
    .A2(\u_multiplier/_1116_ ),
    .ZN(\u_multiplier/_1117_ ));
 NOR2_X1 \u_multiplier/_1995_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_1117_ ),
    .ZN(\u_multiplier/_1118_ ));
 AND2_X1 \u_multiplier/_1996_  (.A1(\u_multiplier/_1112_ ),
    .A2(\u_multiplier/_1118_ ),
    .ZN(\u_multiplier/_1119_ ));
 XNOR2_X2 \u_multiplier/_1997_  (.A(\u_multiplier/_1112_ ),
    .B(\u_multiplier/_1118_ ),
    .ZN(\u_multiplier/_1120_ ));
 AND3_X1 \u_multiplier/_1998_  (.A1(\u_multiplier/_0940_ ),
    .A2(\u_multiplier/_1108_ ),
    .A3(\u_multiplier/_1120_ ),
    .ZN(\u_multiplier/_1121_ ));
 AOI21_X4 \u_multiplier/_1999_  (.A(\u_multiplier/_1120_ ),
    .B1(\u_multiplier/_1108_ ),
    .B2(\u_multiplier/_0940_ ),
    .ZN(\u_multiplier/_1122_ ));
 OR2_X1 \u_multiplier/_2000_  (.A1(\u_multiplier/_1121_ ),
    .A2(\u_multiplier/_1122_ ),
    .ZN(\u_multiplier/_1123_ ));
 AOI211_X2 \u_multiplier/_2001_  (.A(\u_multiplier/_1121_ ),
    .B(\u_multiplier/_1122_ ),
    .C1(\u_multiplier/_1091_ ),
    .C2(\u_multiplier/_1093_ ),
    .ZN(\u_multiplier/_1124_ ));
 OAI211_X1 \u_multiplier/_2002_  (.A(\u_multiplier/_1091_ ),
    .B(\u_multiplier/_1093_ ),
    .C1(\u_multiplier/_1121_ ),
    .C2(\u_multiplier/_1122_ ),
    .ZN(\u_multiplier/_1125_ ));
 XOR2_X2 \u_multiplier/_2003_  (.A(\u_multiplier/_1098_ ),
    .B(\u_multiplier/_1123_ ),
    .Z(\u_multiplier/_1126_ ));
 OAI21_X1 \u_multiplier/_2004_  (.A(\u_multiplier/_1739_ ),
    .B1(\u_multiplier/_1096_ ),
    .B2(\u_multiplier/_1126_ ),
    .ZN(\u_multiplier/_1127_ ));
 AOI21_X1 \u_multiplier/_2005_  (.A(\u_multiplier/_1127_ ),
    .B1(\u_multiplier/_1126_ ),
    .B2(\u_multiplier/_1096_ ),
    .ZN(product[2]));
 AOI21_X2 \u_multiplier/_2006_  (.A(\u_multiplier/_1124_ ),
    .B1(\u_multiplier/_1125_ ),
    .B2(\u_multiplier/_1095_ ),
    .ZN(\u_multiplier/_1128_ ));
 NOR2_X1 \u_multiplier/_2007_  (.A1(\u_multiplier/_1119_ ),
    .A2(\u_multiplier/_1122_ ),
    .ZN(\u_multiplier/_1129_ ));
 MUX2_X1 \u_multiplier/_2008_  (.A(\u_multiplier/_0979_ ),
    .B(\u_multiplier/_0981_ ),
    .S(\u_multiplier/_1059_ ),
    .Z(\u_multiplier/_1130_ ));
 NOR3_X1 \u_multiplier/_2009_  (.A1(\u_multiplier/_0937_ ),
    .A2(\u_multiplier/_1100_ ),
    .A3(\u_multiplier/_1101_ ),
    .ZN(\u_multiplier/_1131_ ));
 MUX2_X1 \u_multiplier/_2010_  (.A(\u_multiplier/_1102_ ),
    .B(\u_multiplier/_1130_ ),
    .S(\u_multiplier/_0937_ ),
    .Z(\u_multiplier/_1132_ ));
 NOR2_X1 \u_multiplier/_2011_  (.A1(\u_multiplier/_0936_ ),
    .A2(\u_multiplier/_1079_ ),
    .ZN(\u_multiplier/_1133_ ));
 AOI211_X2 \u_multiplier/_2012_  (.A(\u_multiplier/K [1]),
    .B(\u_multiplier/_1131_ ),
    .C1(\u_multiplier/_1130_ ),
    .C2(\u_multiplier/_0937_ ),
    .ZN(\u_multiplier/_1134_ ));
 AOI21_X1 \u_multiplier/_2013_  (.A(\u_multiplier/_1133_ ),
    .B1(\u_multiplier/_1132_ ),
    .B2(\u_multiplier/_0936_ ),
    .ZN(\u_multiplier/_1135_ ));
 AOI211_X2 \u_multiplier/_2014_  (.A(\u_multiplier/K [2]),
    .B(\u_multiplier/_1134_ ),
    .C1(\u_multiplier/_1079_ ),
    .C2(\u_multiplier/K [1]),
    .ZN(\u_multiplier/_1136_ ));
 AOI21_X2 \u_multiplier/_2015_  (.A(\u_multiplier/dec_out [3]),
    .B1(\u_multiplier/_1136_ ),
    .B2(\u_multiplier/_0939_ ),
    .ZN(\u_multiplier/_1137_ ));
 MUX2_X1 \u_multiplier/_2016_  (.A(\u_multiplier/_0974_ ),
    .B(\u_multiplier/_0980_ ),
    .S(\u_multiplier/_0934_ ),
    .Z(\u_multiplier/_1138_ ));
 MUX2_X1 \u_multiplier/_2017_  (.A(\u_multiplier/_1138_ ),
    .B(\u_multiplier/_1084_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_1139_ ));
 OR2_X1 \u_multiplier/_2018_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_1139_ ),
    .ZN(\u_multiplier/_1140_ ));
 MUX2_X1 \u_multiplier/_2019_  (.A(\u_multiplier/_0976_ ),
    .B(\u_multiplier/_0982_ ),
    .S(\u_multiplier/_0930_ ),
    .Z(\u_multiplier/_1141_ ));
 MUX2_X1 \u_multiplier/_2020_  (.A(\u_multiplier/_1141_ ),
    .B(\u_multiplier/_1087_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_1142_ ));
 OR2_X1 \u_multiplier/_2021_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_1142_ ),
    .ZN(\u_multiplier/_1143_ ));
 OAI22_X1 \u_multiplier/_2022_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_1140_ ),
    .B1(\u_multiplier/_1143_ ),
    .B2(\u_multiplier/code_y [3]),
    .ZN(\u_multiplier/_1144_ ));
 OR4_X1 \u_multiplier/_2023_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/code_x [3]),
    .A3(\u_multiplier/_1140_ ),
    .A4(\u_multiplier/_1143_ ),
    .ZN(\u_multiplier/_1145_ ));
 NAND2_X1 \u_multiplier/_2024_  (.A1(\u_multiplier/_1144_ ),
    .A2(\u_multiplier/_1145_ ),
    .ZN(\u_multiplier/_1146_ ));
 XOR2_X2 \u_multiplier/_2025_  (.A(\u_multiplier/_1137_ ),
    .B(\u_multiplier/_1146_ ),
    .Z(\u_multiplier/_1147_ ));
 OAI21_X1 \u_multiplier/_2026_  (.A(\u_multiplier/_1147_ ),
    .B1(\u_multiplier/_1122_ ),
    .B2(\u_multiplier/_1119_ ),
    .ZN(\u_multiplier/_1148_ ));
 XOR2_X2 \u_multiplier/_2027_  (.A(\u_multiplier/_1129_ ),
    .B(\u_multiplier/_1147_ ),
    .Z(\u_multiplier/_1149_ ));
 OR2_X1 \u_multiplier/_2028_  (.A1(\u_multiplier/_1128_ ),
    .A2(\u_multiplier/_1149_ ),
    .ZN(\u_multiplier/_1150_ ));
 AOI21_X1 \u_multiplier/_2029_  (.A(\u_multiplier/_0943_ ),
    .B1(\u_multiplier/_1128_ ),
    .B2(\u_multiplier/_1149_ ),
    .ZN(\u_multiplier/_1151_ ));
 AND2_X1 \u_multiplier/_2030_  (.A1(\u_multiplier/_1150_ ),
    .A2(\u_multiplier/_1151_ ),
    .ZN(product[3]));
 AND2_X1 \u_multiplier/_2031_  (.A1(\u_multiplier/_1148_ ),
    .A2(\u_multiplier/_1150_ ),
    .ZN(\u_multiplier/_1152_ ));
 OAI21_X1 \u_multiplier/_2032_  (.A(\u_multiplier/_1148_ ),
    .B1(\u_multiplier/_1149_ ),
    .B2(\u_multiplier/_1128_ ),
    .ZN(\u_multiplier/_1153_ ));
 OAI21_X1 \u_multiplier/_2033_  (.A(\u_multiplier/_1145_ ),
    .B1(\u_multiplier/_1146_ ),
    .B2(\u_multiplier/_1137_ ),
    .ZN(\u_multiplier/_1154_ ));
 MUX2_X1 \u_multiplier/_2034_  (.A(\u_multiplier/_0988_ ),
    .B(\u_multiplier/_0990_ ),
    .S(\u_multiplier/_1059_ ),
    .Z(\u_multiplier/_1155_ ));
 MUX2_X1 \u_multiplier/_2035_  (.A(\u_multiplier/_1130_ ),
    .B(\u_multiplier/_1155_ ),
    .S(\u_multiplier/_0937_ ),
    .Z(\u_multiplier/_1156_ ));
 NOR3_X1 \u_multiplier/_2036_  (.A1(\u_multiplier/_0936_ ),
    .A2(\u_multiplier/_1103_ ),
    .A3(\u_multiplier/_1104_ ),
    .ZN(\u_multiplier/_1157_ ));
 AOI21_X1 \u_multiplier/_2037_  (.A(\u_multiplier/_1157_ ),
    .B1(\u_multiplier/_1156_ ),
    .B2(\u_multiplier/_0936_ ),
    .ZN(\u_multiplier/_1158_ ));
 NOR2_X1 \u_multiplier/_2038_  (.A1(\u_multiplier/_0938_ ),
    .A2(\u_multiplier/_1062_ ),
    .ZN(\u_multiplier/_1159_ ));
 AOI21_X1 \u_multiplier/_2039_  (.A(\u_multiplier/_1159_ ),
    .B1(\u_multiplier/_1158_ ),
    .B2(\u_multiplier/_0938_ ),
    .ZN(\u_multiplier/_1160_ ));
 AOI21_X2 \u_multiplier/_2040_  (.A(\u_multiplier/dec_out [4]),
    .B1(\u_multiplier/_1160_ ),
    .B2(\u_multiplier/_0939_ ),
    .ZN(\u_multiplier/_1161_ ));
 MUX2_X1 \u_multiplier/_2041_  (.A(\u_multiplier/_0979_ ),
    .B(\u_multiplier/_0988_ ),
    .S(\u_multiplier/_0934_ ),
    .Z(\u_multiplier/_1162_ ));
 INV_X1 \u_multiplier/_2042_  (.A(\u_multiplier/_1162_ ),
    .ZN(\u_multiplier/_1163_ ));
 MUX2_X1 \u_multiplier/_2043_  (.A(\u_multiplier/_1162_ ),
    .B(\u_multiplier/_1109_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_1164_ ));
 NOR4_X2 \u_multiplier/_2044_  (.A1(\u_multiplier/code_x [0]),
    .A2(\u_multiplier/code_x [1]),
    .A3(\u_multiplier/_0935_ ),
    .A4(\u_multiplier/_0945_ ),
    .ZN(\u_multiplier/_1165_ ));
 AOI21_X2 \u_multiplier/_2045_  (.A(\u_multiplier/_1165_ ),
    .B1(\u_multiplier/_1164_ ),
    .B2(\u_multiplier/_0935_ ),
    .ZN(\u_multiplier/_1166_ ));
 NOR2_X1 \u_multiplier/_2046_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_1166_ ),
    .ZN(\u_multiplier/_1167_ ));
 MUX2_X1 \u_multiplier/_2047_  (.A(\u_multiplier/_0981_ ),
    .B(\u_multiplier/_0990_ ),
    .S(\u_multiplier/_0930_ ),
    .Z(\u_multiplier/_1168_ ));
 NAND2_X1 \u_multiplier/_2048_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_1114_ ),
    .ZN(\u_multiplier/_1169_ ));
 OAI21_X1 \u_multiplier/_2049_  (.A(\u_multiplier/_1169_ ),
    .B1(\u_multiplier/_1168_ ),
    .B2(\u_multiplier/code_y [1]),
    .ZN(\u_multiplier/_1170_ ));
 NOR2_X1 \u_multiplier/_2050_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_1170_ ),
    .ZN(\u_multiplier/_1171_ ));
 AOI21_X2 \u_multiplier/_2051_  (.A(\u_multiplier/_1171_ ),
    .B1(\u_multiplier/_1068_ ),
    .B2(\u_multiplier/code_y [2]),
    .ZN(\u_multiplier/_1172_ ));
 NOR2_X1 \u_multiplier/_2052_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_1172_ ),
    .ZN(\u_multiplier/_1173_ ));
 NAND2_X1 \u_multiplier/_2053_  (.A1(\u_multiplier/_1167_ ),
    .A2(\u_multiplier/_1173_ ),
    .ZN(\u_multiplier/_1174_ ));
 XOR2_X2 \u_multiplier/_2054_  (.A(\u_multiplier/_1167_ ),
    .B(\u_multiplier/_1173_ ),
    .Z(\u_multiplier/_1175_ ));
 INV_X1 \u_multiplier/_2055_  (.A(\u_multiplier/_1175_ ),
    .ZN(\u_multiplier/_1176_ ));
 XNOR2_X1 \u_multiplier/_2056_  (.A(\u_multiplier/_1161_ ),
    .B(\u_multiplier/_1175_ ),
    .ZN(\u_multiplier/_1177_ ));
 AND2_X1 \u_multiplier/_2057_  (.A1(\u_multiplier/_1154_ ),
    .A2(\u_multiplier/_1177_ ),
    .ZN(\u_multiplier/_1178_ ));
 NAND2_X1 \u_multiplier/_2058_  (.A1(\u_multiplier/_1154_ ),
    .A2(\u_multiplier/_1177_ ),
    .ZN(\u_multiplier/_1179_ ));
 OR2_X1 \u_multiplier/_2059_  (.A1(\u_multiplier/_1154_ ),
    .A2(\u_multiplier/_1177_ ),
    .ZN(\u_multiplier/_1180_ ));
 NAND2_X1 \u_multiplier/_2060_  (.A1(\u_multiplier/_1179_ ),
    .A2(\u_multiplier/_1180_ ),
    .ZN(\u_multiplier/_1181_ ));
 AOI21_X1 \u_multiplier/_2061_  (.A(\u_multiplier/_0943_ ),
    .B1(\u_multiplier/_1152_ ),
    .B2(\u_multiplier/_1181_ ),
    .ZN(\u_multiplier/_1182_ ));
 OAI21_X1 \u_multiplier/_2062_  (.A(\u_multiplier/_1182_ ),
    .B1(\u_multiplier/_1181_ ),
    .B2(\u_multiplier/_1152_ ),
    .ZN(\u_multiplier/_1183_ ));
 INV_X1 \u_multiplier/_2063_  (.A(\u_multiplier/_1183_ ),
    .ZN(product[4]));
 AOI21_X1 \u_multiplier/_2064_  (.A(\u_multiplier/_1178_ ),
    .B1(\u_multiplier/_1180_ ),
    .B2(\u_multiplier/_1153_ ),
    .ZN(\u_multiplier/_1184_ ));
 OAI21_X1 \u_multiplier/_2065_  (.A(\u_multiplier/_1179_ ),
    .B1(\u_multiplier/_1181_ ),
    .B2(\u_multiplier/_1152_ ),
    .ZN(\u_multiplier/_1185_ ));
 OAI21_X2 \u_multiplier/_2066_  (.A(\u_multiplier/_1174_ ),
    .B1(\u_multiplier/_1176_ ),
    .B2(\u_multiplier/_1161_ ),
    .ZN(\u_multiplier/_1186_ ));
 MUX2_X1 \u_multiplier/_2067_  (.A(\u_multiplier/_0991_ ),
    .B(\u_multiplier/_0993_ ),
    .S(\u_multiplier/_1059_ ),
    .Z(\u_multiplier/_1187_ ));
 AND2_X1 \u_multiplier/_2068_  (.A1(\u_multiplier/_0937_ ),
    .A2(\u_multiplier/_1187_ ),
    .ZN(\u_multiplier/_1188_ ));
 AOI21_X1 \u_multiplier/_2069_  (.A(\u_multiplier/_1188_ ),
    .B1(\u_multiplier/_1155_ ),
    .B2(\u_multiplier/K [0]),
    .ZN(\u_multiplier/_1189_ ));
 MUX2_X1 \u_multiplier/_2070_  (.A(\u_multiplier/_1155_ ),
    .B(\u_multiplier/_1187_ ),
    .S(\u_multiplier/_0937_ ),
    .Z(\u_multiplier/_1190_ ));
 MUX2_X1 \u_multiplier/_2071_  (.A(\u_multiplier/_1132_ ),
    .B(\u_multiplier/_1190_ ),
    .S(\u_multiplier/_0936_ ),
    .Z(\u_multiplier/_1191_ ));
 MUX2_X2 \u_multiplier/_2072_  (.A(\u_multiplier/_1080_ ),
    .B(\u_multiplier/_1191_ ),
    .S(\u_multiplier/_0938_ ),
    .Z(\u_multiplier/_1192_ ));
 AOI21_X4 \u_multiplier/_2073_  (.A(\u_multiplier/dec_out [5]),
    .B1(\u_multiplier/_1192_ ),
    .B2(\u_multiplier/_0939_ ),
    .ZN(\u_multiplier/_1193_ ));
 MUX2_X1 \u_multiplier/_2074_  (.A(\u_multiplier/_0988_ ),
    .B(\u_multiplier/_0991_ ),
    .S(\u_multiplier/_0934_ ),
    .Z(\u_multiplier/_1194_ ));
 INV_X1 \u_multiplier/_2075_  (.A(\u_multiplier/_1194_ ),
    .ZN(\u_multiplier/_1195_ ));
 MUX2_X1 \u_multiplier/_2076_  (.A(\u_multiplier/_1195_ ),
    .B(\u_multiplier/_1138_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_1196_ ));
 MUX2_X1 \u_multiplier/_2077_  (.A(\u_multiplier/_1085_ ),
    .B(\u_multiplier/_1196_ ),
    .S(\u_multiplier/_0935_ ),
    .Z(\u_multiplier/_1197_ ));
 MUX2_X1 \u_multiplier/_2078_  (.A(\u_multiplier/_0990_ ),
    .B(\u_multiplier/_0993_ ),
    .S(\u_multiplier/_0930_ ),
    .Z(\u_multiplier/_1198_ ));
 NAND2_X1 \u_multiplier/_2079_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_1141_ ),
    .ZN(\u_multiplier/_1199_ ));
 OAI21_X1 \u_multiplier/_2080_  (.A(\u_multiplier/_1199_ ),
    .B1(\u_multiplier/_1198_ ),
    .B2(\u_multiplier/code_y [1]),
    .ZN(\u_multiplier/_1200_ ));
 MUX2_X1 \u_multiplier/_2081_  (.A(\u_multiplier/_1088_ ),
    .B(\u_multiplier/_1200_ ),
    .S(\u_multiplier/_0931_ ),
    .Z(\u_multiplier/_1201_ ));
 OAI22_X1 \u_multiplier/_2082_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_1197_ ),
    .B1(\u_multiplier/_1201_ ),
    .B2(\u_multiplier/code_y [3]),
    .ZN(\u_multiplier/_1202_ ));
 OR4_X1 \u_multiplier/_2083_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/code_x [3]),
    .A3(\u_multiplier/_1197_ ),
    .A4(\u_multiplier/_1201_ ),
    .ZN(\u_multiplier/_1203_ ));
 AND2_X1 \u_multiplier/_2084_  (.A1(\u_multiplier/_1202_ ),
    .A2(\u_multiplier/_1203_ ),
    .ZN(\u_multiplier/_1204_ ));
 INV_X1 \u_multiplier/_2085_  (.A(\u_multiplier/_1204_ ),
    .ZN(\u_multiplier/_1205_ ));
 XNOR2_X2 \u_multiplier/_2086_  (.A(\u_multiplier/_1193_ ),
    .B(\u_multiplier/_1204_ ),
    .ZN(\u_multiplier/_1206_ ));
 NAND2_X1 \u_multiplier/_2087_  (.A1(\u_multiplier/_1186_ ),
    .A2(\u_multiplier/_1206_ ),
    .ZN(\u_multiplier/_1207_ ));
 XOR2_X2 \u_multiplier/_2088_  (.A(\u_multiplier/_1186_ ),
    .B(\u_multiplier/_1206_ ),
    .Z(\u_multiplier/_1208_ ));
 INV_X1 \u_multiplier/_2089_  (.A(\u_multiplier/_1208_ ),
    .ZN(\u_multiplier/_1209_ ));
 NAND2_X1 \u_multiplier/_2090_  (.A1(\u_multiplier/_1185_ ),
    .A2(\u_multiplier/_1208_ ),
    .ZN(\u_multiplier/_1210_ ));
 OAI21_X1 \u_multiplier/_2091_  (.A(\u_multiplier/_1739_ ),
    .B1(\u_multiplier/_1185_ ),
    .B2(\u_multiplier/_1208_ ),
    .ZN(\u_multiplier/_1211_ ));
 AOI21_X1 \u_multiplier/_2092_  (.A(\u_multiplier/_1211_ ),
    .B1(\u_multiplier/_1208_ ),
    .B2(\u_multiplier/_1185_ ),
    .ZN(product[5]));
 AND2_X1 \u_multiplier/_2093_  (.A1(\u_multiplier/_1207_ ),
    .A2(\u_multiplier/_1210_ ),
    .ZN(\u_multiplier/_1212_ ));
 OAI21_X1 \u_multiplier/_2094_  (.A(\u_multiplier/_1207_ ),
    .B1(\u_multiplier/_1209_ ),
    .B2(\u_multiplier/_1184_ ),
    .ZN(\u_multiplier/_1213_ ));
 OAI21_X2 \u_multiplier/_2095_  (.A(\u_multiplier/_1203_ ),
    .B1(\u_multiplier/_1205_ ),
    .B2(\u_multiplier/_1193_ ),
    .ZN(\u_multiplier/_1214_ ));
 MUX2_X1 \u_multiplier/_2096_  (.A(\u_multiplier/_0960_ ),
    .B(\u_multiplier/_0961_ ),
    .S(\u_multiplier/_1059_ ),
    .Z(\u_multiplier/_1215_ ));
 MUX2_X1 \u_multiplier/_2097_  (.A(\u_multiplier/_1187_ ),
    .B(\u_multiplier/_1215_ ),
    .S(\u_multiplier/_0937_ ),
    .Z(\u_multiplier/_1216_ ));
 MUX2_X1 \u_multiplier/_2098_  (.A(\u_multiplier/_1156_ ),
    .B(\u_multiplier/_1216_ ),
    .S(\u_multiplier/_0936_ ),
    .Z(\u_multiplier/_1217_ ));
 NAND2_X1 \u_multiplier/_2099_  (.A1(\u_multiplier/_0938_ ),
    .A2(\u_multiplier/_1217_ ),
    .ZN(\u_multiplier/_1218_ ));
 OAI21_X2 \u_multiplier/_2100_  (.A(\u_multiplier/_1218_ ),
    .B1(\u_multiplier/_1107_ ),
    .B2(\u_multiplier/_0938_ ),
    .ZN(\u_multiplier/_1219_ ));
 AOI21_X2 \u_multiplier/_2101_  (.A(\u_multiplier/dec_out [6]),
    .B1(\u_multiplier/_1219_ ),
    .B2(\u_multiplier/_0939_ ),
    .ZN(\u_multiplier/_1220_ ));
 MUX2_X1 \u_multiplier/_2102_  (.A(\u_multiplier/_0960_ ),
    .B(\u_multiplier/_0991_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_1221_ ));
 NAND2_X1 \u_multiplier/_2103_  (.A1(\u_multiplier/code_x [1]),
    .A2(\u_multiplier/_1163_ ),
    .ZN(\u_multiplier/_1222_ ));
 OAI21_X1 \u_multiplier/_2104_  (.A(\u_multiplier/_1222_ ),
    .B1(\u_multiplier/_1221_ ),
    .B2(\u_multiplier/code_x [1]),
    .ZN(\u_multiplier/_1223_ ));
 NAND2_X1 \u_multiplier/_2105_  (.A1(\u_multiplier/_0935_ ),
    .A2(\u_multiplier/_1223_ ),
    .ZN(\u_multiplier/_1224_ ));
 OAI21_X2 \u_multiplier/_2106_  (.A(\u_multiplier/_1224_ ),
    .B1(\u_multiplier/_1110_ ),
    .B2(\u_multiplier/_0935_ ),
    .ZN(\u_multiplier/_1225_ ));
 OR2_X1 \u_multiplier/_2107_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_1225_ ),
    .ZN(\u_multiplier/_1226_ ));
 MUX2_X1 \u_multiplier/_2108_  (.A(\u_multiplier/_0962_ ),
    .B(\u_multiplier/_0994_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_1227_ ));
 NOR2_X1 \u_multiplier/_2109_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_1227_ ),
    .ZN(\u_multiplier/_1228_ ));
 AOI21_X1 \u_multiplier/_2110_  (.A(\u_multiplier/_1228_ ),
    .B1(\u_multiplier/_1168_ ),
    .B2(\u_multiplier/code_y [1]),
    .ZN(\u_multiplier/_1229_ ));
 NAND2_X1 \u_multiplier/_2111_  (.A1(\u_multiplier/_0931_ ),
    .A2(\u_multiplier/_1229_ ),
    .ZN(\u_multiplier/_1230_ ));
 OAI21_X2 \u_multiplier/_2112_  (.A(\u_multiplier/_1230_ ),
    .B1(\u_multiplier/_1116_ ),
    .B2(\u_multiplier/_0931_ ),
    .ZN(\u_multiplier/_1231_ ));
 NOR2_X1 \u_multiplier/_2113_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_1231_ ),
    .ZN(\u_multiplier/_1232_ ));
 NOR3_X1 \u_multiplier/_2114_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_1226_ ),
    .A3(\u_multiplier/_1231_ ),
    .ZN(\u_multiplier/_1233_ ));
 XNOR2_X2 \u_multiplier/_2115_  (.A(\u_multiplier/_1226_ ),
    .B(\u_multiplier/_1232_ ),
    .ZN(\u_multiplier/_1234_ ));
 INV_X1 \u_multiplier/_2116_  (.A(\u_multiplier/_1234_ ),
    .ZN(\u_multiplier/_1235_ ));
 NOR2_X1 \u_multiplier/_2117_  (.A1(\u_multiplier/_1220_ ),
    .A2(\u_multiplier/_1235_ ),
    .ZN(\u_multiplier/_1236_ ));
 XNOR2_X2 \u_multiplier/_2118_  (.A(\u_multiplier/_1220_ ),
    .B(\u_multiplier/_1234_ ),
    .ZN(\u_multiplier/_1237_ ));
 AND2_X1 \u_multiplier/_2119_  (.A1(\u_multiplier/_1214_ ),
    .A2(\u_multiplier/_1237_ ),
    .ZN(\u_multiplier/_1238_ ));
 NAND2_X1 \u_multiplier/_2120_  (.A1(\u_multiplier/_1214_ ),
    .A2(\u_multiplier/_1237_ ),
    .ZN(\u_multiplier/_1239_ ));
 XNOR2_X2 \u_multiplier/_2121_  (.A(\u_multiplier/_1214_ ),
    .B(\u_multiplier/_1237_ ),
    .ZN(\u_multiplier/_1240_ ));
 INV_X1 \u_multiplier/_2122_  (.A(\u_multiplier/_1240_ ),
    .ZN(\u_multiplier/_1241_ ));
 AOI21_X1 \u_multiplier/_2123_  (.A(\u_multiplier/_0943_ ),
    .B1(\u_multiplier/_1212_ ),
    .B2(\u_multiplier/_1240_ ),
    .ZN(\u_multiplier/_1242_ ));
 OAI21_X1 \u_multiplier/_2124_  (.A(\u_multiplier/_1242_ ),
    .B1(\u_multiplier/_1240_ ),
    .B2(\u_multiplier/_1212_ ),
    .ZN(\u_multiplier/_1243_ ));
 INV_X1 \u_multiplier/_2125_  (.A(\u_multiplier/_1243_ ),
    .ZN(product[6]));
 AOI21_X1 \u_multiplier/_2126_  (.A(\u_multiplier/_1238_ ),
    .B1(\u_multiplier/_1241_ ),
    .B2(\u_multiplier/_1213_ ),
    .ZN(\u_multiplier/_1244_ ));
 OAI21_X1 \u_multiplier/_2127_  (.A(\u_multiplier/_1239_ ),
    .B1(\u_multiplier/_1240_ ),
    .B2(\u_multiplier/_1212_ ),
    .ZN(\u_multiplier/_1245_ ));
 NOR2_X1 \u_multiplier/_2128_  (.A1(\u_multiplier/_1233_ ),
    .A2(\u_multiplier/_1236_ ),
    .ZN(\u_multiplier/_1246_ ));
 MUX2_X1 \u_multiplier/_2129_  (.A(\u_multiplier/_0956_ ),
    .B(\u_multiplier/_0958_ ),
    .S(\u_multiplier/_1059_ ),
    .Z(\u_multiplier/_1247_ ));
 NAND2_X1 \u_multiplier/_2130_  (.A1(\u_multiplier/_0937_ ),
    .A2(\u_multiplier/_1247_ ),
    .ZN(\u_multiplier/_1248_ ));
 NAND2_X1 \u_multiplier/_2131_  (.A1(\u_multiplier/K [0]),
    .A2(\u_multiplier/_1215_ ),
    .ZN(\u_multiplier/_1249_ ));
 AND2_X1 \u_multiplier/_2132_  (.A1(\u_multiplier/_1248_ ),
    .A2(\u_multiplier/_1249_ ),
    .ZN(\u_multiplier/_1250_ ));
 MUX2_X1 \u_multiplier/_2133_  (.A(\u_multiplier/_1189_ ),
    .B(\u_multiplier/_1250_ ),
    .S(\u_multiplier/_0936_ ),
    .Z(\u_multiplier/_1251_ ));
 MUX2_X1 \u_multiplier/_2134_  (.A(\u_multiplier/_1135_ ),
    .B(\u_multiplier/_1251_ ),
    .S(\u_multiplier/_0938_ ),
    .Z(\u_multiplier/_1252_ ));
 NOR2_X1 \u_multiplier/_2135_  (.A1(\u_multiplier/K [3]),
    .A2(\u_multiplier/_1252_ ),
    .ZN(\u_multiplier/_1253_ ));
 NOR2_X2 \u_multiplier/_2136_  (.A1(\u_multiplier/dec_out [7]),
    .A2(\u_multiplier/_1253_ ),
    .ZN(\u_multiplier/_1254_ ));
 MUX2_X1 \u_multiplier/_2137_  (.A(\u_multiplier/_0956_ ),
    .B(\u_multiplier/_0960_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_1255_ ));
 NAND2_X1 \u_multiplier/_2138_  (.A1(\u_multiplier/code_x [1]),
    .A2(\u_multiplier/_1195_ ),
    .ZN(\u_multiplier/_1256_ ));
 OAI21_X1 \u_multiplier/_2139_  (.A(\u_multiplier/_1256_ ),
    .B1(\u_multiplier/_1255_ ),
    .B2(\u_multiplier/code_x [1]),
    .ZN(\u_multiplier/_1257_ ));
 MUX2_X1 \u_multiplier/_2140_  (.A(\u_multiplier/_1139_ ),
    .B(\u_multiplier/_1257_ ),
    .S(\u_multiplier/_0935_ ),
    .Z(\u_multiplier/_1258_ ));
 NOR2_X2 \u_multiplier/_2141_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_1258_ ),
    .ZN(\u_multiplier/_1259_ ));
 NAND2_X1 \u_multiplier/_2142_  (.A1(\u_multiplier/code_y [0]),
    .A2(\u_multiplier/_0962_ ),
    .ZN(\u_multiplier/_1260_ ));
 OAI21_X1 \u_multiplier/_2143_  (.A(\u_multiplier/_1260_ ),
    .B1(\u_multiplier/_0958_ ),
    .B2(\u_multiplier/code_y [0]),
    .ZN(\u_multiplier/_1261_ ));
 NOR2_X1 \u_multiplier/_2144_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_1261_ ),
    .ZN(\u_multiplier/_1262_ ));
 AOI21_X2 \u_multiplier/_2145_  (.A(\u_multiplier/_1262_ ),
    .B1(\u_multiplier/_1198_ ),
    .B2(\u_multiplier/code_y [1]),
    .ZN(\u_multiplier/_1263_ ));
 MUX2_X2 \u_multiplier/_2146_  (.A(\u_multiplier/_1142_ ),
    .B(\u_multiplier/_1263_ ),
    .S(\u_multiplier/_0931_ ),
    .Z(\u_multiplier/_1264_ ));
 NOR2_X2 \u_multiplier/_2147_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_1264_ ),
    .ZN(\u_multiplier/_1265_ ));
 XNOR2_X2 \u_multiplier/_2148_  (.A(\u_multiplier/_1259_ ),
    .B(\u_multiplier/_1265_ ),
    .ZN(\u_multiplier/_1266_ ));
 NOR2_X1 \u_multiplier/_2149_  (.A1(\u_multiplier/_1254_ ),
    .A2(\u_multiplier/_1266_ ),
    .ZN(\u_multiplier/_1267_ ));
 XOR2_X2 \u_multiplier/_2150_  (.A(\u_multiplier/_1254_ ),
    .B(\u_multiplier/_1266_ ),
    .Z(\u_multiplier/_1268_ ));
 OAI21_X1 \u_multiplier/_2151_  (.A(\u_multiplier/_1268_ ),
    .B1(\u_multiplier/_1236_ ),
    .B2(\u_multiplier/_1233_ ),
    .ZN(\u_multiplier/_1269_ ));
 XNOR2_X2 \u_multiplier/_2152_  (.A(\u_multiplier/_1246_ ),
    .B(\u_multiplier/_1268_ ),
    .ZN(\u_multiplier/_1270_ ));
 INV_X1 \u_multiplier/_2153_  (.A(\u_multiplier/_1270_ ),
    .ZN(\u_multiplier/_1271_ ));
 OAI21_X1 \u_multiplier/_2154_  (.A(\u_multiplier/_1739_ ),
    .B1(\u_multiplier/_1245_ ),
    .B2(\u_multiplier/_1270_ ),
    .ZN(\u_multiplier/_1272_ ));
 AOI21_X1 \u_multiplier/_2155_  (.A(\u_multiplier/_1272_ ),
    .B1(\u_multiplier/_1270_ ),
    .B2(\u_multiplier/_1245_ ),
    .ZN(product[7]));
 OAI21_X2 \u_multiplier/_2156_  (.A(\u_multiplier/_1269_ ),
    .B1(\u_multiplier/_1271_ ),
    .B2(\u_multiplier/_1244_ ),
    .ZN(\u_multiplier/_1273_ ));
 AOI21_X2 \u_multiplier/_2157_  (.A(\u_multiplier/_1267_ ),
    .B1(\u_multiplier/_1265_ ),
    .B2(\u_multiplier/_1259_ ),
    .ZN(\u_multiplier/_1274_ ));
 MUX2_X1 \u_multiplier/_2158_  (.A(\u_multiplier/_0950_ ),
    .B(\u_multiplier/_0952_ ),
    .S(\u_multiplier/_1059_ ),
    .Z(\u_multiplier/_1275_ ));
 MUX2_X1 \u_multiplier/_2159_  (.A(\u_multiplier/_1247_ ),
    .B(\u_multiplier/_1275_ ),
    .S(\u_multiplier/_0937_ ),
    .Z(\u_multiplier/_1276_ ));
 AND2_X1 \u_multiplier/_2160_  (.A1(\u_multiplier/_0936_ ),
    .A2(\u_multiplier/_1276_ ),
    .ZN(\u_multiplier/_1277_ ));
 AOI21_X2 \u_multiplier/_2161_  (.A(\u_multiplier/_1277_ ),
    .B1(\u_multiplier/_1216_ ),
    .B2(\u_multiplier/K [1]),
    .ZN(\u_multiplier/_1278_ ));
 MUX2_X1 \u_multiplier/_2162_  (.A(\u_multiplier/_1158_ ),
    .B(\u_multiplier/_1278_ ),
    .S(\u_multiplier/_0938_ ),
    .Z(\u_multiplier/_1279_ ));
 AOI21_X1 \u_multiplier/_2163_  (.A(\u_multiplier/dec_out [8]),
    .B1(\u_multiplier/_1063_ ),
    .B2(\u_multiplier/K [3]),
    .ZN(\u_multiplier/_1280_ ));
 OAI21_X2 \u_multiplier/_2164_  (.A(\u_multiplier/_1280_ ),
    .B1(\u_multiplier/_1279_ ),
    .B2(\u_multiplier/K [3]),
    .ZN(\u_multiplier/_1281_ ));
 MUX2_X1 \u_multiplier/_2165_  (.A(\u_multiplier/_0950_ ),
    .B(\u_multiplier/_0956_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_1282_ ));
 MUX2_X1 \u_multiplier/_2166_  (.A(\u_multiplier/_1282_ ),
    .B(\u_multiplier/_1221_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_1283_ ));
 MUX2_X1 \u_multiplier/_2167_  (.A(\u_multiplier/_1164_ ),
    .B(\u_multiplier/_1283_ ),
    .S(\u_multiplier/_0935_ ),
    .Z(\u_multiplier/_1284_ ));
 AND2_X1 \u_multiplier/_2168_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_1066_ ),
    .ZN(\u_multiplier/_1285_ ));
 AOI21_X2 \u_multiplier/_2169_  (.A(\u_multiplier/_1285_ ),
    .B1(\u_multiplier/_1284_ ),
    .B2(\u_multiplier/_0933_ ),
    .ZN(\u_multiplier/_1286_ ));
 MUX2_X1 \u_multiplier/_2170_  (.A(\u_multiplier/_0952_ ),
    .B(\u_multiplier/_0958_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_1287_ ));
 NOR2_X1 \u_multiplier/_2171_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_1287_ ),
    .ZN(\u_multiplier/_1288_ ));
 AOI21_X2 \u_multiplier/_2172_  (.A(\u_multiplier/_1288_ ),
    .B1(\u_multiplier/_1227_ ),
    .B2(\u_multiplier/code_y [1]),
    .ZN(\u_multiplier/_1289_ ));
 NAND2_X1 \u_multiplier/_2173_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_1170_ ),
    .ZN(\u_multiplier/_1290_ ));
 OAI21_X2 \u_multiplier/_2174_  (.A(\u_multiplier/_1290_ ),
    .B1(\u_multiplier/_1289_ ),
    .B2(\u_multiplier/code_y [2]),
    .ZN(\u_multiplier/_1291_ ));
 MUX2_X1 \u_multiplier/_2175_  (.A(\u_multiplier/_1069_ ),
    .B(\u_multiplier/_1291_ ),
    .S(\u_multiplier/_0932_ ),
    .Z(\u_multiplier/_1292_ ));
 XOR2_X2 \u_multiplier/_2176_  (.A(\u_multiplier/_1286_ ),
    .B(\u_multiplier/_1292_ ),
    .Z(\u_multiplier/_1293_ ));
 NAND2_X1 \u_multiplier/_2177_  (.A1(\u_multiplier/_1281_ ),
    .A2(\u_multiplier/_1293_ ),
    .ZN(\u_multiplier/_1294_ ));
 XNOR2_X2 \u_multiplier/_2178_  (.A(\u_multiplier/_1281_ ),
    .B(\u_multiplier/_1293_ ),
    .ZN(\u_multiplier/_1295_ ));
 NOR2_X1 \u_multiplier/_2179_  (.A1(\u_multiplier/_1274_ ),
    .A2(\u_multiplier/_1295_ ),
    .ZN(\u_multiplier/_1296_ ));
 XOR2_X2 \u_multiplier/_2180_  (.A(\u_multiplier/_1274_ ),
    .B(\u_multiplier/_1295_ ),
    .Z(\u_multiplier/_1297_ ));
 AND2_X1 \u_multiplier/_2181_  (.A1(\u_multiplier/_1273_ ),
    .A2(\u_multiplier/_1297_ ),
    .ZN(\u_multiplier/_1298_ ));
 OAI21_X1 \u_multiplier/_2182_  (.A(\u_multiplier/_1739_ ),
    .B1(\u_multiplier/_1273_ ),
    .B2(\u_multiplier/_1297_ ),
    .ZN(\u_multiplier/_1299_ ));
 NOR2_X1 \u_multiplier/_2183_  (.A1(\u_multiplier/_1298_ ),
    .A2(\u_multiplier/_1299_ ),
    .ZN(product[8]));
 OAI21_X2 \u_multiplier/_2184_  (.A(\u_multiplier/_1294_ ),
    .B1(\u_multiplier/_1292_ ),
    .B2(\u_multiplier/_1286_ ),
    .ZN(\u_multiplier/_1300_ ));
 MUX2_X1 \u_multiplier/_2185_  (.A(\u_multiplier/_0946_ ),
    .B(\u_multiplier/_0948_ ),
    .S(\u_multiplier/_1059_ ),
    .Z(\u_multiplier/_1301_ ));
 AND2_X1 \u_multiplier/_2186_  (.A1(\u_multiplier/_0937_ ),
    .A2(\u_multiplier/_1301_ ),
    .ZN(\u_multiplier/_1302_ ));
 AOI21_X1 \u_multiplier/_2187_  (.A(\u_multiplier/_1302_ ),
    .B1(\u_multiplier/_1275_ ),
    .B2(\u_multiplier/K [0]),
    .ZN(\u_multiplier/_1303_ ));
 MUX2_X1 \u_multiplier/_2188_  (.A(\u_multiplier/_1250_ ),
    .B(\u_multiplier/_1303_ ),
    .S(\u_multiplier/_0936_ ),
    .Z(\u_multiplier/_1304_ ));
 NOR2_X1 \u_multiplier/_2189_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/_1304_ ),
    .ZN(\u_multiplier/_1305_ ));
 AOI21_X2 \u_multiplier/_2190_  (.A(\u_multiplier/_1305_ ),
    .B1(\u_multiplier/_1191_ ),
    .B2(\u_multiplier/K [2]),
    .ZN(\u_multiplier/_1306_ ));
 NOR2_X1 \u_multiplier/_2191_  (.A1(\u_multiplier/K [3]),
    .A2(\u_multiplier/_1306_ ),
    .ZN(\u_multiplier/_1307_ ));
 AOI211_X2 \u_multiplier/_2192_  (.A(\u_multiplier/dec_out [9]),
    .B(\u_multiplier/_1307_ ),
    .C1(\u_multiplier/_1081_ ),
    .C2(\u_multiplier/K [3]),
    .ZN(\u_multiplier/_1308_ ));
 MUX2_X1 \u_multiplier/_2193_  (.A(\u_multiplier/_0946_ ),
    .B(\u_multiplier/_0950_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_1309_ ));
 MUX2_X1 \u_multiplier/_2194_  (.A(\u_multiplier/_1309_ ),
    .B(\u_multiplier/_1255_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_1310_ ));
 NOR2_X1 \u_multiplier/_2195_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_1310_ ),
    .ZN(\u_multiplier/_1311_ ));
 AOI21_X2 \u_multiplier/_2196_  (.A(\u_multiplier/_1311_ ),
    .B1(\u_multiplier/_1196_ ),
    .B2(\u_multiplier/code_x [2]),
    .ZN(\u_multiplier/_1312_ ));
 NOR2_X1 \u_multiplier/_2197_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_1312_ ),
    .ZN(\u_multiplier/_1313_ ));
 AOI21_X2 \u_multiplier/_2198_  (.A(\u_multiplier/_1313_ ),
    .B1(\u_multiplier/_1086_ ),
    .B2(\u_multiplier/code_x [3]),
    .ZN(\u_multiplier/_1314_ ));
 MUX2_X1 \u_multiplier/_2199_  (.A(\u_multiplier/_0948_ ),
    .B(\u_multiplier/_0952_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_1315_ ));
 NOR2_X1 \u_multiplier/_2200_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_1315_ ),
    .ZN(\u_multiplier/_1316_ ));
 AOI21_X1 \u_multiplier/_2201_  (.A(\u_multiplier/_1316_ ),
    .B1(\u_multiplier/_1261_ ),
    .B2(\u_multiplier/code_y [1]),
    .ZN(\u_multiplier/_1317_ ));
 NOR2_X1 \u_multiplier/_2202_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_1317_ ),
    .ZN(\u_multiplier/_1318_ ));
 AOI21_X2 \u_multiplier/_2203_  (.A(\u_multiplier/_1318_ ),
    .B1(\u_multiplier/_1200_ ),
    .B2(\u_multiplier/code_y [2]),
    .ZN(\u_multiplier/_1319_ ));
 NAND2_X1 \u_multiplier/_2204_  (.A1(\u_multiplier/_0932_ ),
    .A2(\u_multiplier/_1319_ ),
    .ZN(\u_multiplier/_1320_ ));
 OAI21_X1 \u_multiplier/_2205_  (.A(\u_multiplier/_1320_ ),
    .B1(\u_multiplier/_1089_ ),
    .B2(\u_multiplier/_0932_ ),
    .ZN(\u_multiplier/_1321_ ));
 XOR2_X1 \u_multiplier/_2206_  (.A(\u_multiplier/_1314_ ),
    .B(\u_multiplier/_1321_ ),
    .Z(\u_multiplier/_1322_ ));
 INV_X1 \u_multiplier/_2207_  (.A(\u_multiplier/_1322_ ),
    .ZN(\u_multiplier/_1323_ ));
 NOR2_X1 \u_multiplier/_2208_  (.A1(\u_multiplier/_1308_ ),
    .A2(\u_multiplier/_1323_ ),
    .ZN(\u_multiplier/_1324_ ));
 XNOR2_X2 \u_multiplier/_2209_  (.A(\u_multiplier/_1308_ ),
    .B(\u_multiplier/_1323_ ),
    .ZN(\u_multiplier/_1325_ ));
 INV_X1 \u_multiplier/_2210_  (.A(\u_multiplier/_1325_ ),
    .ZN(\u_multiplier/_1326_ ));
 NAND2_X1 \u_multiplier/_2211_  (.A1(\u_multiplier/_1300_ ),
    .A2(\u_multiplier/_1326_ ),
    .ZN(\u_multiplier/_1327_ ));
 XNOR2_X2 \u_multiplier/_2212_  (.A(\u_multiplier/_1300_ ),
    .B(\u_multiplier/_1325_ ),
    .ZN(\u_multiplier/_1328_ ));
 NOR3_X1 \u_multiplier/_2213_  (.A1(\u_multiplier/_1296_ ),
    .A2(\u_multiplier/_1298_ ),
    .A3(\u_multiplier/_1328_ ),
    .ZN(\u_multiplier/_1329_ ));
 NAND3_X2 \u_multiplier/_2214_  (.A1(\u_multiplier/_1273_ ),
    .A2(\u_multiplier/_1297_ ),
    .A3(\u_multiplier/_1328_ ),
    .ZN(\u_multiplier/_1330_ ));
 NAND2_X1 \u_multiplier/_2215_  (.A1(\u_multiplier/_1296_ ),
    .A2(\u_multiplier/_1328_ ),
    .ZN(\u_multiplier/_1331_ ));
 NAND3_X1 \u_multiplier/_2216_  (.A1(\u_multiplier/_1739_ ),
    .A2(\u_multiplier/_1330_ ),
    .A3(\u_multiplier/_1331_ ),
    .ZN(\u_multiplier/_1332_ ));
 NOR2_X1 \u_multiplier/_2217_  (.A1(\u_multiplier/_1329_ ),
    .A2(\u_multiplier/_1332_ ),
    .ZN(product[9]));
 AND2_X1 \u_multiplier/_2218_  (.A1(\u_multiplier/_1327_ ),
    .A2(\u_multiplier/_1331_ ),
    .ZN(\u_multiplier/_1333_ ));
 AOI21_X2 \u_multiplier/_2219_  (.A(\u_multiplier/_1324_ ),
    .B1(\u_multiplier/_1321_ ),
    .B2(\u_multiplier/_1314_ ),
    .ZN(\u_multiplier/_1334_ ));
 MUX2_X1 \u_multiplier/_2220_  (.A(\u_multiplier/_1029_ ),
    .B(\u_multiplier/_1031_ ),
    .S(\u_multiplier/_1059_ ),
    .Z(\u_multiplier/_1335_ ));
 MUX2_X1 \u_multiplier/_2221_  (.A(\u_multiplier/_1301_ ),
    .B(\u_multiplier/_1335_ ),
    .S(\u_multiplier/_0937_ ),
    .Z(\u_multiplier/_1336_ ));
 MUX2_X1 \u_multiplier/_2222_  (.A(\u_multiplier/_1276_ ),
    .B(\u_multiplier/_1336_ ),
    .S(\u_multiplier/_0936_ ),
    .Z(\u_multiplier/_1337_ ));
 MUX2_X1 \u_multiplier/_2223_  (.A(\u_multiplier/_1217_ ),
    .B(\u_multiplier/_1337_ ),
    .S(\u_multiplier/_0938_ ),
    .Z(\u_multiplier/_1338_ ));
 NOR3_X2 \u_multiplier/_2224_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/_0939_ ),
    .A3(\u_multiplier/_1107_ ),
    .ZN(\u_multiplier/_1339_ ));
 AOI211_X2 \u_multiplier/_2225_  (.A(\u_multiplier/dec_out [10]),
    .B(\u_multiplier/_1339_ ),
    .C1(\u_multiplier/_1338_ ),
    .C2(\u_multiplier/_0939_ ),
    .ZN(\u_multiplier/_1340_ ));
 MUX2_X1 \u_multiplier/_2226_  (.A(\u_multiplier/_0946_ ),
    .B(\u_multiplier/_1029_ ),
    .S(\u_multiplier/_0934_ ),
    .Z(\u_multiplier/_1341_ ));
 MUX2_X1 \u_multiplier/_2227_  (.A(\u_multiplier/_1341_ ),
    .B(\u_multiplier/_1282_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_1342_ ));
 NAND2_X1 \u_multiplier/_2228_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_1223_ ),
    .ZN(\u_multiplier/_1343_ ));
 OAI21_X1 \u_multiplier/_2229_  (.A(\u_multiplier/_1343_ ),
    .B1(\u_multiplier/_1342_ ),
    .B2(\u_multiplier/code_x [2]),
    .ZN(\u_multiplier/_1344_ ));
 MUX2_X1 \u_multiplier/_2230_  (.A(\u_multiplier/_1111_ ),
    .B(\u_multiplier/_1344_ ),
    .S(\u_multiplier/_0933_ ),
    .Z(\u_multiplier/_1345_ ));
 MUX2_X1 \u_multiplier/_2231_  (.A(\u_multiplier/_0948_ ),
    .B(\u_multiplier/_1031_ ),
    .S(\u_multiplier/_0930_ ),
    .Z(\u_multiplier/_1346_ ));
 MUX2_X1 \u_multiplier/_2232_  (.A(\u_multiplier/_1346_ ),
    .B(\u_multiplier/_1287_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_1347_ ));
 NAND2_X1 \u_multiplier/_2233_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_1229_ ),
    .ZN(\u_multiplier/_1348_ ));
 OAI21_X1 \u_multiplier/_2234_  (.A(\u_multiplier/_1348_ ),
    .B1(\u_multiplier/_1347_ ),
    .B2(\u_multiplier/code_y [2]),
    .ZN(\u_multiplier/_1349_ ));
 MUX2_X1 \u_multiplier/_2235_  (.A(\u_multiplier/_1117_ ),
    .B(\u_multiplier/_1349_ ),
    .S(\u_multiplier/_0932_ ),
    .Z(\u_multiplier/_1350_ ));
 NOR2_X1 \u_multiplier/_2236_  (.A1(\u_multiplier/_1345_ ),
    .A2(\u_multiplier/_1350_ ),
    .ZN(\u_multiplier/_1351_ ));
 XNOR2_X2 \u_multiplier/_2237_  (.A(\u_multiplier/_1345_ ),
    .B(\u_multiplier/_1350_ ),
    .ZN(\u_multiplier/_1352_ ));
 NOR2_X1 \u_multiplier/_2238_  (.A1(\u_multiplier/_1340_ ),
    .A2(\u_multiplier/_1352_ ),
    .ZN(\u_multiplier/_1353_ ));
 XNOR2_X2 \u_multiplier/_2239_  (.A(\u_multiplier/_1340_ ),
    .B(\u_multiplier/_1352_ ),
    .ZN(\u_multiplier/_1354_ ));
 XNOR2_X2 \u_multiplier/_2240_  (.A(\u_multiplier/_1334_ ),
    .B(\u_multiplier/_1354_ ),
    .ZN(\u_multiplier/_1355_ ));
 AOI21_X1 \u_multiplier/_2241_  (.A(\u_multiplier/_1355_ ),
    .B1(\u_multiplier/_1333_ ),
    .B2(\u_multiplier/_1330_ ),
    .ZN(\u_multiplier/_1356_ ));
 AND3_X1 \u_multiplier/_2242_  (.A1(\u_multiplier/_1330_ ),
    .A2(\u_multiplier/_1333_ ),
    .A3(\u_multiplier/_1355_ ),
    .ZN(\u_multiplier/_1357_ ));
 NOR3_X1 \u_multiplier/_2243_  (.A1(\u_multiplier/_0943_ ),
    .A2(\u_multiplier/_1356_ ),
    .A3(\u_multiplier/_1357_ ),
    .ZN(product[10]));
 NOR2_X1 \u_multiplier/_2244_  (.A1(\u_multiplier/_1351_ ),
    .A2(\u_multiplier/_1353_ ),
    .ZN(\u_multiplier/_1358_ ));
 MUX2_X1 \u_multiplier/_2245_  (.A(\u_multiplier/_1025_ ),
    .B(\u_multiplier/_1027_ ),
    .S(\u_multiplier/_1059_ ),
    .Z(\u_multiplier/_1359_ ));
 MUX2_X1 \u_multiplier/_2246_  (.A(\u_multiplier/_1335_ ),
    .B(\u_multiplier/_1359_ ),
    .S(\u_multiplier/_0937_ ),
    .Z(\u_multiplier/_1360_ ));
 NOR2_X1 \u_multiplier/_2247_  (.A1(\u_multiplier/_0936_ ),
    .A2(\u_multiplier/_1303_ ),
    .ZN(\u_multiplier/_1361_ ));
 AOI21_X2 \u_multiplier/_2248_  (.A(\u_multiplier/_1361_ ),
    .B1(\u_multiplier/_1360_ ),
    .B2(\u_multiplier/_0936_ ),
    .ZN(\u_multiplier/_1362_ ));
 MUX2_X1 \u_multiplier/_2249_  (.A(\u_multiplier/_1251_ ),
    .B(\u_multiplier/_1362_ ),
    .S(\u_multiplier/_0938_ ),
    .Z(\u_multiplier/_1363_ ));
 AOI21_X1 \u_multiplier/_2250_  (.A(\u_multiplier/dec_out [11]),
    .B1(\u_multiplier/_1136_ ),
    .B2(\u_multiplier/K [3]),
    .ZN(\u_multiplier/_1364_ ));
 OAI21_X1 \u_multiplier/_2251_  (.A(\u_multiplier/_1364_ ),
    .B1(\u_multiplier/_1363_ ),
    .B2(\u_multiplier/K [3]),
    .ZN(\u_multiplier/_1365_ ));
 MUX2_X1 \u_multiplier/_2252_  (.A(\u_multiplier/_1025_ ),
    .B(\u_multiplier/_1029_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_1366_ ));
 MUX2_X1 \u_multiplier/_2253_  (.A(\u_multiplier/_1366_ ),
    .B(\u_multiplier/_1309_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_1367_ ));
 NOR2_X1 \u_multiplier/_2254_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_1367_ ),
    .ZN(\u_multiplier/_1368_ ));
 AOI21_X1 \u_multiplier/_2255_  (.A(\u_multiplier/_1368_ ),
    .B1(\u_multiplier/_1257_ ),
    .B2(\u_multiplier/code_x [2]),
    .ZN(\u_multiplier/_1369_ ));
 NOR2_X1 \u_multiplier/_2256_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_1369_ ),
    .ZN(\u_multiplier/_1370_ ));
 AOI21_X2 \u_multiplier/_2257_  (.A(\u_multiplier/_1370_ ),
    .B1(\u_multiplier/_1140_ ),
    .B2(\u_multiplier/code_x [3]),
    .ZN(\u_multiplier/_1371_ ));
 MUX2_X1 \u_multiplier/_2258_  (.A(\u_multiplier/_1027_ ),
    .B(\u_multiplier/_1031_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_1372_ ));
 MUX2_X1 \u_multiplier/_2259_  (.A(\u_multiplier/_1372_ ),
    .B(\u_multiplier/_1315_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_1373_ ));
 NOR2_X1 \u_multiplier/_2260_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_1373_ ),
    .ZN(\u_multiplier/_1374_ ));
 AOI21_X2 \u_multiplier/_2261_  (.A(\u_multiplier/_1374_ ),
    .B1(\u_multiplier/_1263_ ),
    .B2(\u_multiplier/code_y [2]),
    .ZN(\u_multiplier/_1375_ ));
 NAND2_X1 \u_multiplier/_2262_  (.A1(\u_multiplier/_0932_ ),
    .A2(\u_multiplier/_1375_ ),
    .ZN(\u_multiplier/_1376_ ));
 OAI21_X2 \u_multiplier/_2263_  (.A(\u_multiplier/_1376_ ),
    .B1(\u_multiplier/_1143_ ),
    .B2(\u_multiplier/_0932_ ),
    .ZN(\u_multiplier/_1377_ ));
 NAND2_X1 \u_multiplier/_2264_  (.A1(\u_multiplier/_1371_ ),
    .A2(\u_multiplier/_1377_ ),
    .ZN(\u_multiplier/_1378_ ));
 XOR2_X2 \u_multiplier/_2265_  (.A(\u_multiplier/_1371_ ),
    .B(\u_multiplier/_1377_ ),
    .Z(\u_multiplier/_1379_ ));
 NAND2_X1 \u_multiplier/_2266_  (.A1(\u_multiplier/_1365_ ),
    .A2(\u_multiplier/_1379_ ),
    .ZN(\u_multiplier/_1380_ ));
 XNOR2_X1 \u_multiplier/_2267_  (.A(\u_multiplier/_1365_ ),
    .B(\u_multiplier/_1379_ ),
    .ZN(\u_multiplier/_1381_ ));
 NOR2_X1 \u_multiplier/_2268_  (.A1(\u_multiplier/_1358_ ),
    .A2(\u_multiplier/_1381_ ),
    .ZN(\u_multiplier/_1382_ ));
 XOR2_X1 \u_multiplier/_2269_  (.A(\u_multiplier/_1358_ ),
    .B(\u_multiplier/_1381_ ),
    .Z(\u_multiplier/_1383_ ));
 INV_X1 \u_multiplier/_2270_  (.A(\u_multiplier/_1383_ ),
    .ZN(\u_multiplier/_1384_ ));
 OAI21_X1 \u_multiplier/_2271_  (.A(\u_multiplier/_1384_ ),
    .B1(\u_multiplier/_1354_ ),
    .B2(\u_multiplier/_1334_ ),
    .ZN(\u_multiplier/_1385_ ));
 NOR2_X1 \u_multiplier/_2272_  (.A1(\u_multiplier/_1356_ ),
    .A2(\u_multiplier/_1385_ ),
    .ZN(\u_multiplier/_1386_ ));
 AOI211_X2 \u_multiplier/_2273_  (.A(\u_multiplier/_1355_ ),
    .B(\u_multiplier/_1384_ ),
    .C1(\u_multiplier/_1330_ ),
    .C2(\u_multiplier/_1333_ ),
    .ZN(\u_multiplier/_1387_ ));
 NOR3_X1 \u_multiplier/_2274_  (.A1(\u_multiplier/_1334_ ),
    .A2(\u_multiplier/_1354_ ),
    .A3(\u_multiplier/_1384_ ),
    .ZN(\u_multiplier/_1388_ ));
 NOR4_X1 \u_multiplier/_2275_  (.A1(\u_multiplier/_0943_ ),
    .A2(\u_multiplier/_1386_ ),
    .A3(\u_multiplier/_1387_ ),
    .A4(\u_multiplier/_1388_ ),
    .ZN(product[11]));
 OR2_X1 \u_multiplier/_2276_  (.A1(\u_multiplier/_1382_ ),
    .A2(\u_multiplier/_1388_ ),
    .ZN(\u_multiplier/_1389_ ));
 NOR2_X1 \u_multiplier/_2277_  (.A1(\u_multiplier/_1387_ ),
    .A2(\u_multiplier/_1389_ ),
    .ZN(\u_multiplier/_1390_ ));
 NAND2_X1 \u_multiplier/_2278_  (.A1(\u_multiplier/_1378_ ),
    .A2(\u_multiplier/_1380_ ),
    .ZN(\u_multiplier/_1391_ ));
 MUX2_X1 \u_multiplier/_2279_  (.A(\u_multiplier/_1019_ ),
    .B(\u_multiplier/_1021_ ),
    .S(\u_multiplier/_1059_ ),
    .Z(\u_multiplier/_1392_ ));
 MUX2_X1 \u_multiplier/_2280_  (.A(\u_multiplier/_1359_ ),
    .B(\u_multiplier/_1392_ ),
    .S(\u_multiplier/_0937_ ),
    .Z(\u_multiplier/_1393_ ));
 MUX2_X1 \u_multiplier/_2281_  (.A(\u_multiplier/_1336_ ),
    .B(\u_multiplier/_1393_ ),
    .S(\u_multiplier/_0936_ ),
    .Z(\u_multiplier/_1394_ ));
 NAND2_X1 \u_multiplier/_2282_  (.A1(\u_multiplier/_0938_ ),
    .A2(\u_multiplier/_1394_ ),
    .ZN(\u_multiplier/_1395_ ));
 OAI21_X2 \u_multiplier/_2283_  (.A(\u_multiplier/_1395_ ),
    .B1(\u_multiplier/_1278_ ),
    .B2(\u_multiplier/_0938_ ),
    .ZN(\u_multiplier/_1396_ ));
 AND2_X1 \u_multiplier/_2284_  (.A1(\u_multiplier/K [3]),
    .A2(\u_multiplier/_1160_ ),
    .ZN(\u_multiplier/_1397_ ));
 AOI211_X2 \u_multiplier/_2285_  (.A(\u_multiplier/dec_out [12]),
    .B(\u_multiplier/_1397_ ),
    .C1(\u_multiplier/_1396_ ),
    .C2(\u_multiplier/_0939_ ),
    .ZN(\u_multiplier/_1398_ ));
 MUX2_X1 \u_multiplier/_2286_  (.A(\u_multiplier/_1019_ ),
    .B(\u_multiplier/_1025_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_1399_ ));
 MUX2_X1 \u_multiplier/_2287_  (.A(\u_multiplier/_1399_ ),
    .B(\u_multiplier/_1341_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_1400_ ));
 MUX2_X1 \u_multiplier/_2288_  (.A(\u_multiplier/_1283_ ),
    .B(\u_multiplier/_1400_ ),
    .S(\u_multiplier/_0935_ ),
    .Z(\u_multiplier/_1401_ ));
 NOR2_X1 \u_multiplier/_2289_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_1401_ ),
    .ZN(\u_multiplier/_1402_ ));
 AOI21_X2 \u_multiplier/_2290_  (.A(\u_multiplier/_1402_ ),
    .B1(\u_multiplier/_1166_ ),
    .B2(\u_multiplier/code_x [3]),
    .ZN(\u_multiplier/_1403_ ));
 MUX2_X1 \u_multiplier/_2291_  (.A(\u_multiplier/_1021_ ),
    .B(\u_multiplier/_1027_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_1404_ ));
 MUX2_X1 \u_multiplier/_2292_  (.A(\u_multiplier/_1404_ ),
    .B(\u_multiplier/_1346_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_1405_ ));
 MUX2_X1 \u_multiplier/_2293_  (.A(\u_multiplier/_1289_ ),
    .B(\u_multiplier/_1405_ ),
    .S(\u_multiplier/_0931_ ),
    .Z(\u_multiplier/_1406_ ));
 NAND2_X1 \u_multiplier/_2294_  (.A1(\u_multiplier/_0932_ ),
    .A2(\u_multiplier/_1406_ ),
    .ZN(\u_multiplier/_1407_ ));
 OAI21_X2 \u_multiplier/_2295_  (.A(\u_multiplier/_1407_ ),
    .B1(\u_multiplier/_1172_ ),
    .B2(\u_multiplier/_0932_ ),
    .ZN(\u_multiplier/_1408_ ));
 NAND2_X1 \u_multiplier/_2296_  (.A1(\u_multiplier/_1403_ ),
    .A2(\u_multiplier/_1408_ ),
    .ZN(\u_multiplier/_1409_ ));
 NOR2_X1 \u_multiplier/_2297_  (.A1(\u_multiplier/_1403_ ),
    .A2(\u_multiplier/_1408_ ),
    .ZN(\u_multiplier/_1410_ ));
 XOR2_X2 \u_multiplier/_2298_  (.A(\u_multiplier/_1403_ ),
    .B(\u_multiplier/_1408_ ),
    .Z(\u_multiplier/_1411_ ));
 XNOR2_X2 \u_multiplier/_2299_  (.A(\u_multiplier/_1398_ ),
    .B(\u_multiplier/_1411_ ),
    .ZN(\u_multiplier/_1412_ ));
 NAND2_X1 \u_multiplier/_2300_  (.A1(\u_multiplier/_1391_ ),
    .A2(\u_multiplier/_1412_ ),
    .ZN(\u_multiplier/_1413_ ));
 XNOR2_X2 \u_multiplier/_2301_  (.A(\u_multiplier/_1391_ ),
    .B(\u_multiplier/_1412_ ),
    .ZN(\u_multiplier/_1414_ ));
 INV_X1 \u_multiplier/_2302_  (.A(\u_multiplier/_1414_ ),
    .ZN(\u_multiplier/_1415_ ));
 NOR2_X1 \u_multiplier/_2303_  (.A1(\u_multiplier/_1390_ ),
    .A2(\u_multiplier/_1414_ ),
    .ZN(\u_multiplier/_1416_ ));
 NOR3_X1 \u_multiplier/_2304_  (.A1(\u_multiplier/_1387_ ),
    .A2(\u_multiplier/_1389_ ),
    .A3(\u_multiplier/_1415_ ),
    .ZN(\u_multiplier/_1417_ ));
 NOR3_X1 \u_multiplier/_2305_  (.A1(\u_multiplier/_0943_ ),
    .A2(\u_multiplier/_1416_ ),
    .A3(\u_multiplier/_1417_ ),
    .ZN(product[12]));
 OAI21_X1 \u_multiplier/_2306_  (.A(\u_multiplier/_1409_ ),
    .B1(\u_multiplier/_1410_ ),
    .B2(\u_multiplier/_1398_ ),
    .ZN(\u_multiplier/_1418_ ));
 MUX2_X1 \u_multiplier/_2307_  (.A(\u_multiplier/_1015_ ),
    .B(\u_multiplier/_1016_ ),
    .S(\u_multiplier/_1059_ ),
    .Z(\u_multiplier/_1419_ ));
 MUX2_X1 \u_multiplier/_2308_  (.A(\u_multiplier/_1392_ ),
    .B(\u_multiplier/_1419_ ),
    .S(\u_multiplier/_0937_ ),
    .Z(\u_multiplier/_1420_ ));
 MUX2_X1 \u_multiplier/_2309_  (.A(\u_multiplier/_1360_ ),
    .B(\u_multiplier/_1420_ ),
    .S(\u_multiplier/_0936_ ),
    .Z(\u_multiplier/_1421_ ));
 NAND2_X1 \u_multiplier/_2310_  (.A1(\u_multiplier/_0938_ ),
    .A2(\u_multiplier/_1421_ ),
    .ZN(\u_multiplier/_1422_ ));
 OAI21_X1 \u_multiplier/_2311_  (.A(\u_multiplier/_1422_ ),
    .B1(\u_multiplier/_1304_ ),
    .B2(\u_multiplier/_0938_ ),
    .ZN(\u_multiplier/_1423_ ));
 AND2_X1 \u_multiplier/_2312_  (.A1(\u_multiplier/_0939_ ),
    .A2(\u_multiplier/_1423_ ),
    .ZN(\u_multiplier/_1424_ ));
 AOI211_X2 \u_multiplier/_2313_  (.A(\u_multiplier/dec_out [13]),
    .B(\u_multiplier/_1424_ ),
    .C1(\u_multiplier/_1192_ ),
    .C2(\u_multiplier/K [3]),
    .ZN(\u_multiplier/_1425_ ));
 MUX2_X1 \u_multiplier/_2314_  (.A(\u_multiplier/_1015_ ),
    .B(\u_multiplier/_1019_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_1426_ ));
 MUX2_X1 \u_multiplier/_2315_  (.A(\u_multiplier/_1426_ ),
    .B(\u_multiplier/_1366_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_1427_ ));
 OR2_X1 \u_multiplier/_2316_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_1427_ ),
    .ZN(\u_multiplier/_1428_ ));
 OAI21_X1 \u_multiplier/_2317_  (.A(\u_multiplier/_1428_ ),
    .B1(\u_multiplier/_1310_ ),
    .B2(\u_multiplier/_0935_ ),
    .ZN(\u_multiplier/_1429_ ));
 MUX2_X1 \u_multiplier/_2318_  (.A(\u_multiplier/_1197_ ),
    .B(\u_multiplier/_1429_ ),
    .S(\u_multiplier/_0933_ ),
    .Z(\u_multiplier/_1430_ ));
 MUX2_X1 \u_multiplier/_2319_  (.A(\u_multiplier/_1016_ ),
    .B(\u_multiplier/_1021_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_1431_ ));
 MUX2_X1 \u_multiplier/_2320_  (.A(\u_multiplier/_1431_ ),
    .B(\u_multiplier/_1372_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_1432_ ));
 OR2_X1 \u_multiplier/_2321_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_1432_ ),
    .ZN(\u_multiplier/_1433_ ));
 OAI21_X1 \u_multiplier/_2322_  (.A(\u_multiplier/_1433_ ),
    .B1(\u_multiplier/_1317_ ),
    .B2(\u_multiplier/_0931_ ),
    .ZN(\u_multiplier/_1434_ ));
 MUX2_X1 \u_multiplier/_2323_  (.A(\u_multiplier/_1201_ ),
    .B(\u_multiplier/_1434_ ),
    .S(\u_multiplier/_0932_ ),
    .Z(\u_multiplier/_1435_ ));
 OR2_X1 \u_multiplier/_2324_  (.A1(\u_multiplier/_1430_ ),
    .A2(\u_multiplier/_1435_ ),
    .ZN(\u_multiplier/_1436_ ));
 XNOR2_X2 \u_multiplier/_2325_  (.A(\u_multiplier/_1430_ ),
    .B(\u_multiplier/_1435_ ),
    .ZN(\u_multiplier/_1437_ ));
 XOR2_X2 \u_multiplier/_2326_  (.A(\u_multiplier/_1425_ ),
    .B(\u_multiplier/_1437_ ),
    .Z(\u_multiplier/_1438_ ));
 NAND2_X1 \u_multiplier/_2327_  (.A1(\u_multiplier/_1418_ ),
    .A2(\u_multiplier/_1438_ ),
    .ZN(\u_multiplier/_1439_ ));
 XNOR2_X1 \u_multiplier/_2328_  (.A(\u_multiplier/_1418_ ),
    .B(\u_multiplier/_1438_ ),
    .ZN(\u_multiplier/_1440_ ));
 INV_X1 \u_multiplier/_2329_  (.A(\u_multiplier/_1440_ ),
    .ZN(\u_multiplier/_1441_ ));
 OAI211_X1 \u_multiplier/_2330_  (.A(\u_multiplier/_1413_ ),
    .B(\u_multiplier/_1440_ ),
    .C1(\u_multiplier/_1414_ ),
    .C2(\u_multiplier/_1390_ ),
    .ZN(\u_multiplier/_1442_ ));
 OAI211_X2 \u_multiplier/_2331_  (.A(\u_multiplier/_1415_ ),
    .B(\u_multiplier/_1441_ ),
    .C1(\u_multiplier/_1387_ ),
    .C2(\u_multiplier/_1389_ ),
    .ZN(\u_multiplier/_1443_ ));
 OR2_X1 \u_multiplier/_2332_  (.A1(\u_multiplier/_1413_ ),
    .A2(\u_multiplier/_1440_ ),
    .ZN(\u_multiplier/_1444_ ));
 AND4_X1 \u_multiplier/_2333_  (.A1(\u_multiplier/_1739_ ),
    .A2(\u_multiplier/_1442_ ),
    .A3(\u_multiplier/_1443_ ),
    .A4(\u_multiplier/_1444_ ),
    .ZN(product[13]));
 AND2_X1 \u_multiplier/_2334_  (.A1(\u_multiplier/_1439_ ),
    .A2(\u_multiplier/_1444_ ),
    .ZN(\u_multiplier/_1445_ ));
 AND2_X1 \u_multiplier/_2335_  (.A1(\u_multiplier/_1443_ ),
    .A2(\u_multiplier/_1445_ ),
    .ZN(\u_multiplier/_1446_ ));
 OAI21_X2 \u_multiplier/_2336_  (.A(\u_multiplier/_1436_ ),
    .B1(\u_multiplier/_1437_ ),
    .B2(\u_multiplier/_1425_ ),
    .ZN(\u_multiplier/_1447_ ));
 NOR2_X1 \u_multiplier/_2337_  (.A1(\u_multiplier/_1039_ ),
    .A2(\u_multiplier/_1056_ ),
    .ZN(\u_multiplier/_1448_ ));
 NOR2_X1 \u_multiplier/_2338_  (.A1(\u_multiplier/_1042_ ),
    .A2(\u_multiplier/_1448_ ),
    .ZN(\u_multiplier/_1449_ ));
 MUX2_X1 \u_multiplier/_2339_  (.A(\u_multiplier/_1419_ ),
    .B(\u_multiplier/_1449_ ),
    .S(\u_multiplier/_0937_ ),
    .Z(\u_multiplier/_1450_ ));
 MUX2_X1 \u_multiplier/_2340_  (.A(\u_multiplier/_1393_ ),
    .B(\u_multiplier/_1450_ ),
    .S(\u_multiplier/_0936_ ),
    .Z(\u_multiplier/_1451_ ));
 MUX2_X1 \u_multiplier/_2341_  (.A(\u_multiplier/_1337_ ),
    .B(\u_multiplier/_1451_ ),
    .S(\u_multiplier/_0938_ ),
    .Z(\u_multiplier/_1452_ ));
 AND2_X1 \u_multiplier/_2342_  (.A1(\u_multiplier/_0939_ ),
    .A2(\u_multiplier/_1452_ ),
    .ZN(\u_multiplier/_1453_ ));
 AOI211_X2 \u_multiplier/_2343_  (.A(\u_multiplier/dec_out [14]),
    .B(\u_multiplier/_1453_ ),
    .C1(\u_multiplier/_1219_ ),
    .C2(\u_multiplier/K [3]),
    .ZN(\u_multiplier/_1454_ ));
 MUX2_X1 \u_multiplier/_2344_  (.A(\u_multiplier/_1015_ ),
    .B(\u_multiplier/_1039_ ),
    .S(\u_multiplier/_0934_ ),
    .Z(\u_multiplier/_1455_ ));
 MUX2_X1 \u_multiplier/_2345_  (.A(\u_multiplier/_1455_ ),
    .B(\u_multiplier/_1399_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_1456_ ));
 MUX2_X1 \u_multiplier/_2346_  (.A(\u_multiplier/_1342_ ),
    .B(\u_multiplier/_1456_ ),
    .S(\u_multiplier/_0935_ ),
    .Z(\u_multiplier/_1457_ ));
 NOR2_X1 \u_multiplier/_2347_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_1457_ ),
    .ZN(\u_multiplier/_1458_ ));
 AOI21_X2 \u_multiplier/_2348_  (.A(\u_multiplier/_1458_ ),
    .B1(\u_multiplier/_1225_ ),
    .B2(\u_multiplier/code_x [3]),
    .ZN(\u_multiplier/_1459_ ));
 MUX2_X1 \u_multiplier/_2349_  (.A(\u_multiplier/_1016_ ),
    .B(\u_multiplier/_1041_ ),
    .S(\u_multiplier/_0930_ ),
    .Z(\u_multiplier/_1460_ ));
 MUX2_X1 \u_multiplier/_2350_  (.A(\u_multiplier/_1460_ ),
    .B(\u_multiplier/_1404_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_1461_ ));
 MUX2_X1 \u_multiplier/_2351_  (.A(\u_multiplier/_1347_ ),
    .B(\u_multiplier/_1461_ ),
    .S(\u_multiplier/_0931_ ),
    .Z(\u_multiplier/_1462_ ));
 NOR2_X1 \u_multiplier/_2352_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_1462_ ),
    .ZN(\u_multiplier/_1463_ ));
 AOI21_X2 \u_multiplier/_2353_  (.A(\u_multiplier/_1463_ ),
    .B1(\u_multiplier/_1231_ ),
    .B2(\u_multiplier/code_y [3]),
    .ZN(\u_multiplier/_1464_ ));
 NAND2_X1 \u_multiplier/_2354_  (.A1(\u_multiplier/_1459_ ),
    .A2(\u_multiplier/_1464_ ),
    .ZN(\u_multiplier/_1465_ ));
 XNOR2_X2 \u_multiplier/_2355_  (.A(\u_multiplier/_1459_ ),
    .B(\u_multiplier/_1464_ ),
    .ZN(\u_multiplier/_1466_ ));
 XOR2_X2 \u_multiplier/_2356_  (.A(\u_multiplier/_1454_ ),
    .B(\u_multiplier/_1466_ ),
    .Z(\u_multiplier/_1467_ ));
 NAND2_X1 \u_multiplier/_2357_  (.A1(\u_multiplier/_1447_ ),
    .A2(\u_multiplier/_1467_ ),
    .ZN(\u_multiplier/_1468_ ));
 XNOR2_X2 \u_multiplier/_2358_  (.A(\u_multiplier/_1447_ ),
    .B(\u_multiplier/_1467_ ),
    .ZN(\u_multiplier/_1469_ ));
 AOI21_X1 \u_multiplier/_2359_  (.A(\u_multiplier/_0943_ ),
    .B1(\u_multiplier/_1446_ ),
    .B2(\u_multiplier/_1469_ ),
    .ZN(\u_multiplier/_1470_ ));
 OAI21_X1 \u_multiplier/_2360_  (.A(\u_multiplier/_1470_ ),
    .B1(\u_multiplier/_1469_ ),
    .B2(\u_multiplier/_1446_ ),
    .ZN(\u_multiplier/_1471_ ));
 INV_X1 \u_multiplier/_2361_  (.A(\u_multiplier/_1471_ ),
    .ZN(product[14]));
 OAI21_X1 \u_multiplier/_2362_  (.A(\u_multiplier/_1465_ ),
    .B1(\u_multiplier/_1466_ ),
    .B2(\u_multiplier/_1454_ ),
    .ZN(\u_multiplier/_1472_ ));
 NOR3_X2 \u_multiplier/_2363_  (.A1(\u_multiplier/_0937_ ),
    .A2(\u_multiplier/_1042_ ),
    .A3(\u_multiplier/_1448_ ),
    .ZN(\u_multiplier/_1473_ ));
 MUX2_X1 \u_multiplier/_2364_  (.A(\u_multiplier/_1420_ ),
    .B(\u_multiplier/_1473_ ),
    .S(\u_multiplier/_0936_ ),
    .Z(\u_multiplier/_1474_ ));
 NAND2_X1 \u_multiplier/_2365_  (.A1(\u_multiplier/_0938_ ),
    .A2(\u_multiplier/_1474_ ),
    .ZN(\u_multiplier/_1475_ ));
 OAI21_X2 \u_multiplier/_2366_  (.A(\u_multiplier/_1475_ ),
    .B1(\u_multiplier/_1362_ ),
    .B2(\u_multiplier/_0938_ ),
    .ZN(\u_multiplier/_1476_ ));
 NOR2_X1 \u_multiplier/_2367_  (.A1(\u_multiplier/K [3]),
    .A2(\u_multiplier/_1476_ ),
    .ZN(\u_multiplier/_1477_ ));
 AOI21_X1 \u_multiplier/_2368_  (.A(\u_multiplier/_1477_ ),
    .B1(\u_multiplier/_1252_ ),
    .B2(\u_multiplier/K [3]),
    .ZN(\u_multiplier/_1478_ ));
 NOR2_X1 \u_multiplier/_2369_  (.A1(\u_multiplier/dec_out [15]),
    .A2(\u_multiplier/_1478_ ),
    .ZN(\u_multiplier/_1479_ ));
 NOR3_X1 \u_multiplier/_2370_  (.A1(\u_multiplier/_0934_ ),
    .A2(\u_multiplier/code_x [1]),
    .A3(\u_multiplier/_1040_ ),
    .ZN(\u_multiplier/_1480_ ));
 AOI21_X2 \u_multiplier/_2371_  (.A(\u_multiplier/_1480_ ),
    .B1(\u_multiplier/_1426_ ),
    .B2(\u_multiplier/code_x [1]),
    .ZN(\u_multiplier/_1481_ ));
 NOR2_X1 \u_multiplier/_2372_  (.A1(\u_multiplier/_0935_ ),
    .A2(\u_multiplier/_1367_ ),
    .ZN(\u_multiplier/_1482_ ));
 AOI21_X2 \u_multiplier/_2373_  (.A(\u_multiplier/_1482_ ),
    .B1(\u_multiplier/_1481_ ),
    .B2(\u_multiplier/_0935_ ),
    .ZN(\u_multiplier/_1483_ ));
 NAND2_X1 \u_multiplier/_2374_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_1258_ ),
    .ZN(\u_multiplier/_1484_ ));
 OAI21_X2 \u_multiplier/_2375_  (.A(\u_multiplier/_1484_ ),
    .B1(\u_multiplier/_1483_ ),
    .B2(\u_multiplier/code_x [3]),
    .ZN(\u_multiplier/_1485_ ));
 NOR3_X1 \u_multiplier/_2376_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_0930_ ),
    .A3(\u_multiplier/_1042_ ),
    .ZN(\u_multiplier/_1486_ ));
 AOI21_X2 \u_multiplier/_2377_  (.A(\u_multiplier/_1486_ ),
    .B1(\u_multiplier/_1431_ ),
    .B2(\u_multiplier/code_y [1]),
    .ZN(\u_multiplier/_1487_ ));
 NOR2_X1 \u_multiplier/_2378_  (.A1(\u_multiplier/_0931_ ),
    .A2(\u_multiplier/_1373_ ),
    .ZN(\u_multiplier/_1488_ ));
 AOI21_X4 \u_multiplier/_2379_  (.A(\u_multiplier/_1488_ ),
    .B1(\u_multiplier/_1487_ ),
    .B2(\u_multiplier/_0931_ ),
    .ZN(\u_multiplier/_1489_ ));
 NAND2_X1 \u_multiplier/_2380_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_1264_ ),
    .ZN(\u_multiplier/_1490_ ));
 OAI21_X2 \u_multiplier/_2381_  (.A(\u_multiplier/_1490_ ),
    .B1(\u_multiplier/_1489_ ),
    .B2(\u_multiplier/code_y [3]),
    .ZN(\u_multiplier/_1491_ ));
 XOR2_X2 \u_multiplier/_2382_  (.A(\u_multiplier/_1485_ ),
    .B(\u_multiplier/_1491_ ),
    .Z(\u_multiplier/_1492_ ));
 OAI21_X1 \u_multiplier/_2383_  (.A(\u_multiplier/_1492_ ),
    .B1(\u_multiplier/_1478_ ),
    .B2(\u_multiplier/dec_out [15]),
    .ZN(\u_multiplier/_1493_ ));
 XNOR2_X2 \u_multiplier/_2384_  (.A(\u_multiplier/_1479_ ),
    .B(\u_multiplier/_1492_ ),
    .ZN(\u_multiplier/_1494_ ));
 NAND2_X1 \u_multiplier/_2385_  (.A1(\u_multiplier/_1472_ ),
    .A2(\u_multiplier/_1494_ ),
    .ZN(\u_multiplier/_1495_ ));
 XNOR2_X2 \u_multiplier/_2386_  (.A(\u_multiplier/_1472_ ),
    .B(\u_multiplier/_1494_ ),
    .ZN(\u_multiplier/_1496_ ));
 OAI211_X1 \u_multiplier/_2387_  (.A(\u_multiplier/_1468_ ),
    .B(\u_multiplier/_1496_ ),
    .C1(\u_multiplier/_1469_ ),
    .C2(\u_multiplier/_1446_ ),
    .ZN(\u_multiplier/_1497_ ));
 INV_X1 \u_multiplier/_2388_  (.A(\u_multiplier/_1497_ ),
    .ZN(\u_multiplier/_1498_ ));
 AOI211_X2 \u_multiplier/_2389_  (.A(\u_multiplier/_1469_ ),
    .B(\u_multiplier/_1496_ ),
    .C1(\u_multiplier/_1443_ ),
    .C2(\u_multiplier/_1445_ ),
    .ZN(\u_multiplier/_1499_ ));
 OAI21_X1 \u_multiplier/_2390_  (.A(\u_multiplier/_1739_ ),
    .B1(\u_multiplier/_1468_ ),
    .B2(\u_multiplier/_1496_ ),
    .ZN(\u_multiplier/_1500_ ));
 NOR3_X1 \u_multiplier/_2391_  (.A1(\u_multiplier/_1498_ ),
    .A2(\u_multiplier/_1499_ ),
    .A3(\u_multiplier/_1500_ ),
    .ZN(product[15]));
 OAI21_X2 \u_multiplier/_2392_  (.A(\u_multiplier/_1495_ ),
    .B1(\u_multiplier/_1496_ ),
    .B2(\u_multiplier/_1468_ ),
    .ZN(\u_multiplier/_1501_ ));
 NOR2_X1 \u_multiplier/_2393_  (.A1(\u_multiplier/_1499_ ),
    .A2(\u_multiplier/_1501_ ),
    .ZN(\u_multiplier/_1502_ ));
 OAI21_X2 \u_multiplier/_2394_  (.A(\u_multiplier/_1493_ ),
    .B1(\u_multiplier/_1491_ ),
    .B2(\u_multiplier/_1485_ ),
    .ZN(\u_multiplier/_1503_ ));
 AND2_X1 \u_multiplier/_2395_  (.A1(\u_multiplier/K [1]),
    .A2(\u_multiplier/_1450_ ),
    .ZN(\u_multiplier/_1504_ ));
 MUX2_X1 \u_multiplier/_2396_  (.A(\u_multiplier/_1394_ ),
    .B(\u_multiplier/_1504_ ),
    .S(\u_multiplier/_0938_ ),
    .Z(\u_multiplier/_1505_ ));
 NOR2_X1 \u_multiplier/_2397_  (.A1(\u_multiplier/K [3]),
    .A2(\u_multiplier/_1505_ ),
    .ZN(\u_multiplier/_1506_ ));
 AOI21_X1 \u_multiplier/_2398_  (.A(\u_multiplier/_1506_ ),
    .B1(\u_multiplier/_1279_ ),
    .B2(\u_multiplier/K [3]),
    .ZN(\u_multiplier/_1507_ ));
 AND2_X1 \u_multiplier/_2399_  (.A1(\u_multiplier/code_x [1]),
    .A2(\u_multiplier/_1455_ ),
    .ZN(\u_multiplier/_1508_ ));
 MUX2_X1 \u_multiplier/_2400_  (.A(\u_multiplier/_1400_ ),
    .B(\u_multiplier/_1508_ ),
    .S(\u_multiplier/_0935_ ),
    .Z(\u_multiplier/_1509_ ));
 OR2_X1 \u_multiplier/_2401_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_1509_ ),
    .ZN(\u_multiplier/_1510_ ));
 OAI21_X1 \u_multiplier/_2402_  (.A(\u_multiplier/_1510_ ),
    .B1(\u_multiplier/_1284_ ),
    .B2(\u_multiplier/_0933_ ),
    .ZN(\u_multiplier/_1511_ ));
 AND2_X1 \u_multiplier/_2403_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_1460_ ),
    .ZN(\u_multiplier/_1512_ ));
 MUX2_X1 \u_multiplier/_2404_  (.A(\u_multiplier/_1405_ ),
    .B(\u_multiplier/_1512_ ),
    .S(\u_multiplier/_0931_ ),
    .Z(\u_multiplier/_1513_ ));
 NAND2_X1 \u_multiplier/_2405_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_1291_ ),
    .ZN(\u_multiplier/_1514_ ));
 OAI21_X1 \u_multiplier/_2406_  (.A(\u_multiplier/_1514_ ),
    .B1(\u_multiplier/_1513_ ),
    .B2(\u_multiplier/code_y [3]),
    .ZN(\u_multiplier/_1515_ ));
 XOR2_X1 \u_multiplier/_2407_  (.A(\u_multiplier/_1511_ ),
    .B(\u_multiplier/_1515_ ),
    .Z(\u_multiplier/_1516_ ));
 OAI21_X1 \u_multiplier/_2408_  (.A(\u_multiplier/_1516_ ),
    .B1(\u_multiplier/_1507_ ),
    .B2(\u_multiplier/dec_out [16]),
    .ZN(\u_multiplier/_1517_ ));
 OR3_X1 \u_multiplier/_2409_  (.A1(\u_multiplier/dec_out [16]),
    .A2(\u_multiplier/_1507_ ),
    .A3(\u_multiplier/_1516_ ),
    .ZN(\u_multiplier/_1518_ ));
 AND2_X1 \u_multiplier/_2410_  (.A1(\u_multiplier/_1517_ ),
    .A2(\u_multiplier/_1518_ ),
    .ZN(\u_multiplier/_1519_ ));
 NAND2_X1 \u_multiplier/_2411_  (.A1(\u_multiplier/_1503_ ),
    .A2(\u_multiplier/_1519_ ),
    .ZN(\u_multiplier/_1520_ ));
 XNOR2_X2 \u_multiplier/_2412_  (.A(\u_multiplier/_1503_ ),
    .B(\u_multiplier/_1519_ ),
    .ZN(\u_multiplier/_1521_ ));
 INV_X1 \u_multiplier/_2413_  (.A(\u_multiplier/_1521_ ),
    .ZN(\u_multiplier/_1522_ ));
 NOR2_X1 \u_multiplier/_2414_  (.A1(\u_multiplier/_1502_ ),
    .A2(\u_multiplier/_1521_ ),
    .ZN(\u_multiplier/_1523_ ));
 NOR3_X1 \u_multiplier/_2415_  (.A1(\u_multiplier/_1499_ ),
    .A2(\u_multiplier/_1501_ ),
    .A3(\u_multiplier/_1522_ ),
    .ZN(\u_multiplier/_1524_ ));
 NOR3_X1 \u_multiplier/_2416_  (.A1(\u_multiplier/_0943_ ),
    .A2(\u_multiplier/_1523_ ),
    .A3(\u_multiplier/_1524_ ),
    .ZN(product[16]));
 OAI21_X2 \u_multiplier/_2417_  (.A(\u_multiplier/_1517_ ),
    .B1(\u_multiplier/_1515_ ),
    .B2(\u_multiplier/_1511_ ),
    .ZN(\u_multiplier/_1525_ ));
 NAND3_X1 \u_multiplier/_2418_  (.A1(\u_multiplier/K [1]),
    .A2(\u_multiplier/_0938_ ),
    .A3(\u_multiplier/_1473_ ),
    .ZN(\u_multiplier/_1526_ ));
 NAND2_X1 \u_multiplier/_2419_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/_1421_ ),
    .ZN(\u_multiplier/_1527_ ));
 NAND2_X2 \u_multiplier/_2420_  (.A1(\u_multiplier/_1526_ ),
    .A2(\u_multiplier/_1527_ ),
    .ZN(\u_multiplier/_1528_ ));
 NOR2_X1 \u_multiplier/_2421_  (.A1(\u_multiplier/_0939_ ),
    .A2(\u_multiplier/_1306_ ),
    .ZN(\u_multiplier/_1529_ ));
 AOI211_X2 \u_multiplier/_2422_  (.A(\u_multiplier/dec_out [17]),
    .B(\u_multiplier/_1529_ ),
    .C1(\u_multiplier/_1528_ ),
    .C2(\u_multiplier/_0939_ ),
    .ZN(\u_multiplier/_1530_ ));
 INV_X1 \u_multiplier/_2423_  (.A(\u_multiplier/_1530_ ),
    .ZN(\u_multiplier/_1531_ ));
 NAND3_X2 \u_multiplier/_2424_  (.A1(\u_multiplier/code_x [0]),
    .A2(\u_multiplier/code_x [1]),
    .A3(\u_multiplier/_1039_ ),
    .ZN(\u_multiplier/_1532_ ));
 NOR2_X1 \u_multiplier/_2425_  (.A1(\u_multiplier/_0935_ ),
    .A2(\u_multiplier/_1427_ ),
    .ZN(\u_multiplier/_1533_ ));
 AOI21_X2 \u_multiplier/_2426_  (.A(\u_multiplier/_1533_ ),
    .B1(\u_multiplier/_1532_ ),
    .B2(\u_multiplier/_0935_ ),
    .ZN(\u_multiplier/_1534_ ));
 OR2_X1 \u_multiplier/_2427_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_1534_ ),
    .ZN(\u_multiplier/_1535_ ));
 OAI21_X2 \u_multiplier/_2428_  (.A(\u_multiplier/_1535_ ),
    .B1(\u_multiplier/_1312_ ),
    .B2(\u_multiplier/_0933_ ),
    .ZN(\u_multiplier/_1536_ ));
 NAND3_X1 \u_multiplier/_2429_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/code_y [0]),
    .A3(\u_multiplier/_1041_ ),
    .ZN(\u_multiplier/_1537_ ));
 NOR2_X1 \u_multiplier/_2430_  (.A1(\u_multiplier/_0931_ ),
    .A2(\u_multiplier/_1432_ ),
    .ZN(\u_multiplier/_1538_ ));
 AOI21_X2 \u_multiplier/_2431_  (.A(\u_multiplier/_1538_ ),
    .B1(\u_multiplier/_1537_ ),
    .B2(\u_multiplier/_0931_ ),
    .ZN(\u_multiplier/_1539_ ));
 OR2_X1 \u_multiplier/_2432_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_1539_ ),
    .ZN(\u_multiplier/_1540_ ));
 OAI21_X2 \u_multiplier/_2433_  (.A(\u_multiplier/_1540_ ),
    .B1(\u_multiplier/_1319_ ),
    .B2(\u_multiplier/_0932_ ),
    .ZN(\u_multiplier/_1541_ ));
 NOR2_X1 \u_multiplier/_2434_  (.A1(\u_multiplier/_1536_ ),
    .A2(\u_multiplier/_1541_ ),
    .ZN(\u_multiplier/_1542_ ));
 XOR2_X2 \u_multiplier/_2435_  (.A(\u_multiplier/_1536_ ),
    .B(\u_multiplier/_1541_ ),
    .Z(\u_multiplier/_1543_ ));
 XNOR2_X2 \u_multiplier/_2436_  (.A(\u_multiplier/_1530_ ),
    .B(\u_multiplier/_1543_ ),
    .ZN(\u_multiplier/_1544_ ));
 XNOR2_X2 \u_multiplier/_2437_  (.A(\u_multiplier/_1525_ ),
    .B(\u_multiplier/_1544_ ),
    .ZN(\u_multiplier/_1545_ ));
 INV_X1 \u_multiplier/_2438_  (.A(\u_multiplier/_1545_ ),
    .ZN(\u_multiplier/_1546_ ));
 OAI211_X2 \u_multiplier/_2439_  (.A(\u_multiplier/_1522_ ),
    .B(\u_multiplier/_1546_ ),
    .C1(\u_multiplier/_1499_ ),
    .C2(\u_multiplier/_1501_ ),
    .ZN(\u_multiplier/_1547_ ));
 OAI211_X1 \u_multiplier/_2440_  (.A(\u_multiplier/_1520_ ),
    .B(\u_multiplier/_1545_ ),
    .C1(\u_multiplier/_1521_ ),
    .C2(\u_multiplier/_1502_ ),
    .ZN(\u_multiplier/_1548_ ));
 NOR2_X1 \u_multiplier/_2441_  (.A1(\u_multiplier/_1520_ ),
    .A2(\u_multiplier/_1545_ ),
    .ZN(\u_multiplier/_1549_ ));
 NOR2_X1 \u_multiplier/_2442_  (.A1(\u_multiplier/_0943_ ),
    .A2(\u_multiplier/_1549_ ),
    .ZN(\u_multiplier/_1550_ ));
 AND3_X1 \u_multiplier/_2443_  (.A1(\u_multiplier/_1547_ ),
    .A2(\u_multiplier/_1548_ ),
    .A3(\u_multiplier/_1550_ ),
    .ZN(product[17]));
 AOI21_X2 \u_multiplier/_2444_  (.A(\u_multiplier/_1549_ ),
    .B1(\u_multiplier/_1544_ ),
    .B2(\u_multiplier/_1525_ ),
    .ZN(\u_multiplier/_1551_ ));
 AND2_X1 \u_multiplier/_2445_  (.A1(\u_multiplier/_1547_ ),
    .A2(\u_multiplier/_1551_ ),
    .ZN(\u_multiplier/_1552_ ));
 AOI21_X2 \u_multiplier/_2446_  (.A(\u_multiplier/_1542_ ),
    .B1(\u_multiplier/_1543_ ),
    .B2(\u_multiplier/_1531_ ),
    .ZN(\u_multiplier/_1553_ ));
 NAND2_X2 \u_multiplier/_2447_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/_1451_ ),
    .ZN(\u_multiplier/_1554_ ));
 AOI21_X1 \u_multiplier/_2448_  (.A(\u_multiplier/dec_out [18]),
    .B1(\u_multiplier/_1338_ ),
    .B2(\u_multiplier/K [3]),
    .ZN(\u_multiplier/_1555_ ));
 OAI21_X2 \u_multiplier/_2449_  (.A(\u_multiplier/_1555_ ),
    .B1(\u_multiplier/_1554_ ),
    .B2(\u_multiplier/K [3]),
    .ZN(\u_multiplier/_1556_ ));
 AND2_X1 \u_multiplier/_2450_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_1456_ ),
    .ZN(\u_multiplier/_1557_ ));
 NAND2_X1 \u_multiplier/_2451_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_1344_ ),
    .ZN(\u_multiplier/_1558_ ));
 OAI21_X2 \u_multiplier/_2452_  (.A(\u_multiplier/_1558_ ),
    .B1(\u_multiplier/_1557_ ),
    .B2(\u_multiplier/code_x [3]),
    .ZN(\u_multiplier/_1559_ ));
 AND2_X1 \u_multiplier/_2453_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_1461_ ),
    .ZN(\u_multiplier/_1560_ ));
 NAND2_X1 \u_multiplier/_2454_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_1349_ ),
    .ZN(\u_multiplier/_1561_ ));
 OAI21_X2 \u_multiplier/_2455_  (.A(\u_multiplier/_1561_ ),
    .B1(\u_multiplier/_1560_ ),
    .B2(\u_multiplier/code_y [3]),
    .ZN(\u_multiplier/_1562_ ));
 NOR2_X1 \u_multiplier/_2456_  (.A1(\u_multiplier/_1559_ ),
    .A2(\u_multiplier/_1562_ ),
    .ZN(\u_multiplier/_1563_ ));
 XOR2_X2 \u_multiplier/_2457_  (.A(\u_multiplier/_1559_ ),
    .B(\u_multiplier/_1562_ ),
    .Z(\u_multiplier/_1564_ ));
 XNOR2_X2 \u_multiplier/_2458_  (.A(\u_multiplier/_1556_ ),
    .B(\u_multiplier/_1564_ ),
    .ZN(\u_multiplier/_1565_ ));
 NOR2_X1 \u_multiplier/_2459_  (.A1(\u_multiplier/_1553_ ),
    .A2(\u_multiplier/_1565_ ),
    .ZN(\u_multiplier/_1566_ ));
 XNOR2_X2 \u_multiplier/_2460_  (.A(\u_multiplier/_1553_ ),
    .B(\u_multiplier/_1565_ ),
    .ZN(\u_multiplier/_1567_ ));
 NOR2_X1 \u_multiplier/_2461_  (.A1(\u_multiplier/_1552_ ),
    .A2(\u_multiplier/_1567_ ),
    .ZN(\u_multiplier/_1568_ ));
 AND2_X1 \u_multiplier/_2462_  (.A1(\u_multiplier/_1552_ ),
    .A2(\u_multiplier/_1567_ ),
    .ZN(\u_multiplier/_1569_ ));
 NOR3_X1 \u_multiplier/_2463_  (.A1(\u_multiplier/_0943_ ),
    .A2(\u_multiplier/_1568_ ),
    .A3(\u_multiplier/_1569_ ),
    .ZN(product[18]));
 AOI21_X2 \u_multiplier/_2464_  (.A(\u_multiplier/_1563_ ),
    .B1(\u_multiplier/_1564_ ),
    .B2(\u_multiplier/_1556_ ),
    .ZN(\u_multiplier/_1570_ ));
 OR2_X1 \u_multiplier/_2465_  (.A1(\u_multiplier/_0939_ ),
    .A2(\u_multiplier/_1363_ ),
    .ZN(\u_multiplier/_1571_ ));
 AND2_X1 \u_multiplier/_2466_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/_1474_ ),
    .ZN(\u_multiplier/_1572_ ));
 AOI21_X1 \u_multiplier/_2467_  (.A(\u_multiplier/dec_out [19]),
    .B1(\u_multiplier/_1572_ ),
    .B2(\u_multiplier/_0939_ ),
    .ZN(\u_multiplier/_1573_ ));
 NOR2_X1 \u_multiplier/_2468_  (.A1(\u_multiplier/_0935_ ),
    .A2(\u_multiplier/_1481_ ),
    .ZN(\u_multiplier/_1574_ ));
 MUX2_X1 \u_multiplier/_2469_  (.A(\u_multiplier/_1369_ ),
    .B(\u_multiplier/_1574_ ),
    .S(\u_multiplier/_0933_ ),
    .Z(\u_multiplier/_1575_ ));
 NOR2_X1 \u_multiplier/_2470_  (.A1(\u_multiplier/_0931_ ),
    .A2(\u_multiplier/_1487_ ),
    .ZN(\u_multiplier/_1576_ ));
 MUX2_X1 \u_multiplier/_2471_  (.A(\u_multiplier/_1375_ ),
    .B(\u_multiplier/_1576_ ),
    .S(\u_multiplier/_0932_ ),
    .Z(\u_multiplier/_1577_ ));
 XNOR2_X1 \u_multiplier/_2472_  (.A(\u_multiplier/_1575_ ),
    .B(\u_multiplier/_1577_ ),
    .ZN(\u_multiplier/_1578_ ));
 AOI21_X2 \u_multiplier/_2473_  (.A(\u_multiplier/_1578_ ),
    .B1(\u_multiplier/_1573_ ),
    .B2(\u_multiplier/_1571_ ),
    .ZN(\u_multiplier/_1579_ ));
 AND3_X1 \u_multiplier/_2474_  (.A1(\u_multiplier/_1571_ ),
    .A2(\u_multiplier/_1573_ ),
    .A3(\u_multiplier/_1578_ ),
    .ZN(\u_multiplier/_1580_ ));
 OR2_X2 \u_multiplier/_2475_  (.A1(\u_multiplier/_1579_ ),
    .A2(\u_multiplier/_1580_ ),
    .ZN(\u_multiplier/_1581_ ));
 XOR2_X2 \u_multiplier/_2476_  (.A(\u_multiplier/_1570_ ),
    .B(\u_multiplier/_1581_ ),
    .Z(\u_multiplier/_1582_ ));
 INV_X1 \u_multiplier/_2477_  (.A(\u_multiplier/_1582_ ),
    .ZN(\u_multiplier/_1583_ ));
 NOR3_X1 \u_multiplier/_2478_  (.A1(\u_multiplier/_1566_ ),
    .A2(\u_multiplier/_1568_ ),
    .A3(\u_multiplier/_1582_ ),
    .ZN(\u_multiplier/_1584_ ));
 AOI211_X2 \u_multiplier/_2479_  (.A(\u_multiplier/_1567_ ),
    .B(\u_multiplier/_1583_ ),
    .C1(\u_multiplier/_1547_ ),
    .C2(\u_multiplier/_1551_ ),
    .ZN(\u_multiplier/_1585_ ));
 NAND2_X1 \u_multiplier/_2480_  (.A1(\u_multiplier/_1566_ ),
    .A2(\u_multiplier/_1582_ ),
    .ZN(\u_multiplier/_1586_ ));
 NAND2_X1 \u_multiplier/_2481_  (.A1(\u_multiplier/_1739_ ),
    .A2(\u_multiplier/_1586_ ),
    .ZN(\u_multiplier/_1587_ ));
 NOR3_X1 \u_multiplier/_2482_  (.A1(\u_multiplier/_1584_ ),
    .A2(\u_multiplier/_1585_ ),
    .A3(\u_multiplier/_1587_ ),
    .ZN(product[19]));
 OAI21_X1 \u_multiplier/_2483_  (.A(\u_multiplier/_1586_ ),
    .B1(\u_multiplier/_1581_ ),
    .B2(\u_multiplier/_1570_ ),
    .ZN(\u_multiplier/_1588_ ));
 NOR2_X1 \u_multiplier/_2484_  (.A1(\u_multiplier/_1585_ ),
    .A2(\u_multiplier/_1588_ ),
    .ZN(\u_multiplier/_1589_ ));
 AOI21_X2 \u_multiplier/_2485_  (.A(\u_multiplier/_1579_ ),
    .B1(\u_multiplier/_1577_ ),
    .B2(\u_multiplier/_1575_ ),
    .ZN(\u_multiplier/_1590_ ));
 AND2_X1 \u_multiplier/_2486_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/_1504_ ),
    .ZN(\u_multiplier/_1591_ ));
 AND2_X1 \u_multiplier/_2487_  (.A1(\u_multiplier/_0939_ ),
    .A2(\u_multiplier/_1591_ ),
    .ZN(\u_multiplier/_1592_ ));
 AOI211_X2 \u_multiplier/_2488_  (.A(\u_multiplier/dec_out [20]),
    .B(\u_multiplier/_1592_ ),
    .C1(\u_multiplier/_1396_ ),
    .C2(\u_multiplier/K [3]),
    .ZN(\u_multiplier/_1593_ ));
 INV_X1 \u_multiplier/_2489_  (.A(\u_multiplier/_1593_ ),
    .ZN(\u_multiplier/_1594_ ));
 AND2_X1 \u_multiplier/_2490_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_1508_ ),
    .ZN(\u_multiplier/_1595_ ));
 OR2_X1 \u_multiplier/_2491_  (.A1(\u_multiplier/_0933_ ),
    .A2(\u_multiplier/_1401_ ),
    .ZN(\u_multiplier/_1596_ ));
 OAI21_X2 \u_multiplier/_2492_  (.A(\u_multiplier/_1596_ ),
    .B1(\u_multiplier/_1595_ ),
    .B2(\u_multiplier/code_x [3]),
    .ZN(\u_multiplier/_1597_ ));
 AND2_X1 \u_multiplier/_2493_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_1512_ ),
    .ZN(\u_multiplier/_1598_ ));
 OR2_X1 \u_multiplier/_2494_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_1598_ ),
    .ZN(\u_multiplier/_1599_ ));
 OAI21_X2 \u_multiplier/_2495_  (.A(\u_multiplier/_1599_ ),
    .B1(\u_multiplier/_1406_ ),
    .B2(\u_multiplier/_0932_ ),
    .ZN(\u_multiplier/_1600_ ));
 NOR2_X1 \u_multiplier/_2496_  (.A1(\u_multiplier/_1597_ ),
    .A2(\u_multiplier/_1600_ ),
    .ZN(\u_multiplier/_1601_ ));
 XOR2_X2 \u_multiplier/_2497_  (.A(\u_multiplier/_1597_ ),
    .B(\u_multiplier/_1600_ ),
    .Z(\u_multiplier/_1602_ ));
 XNOR2_X1 \u_multiplier/_2498_  (.A(\u_multiplier/_1593_ ),
    .B(\u_multiplier/_1602_ ),
    .ZN(\u_multiplier/_1603_ ));
 INV_X1 \u_multiplier/_2499_  (.A(\u_multiplier/_1603_ ),
    .ZN(\u_multiplier/_1604_ ));
 NOR2_X1 \u_multiplier/_2500_  (.A1(\u_multiplier/_1590_ ),
    .A2(\u_multiplier/_1604_ ),
    .ZN(\u_multiplier/_1605_ ));
 XNOR2_X2 \u_multiplier/_2501_  (.A(\u_multiplier/_1590_ ),
    .B(\u_multiplier/_1604_ ),
    .ZN(\u_multiplier/_1606_ ));
 INV_X1 \u_multiplier/_2502_  (.A(\u_multiplier/_1606_ ),
    .ZN(\u_multiplier/_1607_ ));
 NOR2_X1 \u_multiplier/_2503_  (.A1(\u_multiplier/_1589_ ),
    .A2(\u_multiplier/_1606_ ),
    .ZN(\u_multiplier/_1608_ ));
 AOI21_X1 \u_multiplier/_2504_  (.A(\u_multiplier/_0943_ ),
    .B1(\u_multiplier/_1589_ ),
    .B2(\u_multiplier/_1606_ ),
    .ZN(\u_multiplier/_1609_ ));
 OAI21_X1 \u_multiplier/_2505_  (.A(\u_multiplier/_1609_ ),
    .B1(\u_multiplier/_1606_ ),
    .B2(\u_multiplier/_1589_ ),
    .ZN(\u_multiplier/_1610_ ));
 INV_X2 \u_multiplier/_2506_  (.A(\u_multiplier/_1610_ ),
    .ZN(product[20]));
 AOI21_X2 \u_multiplier/_2507_  (.A(\u_multiplier/_1601_ ),
    .B1(\u_multiplier/_1602_ ),
    .B2(\u_multiplier/_1594_ ),
    .ZN(\u_multiplier/_1611_ ));
 NAND3_X2 \u_multiplier/_2508_  (.A1(\u_multiplier/K [1]),
    .A2(\u_multiplier/K [2]),
    .A3(\u_multiplier/_1473_ ),
    .ZN(\u_multiplier/_1612_ ));
 INV_X1 \u_multiplier/_2509_  (.A(\u_multiplier/_1612_ ),
    .ZN(\u_multiplier/_1613_ ));
 AOI21_X1 \u_multiplier/_2510_  (.A(\u_multiplier/dec_out [21]),
    .B1(\u_multiplier/_1423_ ),
    .B2(\u_multiplier/K [3]),
    .ZN(\u_multiplier/_1614_ ));
 OAI21_X2 \u_multiplier/_2511_  (.A(\u_multiplier/_1614_ ),
    .B1(\u_multiplier/_1612_ ),
    .B2(\u_multiplier/K [3]),
    .ZN(\u_multiplier/_1615_ ));
 NOR2_X2 \u_multiplier/_2512_  (.A1(\u_multiplier/_0935_ ),
    .A2(\u_multiplier/_1532_ ),
    .ZN(\u_multiplier/_1616_ ));
 NAND2_X1 \u_multiplier/_2513_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_1429_ ),
    .ZN(\u_multiplier/_1617_ ));
 OAI21_X2 \u_multiplier/_2514_  (.A(\u_multiplier/_1617_ ),
    .B1(\u_multiplier/_1616_ ),
    .B2(\u_multiplier/code_x [3]),
    .ZN(\u_multiplier/_1618_ ));
 OR2_X1 \u_multiplier/_2515_  (.A1(\u_multiplier/_0931_ ),
    .A2(\u_multiplier/_1537_ ),
    .ZN(\u_multiplier/_1619_ ));
 MUX2_X1 \u_multiplier/_2516_  (.A(\u_multiplier/_1434_ ),
    .B(\u_multiplier/_1619_ ),
    .S(\u_multiplier/_0932_ ),
    .Z(\u_multiplier/_1620_ ));
 NOR2_X1 \u_multiplier/_2517_  (.A1(\u_multiplier/_1618_ ),
    .A2(\u_multiplier/_1620_ ),
    .ZN(\u_multiplier/_1621_ ));
 XOR2_X2 \u_multiplier/_2518_  (.A(\u_multiplier/_1618_ ),
    .B(\u_multiplier/_1620_ ),
    .Z(\u_multiplier/_1622_ ));
 XNOR2_X2 \u_multiplier/_2519_  (.A(\u_multiplier/_1615_ ),
    .B(\u_multiplier/_1622_ ),
    .ZN(\u_multiplier/_1623_ ));
 NOR2_X1 \u_multiplier/_2520_  (.A1(\u_multiplier/_1611_ ),
    .A2(\u_multiplier/_1623_ ),
    .ZN(\u_multiplier/_1624_ ));
 XOR2_X2 \u_multiplier/_2521_  (.A(\u_multiplier/_1611_ ),
    .B(\u_multiplier/_1623_ ),
    .Z(\u_multiplier/_1625_ ));
 NOR3_X1 \u_multiplier/_2522_  (.A1(\u_multiplier/_1605_ ),
    .A2(\u_multiplier/_1608_ ),
    .A3(\u_multiplier/_1625_ ),
    .ZN(\u_multiplier/_1626_ ));
 OAI211_X2 \u_multiplier/_2523_  (.A(\u_multiplier/_1607_ ),
    .B(\u_multiplier/_1625_ ),
    .C1(\u_multiplier/_1585_ ),
    .C2(\u_multiplier/_1588_ ),
    .ZN(\u_multiplier/_1627_ ));
 AND2_X1 \u_multiplier/_2524_  (.A1(\u_multiplier/_1605_ ),
    .A2(\u_multiplier/_1625_ ),
    .ZN(\u_multiplier/_1628_ ));
 OR2_X1 \u_multiplier/_2525_  (.A1(\u_multiplier/_0943_ ),
    .A2(\u_multiplier/_1628_ ),
    .ZN(\u_multiplier/_1629_ ));
 AOI211_X1 \u_multiplier/_2526_  (.A(\u_multiplier/_1626_ ),
    .B(\u_multiplier/_1629_ ),
    .C1(\u_multiplier/_1608_ ),
    .C2(\u_multiplier/_1625_ ),
    .ZN(product[21]));
 NOR2_X1 \u_multiplier/_2527_  (.A1(\u_multiplier/_1624_ ),
    .A2(\u_multiplier/_1628_ ),
    .ZN(\u_multiplier/_1630_ ));
 NAND2_X1 \u_multiplier/_2528_  (.A1(\u_multiplier/_1627_ ),
    .A2(\u_multiplier/_1630_ ),
    .ZN(\u_multiplier/_1631_ ));
 AOI21_X2 \u_multiplier/_2529_  (.A(\u_multiplier/_1621_ ),
    .B1(\u_multiplier/_1622_ ),
    .B2(\u_multiplier/_1615_ ),
    .ZN(\u_multiplier/_1632_ ));
 AOI21_X2 \u_multiplier/_2530_  (.A(\u_multiplier/dec_out [22]),
    .B1(\u_multiplier/_1452_ ),
    .B2(\u_multiplier/K [3]),
    .ZN(\u_multiplier/_1633_ ));
 NAND2_X1 \u_multiplier/_2531_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_1457_ ),
    .ZN(\u_multiplier/_1634_ ));
 NAND2_X1 \u_multiplier/_2532_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_1462_ ),
    .ZN(\u_multiplier/_1635_ ));
 XOR2_X1 \u_multiplier/_2533_  (.A(\u_multiplier/_1634_ ),
    .B(\u_multiplier/_1635_ ),
    .Z(\u_multiplier/_1636_ ));
 INV_X1 \u_multiplier/_2534_  (.A(\u_multiplier/_1636_ ),
    .ZN(\u_multiplier/_1637_ ));
 OR2_X1 \u_multiplier/_2535_  (.A1(\u_multiplier/_1633_ ),
    .A2(\u_multiplier/_1637_ ),
    .ZN(\u_multiplier/_1638_ ));
 XNOR2_X2 \u_multiplier/_2536_  (.A(\u_multiplier/_1633_ ),
    .B(\u_multiplier/_1637_ ),
    .ZN(\u_multiplier/_1639_ ));
 NOR2_X1 \u_multiplier/_2537_  (.A1(\u_multiplier/_1632_ ),
    .A2(\u_multiplier/_1639_ ),
    .ZN(\u_multiplier/_1640_ ));
 XOR2_X2 \u_multiplier/_2538_  (.A(\u_multiplier/_1632_ ),
    .B(\u_multiplier/_1639_ ),
    .Z(\u_multiplier/_1641_ ));
 INV_X1 \u_multiplier/_2539_  (.A(\u_multiplier/_1641_ ),
    .ZN(\u_multiplier/_1642_ ));
 OAI21_X1 \u_multiplier/_2540_  (.A(\u_multiplier/_1739_ ),
    .B1(\u_multiplier/_1631_ ),
    .B2(\u_multiplier/_1641_ ),
    .ZN(\u_multiplier/_1643_ ));
 AOI21_X1 \u_multiplier/_2541_  (.A(\u_multiplier/_1643_ ),
    .B1(\u_multiplier/_1641_ ),
    .B2(\u_multiplier/_1631_ ),
    .ZN(product[22]));
 OAI21_X2 \u_multiplier/_2542_  (.A(\u_multiplier/_1638_ ),
    .B1(\u_multiplier/_1635_ ),
    .B2(\u_multiplier/_1634_ ),
    .ZN(\u_multiplier/_1644_ ));
 AOI21_X2 \u_multiplier/_2543_  (.A(\u_multiplier/dec_out [23]),
    .B1(\u_multiplier/_1476_ ),
    .B2(\u_multiplier/K [3]),
    .ZN(\u_multiplier/_1645_ ));
 NAND2_X1 \u_multiplier/_2544_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_1483_ ),
    .ZN(\u_multiplier/_1646_ ));
 NAND2_X1 \u_multiplier/_2545_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_1489_ ),
    .ZN(\u_multiplier/_1647_ ));
 XNOR2_X2 \u_multiplier/_2546_  (.A(\u_multiplier/_1646_ ),
    .B(\u_multiplier/_1647_ ),
    .ZN(\u_multiplier/_1648_ ));
 OR2_X1 \u_multiplier/_2547_  (.A1(\u_multiplier/_1645_ ),
    .A2(\u_multiplier/_1648_ ),
    .ZN(\u_multiplier/_1649_ ));
 XOR2_X2 \u_multiplier/_2548_  (.A(\u_multiplier/_1645_ ),
    .B(\u_multiplier/_1648_ ),
    .Z(\u_multiplier/_1650_ ));
 NAND2_X1 \u_multiplier/_2549_  (.A1(\u_multiplier/_1644_ ),
    .A2(\u_multiplier/_1650_ ),
    .ZN(\u_multiplier/_1651_ ));
 XOR2_X2 \u_multiplier/_2550_  (.A(\u_multiplier/_1644_ ),
    .B(\u_multiplier/_1650_ ),
    .Z(\u_multiplier/_1652_ ));
 INV_X1 \u_multiplier/_2551_  (.A(\u_multiplier/_1652_ ),
    .ZN(\u_multiplier/_1653_ ));
 AOI211_X1 \u_multiplier/_2552_  (.A(\u_multiplier/_1640_ ),
    .B(\u_multiplier/_1652_ ),
    .C1(\u_multiplier/_1641_ ),
    .C2(\u_multiplier/_1631_ ),
    .ZN(\u_multiplier/_1654_ ));
 AOI211_X2 \u_multiplier/_2553_  (.A(\u_multiplier/_1642_ ),
    .B(\u_multiplier/_1653_ ),
    .C1(\u_multiplier/_1627_ ),
    .C2(\u_multiplier/_1630_ ),
    .ZN(\u_multiplier/_1655_ ));
 NAND2_X1 \u_multiplier/_2554_  (.A1(\u_multiplier/_1640_ ),
    .A2(\u_multiplier/_1652_ ),
    .ZN(\u_multiplier/_1656_ ));
 NAND2_X1 \u_multiplier/_2555_  (.A1(\u_multiplier/_1739_ ),
    .A2(\u_multiplier/_1656_ ),
    .ZN(\u_multiplier/_1657_ ));
 NOR3_X1 \u_multiplier/_2556_  (.A1(\u_multiplier/_1654_ ),
    .A2(\u_multiplier/_1655_ ),
    .A3(\u_multiplier/_1657_ ),
    .ZN(product[23]));
 NAND2_X1 \u_multiplier/_2557_  (.A1(\u_multiplier/_1651_ ),
    .A2(\u_multiplier/_1656_ ),
    .ZN(\u_multiplier/_1658_ ));
 OAI21_X1 \u_multiplier/_2558_  (.A(\u_multiplier/_1649_ ),
    .B1(\u_multiplier/_1647_ ),
    .B2(\u_multiplier/_1646_ ),
    .ZN(\u_multiplier/_1659_ ));
 INV_X1 \u_multiplier/_2559_  (.A(\u_multiplier/_1659_ ),
    .ZN(\u_multiplier/_1660_ ));
 AOI21_X1 \u_multiplier/_2560_  (.A(\u_multiplier/dec_out [24]),
    .B1(\u_multiplier/_1505_ ),
    .B2(\u_multiplier/K [3]),
    .ZN(\u_multiplier/_1661_ ));
 NAND2_X1 \u_multiplier/_2561_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_1509_ ),
    .ZN(\u_multiplier/_1662_ ));
 NAND2_X1 \u_multiplier/_2562_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_1513_ ),
    .ZN(\u_multiplier/_1663_ ));
 XNOR2_X1 \u_multiplier/_2563_  (.A(\u_multiplier/_1662_ ),
    .B(\u_multiplier/_1663_ ),
    .ZN(\u_multiplier/_1664_ ));
 OR2_X1 \u_multiplier/_2564_  (.A1(\u_multiplier/_1661_ ),
    .A2(\u_multiplier/_1664_ ),
    .ZN(\u_multiplier/_1665_ ));
 XNOR2_X1 \u_multiplier/_2565_  (.A(\u_multiplier/_1661_ ),
    .B(\u_multiplier/_1664_ ),
    .ZN(\u_multiplier/_1666_ ));
 NOR2_X1 \u_multiplier/_2566_  (.A1(\u_multiplier/_1660_ ),
    .A2(\u_multiplier/_1666_ ),
    .ZN(\u_multiplier/_1667_ ));
 INV_X1 \u_multiplier/_2567_  (.A(\u_multiplier/_1667_ ),
    .ZN(\u_multiplier/_1668_ ));
 XNOR2_X1 \u_multiplier/_2568_  (.A(\u_multiplier/_1659_ ),
    .B(\u_multiplier/_1666_ ),
    .ZN(\u_multiplier/_1669_ ));
 OAI21_X1 \u_multiplier/_2569_  (.A(\u_multiplier/_1669_ ),
    .B1(\u_multiplier/_1658_ ),
    .B2(\u_multiplier/_1655_ ),
    .ZN(\u_multiplier/_1670_ ));
 NOR3_X1 \u_multiplier/_2570_  (.A1(\u_multiplier/_1655_ ),
    .A2(\u_multiplier/_1658_ ),
    .A3(\u_multiplier/_1669_ ),
    .ZN(\u_multiplier/_1671_ ));
 NOR2_X1 \u_multiplier/_2571_  (.A1(\u_multiplier/_0943_ ),
    .A2(\u_multiplier/_1671_ ),
    .ZN(\u_multiplier/_1672_ ));
 AND2_X1 \u_multiplier/_2572_  (.A1(\u_multiplier/_1670_ ),
    .A2(\u_multiplier/_1672_ ),
    .ZN(product[24]));
 OAI21_X2 \u_multiplier/_2573_  (.A(\u_multiplier/_1665_ ),
    .B1(\u_multiplier/_1663_ ),
    .B2(\u_multiplier/_1662_ ),
    .ZN(\u_multiplier/_1673_ ));
 INV_X1 \u_multiplier/_2574_  (.A(\u_multiplier/_1673_ ),
    .ZN(\u_multiplier/_1674_ ));
 AOI21_X2 \u_multiplier/_2575_  (.A(\u_multiplier/dec_out [25]),
    .B1(\u_multiplier/_1528_ ),
    .B2(\u_multiplier/K [3]),
    .ZN(\u_multiplier/_1675_ ));
 AOI22_X1 \u_multiplier/_2576_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_1534_ ),
    .B1(\u_multiplier/_1539_ ),
    .B2(\u_multiplier/code_y [3]),
    .ZN(\u_multiplier/_1676_ ));
 AND4_X1 \u_multiplier/_2577_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/code_x [3]),
    .A3(\u_multiplier/_1534_ ),
    .A4(\u_multiplier/_1539_ ),
    .ZN(\u_multiplier/_1677_ ));
 OR2_X1 \u_multiplier/_2578_  (.A1(\u_multiplier/_1676_ ),
    .A2(\u_multiplier/_1677_ ),
    .ZN(\u_multiplier/_1678_ ));
 NOR2_X1 \u_multiplier/_2579_  (.A1(\u_multiplier/_1675_ ),
    .A2(\u_multiplier/_1678_ ),
    .ZN(\u_multiplier/_1679_ ));
 XNOR2_X2 \u_multiplier/_2580_  (.A(\u_multiplier/_1675_ ),
    .B(\u_multiplier/_1678_ ),
    .ZN(\u_multiplier/_1680_ ));
 NOR2_X1 \u_multiplier/_2581_  (.A1(\u_multiplier/_1674_ ),
    .A2(\u_multiplier/_1680_ ),
    .ZN(\u_multiplier/_1681_ ));
 XOR2_X2 \u_multiplier/_2582_  (.A(\u_multiplier/_1673_ ),
    .B(\u_multiplier/_1680_ ),
    .Z(\u_multiplier/_1682_ ));
 AOI21_X2 \u_multiplier/_2583_  (.A(\u_multiplier/_1682_ ),
    .B1(\u_multiplier/_1670_ ),
    .B2(\u_multiplier/_1668_ ),
    .ZN(\u_multiplier/_1683_ ));
 AND3_X1 \u_multiplier/_2584_  (.A1(\u_multiplier/_1668_ ),
    .A2(\u_multiplier/_1670_ ),
    .A3(\u_multiplier/_1682_ ),
    .ZN(\u_multiplier/_1684_ ));
 NOR3_X1 \u_multiplier/_2585_  (.A1(\u_multiplier/_0943_ ),
    .A2(\u_multiplier/_1683_ ),
    .A3(\u_multiplier/_1684_ ),
    .ZN(product[25]));
 OR2_X1 \u_multiplier/_2586_  (.A1(\u_multiplier/_1681_ ),
    .A2(\u_multiplier/_1683_ ),
    .ZN(\u_multiplier/_1685_ ));
 NOR2_X1 \u_multiplier/_2587_  (.A1(\u_multiplier/_1677_ ),
    .A2(\u_multiplier/_1679_ ),
    .ZN(\u_multiplier/_1686_ ));
 OAI21_X2 \u_multiplier/_2588_  (.A(\u_multiplier/_0941_ ),
    .B1(\u_multiplier/_1554_ ),
    .B2(\u_multiplier/_0939_ ),
    .ZN(\u_multiplier/_1687_ ));
 AOI22_X2 \u_multiplier/_2589_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_1557_ ),
    .B1(\u_multiplier/_1560_ ),
    .B2(\u_multiplier/code_y [3]),
    .ZN(\u_multiplier/_1688_ ));
 AND4_X1 \u_multiplier/_2590_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/code_x [3]),
    .A3(\u_multiplier/_1557_ ),
    .A4(\u_multiplier/_1560_ ),
    .ZN(\u_multiplier/_1689_ ));
 NOR2_X2 \u_multiplier/_2591_  (.A1(\u_multiplier/_1688_ ),
    .A2(\u_multiplier/_1689_ ),
    .ZN(\u_multiplier/_1690_ ));
 XNOR2_X2 \u_multiplier/_2592_  (.A(\u_multiplier/_1687_ ),
    .B(\u_multiplier/_1690_ ),
    .ZN(\u_multiplier/_1691_ ));
 OR2_X1 \u_multiplier/_2593_  (.A1(\u_multiplier/_1686_ ),
    .A2(\u_multiplier/_1691_ ),
    .ZN(\u_multiplier/_1692_ ));
 XOR2_X2 \u_multiplier/_2594_  (.A(\u_multiplier/_1686_ ),
    .B(\u_multiplier/_1691_ ),
    .Z(\u_multiplier/_1693_ ));
 OAI21_X1 \u_multiplier/_2595_  (.A(\u_multiplier/_1693_ ),
    .B1(\u_multiplier/_1683_ ),
    .B2(\u_multiplier/_1681_ ),
    .ZN(\u_multiplier/_1694_ ));
 OAI21_X1 \u_multiplier/_2596_  (.A(\u_multiplier/_1739_ ),
    .B1(\u_multiplier/_1685_ ),
    .B2(\u_multiplier/_1693_ ),
    .ZN(\u_multiplier/_1695_ ));
 AOI21_X1 \u_multiplier/_2597_  (.A(\u_multiplier/_1695_ ),
    .B1(\u_multiplier/_1693_ ),
    .B2(\u_multiplier/_1685_ ),
    .ZN(product[26]));
 AOI21_X1 \u_multiplier/_2598_  (.A(\u_multiplier/_1689_ ),
    .B1(\u_multiplier/_1690_ ),
    .B2(\u_multiplier/_1687_ ),
    .ZN(\u_multiplier/_1696_ ));
 AOI21_X1 \u_multiplier/_2599_  (.A(\u_multiplier/dec_out [27]),
    .B1(\u_multiplier/_1572_ ),
    .B2(\u_multiplier/K [3]),
    .ZN(\u_multiplier/_1697_ ));
 NAND2_X1 \u_multiplier/_2600_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_1574_ ),
    .ZN(\u_multiplier/_1698_ ));
 NAND2_X1 \u_multiplier/_2601_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/_1576_ ),
    .ZN(\u_multiplier/_1699_ ));
 XOR2_X1 \u_multiplier/_2602_  (.A(\u_multiplier/_1698_ ),
    .B(\u_multiplier/_1699_ ),
    .Z(\u_multiplier/_1700_ ));
 INV_X1 \u_multiplier/_2603_  (.A(\u_multiplier/_1700_ ),
    .ZN(\u_multiplier/_1701_ ));
 OR2_X1 \u_multiplier/_2604_  (.A1(\u_multiplier/_1697_ ),
    .A2(\u_multiplier/_1701_ ),
    .ZN(\u_multiplier/_1702_ ));
 XNOR2_X1 \u_multiplier/_2605_  (.A(\u_multiplier/_1697_ ),
    .B(\u_multiplier/_1701_ ),
    .ZN(\u_multiplier/_1703_ ));
 NOR2_X1 \u_multiplier/_2606_  (.A1(\u_multiplier/_1696_ ),
    .A2(\u_multiplier/_1703_ ),
    .ZN(\u_multiplier/_1704_ ));
 XOR2_X1 \u_multiplier/_2607_  (.A(\u_multiplier/_1696_ ),
    .B(\u_multiplier/_1703_ ),
    .Z(\u_multiplier/_1705_ ));
 INV_X1 \u_multiplier/_2608_  (.A(\u_multiplier/_1705_ ),
    .ZN(\u_multiplier/_1706_ ));
 AOI21_X2 \u_multiplier/_2609_  (.A(\u_multiplier/_1706_ ),
    .B1(\u_multiplier/_1694_ ),
    .B2(\u_multiplier/_1692_ ),
    .ZN(\u_multiplier/_1707_ ));
 NAND3_X1 \u_multiplier/_2610_  (.A1(\u_multiplier/_1692_ ),
    .A2(\u_multiplier/_1694_ ),
    .A3(\u_multiplier/_1706_ ),
    .ZN(\u_multiplier/_1708_ ));
 NAND2_X1 \u_multiplier/_2611_  (.A1(\u_multiplier/_1739_ ),
    .A2(\u_multiplier/_1708_ ),
    .ZN(\u_multiplier/_1709_ ));
 NOR2_X1 \u_multiplier/_2612_  (.A1(\u_multiplier/_1707_ ),
    .A2(\u_multiplier/_1709_ ),
    .ZN(product[27]));
 OAI21_X1 \u_multiplier/_2613_  (.A(\u_multiplier/_1702_ ),
    .B1(\u_multiplier/_1699_ ),
    .B2(\u_multiplier/_1698_ ),
    .ZN(\u_multiplier/_1710_ ));
 AOI21_X1 \u_multiplier/_2614_  (.A(\u_multiplier/dec_out [28]),
    .B1(\u_multiplier/_1591_ ),
    .B2(\u_multiplier/K [3]),
    .ZN(\u_multiplier/_1711_ ));
 INV_X1 \u_multiplier/_2615_  (.A(\u_multiplier/_1711_ ),
    .ZN(\u_multiplier/_1712_ ));
 AOI22_X1 \u_multiplier/_2616_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_1595_ ),
    .B1(\u_multiplier/_1598_ ),
    .B2(\u_multiplier/code_y [3]),
    .ZN(\u_multiplier/_1713_ ));
 AND4_X1 \u_multiplier/_2617_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/code_x [3]),
    .A3(\u_multiplier/_1595_ ),
    .A4(\u_multiplier/_1598_ ),
    .ZN(\u_multiplier/_1714_ ));
 NOR2_X1 \u_multiplier/_2618_  (.A1(\u_multiplier/_1713_ ),
    .A2(\u_multiplier/_1714_ ),
    .ZN(\u_multiplier/_1715_ ));
 XNOR2_X1 \u_multiplier/_2619_  (.A(\u_multiplier/_1711_ ),
    .B(\u_multiplier/_1715_ ),
    .ZN(\u_multiplier/_1716_ ));
 AND2_X1 \u_multiplier/_2620_  (.A1(\u_multiplier/_1710_ ),
    .A2(\u_multiplier/_1716_ ),
    .ZN(\u_multiplier/_1717_ ));
 INV_X1 \u_multiplier/_2621_  (.A(\u_multiplier/_1717_ ),
    .ZN(\u_multiplier/_1718_ ));
 XOR2_X1 \u_multiplier/_2622_  (.A(\u_multiplier/_1710_ ),
    .B(\u_multiplier/_1716_ ),
    .Z(\u_multiplier/_1719_ ));
 OAI21_X1 \u_multiplier/_2623_  (.A(\u_multiplier/_1719_ ),
    .B1(\u_multiplier/_1707_ ),
    .B2(\u_multiplier/_1704_ ),
    .ZN(\u_multiplier/_1720_ ));
 OR3_X1 \u_multiplier/_2624_  (.A1(\u_multiplier/_1704_ ),
    .A2(\u_multiplier/_1707_ ),
    .A3(\u_multiplier/_1719_ ),
    .ZN(\u_multiplier/_1721_ ));
 AND3_X1 \u_multiplier/_2625_  (.A1(\u_multiplier/_1739_ ),
    .A2(\u_multiplier/_1720_ ),
    .A3(\u_multiplier/_1721_ ),
    .ZN(product[28]));
 AOI21_X1 \u_multiplier/_2626_  (.A(\u_multiplier/_1714_ ),
    .B1(\u_multiplier/_1715_ ),
    .B2(\u_multiplier/_1712_ ),
    .ZN(\u_multiplier/_1722_ ));
 AOI21_X2 \u_multiplier/_2627_  (.A(\u_multiplier/dec_out [29]),
    .B1(\u_multiplier/_1613_ ),
    .B2(\u_multiplier/K [3]),
    .ZN(\u_multiplier/_1723_ ));
 NAND2_X1 \u_multiplier/_2628_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_1616_ ),
    .ZN(\u_multiplier/_1724_ ));
 NOR2_X1 \u_multiplier/_2629_  (.A1(\u_multiplier/_0932_ ),
    .A2(\u_multiplier/_1619_ ),
    .ZN(\u_multiplier/_1725_ ));
 NAND3_X1 \u_multiplier/_2630_  (.A1(\u_multiplier/code_x [3]),
    .A2(\u_multiplier/_1616_ ),
    .A3(\u_multiplier/_1725_ ),
    .ZN(\u_multiplier/_1726_ ));
 XOR2_X2 \u_multiplier/_2631_  (.A(\u_multiplier/_1724_ ),
    .B(\u_multiplier/_1725_ ),
    .Z(\u_multiplier/_1727_ ));
 XNOR2_X1 \u_multiplier/_2632_  (.A(\u_multiplier/_1723_ ),
    .B(\u_multiplier/_1727_ ),
    .ZN(\u_multiplier/_1728_ ));
 OR2_X1 \u_multiplier/_2633_  (.A1(\u_multiplier/_1722_ ),
    .A2(\u_multiplier/_1728_ ),
    .ZN(\u_multiplier/_1729_ ));
 INV_X1 \u_multiplier/_2634_  (.A(\u_multiplier/_1729_ ),
    .ZN(\u_multiplier/_1730_ ));
 XNOR2_X1 \u_multiplier/_2635_  (.A(\u_multiplier/_1722_ ),
    .B(\u_multiplier/_1728_ ),
    .ZN(\u_multiplier/_1731_ ));
 AOI21_X2 \u_multiplier/_2636_  (.A(\u_multiplier/_1731_ ),
    .B1(\u_multiplier/_1720_ ),
    .B2(\u_multiplier/_1718_ ),
    .ZN(\u_multiplier/_1732_ ));
 AND3_X1 \u_multiplier/_2637_  (.A1(\u_multiplier/_1718_ ),
    .A2(\u_multiplier/_1720_ ),
    .A3(\u_multiplier/_1731_ ),
    .ZN(\u_multiplier/_1733_ ));
 NOR3_X1 \u_multiplier/_2638_  (.A1(\u_multiplier/_0943_ ),
    .A2(\u_multiplier/_1732_ ),
    .A3(\u_multiplier/_1733_ ),
    .ZN(product[29]));
 OAI21_X2 \u_multiplier/_2639_  (.A(\u_multiplier/_1726_ ),
    .B1(\u_multiplier/_1727_ ),
    .B2(\u_multiplier/_1723_ ),
    .ZN(\u_multiplier/_1734_ ));
 NAND2_X1 \u_multiplier/_2640_  (.A1(\u_multiplier/dec_out [30]),
    .A2(\u_multiplier/_1734_ ),
    .ZN(\u_multiplier/_1735_ ));
 XOR2_X2 \u_multiplier/_2641_  (.A(\u_multiplier/dec_out [30]),
    .B(\u_multiplier/_1734_ ),
    .Z(\u_multiplier/_1736_ ));
 OAI21_X2 \u_multiplier/_2642_  (.A(\u_multiplier/_1736_ ),
    .B1(\u_multiplier/_1732_ ),
    .B2(\u_multiplier/_1730_ ),
    .ZN(\u_multiplier/_1737_ ));
 OR3_X1 \u_multiplier/_2643_  (.A1(\u_multiplier/_1730_ ),
    .A2(\u_multiplier/_1732_ ),
    .A3(\u_multiplier/_1736_ ),
    .ZN(\u_multiplier/_1738_ ));
 AND3_X2 \u_multiplier/_2644_  (.A1(\u_multiplier/_1739_ ),
    .A2(\u_multiplier/_1737_ ),
    .A3(\u_multiplier/_1738_ ),
    .ZN(product[30]));
 AND3_X1 \u_multiplier/_2645_  (.A1(\u_multiplier/_0942_ ),
    .A2(\u_multiplier/_1735_ ),
    .A3(\u_multiplier/_1737_ ),
    .ZN(\u_multiplier/_0917_ ));
 AOI21_X2 \u_multiplier/_2646_  (.A(\u_multiplier/_0942_ ),
    .B1(\u_multiplier/_1735_ ),
    .B2(\u_multiplier/_1737_ ),
    .ZN(\u_multiplier/_0918_ ));
 NOR3_X4 \u_multiplier/_2647_  (.A1(\u_multiplier/_0943_ ),
    .A2(\u_multiplier/_0917_ ),
    .A3(\u_multiplier/_0918_ ),
    .ZN(product[31]));
 MUX2_X2 \u_multiplier/_2648_  (.A(\u_multiplier/_0965_ ),
    .B(\u_multiplier/_0944_ ),
    .S(\u_multiplier/_1059_ ),
    .Z(\u_multiplier/_0827_ ));
 MUX2_X2 \u_multiplier/_2649_  (.A(\u_multiplier/_0969_ ),
    .B(\u_multiplier/_0967_ ),
    .S(\u_multiplier/_1059_ ),
    .Z(\u_multiplier/_0833_ ));
 MUX2_X2 \u_multiplier/_2650_  (.A(\u_multiplier/_0975_ ),
    .B(\u_multiplier/_0973_ ),
    .S(\u_multiplier/_1059_ ),
    .Z(\u_multiplier/_0834_ ));
 MUX2_X2 \u_multiplier/_2651_  (.A(\u_multiplier/_0981_ ),
    .B(\u_multiplier/_0979_ ),
    .S(\u_multiplier/_1059_ ),
    .Z(\u_multiplier/_0835_ ));
 MUX2_X2 \u_multiplier/_2652_  (.A(\u_multiplier/_0990_ ),
    .B(\u_multiplier/_0988_ ),
    .S(\u_multiplier/_1059_ ),
    .Z(\u_multiplier/_0836_ ));
 MUX2_X2 \u_multiplier/_2653_  (.A(\u_multiplier/_0993_ ),
    .B(\u_multiplier/_0991_ ),
    .S(\u_multiplier/_1059_ ),
    .Z(\u_multiplier/_0837_ ));
 MUX2_X2 \u_multiplier/_2654_  (.A(\u_multiplier/_0961_ ),
    .B(\u_multiplier/_0960_ ),
    .S(\u_multiplier/_1059_ ),
    .Z(\u_multiplier/_0838_ ));
 MUX2_X2 \u_multiplier/_2655_  (.A(\u_multiplier/_0958_ ),
    .B(\u_multiplier/_0956_ ),
    .S(\u_multiplier/_1059_ ),
    .Z(\u_multiplier/_0839_ ));
 MUX2_X2 \u_multiplier/_2656_  (.A(\u_multiplier/_0952_ ),
    .B(\u_multiplier/_0950_ ),
    .S(\u_multiplier/_1059_ ),
    .Z(\u_multiplier/_0840_ ));
 MUX2_X2 \u_multiplier/_2657_  (.A(\u_multiplier/_0948_ ),
    .B(\u_multiplier/_0946_ ),
    .S(\u_multiplier/_1059_ ),
    .Z(\u_multiplier/_0841_ ));
 MUX2_X2 \u_multiplier/_2658_  (.A(\u_multiplier/_1031_ ),
    .B(\u_multiplier/_1029_ ),
    .S(\u_multiplier/_1059_ ),
    .Z(\u_multiplier/_0828_ ));
 MUX2_X2 \u_multiplier/_2659_  (.A(\u_multiplier/_1027_ ),
    .B(\u_multiplier/_1025_ ),
    .S(\u_multiplier/_1059_ ),
    .Z(\u_multiplier/_0829_ ));
 MUX2_X2 \u_multiplier/_2660_  (.A(\u_multiplier/_1021_ ),
    .B(\u_multiplier/_1019_ ),
    .S(\u_multiplier/_1059_ ),
    .Z(\u_multiplier/_0830_ ));
 MUX2_X2 \u_multiplier/_2661_  (.A(\u_multiplier/_1016_ ),
    .B(\u_multiplier/_1015_ ),
    .S(\u_multiplier/_1059_ ),
    .Z(\u_multiplier/_0831_ ));
 OAI21_X4 \u_multiplier/_2662_  (.A(\u_multiplier/_1040_ ),
    .B1(\u_multiplier/_1042_ ),
    .B2(\u_multiplier/_1056_ ),
    .ZN(\u_multiplier/_0832_ ));
 NAND2_X1 \u_multiplier/_2663_  (.A1(\u_multiplier/code_y [0]),
    .A2(\u_multiplier/code_x [0]),
    .ZN(\u_multiplier/_0919_ ));
 NAND2_X1 \u_multiplier/_2664_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/code_x [1]),
    .ZN(\u_multiplier/_0920_ ));
 XOR2_X2 \u_multiplier/_2665_  (.A(\u_multiplier/code_y [1]),
    .B(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_0921_ ));
 NAND3_X2 \u_multiplier/_2666_  (.A1(\u_multiplier/code_y [0]),
    .A2(\u_multiplier/code_x [0]),
    .A3(\u_multiplier/_0921_ ),
    .ZN(\u_multiplier/_0922_ ));
 XNOR2_X2 \u_multiplier/_2667_  (.A(\u_multiplier/_0919_ ),
    .B(\u_multiplier/_0921_ ),
    .ZN(\u_multiplier/_0843_ ));
 XNOR2_X2 \u_multiplier/_2668_  (.A(\u_multiplier/code_y [2]),
    .B(\u_multiplier/code_x [2]),
    .ZN(\u_multiplier/_0923_ ));
 AOI21_X4 \u_multiplier/_2669_  (.A(\u_multiplier/_0923_ ),
    .B1(\u_multiplier/_0922_ ),
    .B2(\u_multiplier/_0920_ ),
    .ZN(\u_multiplier/_0924_ ));
 AND3_X1 \u_multiplier/_2670_  (.A1(\u_multiplier/_0920_ ),
    .A2(\u_multiplier/_0922_ ),
    .A3(\u_multiplier/_0923_ ),
    .ZN(\u_multiplier/_0925_ ));
 NOR2_X4 \u_multiplier/_2671_  (.A1(\u_multiplier/_0924_ ),
    .A2(\u_multiplier/_0925_ ),
    .ZN(\u_multiplier/_0844_ ));
 AOI21_X4 \u_multiplier/_2672_  (.A(\u_multiplier/_0924_ ),
    .B1(\u_multiplier/code_x [2]),
    .B2(\u_multiplier/code_y [2]),
    .ZN(\u_multiplier/_0926_ ));
 NOR2_X1 \u_multiplier/_2673_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/code_x [3]),
    .ZN(\u_multiplier/_0927_ ));
 NAND2_X1 \u_multiplier/_2674_  (.A1(\u_multiplier/code_y [3]),
    .A2(\u_multiplier/code_x [3]),
    .ZN(\u_multiplier/_0928_ ));
 XOR2_X2 \u_multiplier/_2675_  (.A(\u_multiplier/code_y [3]),
    .B(\u_multiplier/code_x [3]),
    .Z(\u_multiplier/_0929_ ));
 XNOR2_X2 \u_multiplier/_2676_  (.A(\u_multiplier/_0926_ ),
    .B(\u_multiplier/_0929_ ),
    .ZN(\u_multiplier/_0845_ ));
 XOR2_X2 \u_multiplier/_2677_  (.A(\u_multiplier/code_y [0]),
    .B(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_0842_ ));
 AOI21_X4 \u_multiplier/_2678_  (.A(\u_multiplier/_0927_ ),
    .B1(\u_multiplier/_0928_ ),
    .B2(\u_multiplier/_0926_ ),
    .ZN(\u_multiplier/_0846_ ));
 INV_X4 \u_multiplier/dec/_089_  (.A(\u_multiplier/_0846_ ),
    .ZN(\u_multiplier/dec/_068_ ));
 INV_X1 \u_multiplier/dec/_090_  (.A(\u_multiplier/_0842_ ),
    .ZN(\u_multiplier/dec/_069_ ));
 INV_X1 \u_multiplier/dec/_091_  (.A(\u_multiplier/_0843_ ),
    .ZN(\u_multiplier/dec/_070_ ));
 INV_X1 \u_multiplier/dec/_092_  (.A(\u_multiplier/_0844_ ),
    .ZN(\u_multiplier/dec/_071_ ));
 INV_X1 \u_multiplier/dec/_093_  (.A(\u_multiplier/_0845_ ),
    .ZN(\u_multiplier/dec/_072_ ));
 NOR2_X1 \u_multiplier/dec/_094_  (.A1(\u_multiplier/_0842_ ),
    .A2(\u_multiplier/_0843_ ),
    .ZN(\u_multiplier/dec/_073_ ));
 OR3_X1 \u_multiplier/dec/_095_  (.A1(\u_multiplier/_0842_ ),
    .A2(\u_multiplier/_0843_ ),
    .A3(\u_multiplier/_0844_ ),
    .ZN(\u_multiplier/dec/_074_ ));
 NOR3_X1 \u_multiplier/dec/_096_  (.A1(\u_multiplier/_0846_ ),
    .A2(\u_multiplier/_0845_ ),
    .A3(\u_multiplier/dec/_074_ ),
    .ZN(\u_multiplier/dec_out [0]));
 NAND2_X2 \u_multiplier/dec/_097_  (.A1(\u_multiplier/_0842_ ),
    .A2(\u_multiplier/dec/_070_ ),
    .ZN(\u_multiplier/dec/_075_ ));
 NOR4_X2 \u_multiplier/dec/_098_  (.A1(\u_multiplier/_0846_ ),
    .A2(\u_multiplier/_0844_ ),
    .A3(\u_multiplier/_0845_ ),
    .A4(\u_multiplier/dec/_075_ ),
    .ZN(\u_multiplier/dec_out [1]));
 NAND2_X1 \u_multiplier/dec/_099_  (.A1(\u_multiplier/dec/_069_ ),
    .A2(\u_multiplier/_0843_ ),
    .ZN(\u_multiplier/dec/_076_ ));
 NOR4_X1 \u_multiplier/dec/_100_  (.A1(\u_multiplier/_0846_ ),
    .A2(\u_multiplier/_0844_ ),
    .A3(\u_multiplier/_0845_ ),
    .A4(\u_multiplier/dec/_076_ ),
    .ZN(\u_multiplier/dec_out [2]));
 NAND2_X2 \u_multiplier/dec/_101_  (.A1(\u_multiplier/_0842_ ),
    .A2(\u_multiplier/_0843_ ),
    .ZN(\u_multiplier/dec/_077_ ));
 NOR4_X2 \u_multiplier/dec/_102_  (.A1(\u_multiplier/_0846_ ),
    .A2(\u_multiplier/_0844_ ),
    .A3(\u_multiplier/_0845_ ),
    .A4(\u_multiplier/dec/_077_ ),
    .ZN(\u_multiplier/dec_out [3]));
 NAND2_X1 \u_multiplier/dec/_103_  (.A1(\u_multiplier/_0844_ ),
    .A2(\u_multiplier/dec/_073_ ),
    .ZN(\u_multiplier/dec/_078_ ));
 NOR3_X1 \u_multiplier/dec/_104_  (.A1(\u_multiplier/_0846_ ),
    .A2(\u_multiplier/_0845_ ),
    .A3(\u_multiplier/dec/_078_ ),
    .ZN(\u_multiplier/dec_out [4]));
 NAND3_X1 \u_multiplier/dec/_105_  (.A1(\u_multiplier/_0842_ ),
    .A2(\u_multiplier/dec/_070_ ),
    .A3(\u_multiplier/_0844_ ),
    .ZN(\u_multiplier/dec/_079_ ));
 NOR3_X2 \u_multiplier/dec/_106_  (.A1(\u_multiplier/_0846_ ),
    .A2(\u_multiplier/_0845_ ),
    .A3(\u_multiplier/dec/_079_ ),
    .ZN(\u_multiplier/dec_out [5]));
 NAND3_X1 \u_multiplier/dec/_107_  (.A1(\u_multiplier/dec/_069_ ),
    .A2(\u_multiplier/_0843_ ),
    .A3(\u_multiplier/_0844_ ),
    .ZN(\u_multiplier/dec/_080_ ));
 NOR3_X1 \u_multiplier/dec/_108_  (.A1(\u_multiplier/_0846_ ),
    .A2(\u_multiplier/_0845_ ),
    .A3(\u_multiplier/dec/_080_ ),
    .ZN(\u_multiplier/dec_out [6]));
 NAND3_X1 \u_multiplier/dec/_109_  (.A1(\u_multiplier/_0842_ ),
    .A2(\u_multiplier/_0843_ ),
    .A3(\u_multiplier/_0844_ ),
    .ZN(\u_multiplier/dec/_081_ ));
 NOR3_X1 \u_multiplier/dec/_110_  (.A1(\u_multiplier/_0846_ ),
    .A2(\u_multiplier/_0845_ ),
    .A3(\u_multiplier/dec/_081_ ),
    .ZN(\u_multiplier/dec_out [7]));
 OR2_X1 \u_multiplier/dec/_111_  (.A1(\u_multiplier/dec/_072_ ),
    .A2(\u_multiplier/dec/_074_ ),
    .ZN(\u_multiplier/dec/_082_ ));
 NOR2_X1 \u_multiplier/dec/_112_  (.A1(\u_multiplier/_0846_ ),
    .A2(\u_multiplier/dec/_082_ ),
    .ZN(\u_multiplier/dec_out [8]));
 NAND4_X1 \u_multiplier/dec/_113_  (.A1(\u_multiplier/_0842_ ),
    .A2(\u_multiplier/dec/_070_ ),
    .A3(\u_multiplier/dec/_071_ ),
    .A4(\u_multiplier/_0845_ ),
    .ZN(\u_multiplier/dec/_083_ ));
 NOR2_X1 \u_multiplier/dec/_114_  (.A1(\u_multiplier/_0846_ ),
    .A2(\u_multiplier/dec/_083_ ),
    .ZN(\u_multiplier/dec_out [9]));
 NAND4_X1 \u_multiplier/dec/_115_  (.A1(\u_multiplier/dec/_069_ ),
    .A2(\u_multiplier/_0843_ ),
    .A3(\u_multiplier/dec/_071_ ),
    .A4(\u_multiplier/_0845_ ),
    .ZN(\u_multiplier/dec/_084_ ));
 NOR2_X1 \u_multiplier/dec/_116_  (.A1(\u_multiplier/_0846_ ),
    .A2(\u_multiplier/dec/_084_ ),
    .ZN(\u_multiplier/dec_out [10]));
 NOR4_X1 \u_multiplier/dec/_117_  (.A1(\u_multiplier/_0846_ ),
    .A2(\u_multiplier/_0844_ ),
    .A3(\u_multiplier/dec/_072_ ),
    .A4(\u_multiplier/dec/_077_ ),
    .ZN(\u_multiplier/dec_out [11]));
 NAND3_X1 \u_multiplier/dec/_118_  (.A1(\u_multiplier/_0844_ ),
    .A2(\u_multiplier/_0845_ ),
    .A3(\u_multiplier/dec/_073_ ),
    .ZN(\u_multiplier/dec/_085_ ));
 NOR2_X1 \u_multiplier/dec/_119_  (.A1(\u_multiplier/_0846_ ),
    .A2(\u_multiplier/dec/_085_ ),
    .ZN(\u_multiplier/dec_out [12]));
 NAND4_X1 \u_multiplier/dec/_120_  (.A1(\u_multiplier/_0842_ ),
    .A2(\u_multiplier/dec/_070_ ),
    .A3(\u_multiplier/_0844_ ),
    .A4(\u_multiplier/_0845_ ),
    .ZN(\u_multiplier/dec/_086_ ));
 NOR2_X1 \u_multiplier/dec/_121_  (.A1(\u_multiplier/_0846_ ),
    .A2(\u_multiplier/dec/_086_ ),
    .ZN(\u_multiplier/dec_out [13]));
 NAND4_X1 \u_multiplier/dec/_122_  (.A1(\u_multiplier/dec/_069_ ),
    .A2(\u_multiplier/_0843_ ),
    .A3(\u_multiplier/_0844_ ),
    .A4(\u_multiplier/_0845_ ),
    .ZN(\u_multiplier/dec/_087_ ));
 NOR2_X1 \u_multiplier/dec/_123_  (.A1(\u_multiplier/_0846_ ),
    .A2(\u_multiplier/dec/_087_ ),
    .ZN(\u_multiplier/dec_out [14]));
 OR2_X1 \u_multiplier/dec/_124_  (.A1(\u_multiplier/dec/_072_ ),
    .A2(\u_multiplier/dec/_081_ ),
    .ZN(\u_multiplier/dec/_088_ ));
 NOR2_X1 \u_multiplier/dec/_125_  (.A1(\u_multiplier/_0846_ ),
    .A2(\u_multiplier/dec/_088_ ),
    .ZN(\u_multiplier/dec_out [15]));
 NOR3_X1 \u_multiplier/dec/_126_  (.A1(\u_multiplier/dec/_068_ ),
    .A2(\u_multiplier/_0845_ ),
    .A3(\u_multiplier/dec/_074_ ),
    .ZN(\u_multiplier/dec_out [16]));
 NOR4_X2 \u_multiplier/dec/_127_  (.A1(\u_multiplier/dec/_068_ ),
    .A2(\u_multiplier/_0844_ ),
    .A3(\u_multiplier/_0845_ ),
    .A4(\u_multiplier/dec/_075_ ),
    .ZN(\u_multiplier/dec_out [17]));
 NOR4_X1 \u_multiplier/dec/_128_  (.A1(\u_multiplier/dec/_068_ ),
    .A2(\u_multiplier/_0844_ ),
    .A3(\u_multiplier/_0845_ ),
    .A4(\u_multiplier/dec/_076_ ),
    .ZN(\u_multiplier/dec_out [18]));
 NOR4_X1 \u_multiplier/dec/_129_  (.A1(\u_multiplier/dec/_068_ ),
    .A2(\u_multiplier/_0844_ ),
    .A3(\u_multiplier/_0845_ ),
    .A4(\u_multiplier/dec/_077_ ),
    .ZN(\u_multiplier/dec_out [19]));
 NOR3_X1 \u_multiplier/dec/_130_  (.A1(\u_multiplier/dec/_068_ ),
    .A2(\u_multiplier/_0845_ ),
    .A3(\u_multiplier/dec/_078_ ),
    .ZN(\u_multiplier/dec_out [20]));
 NOR3_X1 \u_multiplier/dec/_131_  (.A1(\u_multiplier/dec/_068_ ),
    .A2(\u_multiplier/_0845_ ),
    .A3(\u_multiplier/dec/_079_ ),
    .ZN(\u_multiplier/dec_out [21]));
 NOR3_X1 \u_multiplier/dec/_132_  (.A1(\u_multiplier/dec/_068_ ),
    .A2(\u_multiplier/_0845_ ),
    .A3(\u_multiplier/dec/_080_ ),
    .ZN(\u_multiplier/dec_out [22]));
 NOR3_X1 \u_multiplier/dec/_133_  (.A1(\u_multiplier/dec/_068_ ),
    .A2(\u_multiplier/_0845_ ),
    .A3(\u_multiplier/dec/_081_ ),
    .ZN(\u_multiplier/dec_out [23]));
 NOR2_X1 \u_multiplier/dec/_134_  (.A1(\u_multiplier/dec/_068_ ),
    .A2(\u_multiplier/dec/_082_ ),
    .ZN(\u_multiplier/dec_out [24]));
 NOR2_X1 \u_multiplier/dec/_135_  (.A1(\u_multiplier/dec/_068_ ),
    .A2(\u_multiplier/dec/_083_ ),
    .ZN(\u_multiplier/dec_out [25]));
 NOR2_X1 \u_multiplier/dec/_136_  (.A1(\u_multiplier/dec/_068_ ),
    .A2(\u_multiplier/dec/_084_ ),
    .ZN(\u_multiplier/dec_out [26]));
 NOR4_X1 \u_multiplier/dec/_137_  (.A1(\u_multiplier/dec/_068_ ),
    .A2(\u_multiplier/_0844_ ),
    .A3(\u_multiplier/dec/_072_ ),
    .A4(\u_multiplier/dec/_077_ ),
    .ZN(\u_multiplier/dec_out [27]));
 NOR2_X1 \u_multiplier/dec/_138_  (.A1(\u_multiplier/dec/_068_ ),
    .A2(\u_multiplier/dec/_085_ ),
    .ZN(\u_multiplier/dec_out [28]));
 NOR2_X1 \u_multiplier/dec/_139_  (.A1(\u_multiplier/dec/_068_ ),
    .A2(\u_multiplier/dec/_086_ ),
    .ZN(\u_multiplier/dec_out [29]));
 NOR2_X1 \u_multiplier/dec/_140_  (.A1(\u_multiplier/dec/_068_ ),
    .A2(\u_multiplier/dec/_087_ ),
    .ZN(\u_multiplier/dec_out [30]));
 NOR2_X1 \u_multiplier/dec/_141_  (.A1(\u_multiplier/dec/_068_ ),
    .A2(\u_multiplier/dec/_088_ ),
    .ZN(\u_multiplier/dec_out [31]));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_2_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_2_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_2_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_2_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_2_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_2_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_2_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_2_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_2_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_2_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_2_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_2_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_2_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_2_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_2_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_2_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_2_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_2_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_2_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_2_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_2_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_2_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_2_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_2_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_2_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_2_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_2_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_2_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_2_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_2_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_2_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_2_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_2_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_2_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_2_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_2_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_2_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_2_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_2_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_2_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_2_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_2_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_2_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_2_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_2_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_2_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_2_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_2_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_2_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_2_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_2_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_2_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_2_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_2_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_2_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_2_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_2_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_2_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_2_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_2_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_2_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_2_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_2_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_2_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_2_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_2_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_2_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_2_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_2_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_2_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_2_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_2_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_2_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_2_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_2_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_2_Right_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_2_Right_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_2_Right_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_2_Right_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_2_Right_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_2_Right_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_2_Right_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_2_Right_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_2_Right_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_2_Right_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_2_Right_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_2_Right_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_2_Right_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_2_Right_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_2_Right_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_2_Right_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_2_Right_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_2_Right_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_2_Right_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_2_Right_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_2_Right_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_2_Right_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_2_Right_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_2_Right_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_2_Right_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_2_Right_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_2_Right_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_2_Right_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_2_Right_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_2_Right_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_1_Left_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_1_Left_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_1_Left_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_1_Left_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_1_Left_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_1_Left_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_1_Left_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_1_Left_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_1_Left_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_1_Left_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_1_Left_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_1_Left_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_1_Left_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_1_Left_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_1_Left_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_1_Left_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_1_Left_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_1_Left_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_1_Left_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_1_Left_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_1_Left_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_1_Left_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_1_Left_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_1_Left_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_1_Left_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_1_Left_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_1_Left_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_1_Left_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_1_Left_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_1_Left_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_1_Left_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_1_Left_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_1_Left_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_1_Left_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_1_Left_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_1_Left_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_1_Left_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_1_Left_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_1_Left_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_1_Left_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_1_Left_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_1_Left_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_1_Left_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_1_Left_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_1_Left_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_1_Left_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_1_Left_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_1_Left_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_1_Left_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_1_Left_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_1_Left_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_1_Left_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_1_Left_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_1_Left_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_1_Left_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_1_Left_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_1_Left_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_1_Left_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_1_Left_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_1_Left_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_1_Left_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_1_Left_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_1_Left_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_1_Left_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_1_Left_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_1_Left_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_1_Left_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_1_Left_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_1_Left_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_1_Left_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_1_Left_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_1_Left_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_1_Left_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_1_Left_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_1_Left_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_1_Left_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_1_Left_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_1_Left_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_1_Left_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_1_Left_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_1_Left_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_1_Left_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_1_Left_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_1_Left_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_1_Left_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_1_Left_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_1_Left_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_1_Left_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_1_Left_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_1_Left_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_1_Left_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_1_Left_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_1_Left_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_1_Left_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_1_Left_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_1_Left_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_1_Left_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_1_Left_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_1_Left_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_1_Left_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_1_Left_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_1_Left_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_1_Left_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_1_Left_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Left_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Left_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Left_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Left_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Left_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Left_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Left_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Left_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Left_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Left_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Left_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Left_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Left_265 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Left_266 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Left_267 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Left_268 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Left_269 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Left_270 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Left_271 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Left_272 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_1_Left_273 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_2_Left_274 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_2_Left_275 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_2_Left_276 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_2_Left_277 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_2_Left_278 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_2_Left_279 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_2_Left_280 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_2_Left_281 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_2_Left_282 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_2_Left_283 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_2_Left_284 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_2_Left_285 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_2_Left_286 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_2_Left_287 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_2_Left_288 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_2_Left_289 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_2_Left_290 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_2_Left_291 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_2_Left_292 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_2_Left_293 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_2_Left_294 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_2_Left_295 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_2_Left_296 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_2_Left_297 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_2_Left_298 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_2_Left_299 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_2_Left_300 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_2_Left_301 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_2_Left_302 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_2_Left_303 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_2_Left_304 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_2_Left_305 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_2_Left_306 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_2_Left_307 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_2_Left_308 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_2_Left_309 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_2_Left_310 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_2_Left_311 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_2_Left_312 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_2_Left_313 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_2_Left_314 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_2_Left_315 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_2_Left_316 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_2_Left_317 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_2_Left_318 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_2_Left_319 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_2_Left_320 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_2_Left_321 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_2_Left_322 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_2_Left_323 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_2_Left_324 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_2_Left_325 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_2_Left_326 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_2_Left_327 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_2_Left_328 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_2_Left_329 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_2_Left_330 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_2_Left_331 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_2_Left_332 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_2_Left_333 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_2_Left_334 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_2_Left_335 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_2_Left_336 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_2_Left_337 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_2_Left_338 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_2_Left_339 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_2_Left_340 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_2_Left_341 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_2_Left_342 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_2_Left_343 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_2_Left_344 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_2_Left_345 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_2_Left_346 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_2_Left_347 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_2_Left_348 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_2_Left_349 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_2_Left_350 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_2_Left_351 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_2_Left_352 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_2_Left_353 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_2_Left_354 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_2_Left_355 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_2_Left_356 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_2_Left_357 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_2_Left_358 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_2_Left_359 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_2_Left_360 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_2_Left_361 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_2_Left_362 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_2_Left_363 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_2_Left_364 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_2_Left_365 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_2_Left_366 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_2_Left_367 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_2_Left_368 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_2_Left_369 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_2_Left_370 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_2_Left_371 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_2_Left_372 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_2_Left_373 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_2_Left_374 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_2_Left_375 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_2_Left_376 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_2_Left_377 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_2_Left_378 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_1_Right_379 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_1_Right_380 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_1_Right_381 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_1_Right_382 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_1_Right_383 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_1_Right_384 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_1_Right_385 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_1_Right_386 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_1_Right_387 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_1_Right_388 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_1_Right_389 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_1_Right_390 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_1_Right_391 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_1_Right_392 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_1_Right_393 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_1_Right_394 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_1_Right_395 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_1_Right_396 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_1_Right_397 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_1_Right_398 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_1_Right_399 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_1_Right_400 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_1_Right_401 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_1_Right_402 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_1_Right_403 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_1_Right_404 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_1_Right_405 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_1_Right_406 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_1_Right_407 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_1_Right_408 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_1_Right_409 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_1_Right_410 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_1_Right_411 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_1_Right_412 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_1_Right_413 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_1_Right_414 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_1_Right_415 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_1_Right_416 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_1_Right_417 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_1_Right_418 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_1_Right_419 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_1_Right_420 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_1_Right_421 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_1_Right_422 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_1_Right_423 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_1_Right_424 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_1_Right_425 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_1_Right_426 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_1_Right_427 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_1_Right_428 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_1_Right_429 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_1_Right_430 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_1_Right_431 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_1_Right_432 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_1_Right_433 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_1_Right_434 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_1_Right_435 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_1_Right_436 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_1_Right_437 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_1_Right_438 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_1_Right_439 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_1_Right_440 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_1_Right_441 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_1_Right_442 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_1_Right_443 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_1_Right_444 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_1_Right_445 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_1_Right_446 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_1_Right_447 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_1_Right_448 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_1_Right_449 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_1_Right_450 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_1_Right_451 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_1_Right_452 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_1_Right_453 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_1_Right_454 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_1_Right_455 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_1_Right_456 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_1_Right_457 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_1_Right_458 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_1_Right_459 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_1_Right_460 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_1_Right_461 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_1_Right_462 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_1_Right_463 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_1_Right_464 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_1_Right_465 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_1_Right_466 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_1_Right_467 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_1_Right_468 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_1_Right_469 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_1_Right_470 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_1_Right_471 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_1_Right_472 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_1_Right_473 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_1_Right_474 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_1_Right_475 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_1_Right_476 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_1_Right_477 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_1_Right_478 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_1_Right_479 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_1_Right_480 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_1_Right_481 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_1_Right_482 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_1_Right_483 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_484 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_485 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_486 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_487 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_488 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_489 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_490 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_117_491 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_492 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_493 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_494 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_495 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_496 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_497 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_498 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_499 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_500 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_501 ();
 LOGIC1_X1 \u_multiplier/NOD/nod_cels[13].Nod_bits/_07__55  (.Z(net55));
 CLKBUF_X1 hold56 (.A(net130),
    .Z(net56));
 BUF_X1 input2 (.A(data_in[0]),
    .Z(net2));
 BUF_X2 input3 (.A(data_in[10]),
    .Z(net3));
 BUF_X1 input4 (.A(data_in[11]),
    .Z(net4));
 BUF_X2 input5 (.A(data_in[12]),
    .Z(net5));
 BUF_X1 input6 (.A(data_in[13]),
    .Z(net6));
 BUF_X2 input7 (.A(data_in[14]),
    .Z(net7));
 CLKBUF_X3 input8 (.A(data_in[15]),
    .Z(net8));
 CLKBUF_X3 input9 (.A(data_in[1]),
    .Z(net9));
 BUF_X1 input10 (.A(data_in[2]),
    .Z(net10));
 BUF_X2 input11 (.A(data_in[3]),
    .Z(net11));
 BUF_X2 input12 (.A(data_in[4]),
    .Z(net12));
 BUF_X1 input13 (.A(data_in[5]),
    .Z(net13));
 BUF_X1 input14 (.A(data_in[6]),
    .Z(net14));
 BUF_X1 input15 (.A(data_in[7]),
    .Z(net15));
 CLKBUF_X3 input16 (.A(data_in[8]),
    .Z(net16));
 BUF_X2 input17 (.A(data_in[9]),
    .Z(net17));
 CLKBUF_X3 input18 (.A(init_enable),
    .Z(net18));
 CLKBUF_X3 input19 (.A(pe_ce),
    .Z(net19));
 BUF_X8 input20 (.A(rst_n),
    .Z(net20));
 BUF_X1 output21 (.A(net21),
    .Z(curr_state[1]));
 BUF_X1 output22 (.A(net22),
    .Z(data_out[0]));
 BUF_X1 output23 (.A(net23),
    .Z(data_out[10]));
 BUF_X1 output24 (.A(net24),
    .Z(data_out[11]));
 BUF_X1 output25 (.A(net25),
    .Z(data_out[12]));
 BUF_X1 output26 (.A(net26),
    .Z(data_out[13]));
 BUF_X1 output27 (.A(net27),
    .Z(data_out[14]));
 BUF_X1 output28 (.A(net28),
    .Z(data_out[15]));
 BUF_X1 output29 (.A(net29),
    .Z(data_out[16]));
 BUF_X1 output30 (.A(net30),
    .Z(data_out[17]));
 BUF_X1 output31 (.A(net31),
    .Z(data_out[18]));
 BUF_X1 output32 (.A(net32),
    .Z(data_out[19]));
 BUF_X1 output33 (.A(net33),
    .Z(data_out[1]));
 BUF_X1 output34 (.A(net34),
    .Z(data_out[20]));
 BUF_X1 output35 (.A(net35),
    .Z(data_out[21]));
 BUF_X1 output36 (.A(net36),
    .Z(data_out[22]));
 BUF_X1 output37 (.A(net37),
    .Z(data_out[23]));
 BUF_X1 output38 (.A(net38),
    .Z(data_out[24]));
 BUF_X1 output39 (.A(net39),
    .Z(data_out[25]));
 BUF_X1 output40 (.A(net40),
    .Z(data_out[26]));
 BUF_X1 output41 (.A(net41),
    .Z(data_out[27]));
 BUF_X1 output42 (.A(net42),
    .Z(data_out[28]));
 BUF_X1 output43 (.A(net43),
    .Z(data_out[29]));
 BUF_X1 output44 (.A(net44),
    .Z(data_out[2]));
 BUF_X1 output45 (.A(net45),
    .Z(data_out[30]));
 BUF_X1 output46 (.A(net46),
    .Z(data_out[31]));
 BUF_X1 output47 (.A(net47),
    .Z(data_out[3]));
 BUF_X1 output48 (.A(net48),
    .Z(data_out[4]));
 BUF_X1 output49 (.A(net49),
    .Z(data_out[5]));
 BUF_X1 output50 (.A(net50),
    .Z(data_out[6]));
 BUF_X1 output51 (.A(net51),
    .Z(data_out[7]));
 BUF_X1 output52 (.A(net52),
    .Z(data_out[8]));
 BUF_X1 output53 (.A(net53),
    .Z(data_out[9]));
 BUF_X1 output54 (.A(net54),
    .Z(valid_reg_out));
 CLKBUF_X1 hold57 (.A(_174_),
    .Z(net57));
 CLKBUF_X1 hold58 (.A(net77),
    .Z(net58));
 CLKBUF_X1 hold59 (.A(net83),
    .Z(net59));
 CLKBUF_X1 hold60 (.A(net105),
    .Z(net60));
 CLKBUF_X1 hold61 (.A(net102),
    .Z(net61));
 CLKBUF_X1 hold62 (.A(net80),
    .Z(net62));
 CLKBUF_X1 hold63 (.A(net87),
    .Z(net63));
 CLKBUF_X1 hold64 (.A(net100),
    .Z(net64));
 CLKBUF_X1 hold65 (.A(net108),
    .Z(net65));
 CLKBUF_X1 hold66 (.A(net111),
    .Z(net66));
 CLKBUF_X1 hold67 (.A(net116),
    .Z(net67));
 CLKBUF_X1 hold68 (.A(net119),
    .Z(net68));
 CLKBUF_X1 hold69 (.A(net124),
    .Z(net69));
 CLKBUF_X1 hold70 (.A(net122),
    .Z(net70));
 CLKBUF_X1 hold71 (.A(net127),
    .Z(net71));
 CLKBUF_X1 hold72 (.A(net132),
    .Z(net72));
 CLKBUF_X1 hold73 (.A(net133),
    .Z(net73));
 CLKBUF_X1 hold74 (.A(net131),
    .Z(net74));
 CLKBUF_X1 hold75 (.A(net129),
    .Z(net75));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_2_0_0_clk));
 CLKBUF_X3 clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_2_1_0_clk));
 CLKBUF_X3 clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .Z(clknet_2_2_0_clk));
 CLKBUF_X3 clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .Z(clknet_2_3_0_clk));
 CLKBUF_X3 clkbuf_3_0_0_clk (.A(clknet_2_0_0_clk),
    .Z(clknet_3_0_0_clk));
 CLKBUF_X3 clkbuf_3_1_0_clk (.A(clknet_2_0_0_clk),
    .Z(clknet_3_1_0_clk));
 CLKBUF_X3 clkbuf_3_2_0_clk (.A(clknet_2_1_0_clk),
    .Z(clknet_3_2_0_clk));
 CLKBUF_X3 clkbuf_3_3_0_clk (.A(clknet_2_1_0_clk),
    .Z(clknet_3_3_0_clk));
 CLKBUF_X3 clkbuf_3_4_0_clk (.A(clknet_2_2_0_clk),
    .Z(clknet_3_4_0_clk));
 CLKBUF_X3 clkbuf_3_5_0_clk (.A(clknet_2_2_0_clk),
    .Z(clknet_3_5_0_clk));
 CLKBUF_X3 clkbuf_3_6_0_clk (.A(clknet_2_3_0_clk),
    .Z(clknet_3_6_0_clk));
 CLKBUF_X3 clkbuf_3_7_0_clk (.A(clknet_2_3_0_clk),
    .Z(clknet_3_7_0_clk));
 INV_X2 clkload0 (.A(clknet_3_0_0_clk));
 INV_X2 clkload1 (.A(clknet_3_2_0_clk));
 INV_X1 clkload2 (.A(clknet_3_4_0_clk));
 INV_X2 clkload3 (.A(clknet_3_6_0_clk));
 CLKBUF_X1 hold1 (.A(net134),
    .Z(net1));
 CLKBUF_X1 hold2 (.A(net135),
    .Z(net76));
 CLKBUF_X1 hold3 (.A(_401_),
    .Z(net77));
 CLKBUF_X1 hold4 (.A(net58),
    .Z(net78));
 CLKBUF_X1 hold5 (.A(_119_),
    .Z(net79));
 CLKBUF_X1 hold6 (.A(addr_ptr[4]),
    .Z(net80));
 CLKBUF_X1 hold7 (.A(net62),
    .Z(net81));
 CLKBUF_X1 hold8 (.A(net137),
    .Z(net82));
 CLKBUF_X1 hold9 (.A(_400_),
    .Z(net83));
 CLKBUF_X1 hold10 (.A(net59),
    .Z(net84));
 CLKBUF_X1 hold11 (.A(_118_),
    .Z(net85));
 CLKBUF_X1 hold12 (.A(net136),
    .Z(net86));
 CLKBUF_X1 hold13 (.A(addr_ptr[1]),
    .Z(net87));
 CLKBUF_X1 hold14 (.A(net63),
    .Z(net88));
 CLKBUF_X1 hold15 (.A(net141),
    .Z(net89));
 CLKBUF_X1 hold16 (.A(_403_),
    .Z(net90));
 CLKBUF_X1 hold17 (.A(_279_),
    .Z(net91));
 CLKBUF_X1 hold18 (.A(_121_),
    .Z(net92));
 CLKBUF_X1 hold19 (.A(curr_state[0]),
    .Z(net93));
 CLKBUF_X1 hold20 (.A(_240_),
    .Z(net94));
 CLKBUF_X1 hold21 (.A(net138),
    .Z(net95));
 CLKBUF_X1 hold22 (.A(net140),
    .Z(net96));
 CLKBUF_X1 hold23 (.A(_404_),
    .Z(net97));
 CLKBUF_X1 hold24 (.A(_281_),
    .Z(net98));
 CLKBUF_X1 hold25 (.A(net139),
    .Z(net99));
 CLKBUF_X1 hold26 (.A(addr_ptr[3]),
    .Z(net100));
 CLKBUF_X1 hold27 (.A(net64),
    .Z(net101));
 CLKBUF_X1 hold28 (.A(_407_),
    .Z(net102));
 CLKBUF_X1 hold29 (.A(net61),
    .Z(net103));
 CLKBUF_X1 hold30 (.A(_173_),
    .Z(net104));
 CLKBUF_X1 hold31 (.A(_406_),
    .Z(net105));
 CLKBUF_X1 hold32 (.A(net60),
    .Z(net106));
 CLKBUF_X1 hold33 (.A(_172_),
    .Z(net107));
 CLKBUF_X1 hold34 (.A(addr_ptr[2]),
    .Z(net108));
 CLKBUF_X1 hold35 (.A(net65),
    .Z(net109));
 CLKBUF_X1 hold36 (.A(\u_multiplier/LODx/z [7]),
    .Z(net110));
 CLKBUF_X1 hold37 (.A(addr_ptr[0]),
    .Z(net111));
 CLKBUF_X1 hold38 (.A(net66),
    .Z(net112));
 CLKBUF_X1 hold39 (.A(data_in_reg[0]),
    .Z(net113));
 CLKBUF_X1 hold40 (.A(curr_state[2]),
    .Z(net114));
 CLKBUF_X1 hold41 (.A(_195_),
    .Z(net115));
 CLKBUF_X1 hold42 (.A(_405_),
    .Z(net116));
 CLKBUF_X1 hold43 (.A(net67),
    .Z(net117));
 CLKBUF_X1 hold44 (.A(_171_),
    .Z(net118));
 CLKBUF_X1 hold45 (.A(_402_),
    .Z(net119));
 CLKBUF_X1 hold46 (.A(net68),
    .Z(net120));
 CLKBUF_X1 hold47 (.A(_120_),
    .Z(net121));
 CLKBUF_X1 hold48 (.A(\u_multiplier/LODx/z [15]),
    .Z(net122));
 CLKBUF_X1 hold49 (.A(net70),
    .Z(net123));
 CLKBUF_X1 hold50 (.A(_409_),
    .Z(net124));
 CLKBUF_X1 hold51 (.A(net69),
    .Z(net125));
 CLKBUF_X1 hold52 (.A(_175_),
    .Z(net126));
 CLKBUF_X1 hold53 (.A(data_in_reg[13]),
    .Z(net127));
 CLKBUF_X1 hold54 (.A(net71),
    .Z(net128));
 CLKBUF_X1 hold55 (.A(data_in_reg[5]),
    .Z(net129));
 CLKBUF_X1 hold76 (.A(_408_),
    .Z(net130));
 CLKBUF_X1 hold77 (.A(data_in_reg[10]),
    .Z(net131));
 CLKBUF_X1 hold78 (.A(data_in_reg[4]),
    .Z(net132));
 CLKBUF_X1 hold79 (.A(data_in_reg[12]),
    .Z(net133));
 CLKBUF_X1 hold80 (.A(data_in_reg[14]),
    .Z(net134));
 CLKBUF_X1 hold81 (.A(\u_multiplier/LODx/z [3]),
    .Z(net135));
 CLKBUF_X1 hold82 (.A(data_in_reg[1]),
    .Z(net136));
 CLKBUF_X1 hold83 (.A(\u_multiplier/LODx/z [11]),
    .Z(net137));
 CLKBUF_X1 hold84 (.A(data_in_reg[8]),
    .Z(net138));
 CLKBUF_X1 hold85 (.A(data_in_reg[9]),
    .Z(net139));
 CLKBUF_X1 hold86 (.A(data_in_reg[2]),
    .Z(net140));
 CLKBUF_X1 hold87 (.A(data_in_reg[6]),
    .Z(net141));
 assign init_done = curr_state[1];
 assign valid_out = valid_reg_out;
endmodule
