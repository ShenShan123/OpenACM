module sram_multiplier_system (clk,
    init_done,
    init_enable,
    pe_ce,
    rst_n,
    valid_out,
    data_in,
    data_out);
 input clk;
 output init_done;
 input init_enable;
 input pe_ce;
 input rst_n;
 output valid_out;
 input [31:0] data_in;
 output [63:0] data_out;

 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net142;
 wire net150;
 wire u_multiplier_pp1_0 ;
 wire u_multiplier_pp1_62 ;
 wire u_multiplier_pp2_0 ;
 wire u_multiplier_pp2_62 ;
 wire u_multiplier_pp3_0 ;
 wire u_multiplier_pp3_62 ;
 wire u_multiplier_Final_add_Cout ;
 wire u_multiplier_Final_add_c1 ;
 wire u_multiplier_Final_add_cla1_c1 ;
 wire u_multiplier_Final_add_cla1_cla1_c1 ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_c1 ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__25_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__26_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__27_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__28_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__29_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__30_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__31_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__32_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__33_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__34_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__35_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__36_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__37_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__38_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla1__39_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__25_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__26_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__27_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__28_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__29_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__30_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__31_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__32_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__33_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__34_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__35_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__36_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__37_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__38_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla1_cla2__39_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_c1 ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__25_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__26_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__27_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__28_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__29_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__30_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__31_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__32_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__33_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__34_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__35_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__36_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__37_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__38_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla1__39_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__25_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__26_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__27_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__28_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__29_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__30_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__31_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__32_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__33_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__34_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__35_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__36_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__37_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__38_ ;
 wire u_multiplier_Final_add_cla1_cla1_cla2_cla2__39_ ;
 wire u_multiplier_Final_add_cla1_cla2_c1 ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_c1 ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__25_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__26_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__27_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__28_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__29_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__30_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__31_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__32_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__33_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__34_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__35_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__36_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__37_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__38_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla1__39_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__25_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__26_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__27_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__28_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__29_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__30_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__31_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__32_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__33_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__34_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__35_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__36_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__37_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__38_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla1_cla2__39_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_c1 ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__25_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__26_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__27_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__28_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__29_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__30_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__31_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__32_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__33_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__34_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__35_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__36_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__37_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__38_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla1__39_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__25_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__26_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__27_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__28_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__29_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__30_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__31_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__32_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__33_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__34_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__35_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__36_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__37_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__38_ ;
 wire u_multiplier_Final_add_cla1_cla2_cla2_cla2__39_ ;
 wire u_multiplier_Final_add_cla2_c1 ;
 wire u_multiplier_Final_add_cla2_cla1_c1 ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_c1 ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__25_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__26_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__27_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__28_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__29_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__30_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__31_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__32_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__33_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__34_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__35_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__36_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__37_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__38_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla1__39_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__25_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__26_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__27_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__28_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__29_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__30_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__31_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__32_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__33_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__34_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__35_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__36_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__37_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__38_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla1_cla2__39_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_c1 ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__25_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__26_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__27_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__28_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__29_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__30_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__31_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__32_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__33_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__34_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__35_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__36_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__37_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__38_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla1__39_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__25_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__26_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__27_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__28_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__29_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__30_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__31_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__32_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__33_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__34_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__35_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__36_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__37_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__38_ ;
 wire u_multiplier_Final_add_cla2_cla1_cla2_cla2__39_ ;
 wire u_multiplier_Final_add_cla2_cla2_c1 ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_c1 ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__25_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__26_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__27_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__28_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__29_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__30_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__31_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__32_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__33_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__34_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__35_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__36_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__37_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__38_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla1__39_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__25_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__26_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__27_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__28_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__29_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__30_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__31_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__32_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__33_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__34_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__35_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__36_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__37_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__38_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla1_cla2__39_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_c1 ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__25_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__26_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__27_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__28_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__29_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__30_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__31_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__32_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__33_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__34_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__35_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__36_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__37_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__38_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla1__39_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__25_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__26_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__27_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__28_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__29_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__30_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__31_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__32_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__33_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__34_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__35_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__36_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__37_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__38_ ;
 wire u_multiplier_Final_add_cla2_cla2_cla2_cla2__39_ ;
 wire u_multiplier_STAGE1__0607_ ;
 wire u_multiplier_STAGE1__0608_ ;
 wire u_multiplier_STAGE1__0609_ ;
 wire u_multiplier_STAGE1__0610_ ;
 wire u_multiplier_STAGE1__0611_ ;
 wire u_multiplier_STAGE1__0612_ ;
 wire u_multiplier_STAGE1__0613_ ;
 wire u_multiplier_STAGE1__0614_ ;
 wire u_multiplier_STAGE1__0615_ ;
 wire u_multiplier_STAGE1__0616_ ;
 wire u_multiplier_STAGE1__0617_ ;
 wire u_multiplier_STAGE1__0618_ ;
 wire u_multiplier_STAGE1__0619_ ;
 wire u_multiplier_STAGE1__0620_ ;
 wire u_multiplier_STAGE1__0621_ ;
 wire u_multiplier_STAGE1__0622_ ;
 wire u_multiplier_STAGE1__0623_ ;
 wire u_multiplier_STAGE1__0624_ ;
 wire u_multiplier_STAGE1__0625_ ;
 wire u_multiplier_STAGE1__0626_ ;
 wire u_multiplier_STAGE1__0627_ ;
 wire u_multiplier_STAGE1__0628_ ;
 wire u_multiplier_STAGE1__0629_ ;
 wire u_multiplier_STAGE1__0630_ ;
 wire u_multiplier_STAGE1__0631_ ;
 wire u_multiplier_STAGE1__0632_ ;
 wire u_multiplier_STAGE1__0633_ ;
 wire u_multiplier_STAGE1__0634_ ;
 wire u_multiplier_STAGE1__0635_ ;
 wire u_multiplier_STAGE1__0636_ ;
 wire u_multiplier_STAGE1__0637_ ;
 wire u_multiplier_STAGE1__0638_ ;
 wire u_multiplier_STAGE1__0639_ ;
 wire u_multiplier_STAGE1__0640_ ;
 wire u_multiplier_STAGE1__0641_ ;
 wire u_multiplier_STAGE1__0642_ ;
 wire u_multiplier_STAGE1__0643_ ;
 wire u_multiplier_STAGE1__0644_ ;
 wire u_multiplier_STAGE1__0645_ ;
 wire u_multiplier_STAGE1__0646_ ;
 wire u_multiplier_STAGE1__0647_ ;
 wire u_multiplier_STAGE1__0648_ ;
 wire u_multiplier_STAGE1__0649_ ;
 wire u_multiplier_STAGE1__0650_ ;
 wire u_multiplier_STAGE1__0651_ ;
 wire u_multiplier_STAGE1__0652_ ;
 wire u_multiplier_STAGE1__0653_ ;
 wire u_multiplier_STAGE1__0654_ ;
 wire u_multiplier_STAGE1__0655_ ;
 wire u_multiplier_STAGE1__0656_ ;
 wire u_multiplier_STAGE1__0657_ ;
 wire u_multiplier_STAGE1__0658_ ;
 wire u_multiplier_STAGE1__0659_ ;
 wire u_multiplier_STAGE1__0660_ ;
 wire u_multiplier_STAGE1__0661_ ;
 wire u_multiplier_STAGE1__0662_ ;
 wire u_multiplier_STAGE1__0663_ ;
 wire u_multiplier_STAGE1__0664_ ;
 wire u_multiplier_STAGE1__0665_ ;
 wire u_multiplier_STAGE1__0666_ ;
 wire u_multiplier_STAGE1__0667_ ;
 wire u_multiplier_STAGE1__0668_ ;
 wire u_multiplier_STAGE1__0669_ ;
 wire u_multiplier_STAGE1__0670_ ;
 wire u_multiplier_STAGE1__0671_ ;
 wire u_multiplier_STAGE1__0672_ ;
 wire u_multiplier_STAGE1__0673_ ;
 wire u_multiplier_STAGE1__0674_ ;
 wire u_multiplier_STAGE1__0675_ ;
 wire u_multiplier_STAGE1__0676_ ;
 wire u_multiplier_STAGE1__0677_ ;
 wire u_multiplier_STAGE1__0678_ ;
 wire u_multiplier_STAGE1__0679_ ;
 wire u_multiplier_STAGE1__0680_ ;
 wire u_multiplier_STAGE1__0681_ ;
 wire u_multiplier_STAGE1__0682_ ;
 wire u_multiplier_STAGE1__0683_ ;
 wire u_multiplier_STAGE1__0684_ ;
 wire u_multiplier_STAGE1__0685_ ;
 wire u_multiplier_STAGE1__0686_ ;
 wire u_multiplier_STAGE1__0687_ ;
 wire u_multiplier_STAGE1__0688_ ;
 wire u_multiplier_STAGE1__0689_ ;
 wire u_multiplier_STAGE1__0690_ ;
 wire u_multiplier_STAGE1__0691_ ;
 wire u_multiplier_STAGE1__0692_ ;
 wire u_multiplier_STAGE1__0693_ ;
 wire u_multiplier_STAGE1__0694_ ;
 wire u_multiplier_STAGE1__0695_ ;
 wire u_multiplier_STAGE1__0696_ ;
 wire u_multiplier_STAGE1__0697_ ;
 wire u_multiplier_STAGE1__0698_ ;
 wire u_multiplier_STAGE1__0699_ ;
 wire u_multiplier_STAGE1__0700_ ;
 wire u_multiplier_STAGE1__0701_ ;
 wire u_multiplier_STAGE1__0702_ ;
 wire u_multiplier_STAGE1__0703_ ;
 wire u_multiplier_STAGE1__0704_ ;
 wire u_multiplier_STAGE1__0705_ ;
 wire u_multiplier_STAGE1__0706_ ;
 wire u_multiplier_STAGE1__0707_ ;
 wire u_multiplier_STAGE1__0708_ ;
 wire u_multiplier_STAGE1__0709_ ;
 wire u_multiplier_STAGE1__0710_ ;
 wire u_multiplier_STAGE1__0711_ ;
 wire u_multiplier_STAGE1__0712_ ;
 wire u_multiplier_STAGE1__0713_ ;
 wire u_multiplier_STAGE1__0714_ ;
 wire u_multiplier_STAGE1__0715_ ;
 wire u_multiplier_STAGE1__0716_ ;
 wire u_multiplier_STAGE1__0717_ ;
 wire u_multiplier_STAGE1__0718_ ;
 wire u_multiplier_STAGE1__0719_ ;
 wire u_multiplier_STAGE1__0720_ ;
 wire u_multiplier_STAGE1__0721_ ;
 wire u_multiplier_STAGE1__0722_ ;
 wire u_multiplier_STAGE1__0723_ ;
 wire u_multiplier_STAGE1__0724_ ;
 wire u_multiplier_STAGE1__0725_ ;
 wire u_multiplier_STAGE1__0726_ ;
 wire u_multiplier_STAGE1__0727_ ;
 wire u_multiplier_STAGE1__0728_ ;
 wire u_multiplier_STAGE1__0729_ ;
 wire u_multiplier_STAGE1__0730_ ;
 wire u_multiplier_STAGE1__0731_ ;
 wire u_multiplier_STAGE1__0732_ ;
 wire u_multiplier_STAGE1__0733_ ;
 wire u_multiplier_STAGE1__0734_ ;
 wire u_multiplier_STAGE1__0735_ ;
 wire u_multiplier_STAGE1__0736_ ;
 wire u_multiplier_STAGE1__0737_ ;
 wire u_multiplier_STAGE1__0738_ ;
 wire u_multiplier_STAGE1__0739_ ;
 wire u_multiplier_STAGE1__0740_ ;
 wire u_multiplier_STAGE1__0741_ ;
 wire u_multiplier_STAGE1__0742_ ;
 wire u_multiplier_STAGE1__0743_ ;
 wire u_multiplier_STAGE1__0744_ ;
 wire u_multiplier_STAGE1__0745_ ;
 wire u_multiplier_STAGE1__0746_ ;
 wire u_multiplier_STAGE1__0747_ ;
 wire u_multiplier_STAGE1__0748_ ;
 wire u_multiplier_STAGE1__0749_ ;
 wire u_multiplier_STAGE1__0750_ ;
 wire u_multiplier_STAGE1__0751_ ;
 wire u_multiplier_STAGE1__0752_ ;
 wire u_multiplier_STAGE1__0753_ ;
 wire u_multiplier_STAGE1__0754_ ;
 wire u_multiplier_STAGE1__0755_ ;
 wire u_multiplier_STAGE1__0756_ ;
 wire u_multiplier_STAGE1__0757_ ;
 wire u_multiplier_STAGE1__0758_ ;
 wire u_multiplier_STAGE1__0759_ ;
 wire u_multiplier_STAGE1__0760_ ;
 wire u_multiplier_STAGE1__0761_ ;
 wire u_multiplier_STAGE1__0762_ ;
 wire u_multiplier_STAGE1__0763_ ;
 wire u_multiplier_STAGE1__0764_ ;
 wire u_multiplier_STAGE1__0765_ ;
 wire u_multiplier_STAGE1__0766_ ;
 wire u_multiplier_STAGE1__0767_ ;
 wire u_multiplier_STAGE1__0768_ ;
 wire u_multiplier_STAGE1__0769_ ;
 wire u_multiplier_STAGE1__0770_ ;
 wire u_multiplier_STAGE1__0771_ ;
 wire u_multiplier_STAGE1__0772_ ;
 wire u_multiplier_STAGE1__0773_ ;
 wire u_multiplier_STAGE1__0774_ ;
 wire u_multiplier_STAGE1__0775_ ;
 wire u_multiplier_STAGE1__0776_ ;
 wire u_multiplier_STAGE1__0777_ ;
 wire u_multiplier_STAGE1__0778_ ;
 wire u_multiplier_STAGE1__0779_ ;
 wire u_multiplier_STAGE1__0780_ ;
 wire u_multiplier_STAGE1__0781_ ;
 wire u_multiplier_STAGE1__0782_ ;
 wire u_multiplier_STAGE1__0783_ ;
 wire u_multiplier_STAGE1__0784_ ;
 wire u_multiplier_STAGE1__0785_ ;
 wire u_multiplier_STAGE1__0786_ ;
 wire u_multiplier_STAGE1__0787_ ;
 wire u_multiplier_STAGE1__0788_ ;
 wire u_multiplier_STAGE1__0789_ ;
 wire u_multiplier_STAGE1__0790_ ;
 wire u_multiplier_STAGE1__0791_ ;
 wire u_multiplier_STAGE1__0792_ ;
 wire u_multiplier_STAGE1__0793_ ;
 wire u_multiplier_STAGE1__0794_ ;
 wire u_multiplier_STAGE1__0795_ ;
 wire u_multiplier_STAGE1__0796_ ;
 wire u_multiplier_STAGE1__0797_ ;
 wire u_multiplier_STAGE1__0798_ ;
 wire u_multiplier_STAGE1__0799_ ;
 wire u_multiplier_STAGE1__0800_ ;
 wire u_multiplier_STAGE1__0801_ ;
 wire u_multiplier_STAGE1__0802_ ;
 wire u_multiplier_STAGE1__0803_ ;
 wire u_multiplier_STAGE1__0804_ ;
 wire u_multiplier_STAGE1__0805_ ;
 wire u_multiplier_STAGE1__0806_ ;
 wire u_multiplier_STAGE1__0807_ ;
 wire u_multiplier_STAGE1__0808_ ;
 wire u_multiplier_STAGE1__0809_ ;
 wire u_multiplier_STAGE1__0810_ ;
 wire u_multiplier_STAGE1__0811_ ;
 wire u_multiplier_STAGE1__0812_ ;
 wire u_multiplier_STAGE1__0813_ ;
 wire u_multiplier_STAGE1__0814_ ;
 wire u_multiplier_STAGE1__0815_ ;
 wire u_multiplier_STAGE1__0816_ ;
 wire u_multiplier_STAGE1__0817_ ;
 wire u_multiplier_STAGE1__0818_ ;
 wire u_multiplier_STAGE1__0819_ ;
 wire u_multiplier_STAGE1__0820_ ;
 wire u_multiplier_STAGE1__0821_ ;
 wire u_multiplier_STAGE1__0822_ ;
 wire u_multiplier_STAGE1__0823_ ;
 wire u_multiplier_STAGE1__0824_ ;
 wire u_multiplier_STAGE1__0825_ ;
 wire u_multiplier_STAGE1__0826_ ;
 wire u_multiplier_STAGE1__0827_ ;
 wire u_multiplier_STAGE1__0828_ ;
 wire u_multiplier_STAGE1__0829_ ;
 wire u_multiplier_STAGE1__0830_ ;
 wire u_multiplier_STAGE1__0831_ ;
 wire u_multiplier_STAGE1__0832_ ;
 wire u_multiplier_STAGE1__0833_ ;
 wire u_multiplier_STAGE1__0834_ ;
 wire u_multiplier_STAGE1__0835_ ;
 wire u_multiplier_STAGE1__0836_ ;
 wire u_multiplier_STAGE1__0837_ ;
 wire u_multiplier_STAGE1__0838_ ;
 wire u_multiplier_STAGE1__0839_ ;
 wire u_multiplier_STAGE1__0840_ ;
 wire u_multiplier_STAGE1__0841_ ;
 wire u_multiplier_STAGE1__0842_ ;
 wire u_multiplier_STAGE1__0843_ ;
 wire u_multiplier_STAGE1__0844_ ;
 wire u_multiplier_STAGE1__0845_ ;
 wire u_multiplier_STAGE1__0846_ ;
 wire u_multiplier_STAGE1__0847_ ;
 wire u_multiplier_STAGE1__0848_ ;
 wire u_multiplier_STAGE1__0849_ ;
 wire u_multiplier_STAGE1__0850_ ;
 wire u_multiplier_STAGE1__0851_ ;
 wire u_multiplier_STAGE1__0852_ ;
 wire u_multiplier_STAGE1__0853_ ;
 wire u_multiplier_STAGE1__0854_ ;
 wire u_multiplier_STAGE1__0855_ ;
 wire u_multiplier_STAGE1__0856_ ;
 wire u_multiplier_STAGE1__0857_ ;
 wire u_multiplier_STAGE1__0858_ ;
 wire u_multiplier_STAGE1__0859_ ;
 wire u_multiplier_STAGE1__0860_ ;
 wire u_multiplier_STAGE1__0861_ ;
 wire u_multiplier_STAGE1__0862_ ;
 wire u_multiplier_STAGE1__0863_ ;
 wire u_multiplier_STAGE1__0864_ ;
 wire u_multiplier_STAGE1__0865_ ;
 wire u_multiplier_STAGE1__0866_ ;
 wire u_multiplier_STAGE1__0867_ ;
 wire u_multiplier_STAGE1__0868_ ;
 wire u_multiplier_STAGE1__0869_ ;
 wire u_multiplier_STAGE1__0870_ ;
 wire u_multiplier_STAGE1__0871_ ;
 wire u_multiplier_STAGE1__0872_ ;
 wire u_multiplier_STAGE1__0873_ ;
 wire u_multiplier_STAGE1__0874_ ;
 wire u_multiplier_STAGE1__0875_ ;
 wire u_multiplier_STAGE1__0876_ ;
 wire u_multiplier_STAGE1__0877_ ;
 wire u_multiplier_STAGE1__0878_ ;
 wire u_multiplier_STAGE1__0879_ ;
 wire u_multiplier_STAGE1__0880_ ;
 wire u_multiplier_STAGE1__0881_ ;
 wire u_multiplier_STAGE1__0882_ ;
 wire u_multiplier_STAGE1__0883_ ;
 wire u_multiplier_STAGE1__0884_ ;
 wire u_multiplier_STAGE1__0885_ ;
 wire u_multiplier_STAGE1__0886_ ;
 wire u_multiplier_STAGE1__0887_ ;
 wire u_multiplier_STAGE1__0888_ ;
 wire u_multiplier_STAGE1__0889_ ;
 wire u_multiplier_STAGE1__0890_ ;
 wire u_multiplier_STAGE1__0891_ ;
 wire u_multiplier_STAGE1__0892_ ;
 wire u_multiplier_STAGE1__0893_ ;
 wire u_multiplier_STAGE1__0894_ ;
 wire u_multiplier_STAGE1__0895_ ;
 wire u_multiplier_STAGE1__0896_ ;
 wire u_multiplier_STAGE1__0897_ ;
 wire u_multiplier_STAGE1__0898_ ;
 wire u_multiplier_STAGE1__0899_ ;
 wire u_multiplier_STAGE1__0900_ ;
 wire u_multiplier_STAGE1__0901_ ;
 wire u_multiplier_STAGE1__0902_ ;
 wire u_multiplier_STAGE1__0903_ ;
 wire u_multiplier_STAGE1__0904_ ;
 wire u_multiplier_STAGE1__0905_ ;
 wire u_multiplier_STAGE1__0906_ ;
 wire u_multiplier_STAGE1__0907_ ;
 wire u_multiplier_STAGE1__0908_ ;
 wire u_multiplier_STAGE1__0909_ ;
 wire u_multiplier_STAGE1__0910_ ;
 wire u_multiplier_STAGE1__0911_ ;
 wire u_multiplier_STAGE1__0912_ ;
 wire u_multiplier_STAGE1__0913_ ;
 wire u_multiplier_STAGE1__0914_ ;
 wire u_multiplier_STAGE1__0915_ ;
 wire u_multiplier_STAGE1__0916_ ;
 wire u_multiplier_STAGE1__0917_ ;
 wire u_multiplier_STAGE1__0918_ ;
 wire u_multiplier_STAGE1__0919_ ;
 wire u_multiplier_STAGE1__0920_ ;
 wire u_multiplier_STAGE1__0921_ ;
 wire u_multiplier_STAGE1__0922_ ;
 wire u_multiplier_STAGE1__0923_ ;
 wire u_multiplier_STAGE1__0924_ ;
 wire u_multiplier_STAGE1__0925_ ;
 wire u_multiplier_STAGE1__0926_ ;
 wire u_multiplier_STAGE1__0927_ ;
 wire u_multiplier_STAGE1__0928_ ;
 wire u_multiplier_STAGE1__0929_ ;
 wire u_multiplier_STAGE1__0930_ ;
 wire u_multiplier_STAGE1__0931_ ;
 wire u_multiplier_STAGE1__0932_ ;
 wire u_multiplier_STAGE1__0933_ ;
 wire u_multiplier_STAGE1__0934_ ;
 wire u_multiplier_STAGE1__0935_ ;
 wire u_multiplier_STAGE1__0936_ ;
 wire u_multiplier_STAGE1__0937_ ;
 wire u_multiplier_STAGE1__0938_ ;
 wire u_multiplier_STAGE1__0939_ ;
 wire u_multiplier_STAGE1__0940_ ;
 wire u_multiplier_STAGE1__0941_ ;
 wire u_multiplier_STAGE1__0942_ ;
 wire u_multiplier_STAGE1__0943_ ;
 wire u_multiplier_STAGE1__0944_ ;
 wire u_multiplier_STAGE1__0945_ ;
 wire u_multiplier_STAGE1__0946_ ;
 wire u_multiplier_STAGE1__0947_ ;
 wire u_multiplier_STAGE1__0948_ ;
 wire u_multiplier_STAGE1__0949_ ;
 wire u_multiplier_STAGE1__0950_ ;
 wire u_multiplier_STAGE1__0951_ ;
 wire u_multiplier_STAGE1__0952_ ;
 wire u_multiplier_STAGE1__0953_ ;
 wire u_multiplier_STAGE1__0954_ ;
 wire u_multiplier_STAGE1__0955_ ;
 wire u_multiplier_STAGE1__0956_ ;
 wire u_multiplier_STAGE1__0957_ ;
 wire u_multiplier_STAGE1__0958_ ;
 wire u_multiplier_STAGE1__0959_ ;
 wire u_multiplier_STAGE1__0960_ ;
 wire u_multiplier_STAGE1__0961_ ;
 wire u_multiplier_STAGE1__0962_ ;
 wire u_multiplier_STAGE1__0963_ ;
 wire u_multiplier_STAGE1__0964_ ;
 wire u_multiplier_STAGE1__0965_ ;
 wire u_multiplier_STAGE1__0966_ ;
 wire u_multiplier_STAGE1__0967_ ;
 wire u_multiplier_STAGE1__0968_ ;
 wire u_multiplier_STAGE1__0969_ ;
 wire u_multiplier_STAGE1__0970_ ;
 wire u_multiplier_STAGE1__0971_ ;
 wire u_multiplier_STAGE1__0972_ ;
 wire u_multiplier_STAGE1__0973_ ;
 wire u_multiplier_STAGE1__0974_ ;
 wire u_multiplier_STAGE1__0975_ ;
 wire u_multiplier_STAGE1__0976_ ;
 wire u_multiplier_STAGE1__0977_ ;
 wire u_multiplier_STAGE1__0978_ ;
 wire u_multiplier_STAGE1__0979_ ;
 wire u_multiplier_STAGE1__0980_ ;
 wire u_multiplier_STAGE1__0981_ ;
 wire u_multiplier_STAGE1__0982_ ;
 wire u_multiplier_STAGE1__0983_ ;
 wire u_multiplier_STAGE1__0984_ ;
 wire u_multiplier_STAGE1__0985_ ;
 wire u_multiplier_STAGE1__0986_ ;
 wire u_multiplier_STAGE1__0987_ ;
 wire u_multiplier_STAGE1__0988_ ;
 wire u_multiplier_STAGE1__0989_ ;
 wire u_multiplier_STAGE1__0990_ ;
 wire u_multiplier_STAGE1__0991_ ;
 wire u_multiplier_STAGE1__0992_ ;
 wire u_multiplier_STAGE1__0993_ ;
 wire u_multiplier_STAGE1__0994_ ;
 wire u_multiplier_STAGE1__0995_ ;
 wire u_multiplier_STAGE1__0996_ ;
 wire u_multiplier_STAGE1__0997_ ;
 wire u_multiplier_STAGE1__0998_ ;
 wire u_multiplier_STAGE1__0999_ ;
 wire u_multiplier_STAGE1__1000_ ;
 wire u_multiplier_STAGE1__1001_ ;
 wire u_multiplier_STAGE1__1002_ ;
 wire u_multiplier_STAGE1__1003_ ;
 wire u_multiplier_STAGE1__1004_ ;
 wire u_multiplier_STAGE1__1005_ ;
 wire u_multiplier_STAGE1__1006_ ;
 wire u_multiplier_STAGE1__1007_ ;
 wire u_multiplier_STAGE1__1008_ ;
 wire u_multiplier_STAGE1__1009_ ;
 wire u_multiplier_STAGE1__1010_ ;
 wire u_multiplier_STAGE1__1011_ ;
 wire u_multiplier_STAGE1__1012_ ;
 wire u_multiplier_STAGE1__1013_ ;
 wire u_multiplier_STAGE1__1014_ ;
 wire u_multiplier_STAGE1__1015_ ;
 wire u_multiplier_STAGE1__1016_ ;
 wire u_multiplier_STAGE1__1017_ ;
 wire u_multiplier_STAGE1__1018_ ;
 wire u_multiplier_STAGE1__1019_ ;
 wire u_multiplier_STAGE1__1020_ ;
 wire u_multiplier_STAGE1__1021_ ;
 wire u_multiplier_STAGE1__1022_ ;
 wire u_multiplier_STAGE1__1023_ ;
 wire u_multiplier_STAGE1__1024_ ;
 wire u_multiplier_STAGE1__1025_ ;
 wire u_multiplier_STAGE1__1026_ ;
 wire u_multiplier_STAGE1__1027_ ;
 wire u_multiplier_STAGE1__1028_ ;
 wire u_multiplier_STAGE1__1029_ ;
 wire u_multiplier_STAGE1__1030_ ;
 wire u_multiplier_STAGE1__1031_ ;
 wire u_multiplier_STAGE1__1032_ ;
 wire u_multiplier_STAGE1__1033_ ;
 wire u_multiplier_STAGE1__1034_ ;
 wire u_multiplier_STAGE1__1035_ ;
 wire u_multiplier_STAGE1__1036_ ;
 wire u_multiplier_STAGE1__1037_ ;
 wire u_multiplier_STAGE1__1038_ ;
 wire u_multiplier_STAGE1__1039_ ;
 wire u_multiplier_STAGE1__1040_ ;
 wire u_multiplier_STAGE1__1041_ ;
 wire u_multiplier_STAGE1__1042_ ;
 wire u_multiplier_STAGE1__1043_ ;
 wire u_multiplier_STAGE1__1044_ ;
 wire u_multiplier_STAGE1__1045_ ;
 wire u_multiplier_STAGE1__1046_ ;
 wire u_multiplier_STAGE1__1047_ ;
 wire u_multiplier_STAGE1__1048_ ;
 wire u_multiplier_STAGE1__1049_ ;
 wire u_multiplier_STAGE1__1050_ ;
 wire u_multiplier_STAGE1__1051_ ;
 wire u_multiplier_STAGE1__1052_ ;
 wire u_multiplier_STAGE1__1053_ ;
 wire u_multiplier_STAGE1__1054_ ;
 wire u_multiplier_STAGE1__1055_ ;
 wire u_multiplier_STAGE1__1056_ ;
 wire u_multiplier_STAGE1__1057_ ;
 wire u_multiplier_STAGE1__1058_ ;
 wire u_multiplier_STAGE1__1059_ ;
 wire u_multiplier_STAGE1__1060_ ;
 wire u_multiplier_STAGE1__1061_ ;
 wire u_multiplier_STAGE1__1062_ ;
 wire u_multiplier_STAGE1__1063_ ;
 wire u_multiplier_STAGE1__1064_ ;
 wire u_multiplier_STAGE1__1065_ ;
 wire u_multiplier_STAGE1__1066_ ;
 wire u_multiplier_STAGE1__1067_ ;
 wire u_multiplier_STAGE1__1068_ ;
 wire u_multiplier_STAGE1__1069_ ;
 wire u_multiplier_STAGE1__1070_ ;
 wire u_multiplier_STAGE1__1071_ ;
 wire u_multiplier_STAGE1__1072_ ;
 wire u_multiplier_STAGE1__1073_ ;
 wire u_multiplier_STAGE1__1074_ ;
 wire u_multiplier_STAGE1__1075_ ;
 wire u_multiplier_STAGE1__1076_ ;
 wire u_multiplier_STAGE1__1077_ ;
 wire u_multiplier_STAGE1__1078_ ;
 wire u_multiplier_STAGE1__1079_ ;
 wire u_multiplier_STAGE1__1080_ ;
 wire u_multiplier_STAGE1__1081_ ;
 wire u_multiplier_STAGE1__1082_ ;
 wire u_multiplier_STAGE1__1083_ ;
 wire u_multiplier_STAGE1__1084_ ;
 wire u_multiplier_STAGE1__1085_ ;
 wire u_multiplier_STAGE1__1086_ ;
 wire u_multiplier_STAGE1__1087_ ;
 wire u_multiplier_STAGE1__1088_ ;
 wire u_multiplier_STAGE1__1089_ ;
 wire u_multiplier_STAGE1__1090_ ;
 wire u_multiplier_STAGE1__1091_ ;
 wire u_multiplier_STAGE1__1092_ ;
 wire u_multiplier_STAGE1__1093_ ;
 wire u_multiplier_STAGE1__1094_ ;
 wire u_multiplier_STAGE1__1095_ ;
 wire u_multiplier_STAGE1__1096_ ;
 wire u_multiplier_STAGE1__1097_ ;
 wire u_multiplier_STAGE1__1098_ ;
 wire u_multiplier_STAGE1__1099_ ;
 wire u_multiplier_STAGE1__1100_ ;
 wire u_multiplier_STAGE1__1101_ ;
 wire u_multiplier_STAGE1__1102_ ;
 wire u_multiplier_STAGE1__1103_ ;
 wire u_multiplier_STAGE1__1104_ ;
 wire u_multiplier_STAGE1__1105_ ;
 wire u_multiplier_STAGE1__1106_ ;
 wire u_multiplier_STAGE1__1107_ ;
 wire u_multiplier_STAGE1__1108_ ;
 wire u_multiplier_STAGE1__1109_ ;
 wire u_multiplier_STAGE1__1110_ ;
 wire u_multiplier_STAGE1__1111_ ;
 wire u_multiplier_STAGE1__1112_ ;
 wire u_multiplier_STAGE1__1113_ ;
 wire u_multiplier_STAGE1__1114_ ;
 wire u_multiplier_STAGE1__1115_ ;
 wire u_multiplier_STAGE1__1116_ ;
 wire u_multiplier_STAGE1__1117_ ;
 wire u_multiplier_STAGE1__1118_ ;
 wire u_multiplier_STAGE1__1119_ ;
 wire u_multiplier_STAGE1__1120_ ;
 wire u_multiplier_STAGE1__1121_ ;
 wire u_multiplier_STAGE1__1122_ ;
 wire u_multiplier_STAGE1__1123_ ;
 wire u_multiplier_STAGE1__1124_ ;
 wire u_multiplier_STAGE1__1125_ ;
 wire u_multiplier_STAGE1__1126_ ;
 wire u_multiplier_STAGE1__1127_ ;
 wire u_multiplier_STAGE1__1128_ ;
 wire u_multiplier_STAGE1__1129_ ;
 wire u_multiplier_STAGE1__1130_ ;
 wire u_multiplier_STAGE1__1131_ ;
 wire u_multiplier_STAGE1__1132_ ;
 wire u_multiplier_STAGE1__1133_ ;
 wire u_multiplier_STAGE1__1134_ ;
 wire u_multiplier_STAGE1__1135_ ;
 wire u_multiplier_STAGE1__1136_ ;
 wire u_multiplier_STAGE1__1137_ ;
 wire u_multiplier_STAGE1__1138_ ;
 wire u_multiplier_STAGE1__1139_ ;
 wire u_multiplier_STAGE1__1140_ ;
 wire u_multiplier_STAGE1__1141_ ;
 wire u_multiplier_STAGE1__1142_ ;
 wire u_multiplier_STAGE1__1143_ ;
 wire u_multiplier_STAGE1__1144_ ;
 wire u_multiplier_STAGE1__1145_ ;
 wire u_multiplier_STAGE1__1146_ ;
 wire u_multiplier_STAGE1__1147_ ;
 wire u_multiplier_STAGE1__1148_ ;
 wire u_multiplier_STAGE1__1149_ ;
 wire net125;
 wire u_multiplier_STAGE1_pp1_32_1_cout ;
 wire u_multiplier_STAGE1_pp1_32_2_cout ;
 wire u_multiplier_STAGE1_pp1_32_3_cout ;
 wire u_multiplier_STAGE1_pp1_32_4_cout ;
 wire u_multiplier_STAGE1_pp1_32_5_cout ;
 wire u_multiplier_STAGE1_pp1_32_6_cout ;
 wire u_multiplier_STAGE1_pp1_32_7_cout ;
 wire u_multiplier_STAGE1_pp1_33_1_cout ;
 wire u_multiplier_STAGE1_pp1_33_2_cout ;
 wire u_multiplier_STAGE1_pp1_33_3_cout ;
 wire u_multiplier_STAGE1_pp1_33_4_cout ;
 wire u_multiplier_STAGE1_pp1_33_5_cout ;
 wire u_multiplier_STAGE1_pp1_33_6_cout ;
 wire u_multiplier_STAGE1_pp1_33_7_cout ;
 wire u_multiplier_STAGE1_pp1_34_1_cout ;
 wire u_multiplier_STAGE1_pp1_34_2_cout ;
 wire u_multiplier_STAGE1_pp1_34_3_cout ;
 wire u_multiplier_STAGE1_pp1_34_4_cout ;
 wire u_multiplier_STAGE1_pp1_34_5_cout ;
 wire u_multiplier_STAGE1_pp1_34_6_cout ;
 wire u_multiplier_STAGE1_pp1_34_7_cout ;
 wire u_multiplier_STAGE1_pp1_35_1_cout ;
 wire u_multiplier_STAGE1_pp1_35_2_cout ;
 wire u_multiplier_STAGE1_pp1_35_3_cout ;
 wire u_multiplier_STAGE1_pp1_35_4_cout ;
 wire u_multiplier_STAGE1_pp1_35_5_cout ;
 wire u_multiplier_STAGE1_pp1_35_6_cout ;
 wire u_multiplier_STAGE1_pp1_36_1_cout ;
 wire u_multiplier_STAGE1_pp1_36_2_cout ;
 wire u_multiplier_STAGE1_pp1_36_3_cout ;
 wire u_multiplier_STAGE1_pp1_36_4_cout ;
 wire u_multiplier_STAGE1_pp1_36_5_cout ;
 wire u_multiplier_STAGE1_pp1_36_6_cout ;
 wire u_multiplier_STAGE1_pp1_37_1_cout ;
 wire u_multiplier_STAGE1_pp1_37_2_cout ;
 wire u_multiplier_STAGE1_pp1_37_3_cout ;
 wire u_multiplier_STAGE1_pp1_37_4_cout ;
 wire u_multiplier_STAGE1_pp1_37_5_cout ;
 wire u_multiplier_STAGE1_pp1_38_1_cout ;
 wire u_multiplier_STAGE1_pp1_38_2_cout ;
 wire u_multiplier_STAGE1_pp1_38_3_cout ;
 wire u_multiplier_STAGE1_pp1_38_4_cout ;
 wire u_multiplier_STAGE1_pp1_38_5_cout ;
 wire u_multiplier_STAGE1_pp1_39_1_cout ;
 wire u_multiplier_STAGE1_pp1_39_2_cout ;
 wire u_multiplier_STAGE1_pp1_39_3_cout ;
 wire u_multiplier_STAGE1_pp1_39_4_cout ;
 wire u_multiplier_STAGE1_pp1_40_1_cout ;
 wire u_multiplier_STAGE1_pp1_40_2_cout ;
 wire u_multiplier_STAGE1_pp1_40_3_cout ;
 wire u_multiplier_STAGE1_pp1_40_4_cout ;
 wire u_multiplier_STAGE1_pp1_41_1_cout ;
 wire u_multiplier_STAGE1_pp1_41_2_cout ;
 wire u_multiplier_STAGE1_pp1_41_3_cout ;
 wire u_multiplier_STAGE1_pp1_42_1_cout ;
 wire u_multiplier_STAGE1_pp1_42_2_cout ;
 wire u_multiplier_STAGE1_pp1_42_3_cout ;
 wire u_multiplier_STAGE1_pp1_43_1_cout ;
 wire u_multiplier_STAGE1_pp1_43_2_cout ;
 wire u_multiplier_STAGE1_pp1_44_1_cout ;
 wire u_multiplier_STAGE1_pp1_44_2_cout ;
 wire u_multiplier_STAGE1_pp1_45_1_cout ;
 wire u_multiplier_STAGE1_pp1_46_1_cout ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_4__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_4__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_4__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_4__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_4__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_4__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_4__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_5__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_5__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_5__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_5__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_5__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_5__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_5__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_6__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_6__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_6__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_6__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_6__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_6__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_6__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_7__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_7__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_7__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_7__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_7__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_7__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_32_7__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_4__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_4__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_4__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_4__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_4__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_4__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_4__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_5__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_5__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_5__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_5__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_5__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_5__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_5__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_6__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_6__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_6__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_6__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_6__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_6__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_6__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_7__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_7__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_7__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_7__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_7__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_7__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_33_7__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_4__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_4__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_4__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_4__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_4__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_4__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_4__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_5__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_5__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_5__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_5__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_5__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_5__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_5__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_6__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_6__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_6__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_6__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_6__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_6__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_6__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_7__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_7__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_7__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_7__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_7__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_7__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_34_7__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_4__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_4__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_4__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_4__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_4__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_4__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_4__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_5__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_5__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_5__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_5__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_5__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_5__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_5__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_6__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_6__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_6__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_6__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_6__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_6__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_35_6__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_4__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_4__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_4__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_4__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_4__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_4__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_4__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_5__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_5__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_5__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_5__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_5__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_5__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_5__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_6__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_6__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_6__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_6__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_6__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_6__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_36_6__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_4__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_4__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_4__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_4__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_4__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_4__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_4__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_5__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_5__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_5__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_5__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_5__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_5__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_37_5__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_4__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_4__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_4__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_4__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_4__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_4__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_4__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_5__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_5__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_5__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_5__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_5__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_5__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_38_5__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_4__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_4__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_4__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_4__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_4__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_4__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_39_4__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_4__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_4__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_4__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_4__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_4__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_4__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_40_4__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_41_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_3__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_3__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_3__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_3__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_3__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_3__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_42_3__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_43_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_2__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_2__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_2__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_2__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_2__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_2__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_44_2__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_45_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_45_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_45_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_45_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_45_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_45_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_45_1__17_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_46_1__11_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_46_1__12_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_46_1__13_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_46_1__14_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_46_1__15_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_46_1__16_ ;
 wire u_multiplier_STAGE1_E_4_2_pp_46_1__17_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_32_1__08_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_32_1__09_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_32_1__10_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_32_1__11_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_35_1__08_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_35_1__09_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_35_1__10_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_35_1__11_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_37_1__08_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_37_1__09_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_37_1__10_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_37_1__11_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_39_1__08_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_39_1__09_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_39_1__10_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_39_1__11_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_41_1__08_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_41_1__09_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_41_1__10_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_41_1__11_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_43_1__08_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_43_1__09_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_43_1__10_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_43_1__11_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_45_1__08_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_45_1__09_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_45_1__10_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_45_1__11_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_47_1__08_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_47_1__09_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_47_1__10_ ;
 wire u_multiplier_STAGE1_Full_adder_pp_47_1__11_ ;
 wire u_multiplier_STAGE1_acci1_pp_17_0__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_17_0__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_17_0__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_17_0__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_17_0__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_17_0__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_18_0__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_18_0__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_18_0__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_18_0__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_18_0__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_18_0__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_19_0__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_19_0__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_19_0__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_19_0__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_19_0__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_19_0__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_19_1__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_19_1__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_19_1__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_19_1__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_19_1__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_19_1__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_20_0__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_20_0__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_20_0__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_20_0__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_20_0__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_20_0__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_20_1__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_20_1__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_20_1__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_20_1__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_20_1__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_20_1__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_21_0__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_21_0__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_21_0__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_21_0__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_21_0__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_21_0__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_21_1__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_21_1__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_21_1__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_21_1__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_21_1__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_21_1__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_21_2__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_21_2__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_21_2__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_21_2__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_21_2__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_21_2__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_22_0__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_22_0__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_22_0__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_22_0__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_22_0__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_22_0__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_22_1__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_22_1__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_22_1__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_22_1__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_22_1__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_22_1__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_22_2__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_22_2__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_22_2__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_22_2__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_22_2__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_22_2__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_23_0__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_23_0__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_23_0__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_23_0__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_23_0__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_23_0__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_23_1__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_23_1__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_23_1__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_23_1__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_23_1__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_23_1__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_23_2__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_23_2__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_23_2__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_23_2__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_23_2__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_23_2__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_23_3__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_23_3__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_23_3__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_23_3__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_23_3__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_23_3__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_24_0__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_24_0__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_24_0__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_24_0__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_24_0__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_24_0__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_24_1__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_24_1__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_24_1__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_24_1__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_24_1__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_24_1__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_24_2__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_24_2__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_24_2__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_24_2__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_24_2__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_24_2__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_24_3__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_24_3__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_24_3__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_24_3__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_24_3__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_24_3__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_0__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_0__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_0__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_0__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_0__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_0__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_1__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_1__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_1__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_1__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_1__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_1__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_2__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_2__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_2__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_2__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_2__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_2__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_3__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_3__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_3__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_3__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_3__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_3__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_4__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_4__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_4__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_4__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_4__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_25_4__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_0__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_0__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_0__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_0__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_0__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_0__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_1__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_1__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_1__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_1__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_1__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_1__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_2__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_2__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_2__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_2__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_2__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_2__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_3__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_3__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_3__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_3__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_3__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_3__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_4__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_4__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_4__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_4__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_4__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_26_4__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_0__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_0__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_0__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_0__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_0__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_0__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_1__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_1__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_1__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_1__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_1__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_1__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_2__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_2__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_2__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_2__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_2__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_2__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_3__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_3__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_3__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_3__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_3__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_3__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_4__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_4__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_4__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_4__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_4__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_4__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_5__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_5__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_5__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_5__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_5__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_27_5__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_0__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_0__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_0__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_0__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_0__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_0__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_1__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_1__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_1__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_1__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_1__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_1__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_2__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_2__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_2__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_2__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_2__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_2__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_3__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_3__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_3__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_3__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_3__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_3__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_4__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_4__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_4__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_4__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_4__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_4__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_5__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_5__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_5__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_5__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_5__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_28_5__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_0__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_0__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_0__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_0__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_0__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_0__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_1__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_1__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_1__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_1__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_1__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_1__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_2__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_2__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_2__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_2__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_2__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_2__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_3__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_3__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_3__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_3__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_3__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_3__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_4__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_4__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_4__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_4__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_4__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_4__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_5__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_5__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_5__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_5__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_5__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_5__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_6__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_6__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_6__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_6__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_6__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_29_6__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_0__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_0__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_0__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_0__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_0__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_0__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_1__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_1__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_1__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_1__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_1__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_1__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_2__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_2__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_2__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_2__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_2__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_2__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_3__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_3__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_3__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_3__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_3__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_3__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_4__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_4__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_4__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_4__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_4__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_4__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_5__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_5__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_5__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_5__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_5__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_5__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_6__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_6__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_6__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_6__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_6__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_30_6__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_0__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_0__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_0__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_0__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_0__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_0__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_1__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_1__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_1__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_1__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_1__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_1__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_2__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_2__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_2__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_2__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_2__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_2__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_3__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_3__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_3__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_3__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_3__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_3__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_4__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_4__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_4__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_4__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_4__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_4__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_5__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_5__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_5__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_5__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_5__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_5__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_6__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_6__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_6__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_6__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_6__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_6__20_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_7__15_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_7__16_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_7__17_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_7__18_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_7__19_ ;
 wire u_multiplier_STAGE1_acci1_pp_31_7__20_ ;
 wire net133;
 wire u_multiplier_STAGE2_pp2_32_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_32_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_32_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_32_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_33_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_33_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_33_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_33_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_34_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_34_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_34_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_34_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_35_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_35_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_35_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_35_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_36_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_36_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_36_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_36_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_37_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_37_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_37_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_37_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_38_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_38_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_38_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_38_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_39_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_39_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_39_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_39_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_40_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_40_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_40_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_40_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_41_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_41_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_41_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_41_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_42_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_42_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_42_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_42_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_43_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_43_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_43_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_43_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_44_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_44_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_44_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_44_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_45_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_45_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_45_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_45_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_46_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_46_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_46_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_46_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_47_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_47_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_47_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_47_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_48_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_48_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_48_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_48_e42_4_cout ;
 wire u_multiplier_STAGE2_pp2_49_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_49_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_49_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_50_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_50_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_50_e42_3_cout ;
 wire u_multiplier_STAGE2_pp2_51_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_51_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_52_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_52_e42_2_cout ;
 wire u_multiplier_STAGE2_pp2_53_e42_1_cout ;
 wire u_multiplier_STAGE2_pp2_54_e42_1_cout ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_32_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_33_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_34_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_35_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_36_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_37_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_38_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_39_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_40_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_41_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_42_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_43_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_44_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_45_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_46_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_47_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_4__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_4__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_4__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_4__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_4__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_4__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_48_4__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_49_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_3__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_3__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_3__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_3__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_3__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_3__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_50_3__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_51_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_2__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_2__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_2__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_2__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_2__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_2__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_52_2__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_53_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_53_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_53_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_53_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_53_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_53_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_53_1__17_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_54_1__11_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_54_1__12_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_54_1__13_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_54_1__14_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_54_1__15_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_54_1__16_ ;
 wire u_multiplier_STAGE2_E_4_2_pp2_54_1__17_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_49_1__08_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_49_1__09_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_49_1__10_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_49_1__11_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_51_1__08_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_51_1__09_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_51_1__10_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_51_1__11_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_53_1__08_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_53_1__09_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_53_1__10_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_53_1__11_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_55_1__08_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_55_1__09_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_55_1__10_ ;
 wire u_multiplier_STAGE2_Full_adder_pp2_55_1__11_ ;
 wire u_multiplier_STAGE2_acci_pp2_10_0__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_10_0__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_10_0__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_10_0__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_10_0__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_10_0__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_11_0__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_11_0__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_11_0__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_11_0__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_11_0__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_11_0__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_11_1__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_11_1__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_11_1__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_11_1__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_11_1__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_11_1__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_12_0__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_12_0__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_12_0__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_12_0__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_12_0__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_12_0__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_12_1__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_12_1__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_12_1__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_12_1__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_12_1__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_12_1__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_13_0__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_13_0__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_13_0__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_13_0__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_13_0__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_13_0__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_13_1__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_13_1__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_13_1__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_13_1__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_13_1__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_13_1__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_13_2__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_13_2__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_13_2__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_13_2__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_13_2__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_13_2__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_14_0__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_14_0__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_14_0__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_14_0__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_14_0__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_14_0__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_14_1__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_14_1__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_14_1__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_14_1__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_14_1__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_14_1__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_14_2__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_14_2__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_14_2__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_14_2__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_14_2__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_14_2__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_15_0__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_15_0__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_15_0__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_15_0__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_15_0__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_15_0__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_15_1__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_15_1__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_15_1__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_15_1__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_15_1__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_15_1__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_15_2__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_15_2__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_15_2__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_15_2__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_15_2__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_15_2__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_15_3__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_15_3__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_15_3__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_15_3__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_15_3__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_15_3__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_16_0__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_16_0__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_16_0__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_16_0__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_16_0__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_16_0__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_16_1__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_16_1__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_16_1__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_16_1__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_16_1__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_16_1__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_16_2__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_16_2__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_16_2__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_16_2__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_16_2__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_16_2__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_16_3__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_16_3__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_16_3__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_16_3__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_16_3__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_16_3__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_17_0__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_17_0__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_17_0__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_17_0__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_17_0__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_17_0__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_17_1__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_17_1__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_17_1__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_17_1__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_17_1__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_17_1__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_17_2__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_17_2__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_17_2__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_17_2__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_17_2__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_17_2__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_17_3__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_17_3__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_17_3__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_17_3__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_17_3__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_17_3__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_18_0__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_18_0__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_18_0__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_18_0__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_18_0__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_18_0__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_18_1__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_18_1__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_18_1__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_18_1__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_18_1__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_18_1__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_18_2__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_18_2__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_18_2__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_18_2__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_18_2__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_18_2__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_18_3__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_18_3__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_18_3__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_18_3__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_18_3__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_18_3__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_19_0__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_19_0__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_19_0__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_19_0__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_19_0__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_19_0__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_19_1__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_19_1__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_19_1__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_19_1__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_19_1__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_19_1__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_19_2__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_19_2__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_19_2__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_19_2__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_19_2__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_19_2__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_19_3__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_19_3__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_19_3__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_19_3__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_19_3__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_19_3__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_20_0__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_20_0__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_20_0__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_20_0__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_20_0__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_20_0__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_20_1__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_20_1__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_20_1__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_20_1__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_20_1__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_20_1__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_20_2__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_20_2__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_20_2__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_20_2__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_20_2__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_20_2__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_20_3__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_20_3__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_20_3__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_20_3__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_20_3__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_20_3__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_21_0__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_21_0__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_21_0__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_21_0__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_21_0__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_21_0__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_21_1__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_21_1__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_21_1__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_21_1__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_21_1__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_21_1__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_21_2__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_21_2__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_21_2__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_21_2__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_21_2__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_21_2__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_21_3__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_21_3__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_21_3__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_21_3__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_21_3__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_21_3__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_22_0__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_22_0__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_22_0__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_22_0__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_22_0__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_22_0__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_22_1__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_22_1__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_22_1__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_22_1__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_22_1__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_22_1__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_22_2__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_22_2__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_22_2__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_22_2__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_22_2__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_22_2__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_22_3__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_22_3__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_22_3__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_22_3__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_22_3__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_22_3__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_23_0__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_23_0__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_23_0__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_23_0__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_23_0__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_23_0__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_23_1__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_23_1__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_23_1__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_23_1__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_23_1__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_23_1__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_23_2__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_23_2__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_23_2__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_23_2__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_23_2__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_23_2__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_23_3__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_23_3__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_23_3__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_23_3__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_23_3__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_23_3__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_24_0__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_24_0__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_24_0__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_24_0__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_24_0__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_24_0__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_24_1__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_24_1__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_24_1__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_24_1__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_24_1__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_24_1__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_24_2__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_24_2__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_24_2__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_24_2__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_24_2__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_24_2__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_24_3__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_24_3__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_24_3__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_24_3__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_24_3__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_24_3__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_25_0__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_25_0__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_25_0__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_25_0__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_25_0__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_25_0__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_25_1__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_25_1__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_25_1__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_25_1__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_25_1__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_25_1__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_25_2__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_25_2__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_25_2__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_25_2__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_25_2__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_25_2__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_25_3__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_25_3__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_25_3__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_25_3__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_25_3__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_25_3__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_26_0__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_26_0__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_26_0__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_26_0__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_26_0__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_26_0__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_26_1__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_26_1__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_26_1__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_26_1__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_26_1__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_26_1__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_26_2__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_26_2__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_26_2__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_26_2__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_26_2__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_26_2__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_26_3__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_26_3__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_26_3__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_26_3__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_26_3__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_26_3__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_27_0__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_27_0__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_27_0__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_27_0__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_27_0__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_27_0__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_27_1__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_27_1__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_27_1__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_27_1__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_27_1__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_27_1__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_27_2__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_27_2__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_27_2__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_27_2__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_27_2__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_27_2__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_27_3__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_27_3__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_27_3__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_27_3__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_27_3__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_27_3__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_28_0__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_28_0__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_28_0__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_28_0__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_28_0__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_28_0__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_28_1__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_28_1__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_28_1__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_28_1__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_28_1__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_28_1__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_28_2__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_28_2__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_28_2__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_28_2__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_28_2__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_28_2__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_28_3__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_28_3__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_28_3__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_28_3__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_28_3__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_28_3__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_29_0__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_29_0__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_29_0__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_29_0__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_29_0__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_29_0__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_29_1__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_29_1__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_29_1__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_29_1__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_29_1__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_29_1__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_29_2__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_29_2__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_29_2__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_29_2__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_29_2__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_29_2__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_29_3__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_29_3__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_29_3__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_29_3__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_29_3__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_29_3__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_30_0__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_30_0__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_30_0__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_30_0__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_30_0__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_30_0__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_30_1__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_30_1__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_30_1__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_30_1__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_30_1__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_30_1__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_30_2__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_30_2__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_30_2__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_30_2__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_30_2__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_30_2__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_30_3__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_30_3__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_30_3__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_30_3__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_30_3__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_30_3__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_31_0__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_31_0__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_31_0__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_31_0__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_31_0__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_31_0__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_31_1__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_31_1__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_31_1__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_31_1__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_31_1__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_31_1__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_31_2__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_31_2__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_31_2__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_31_2__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_31_2__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_31_2__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_31_3__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_31_3__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_31_3__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_31_3__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_31_3__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_31_3__20_ ;
 wire u_multiplier_STAGE2_acci_pp2_9_0__15_ ;
 wire u_multiplier_STAGE2_acci_pp2_9_0__16_ ;
 wire u_multiplier_STAGE2_acci_pp2_9_0__17_ ;
 wire u_multiplier_STAGE2_acci_pp2_9_0__18_ ;
 wire u_multiplier_STAGE2_acci_pp2_9_0__19_ ;
 wire u_multiplier_STAGE2_acci_pp2_9_0__20_ ;
 wire net137;
 wire u_multiplier_STAGE3_pp3_32_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_32_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_33_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_33_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_34_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_34_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_35_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_35_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_36_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_36_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_37_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_37_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_38_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_38_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_39_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_39_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_40_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_40_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_41_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_41_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_42_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_42_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_43_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_43_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_44_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_44_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_45_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_45_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_46_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_46_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_47_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_47_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_48_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_48_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_49_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_49_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_50_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_50_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_51_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_51_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_52_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_52_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_53_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_53_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_54_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_54_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_55_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_55_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_56_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_56_e42_2_cout ;
 wire u_multiplier_STAGE3_pp3_57_e42_1_cout ;
 wire u_multiplier_STAGE3_pp3_58_e42_1_cout ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_32_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_33_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_34_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_35_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_36_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_37_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_38_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_39_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_40_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_41_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_42_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_43_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_44_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_45_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_46_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_47_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_48_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_49_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_50_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_51_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_52_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_53_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_54_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_55_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_2__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_2__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_2__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_2__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_2__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_2__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_56_2__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_57_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_57_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_57_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_57_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_57_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_57_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_57_1__17_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_58_1__11_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_58_1__12_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_58_1__13_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_58_1__14_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_58_1__15_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_58_1__16_ ;
 wire u_multiplier_STAGE3_E_4_2_pp3_58_1__17_ ;
 wire u_multiplier_STAGE3_Full_adder_pp3_57_1__08_ ;
 wire u_multiplier_STAGE3_Full_adder_pp3_57_1__09_ ;
 wire u_multiplier_STAGE3_Full_adder_pp3_57_1__10_ ;
 wire u_multiplier_STAGE3_Full_adder_pp3_57_1__11_ ;
 wire u_multiplier_STAGE3_Full_adder_pp3_59_1__08_ ;
 wire u_multiplier_STAGE3_Full_adder_pp3_59_1__09_ ;
 wire u_multiplier_STAGE3_Full_adder_pp3_59_1__10_ ;
 wire u_multiplier_STAGE3_Full_adder_pp3_59_1__11_ ;
 wire u_multiplier_STAGE3_acci_pp3_10_0__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_10_0__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_10_0__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_10_0__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_10_0__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_10_0__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_10_1__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_10_1__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_10_1__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_10_1__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_10_1__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_10_1__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_11_0__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_11_0__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_11_0__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_11_0__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_11_0__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_11_0__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_11_1__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_11_1__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_11_1__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_11_1__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_11_1__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_11_1__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_12_0__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_12_0__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_12_0__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_12_0__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_12_0__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_12_0__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_12_1__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_12_1__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_12_1__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_12_1__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_12_1__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_12_1__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_13_0__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_13_0__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_13_0__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_13_0__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_13_0__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_13_0__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_13_1__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_13_1__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_13_1__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_13_1__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_13_1__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_13_1__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_14_0__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_14_0__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_14_0__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_14_0__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_14_0__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_14_0__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_14_1__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_14_1__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_14_1__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_14_1__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_14_1__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_14_1__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_15_0__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_15_0__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_15_0__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_15_0__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_15_0__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_15_0__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_15_1__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_15_1__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_15_1__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_15_1__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_15_1__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_15_1__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_16_0__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_16_0__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_16_0__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_16_0__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_16_0__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_16_0__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_16_1__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_16_1__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_16_1__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_16_1__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_16_1__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_16_1__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_17_0__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_17_0__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_17_0__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_17_0__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_17_0__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_17_0__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_17_1__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_17_1__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_17_1__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_17_1__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_17_1__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_17_1__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_18_0__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_18_0__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_18_0__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_18_0__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_18_0__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_18_0__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_18_1__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_18_1__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_18_1__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_18_1__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_18_1__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_18_1__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_19_0__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_19_0__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_19_0__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_19_0__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_19_0__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_19_0__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_19_1__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_19_1__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_19_1__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_19_1__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_19_1__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_19_1__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_20_0__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_20_0__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_20_0__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_20_0__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_20_0__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_20_0__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_20_1__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_20_1__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_20_1__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_20_1__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_20_1__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_20_1__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_21_0__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_21_0__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_21_0__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_21_0__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_21_0__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_21_0__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_21_1__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_21_1__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_21_1__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_21_1__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_21_1__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_21_1__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_22_0__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_22_0__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_22_0__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_22_0__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_22_0__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_22_0__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_22_1__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_22_1__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_22_1__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_22_1__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_22_1__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_22_1__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_23_0__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_23_0__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_23_0__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_23_0__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_23_0__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_23_0__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_23_1__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_23_1__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_23_1__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_23_1__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_23_1__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_23_1__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_24_0__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_24_0__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_24_0__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_24_0__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_24_0__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_24_0__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_24_1__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_24_1__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_24_1__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_24_1__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_24_1__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_24_1__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_25_0__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_25_0__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_25_0__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_25_0__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_25_0__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_25_0__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_25_1__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_25_1__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_25_1__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_25_1__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_25_1__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_25_1__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_26_0__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_26_0__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_26_0__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_26_0__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_26_0__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_26_0__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_26_1__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_26_1__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_26_1__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_26_1__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_26_1__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_26_1__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_27_0__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_27_0__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_27_0__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_27_0__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_27_0__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_27_0__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_27_1__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_27_1__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_27_1__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_27_1__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_27_1__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_27_1__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_28_0__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_28_0__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_28_0__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_28_0__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_28_0__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_28_0__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_28_1__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_28_1__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_28_1__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_28_1__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_28_1__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_28_1__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_29_0__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_29_0__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_29_0__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_29_0__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_29_0__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_29_0__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_29_1__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_29_1__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_29_1__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_29_1__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_29_1__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_29_1__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_30_0__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_30_0__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_30_0__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_30_0__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_30_0__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_30_0__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_30_1__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_30_1__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_30_1__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_30_1__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_30_1__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_30_1__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_31_0__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_31_0__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_31_0__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_31_0__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_31_0__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_31_0__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_31_1__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_31_1__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_31_1__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_31_1__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_31_1__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_31_1__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_5_0__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_5_0__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_5_0__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_5_0__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_5_0__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_5_0__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_6_0__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_6_0__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_6_0__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_6_0__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_6_0__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_6_0__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_7_0__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_7_0__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_7_0__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_7_0__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_7_0__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_7_0__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_7_1__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_7_1__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_7_1__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_7_1__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_7_1__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_7_1__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_8_0__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_8_0__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_8_0__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_8_0__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_8_0__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_8_0__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_8_1__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_8_1__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_8_1__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_8_1__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_8_1__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_8_1__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_9_0__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_9_0__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_9_0__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_9_0__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_9_0__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_9_0__20_ ;
 wire u_multiplier_STAGE3_acci_pp3_9_1__15_ ;
 wire u_multiplier_STAGE3_acci_pp3_9_1__16_ ;
 wire u_multiplier_STAGE3_acci_pp3_9_1__17_ ;
 wire u_multiplier_STAGE3_acci_pp3_9_1__18_ ;
 wire u_multiplier_STAGE3_acci_pp3_9_1__19_ ;
 wire u_multiplier_STAGE3_acci_pp3_9_1__20_ ;
 wire u_multiplier_STAGE4_pp4_32_c2 ;
 wire u_multiplier_STAGE4_pp4_33_c2 ;
 wire u_multiplier_STAGE4_pp4_34_c2 ;
 wire u_multiplier_STAGE4_pp4_35_c2 ;
 wire u_multiplier_STAGE4_pp4_36_c2 ;
 wire u_multiplier_STAGE4_pp4_37_c2 ;
 wire u_multiplier_STAGE4_pp4_38_c2 ;
 wire u_multiplier_STAGE4_pp4_39_c2 ;
 wire u_multiplier_STAGE4_pp4_40_c2 ;
 wire u_multiplier_STAGE4_pp4_41_c2 ;
 wire u_multiplier_STAGE4_pp4_42_c2 ;
 wire u_multiplier_STAGE4_pp4_43_c2 ;
 wire u_multiplier_STAGE4_pp4_44_c2 ;
 wire u_multiplier_STAGE4_pp4_45_c2 ;
 wire u_multiplier_STAGE4_pp4_46_c2 ;
 wire u_multiplier_STAGE4_pp4_47_c2 ;
 wire u_multiplier_STAGE4_pp4_48_c2 ;
 wire u_multiplier_STAGE4_pp4_49_c2 ;
 wire u_multiplier_STAGE4_pp4_50_c2 ;
 wire u_multiplier_STAGE4_pp4_51_c2 ;
 wire u_multiplier_STAGE4_pp4_52_c2 ;
 wire u_multiplier_STAGE4_pp4_53_c2 ;
 wire u_multiplier_STAGE4_pp4_54_c2 ;
 wire u_multiplier_STAGE4_pp4_55_c2 ;
 wire u_multiplier_STAGE4_pp4_56_c2 ;
 wire u_multiplier_STAGE4_pp4_57_c2 ;
 wire u_multiplier_STAGE4_pp4_58_c2 ;
 wire u_multiplier_STAGE4_pp4_59_c2 ;
 wire u_multiplier_STAGE4_pp4_60_c2 ;
 wire u_multiplier_STAGE4_ACCI_pp4_10__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_10__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_10__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_10__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_10__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_10__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_11__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_11__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_11__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_11__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_11__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_11__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_12__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_12__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_12__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_12__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_12__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_12__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_13__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_13__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_13__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_13__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_13__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_13__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_14__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_14__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_14__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_14__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_14__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_14__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_15__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_15__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_15__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_15__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_15__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_15__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_16__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_16__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_16__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_16__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_16__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_16__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_17__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_17__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_17__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_17__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_17__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_17__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_18__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_18__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_18__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_18__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_18__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_18__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_19__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_19__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_19__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_19__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_19__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_19__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_20__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_20__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_20__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_20__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_20__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_20__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_21__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_21__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_21__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_21__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_21__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_21__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_22__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_22__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_22__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_22__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_22__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_22__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_23__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_23__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_23__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_23__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_23__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_23__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_24__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_24__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_24__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_24__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_24__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_24__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_25__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_25__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_25__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_25__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_25__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_25__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_26__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_26__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_26__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_26__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_26__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_26__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_27__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_27__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_27__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_27__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_27__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_27__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_28__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_28__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_28__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_28__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_28__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_28__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_29__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_29__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_29__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_29__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_29__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_29__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_3__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_3__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_3__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_3__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_3__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_3__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_30__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_30__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_30__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_30__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_30__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_30__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_31__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_31__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_31__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_31__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_31__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_31__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_4__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_4__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_4__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_4__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_4__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_4__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_5__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_5__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_5__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_5__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_5__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_5__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_6__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_6__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_6__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_6__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_6__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_6__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_7__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_7__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_7__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_7__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_7__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_7__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_8__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_8__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_8__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_8__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_8__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_8__20_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_9__15_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_9__16_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_9__17_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_9__18_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_9__19_ ;
 wire u_multiplier_STAGE4_ACCI_pp4_9__20_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_32__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_32__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_32__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_32__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_32__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_32__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_32__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_33__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_33__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_33__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_33__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_33__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_33__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_33__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_34__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_34__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_34__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_34__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_34__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_34__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_34__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_35__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_35__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_35__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_35__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_35__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_35__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_35__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_36__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_36__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_36__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_36__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_36__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_36__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_36__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_37__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_37__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_37__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_37__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_37__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_37__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_37__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_38__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_38__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_38__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_38__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_38__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_38__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_38__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_39__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_39__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_39__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_39__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_39__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_39__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_39__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_40__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_40__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_40__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_40__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_40__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_40__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_40__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_41__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_41__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_41__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_41__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_41__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_41__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_41__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_42__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_42__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_42__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_42__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_42__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_42__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_42__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_43__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_43__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_43__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_43__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_43__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_43__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_43__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_44__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_44__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_44__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_44__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_44__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_44__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_44__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_45__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_45__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_45__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_45__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_45__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_45__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_45__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_46__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_46__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_46__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_46__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_46__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_46__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_46__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_47__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_47__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_47__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_47__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_47__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_47__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_47__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_48__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_48__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_48__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_48__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_48__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_48__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_48__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_49__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_49__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_49__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_49__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_49__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_49__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_49__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_50__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_50__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_50__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_50__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_50__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_50__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_50__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_51__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_51__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_51__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_51__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_51__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_51__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_51__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_52__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_52__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_52__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_52__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_52__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_52__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_52__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_53__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_53__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_53__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_53__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_53__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_53__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_53__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_54__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_54__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_54__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_54__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_54__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_54__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_54__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_55__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_55__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_55__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_55__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_55__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_55__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_55__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_56__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_56__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_56__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_56__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_56__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_56__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_56__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_57__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_57__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_57__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_57__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_57__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_57__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_57__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_58__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_58__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_58__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_58__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_58__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_58__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_58__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_59__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_59__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_59__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_59__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_59__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_59__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_59__17_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_60__11_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_60__12_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_60__13_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_60__14_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_60__15_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_60__16_ ;
 wire u_multiplier_STAGE4_E_4_2_pp4_60__17_ ;
 wire u_multiplier_STAGE4_Full_adder_pp4_61__08_ ;
 wire u_multiplier_STAGE4_Full_adder_pp4_61__09_ ;
 wire u_multiplier_STAGE4_Full_adder_pp4_61__10_ ;
 wire u_multiplier_STAGE4_Full_adder_pp4_61__11_ ;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire valid_reg_out;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net134;
 wire net135;
 wire net136;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire clknet_0_clk;
 wire clknet_1_0_0_clk;
 wire clknet_1_1_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_4_0__leaf_clk;
 wire clknet_4_1__leaf_clk;
 wire clknet_4_2__leaf_clk;
 wire clknet_4_3__leaf_clk;
 wire clknet_4_4__leaf_clk;
 wire clknet_4_5__leaf_clk;
 wire clknet_4_6__leaf_clk;
 wire clknet_4_7__leaf_clk;
 wire clknet_4_8__leaf_clk;
 wire clknet_4_9__leaf_clk;
 wire clknet_4_10__leaf_clk;
 wire clknet_4_11__leaf_clk;
 wire clknet_4_12__leaf_clk;
 wire clknet_4_13__leaf_clk;
 wire clknet_4_14__leaf_clk;
 wire clknet_4_15__leaf_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire [5:0] addr_ptr;
 wire [2:0] curr_state;
 wire [31:0] data_in_reg;
 wire [5:0] init_count;
 wire [63:0] product;
 wire [31:0] sram_rdata;
 wire [31:0] sram_rdata_reg;
 wire [62:0] u_multiplier_A ;
 wire [62:0] u_multiplier_B ;
 wire [1:0] u_multiplier_pp1_1 ;
 wire [10:0] u_multiplier_pp1_10 ;
 wire [11:0] u_multiplier_pp1_11 ;
 wire [12:0] u_multiplier_pp1_12 ;
 wire [13:0] u_multiplier_pp1_13 ;
 wire [14:0] u_multiplier_pp1_14 ;
 wire [15:0] u_multiplier_pp1_15 ;
 wire [15:0] u_multiplier_pp1_16 ;
 wire [15:0] u_multiplier_pp1_17 ;
 wire [15:0] u_multiplier_pp1_18 ;
 wire [15:0] u_multiplier_pp1_19 ;
 wire [2:0] u_multiplier_pp1_2 ;
 wire [15:0] u_multiplier_pp1_20 ;
 wire [15:0] u_multiplier_pp1_21 ;
 wire [15:0] u_multiplier_pp1_22 ;
 wire [15:0] u_multiplier_pp1_23 ;
 wire [15:0] u_multiplier_pp1_24 ;
 wire [15:0] u_multiplier_pp1_25 ;
 wire [15:0] u_multiplier_pp1_26 ;
 wire [15:0] u_multiplier_pp1_27 ;
 wire [15:0] u_multiplier_pp1_28 ;
 wire [15:0] u_multiplier_pp1_29 ;
 wire [3:0] u_multiplier_pp1_3 ;
 wire [15:0] u_multiplier_pp1_30 ;
 wire [15:0] u_multiplier_pp1_31 ;
 wire [15:0] u_multiplier_pp1_32 ;
 wire [15:0] u_multiplier_pp1_33 ;
 wire [15:0] u_multiplier_pp1_34 ;
 wire [15:0] u_multiplier_pp1_35 ;
 wire [15:0] u_multiplier_pp1_36 ;
 wire [15:0] u_multiplier_pp1_37 ;
 wire [15:0] u_multiplier_pp1_38 ;
 wire [15:0] u_multiplier_pp1_39 ;
 wire [4:0] u_multiplier_pp1_4 ;
 wire [15:0] u_multiplier_pp1_40 ;
 wire [15:0] u_multiplier_pp1_41 ;
 wire [15:0] u_multiplier_pp1_42 ;
 wire [15:0] u_multiplier_pp1_43 ;
 wire [15:0] u_multiplier_pp1_44 ;
 wire [15:0] u_multiplier_pp1_45 ;
 wire [15:0] u_multiplier_pp1_46 ;
 wire [15:0] u_multiplier_pp1_47 ;
 wire [15:0] u_multiplier_pp1_48 ;
 wire [13:0] u_multiplier_pp1_49 ;
 wire [5:0] u_multiplier_pp1_5 ;
 wire [12:0] u_multiplier_pp1_50 ;
 wire [11:0] u_multiplier_pp1_51 ;
 wire [10:0] u_multiplier_pp1_52 ;
 wire [9:0] u_multiplier_pp1_53 ;
 wire [8:0] u_multiplier_pp1_54 ;
 wire [7:0] u_multiplier_pp1_55 ;
 wire [6:0] u_multiplier_pp1_56 ;
 wire [5:0] u_multiplier_pp1_57 ;
 wire [4:0] u_multiplier_pp1_58 ;
 wire [3:0] u_multiplier_pp1_59 ;
 wire [6:0] u_multiplier_pp1_6 ;
 wire [2:0] u_multiplier_pp1_60 ;
 wire [1:0] u_multiplier_pp1_61 ;
 wire [7:0] u_multiplier_pp1_7 ;
 wire [8:0] u_multiplier_pp1_8 ;
 wire [9:0] u_multiplier_pp1_9 ;
 wire [1:0] u_multiplier_pp2_1 ;
 wire [7:0] u_multiplier_pp2_10 ;
 wire [7:0] u_multiplier_pp2_11 ;
 wire [7:0] u_multiplier_pp2_12 ;
 wire [7:0] u_multiplier_pp2_13 ;
 wire [7:0] u_multiplier_pp2_14 ;
 wire [7:0] u_multiplier_pp2_15 ;
 wire [7:0] u_multiplier_pp2_16 ;
 wire [7:0] u_multiplier_pp2_17 ;
 wire [7:0] u_multiplier_pp2_18 ;
 wire [7:0] u_multiplier_pp2_19 ;
 wire [2:0] u_multiplier_pp2_2 ;
 wire [7:0] u_multiplier_pp2_20 ;
 wire [7:0] u_multiplier_pp2_21 ;
 wire [7:0] u_multiplier_pp2_22 ;
 wire [7:0] u_multiplier_pp2_23 ;
 wire [7:0] u_multiplier_pp2_24 ;
 wire [7:0] u_multiplier_pp2_25 ;
 wire [7:0] u_multiplier_pp2_26 ;
 wire [7:0] u_multiplier_pp2_27 ;
 wire [7:0] u_multiplier_pp2_28 ;
 wire [7:0] u_multiplier_pp2_29 ;
 wire [3:0] u_multiplier_pp2_3 ;
 wire [7:0] u_multiplier_pp2_30 ;
 wire [7:0] u_multiplier_pp2_31 ;
 wire [7:0] u_multiplier_pp2_32 ;
 wire [7:0] u_multiplier_pp2_33 ;
 wire [7:0] u_multiplier_pp2_34 ;
 wire [7:0] u_multiplier_pp2_35 ;
 wire [7:0] u_multiplier_pp2_36 ;
 wire [7:0] u_multiplier_pp2_37 ;
 wire [7:0] u_multiplier_pp2_38 ;
 wire [7:0] u_multiplier_pp2_39 ;
 wire [4:0] u_multiplier_pp2_4 ;
 wire [7:0] u_multiplier_pp2_40 ;
 wire [7:0] u_multiplier_pp2_41 ;
 wire [7:0] u_multiplier_pp2_42 ;
 wire [7:0] u_multiplier_pp2_43 ;
 wire [7:0] u_multiplier_pp2_44 ;
 wire [7:0] u_multiplier_pp2_45 ;
 wire [7:0] u_multiplier_pp2_46 ;
 wire [7:0] u_multiplier_pp2_47 ;
 wire [7:0] u_multiplier_pp2_48 ;
 wire [7:0] u_multiplier_pp2_49 ;
 wire [5:0] u_multiplier_pp2_5 ;
 wire [7:0] u_multiplier_pp2_50 ;
 wire [7:0] u_multiplier_pp2_51 ;
 wire [7:0] u_multiplier_pp2_52 ;
 wire [7:0] u_multiplier_pp2_53 ;
 wire [7:0] u_multiplier_pp2_54 ;
 wire [7:0] u_multiplier_pp2_55 ;
 wire [7:0] u_multiplier_pp2_56 ;
 wire [5:0] u_multiplier_pp2_57 ;
 wire [4:0] u_multiplier_pp2_58 ;
 wire [3:0] u_multiplier_pp2_59 ;
 wire [6:0] u_multiplier_pp2_6 ;
 wire [2:0] u_multiplier_pp2_60 ;
 wire [1:0] u_multiplier_pp2_61 ;
 wire [7:0] u_multiplier_pp2_7 ;
 wire [7:0] u_multiplier_pp2_8 ;
 wire [7:0] u_multiplier_pp2_9 ;
 wire [1:0] u_multiplier_pp3_1 ;
 wire [3:0] u_multiplier_pp3_10 ;
 wire [3:0] u_multiplier_pp3_11 ;
 wire [3:0] u_multiplier_pp3_12 ;
 wire [3:0] u_multiplier_pp3_13 ;
 wire [3:0] u_multiplier_pp3_14 ;
 wire [3:0] u_multiplier_pp3_15 ;
 wire [3:0] u_multiplier_pp3_16 ;
 wire [3:0] u_multiplier_pp3_17 ;
 wire [3:0] u_multiplier_pp3_18 ;
 wire [3:0] u_multiplier_pp3_19 ;
 wire [2:0] u_multiplier_pp3_2 ;
 wire [3:0] u_multiplier_pp3_20 ;
 wire [3:0] u_multiplier_pp3_21 ;
 wire [3:0] u_multiplier_pp3_22 ;
 wire [3:0] u_multiplier_pp3_23 ;
 wire [3:0] u_multiplier_pp3_24 ;
 wire [3:0] u_multiplier_pp3_25 ;
 wire [3:0] u_multiplier_pp3_26 ;
 wire [3:0] u_multiplier_pp3_27 ;
 wire [3:0] u_multiplier_pp3_28 ;
 wire [3:0] u_multiplier_pp3_29 ;
 wire [3:0] u_multiplier_pp3_3 ;
 wire [3:0] u_multiplier_pp3_30 ;
 wire [3:0] u_multiplier_pp3_31 ;
 wire [3:0] u_multiplier_pp3_32 ;
 wire [3:0] u_multiplier_pp3_33 ;
 wire [3:0] u_multiplier_pp3_34 ;
 wire [3:0] u_multiplier_pp3_35 ;
 wire [3:0] u_multiplier_pp3_36 ;
 wire [3:0] u_multiplier_pp3_37 ;
 wire [3:0] u_multiplier_pp3_38 ;
 wire [3:0] u_multiplier_pp3_39 ;
 wire [3:0] u_multiplier_pp3_4 ;
 wire [3:0] u_multiplier_pp3_40 ;
 wire [3:0] u_multiplier_pp3_41 ;
 wire [3:0] u_multiplier_pp3_42 ;
 wire [3:0] u_multiplier_pp3_43 ;
 wire [3:0] u_multiplier_pp3_44 ;
 wire [3:0] u_multiplier_pp3_45 ;
 wire [3:0] u_multiplier_pp3_46 ;
 wire [3:0] u_multiplier_pp3_47 ;
 wire [3:0] u_multiplier_pp3_48 ;
 wire [3:0] u_multiplier_pp3_49 ;
 wire [3:0] u_multiplier_pp3_5 ;
 wire [3:0] u_multiplier_pp3_50 ;
 wire [3:0] u_multiplier_pp3_51 ;
 wire [3:0] u_multiplier_pp3_52 ;
 wire [3:0] u_multiplier_pp3_53 ;
 wire [3:0] u_multiplier_pp3_54 ;
 wire [3:0] u_multiplier_pp3_55 ;
 wire [3:0] u_multiplier_pp3_56 ;
 wire [3:0] u_multiplier_pp3_57 ;
 wire [3:0] u_multiplier_pp3_58 ;
 wire [3:0] u_multiplier_pp3_59 ;
 wire [3:0] u_multiplier_pp3_6 ;
 wire [3:0] u_multiplier_pp3_60 ;
 wire [1:0] u_multiplier_pp3_61 ;
 wire [3:0] u_multiplier_pp3_7 ;
 wire [3:0] u_multiplier_pp3_8 ;
 wire [3:0] u_multiplier_pp3_9 ;

 INV_X2 _0675_ (.A(net9),
    .ZN(_0370_));
 INV_X2 _0676_ (.A(net43),
    .ZN(_0307_));
 INV_X1 _0677_ (.A(init_count[5]),
    .ZN(_0371_));
 INV_X1 _0678_ (.A(curr_state[2]),
    .ZN(_0372_));
 INV_X1 _0679_ (.A(net45),
    .ZN(_0373_));
 INV_X1 _0680_ (.A(net168),
    .ZN(_0374_));
 NOR2_X4 _0681_ (.A1(_0370_),
    .A2(_0373_),
    .ZN(_0303_));
 NAND2_X2 _0682_ (.A1(net9),
    .A2(net218),
    .ZN(_0308_));
 NAND2_X1 _0683_ (.A1(init_count[1]),
    .A2(init_count[0]),
    .ZN(_0375_));
 AND4_X2 _0684_ (.A1(init_count[1]),
    .A2(init_count[0]),
    .A3(init_count[3]),
    .A4(init_count[2]),
    .ZN(_0376_));
 INV_X1 _0685_ (.A(_0376_),
    .ZN(_0377_));
 AND2_X1 _0686_ (.A1(init_count[5]),
    .A2(init_count[4]),
    .ZN(_0378_));
 AND3_X1 _0687_ (.A1(net43),
    .A2(_0376_),
    .A3(_0378_),
    .ZN(_0379_));
 NOR2_X2 _0688_ (.A1(_0370_),
    .A2(_0307_),
    .ZN(_0380_));
 NAND2_X2 _0689_ (.A1(net9),
    .A2(net43),
    .ZN(_0381_));
 AND3_X1 _0690_ (.A1(curr_state[2]),
    .A2(_0376_),
    .A3(_0378_),
    .ZN(_0382_));
 NAND2_X1 _0691_ (.A1(_0380_),
    .A2(_0382_),
    .ZN(_0383_));
 OAI21_X1 _0692_ (.A(_0383_),
    .B1(_0373_),
    .B2(_0370_),
    .ZN(_0305_));
 NAND3_X1 _0693_ (.A1(net42),
    .A2(net192),
    .A3(_0380_),
    .ZN(_0384_));
 OAI21_X1 _0694_ (.A(net193),
    .B1(_0379_),
    .B2(_0308_),
    .ZN(_0306_));
 AOI22_X1 _0695_ (.A1(net9),
    .A2(net152),
    .B1(_0380_),
    .B2(net42),
    .ZN(_0304_));
 AND2_X1 _0696_ (.A1(net9),
    .A2(sram_rdata[0]),
    .ZN(_0271_));
 AND2_X1 _0697_ (.A1(net9),
    .A2(sram_rdata[1]),
    .ZN(_0282_));
 AND2_X1 _0698_ (.A1(net9),
    .A2(sram_rdata[2]),
    .ZN(_0293_));
 AND2_X1 _0699_ (.A1(net9),
    .A2(sram_rdata[3]),
    .ZN(_0296_));
 AND2_X1 _0700_ (.A1(net9),
    .A2(sram_rdata[4]),
    .ZN(_0297_));
 AND2_X1 _0701_ (.A1(net9),
    .A2(sram_rdata[5]),
    .ZN(_0298_));
 AND2_X1 _0702_ (.A1(net9),
    .A2(sram_rdata[6]),
    .ZN(_0299_));
 AND2_X1 _0703_ (.A1(net9),
    .A2(sram_rdata[7]),
    .ZN(_0300_));
 AND2_X1 _0704_ (.A1(net9),
    .A2(sram_rdata[8]),
    .ZN(_0301_));
 AND2_X1 _0705_ (.A1(net9),
    .A2(sram_rdata[9]),
    .ZN(_0302_));
 AND2_X1 _0706_ (.A1(net9),
    .A2(sram_rdata[10]),
    .ZN(_0272_));
 AND2_X1 _0707_ (.A1(net9),
    .A2(sram_rdata[11]),
    .ZN(_0273_));
 AND2_X1 _0708_ (.A1(net9),
    .A2(sram_rdata[12]),
    .ZN(_0274_));
 AND2_X1 _0709_ (.A1(net9),
    .A2(sram_rdata[13]),
    .ZN(_0275_));
 AND2_X1 _0710_ (.A1(net9),
    .A2(sram_rdata[14]),
    .ZN(_0276_));
 AND2_X1 _0711_ (.A1(net9),
    .A2(sram_rdata[15]),
    .ZN(_0277_));
 AND2_X1 _0712_ (.A1(net9),
    .A2(sram_rdata[16]),
    .ZN(_0278_));
 AND2_X1 _0713_ (.A1(net9),
    .A2(sram_rdata[17]),
    .ZN(_0279_));
 AND2_X1 _0714_ (.A1(net9),
    .A2(sram_rdata[18]),
    .ZN(_0280_));
 AND2_X1 _0715_ (.A1(net9),
    .A2(sram_rdata[19]),
    .ZN(_0281_));
 AND2_X1 _0716_ (.A1(net9),
    .A2(sram_rdata[20]),
    .ZN(_0283_));
 AND2_X1 _0717_ (.A1(net9),
    .A2(sram_rdata[21]),
    .ZN(_0284_));
 AND2_X1 _0718_ (.A1(net9),
    .A2(sram_rdata[22]),
    .ZN(_0285_));
 AND2_X1 _0719_ (.A1(net9),
    .A2(sram_rdata[23]),
    .ZN(_0286_));
 AND2_X1 _0720_ (.A1(net9),
    .A2(sram_rdata[24]),
    .ZN(_0287_));
 AND2_X1 _0721_ (.A1(net9),
    .A2(sram_rdata[25]),
    .ZN(_0288_));
 AND2_X1 _0722_ (.A1(net9),
    .A2(sram_rdata[26]),
    .ZN(_0289_));
 AND2_X1 _0723_ (.A1(net9),
    .A2(sram_rdata[27]),
    .ZN(_0290_));
 AND2_X1 _0724_ (.A1(net9),
    .A2(sram_rdata[28]),
    .ZN(_0291_));
 AND2_X1 _0725_ (.A1(net9),
    .A2(sram_rdata[29]),
    .ZN(_0292_));
 AND2_X1 _0726_ (.A1(net9),
    .A2(sram_rdata[30]),
    .ZN(_0294_));
 AND2_X1 _0727_ (.A1(net9),
    .A2(sram_rdata[31]),
    .ZN(_0295_));
 AND2_X1 _0728_ (.A1(product[0]),
    .A2(net7),
    .ZN(_0201_));
 AND2_X1 _0729_ (.A1(product[1]),
    .A2(net7),
    .ZN(_0212_));
 AND2_X1 _0730_ (.A1(product[2]),
    .A2(net7),
    .ZN(_0223_));
 AND2_X1 _0731_ (.A1(product[3]),
    .A2(net7),
    .ZN(_0234_));
 AND2_X1 _0732_ (.A1(product[4]),
    .A2(_0303_),
    .ZN(_0245_));
 AND2_X1 _0733_ (.A1(product[5]),
    .A2(_0303_),
    .ZN(_0256_));
 AND2_X1 _0734_ (.A1(product[6]),
    .A2(net7),
    .ZN(_0261_));
 AND2_X1 _0735_ (.A1(product[7]),
    .A2(net7),
    .ZN(_0262_));
 AND2_X1 _0736_ (.A1(product[8]),
    .A2(_0303_),
    .ZN(_0263_));
 AND2_X1 _0737_ (.A1(product[9]),
    .A2(_0303_),
    .ZN(_0264_));
 AND2_X1 _0738_ (.A1(product[10]),
    .A2(net7),
    .ZN(_0202_));
 AND2_X1 _0739_ (.A1(product[11]),
    .A2(_0303_),
    .ZN(_0203_));
 AND2_X1 _0740_ (.A1(product[12]),
    .A2(_0303_),
    .ZN(_0204_));
 AND2_X1 _0741_ (.A1(product[13]),
    .A2(net7),
    .ZN(_0205_));
 AND2_X1 _0742_ (.A1(product[14]),
    .A2(net7),
    .ZN(_0206_));
 AND2_X1 _0743_ (.A1(product[15]),
    .A2(net7),
    .ZN(_0207_));
 AND2_X1 _0744_ (.A1(product[16]),
    .A2(net7),
    .ZN(_0208_));
 AND2_X1 _0745_ (.A1(product[17]),
    .A2(net7),
    .ZN(_0209_));
 AND2_X1 _0746_ (.A1(product[18]),
    .A2(net7),
    .ZN(_0210_));
 AND2_X1 _0747_ (.A1(product[19]),
    .A2(_0303_),
    .ZN(_0211_));
 AND2_X1 _0748_ (.A1(product[20]),
    .A2(net7),
    .ZN(_0213_));
 AND2_X1 _0749_ (.A1(product[21]),
    .A2(net7),
    .ZN(_0214_));
 AND2_X1 _0750_ (.A1(product[22]),
    .A2(_0303_),
    .ZN(_0215_));
 AND2_X1 _0751_ (.A1(product[23]),
    .A2(_0303_),
    .ZN(_0216_));
 AND2_X1 _0752_ (.A1(product[24]),
    .A2(net7),
    .ZN(_0217_));
 AND2_X1 _0753_ (.A1(product[25]),
    .A2(_0303_),
    .ZN(_0218_));
 AND2_X1 _0754_ (.A1(product[26]),
    .A2(_0303_),
    .ZN(_0219_));
 AND2_X1 _0755_ (.A1(product[27]),
    .A2(_0303_),
    .ZN(_0220_));
 AND2_X1 _0756_ (.A1(product[28]),
    .A2(_0303_),
    .ZN(_0221_));
 AND2_X1 _0757_ (.A1(product[29]),
    .A2(net7),
    .ZN(_0222_));
 AND2_X1 _0758_ (.A1(product[30]),
    .A2(_0303_),
    .ZN(_0224_));
 AND2_X1 _0759_ (.A1(product[31]),
    .A2(_0303_),
    .ZN(_0225_));
 AND2_X1 _0760_ (.A1(product[32]),
    .A2(_0303_),
    .ZN(_0226_));
 AND2_X1 _0761_ (.A1(product[33]),
    .A2(net7),
    .ZN(_0227_));
 AND2_X1 _0762_ (.A1(product[34]),
    .A2(net7),
    .ZN(_0228_));
 AND2_X1 _0763_ (.A1(product[35]),
    .A2(net7),
    .ZN(_0229_));
 AND2_X1 _0764_ (.A1(product[36]),
    .A2(_0303_),
    .ZN(_0230_));
 AND2_X1 _0765_ (.A1(product[37]),
    .A2(_0303_),
    .ZN(_0231_));
 AND2_X1 _0766_ (.A1(product[38]),
    .A2(net7),
    .ZN(_0232_));
 AND2_X1 _0767_ (.A1(product[39]),
    .A2(_0303_),
    .ZN(_0233_));
 AND2_X1 _0768_ (.A1(product[40]),
    .A2(net7),
    .ZN(_0235_));
 AND2_X1 _0769_ (.A1(product[41]),
    .A2(net7),
    .ZN(_0236_));
 AND2_X1 _0770_ (.A1(product[42]),
    .A2(net7),
    .ZN(_0237_));
 AND2_X1 _0771_ (.A1(product[43]),
    .A2(_0303_),
    .ZN(_0238_));
 AND2_X1 _0772_ (.A1(product[44]),
    .A2(_0303_),
    .ZN(_0239_));
 AND2_X1 _0773_ (.A1(product[45]),
    .A2(_0303_),
    .ZN(_0240_));
 AND2_X1 _0774_ (.A1(product[46]),
    .A2(_0303_),
    .ZN(_0241_));
 AND2_X1 _0775_ (.A1(product[47]),
    .A2(_0303_),
    .ZN(_0242_));
 AND2_X1 _0776_ (.A1(product[48]),
    .A2(_0303_),
    .ZN(_0243_));
 AND2_X1 _0777_ (.A1(product[49]),
    .A2(_0303_),
    .ZN(_0244_));
 AND2_X1 _0778_ (.A1(product[50]),
    .A2(_0303_),
    .ZN(_0246_));
 AND2_X1 _0779_ (.A1(product[51]),
    .A2(_0303_),
    .ZN(_0247_));
 AND2_X1 _0780_ (.A1(product[52]),
    .A2(_0303_),
    .ZN(_0248_));
 AND2_X1 _0781_ (.A1(product[53]),
    .A2(net7),
    .ZN(_0249_));
 AND2_X1 _0782_ (.A1(product[54]),
    .A2(net7),
    .ZN(_0250_));
 AND2_X1 _0783_ (.A1(product[55]),
    .A2(net7),
    .ZN(_0251_));
 AND2_X1 _0784_ (.A1(product[56]),
    .A2(net7),
    .ZN(_0252_));
 AND2_X1 _0785_ (.A1(product[57]),
    .A2(net7),
    .ZN(_0253_));
 AND2_X1 _0786_ (.A1(product[58]),
    .A2(_0303_),
    .ZN(_0254_));
 AND2_X1 _0787_ (.A1(product[59]),
    .A2(net7),
    .ZN(_0255_));
 AND2_X1 _0788_ (.A1(product[60]),
    .A2(net7),
    .ZN(_0257_));
 AND2_X1 _0789_ (.A1(product[61]),
    .A2(_0303_),
    .ZN(_0258_));
 AND2_X1 _0790_ (.A1(product[62]),
    .A2(net7),
    .ZN(_0259_));
 AND2_X1 _0791_ (.A1(product[63]),
    .A2(net7),
    .ZN(_0260_));
 AND2_X1 _0792_ (.A1(net9),
    .A2(net10),
    .ZN(_0169_));
 AND2_X1 _0793_ (.A1(net8),
    .A2(net21),
    .ZN(_0180_));
 AND2_X1 _0794_ (.A1(net8),
    .A2(net32),
    .ZN(_0191_));
 AND2_X1 _0795_ (.A1(net9),
    .A2(net35),
    .ZN(_0194_));
 AND2_X1 _0796_ (.A1(net9),
    .A2(net36),
    .ZN(_0195_));
 AND2_X1 _0797_ (.A1(net8),
    .A2(net37),
    .ZN(_0196_));
 AND2_X1 _0798_ (.A1(net8),
    .A2(net38),
    .ZN(_0197_));
 AND2_X1 _0799_ (.A1(net8),
    .A2(net39),
    .ZN(_0198_));
 AND2_X1 _0800_ (.A1(net44),
    .A2(net40),
    .ZN(_0199_));
 AND2_X1 _0801_ (.A1(net9),
    .A2(net41),
    .ZN(_0200_));
 AND2_X1 _0802_ (.A1(net8),
    .A2(net11),
    .ZN(_0170_));
 AND2_X1 _0803_ (.A1(net8),
    .A2(net12),
    .ZN(_0171_));
 AND2_X1 _0804_ (.A1(net8),
    .A2(net13),
    .ZN(_0172_));
 AND2_X1 _0805_ (.A1(net9),
    .A2(net14),
    .ZN(_0173_));
 AND2_X1 _0806_ (.A1(net8),
    .A2(net15),
    .ZN(_0174_));
 AND2_X1 _0807_ (.A1(net8),
    .A2(net16),
    .ZN(_0175_));
 AND2_X1 _0808_ (.A1(net8),
    .A2(net17),
    .ZN(_0176_));
 AND2_X1 _0809_ (.A1(net9),
    .A2(net18),
    .ZN(_0177_));
 AND2_X1 _0810_ (.A1(net8),
    .A2(net19),
    .ZN(_0178_));
 AND2_X1 _0811_ (.A1(net9),
    .A2(net20),
    .ZN(_0179_));
 AND2_X1 _0812_ (.A1(net8),
    .A2(net22),
    .ZN(_0181_));
 AND2_X1 _0813_ (.A1(net8),
    .A2(net23),
    .ZN(_0182_));
 AND2_X1 _0814_ (.A1(net44),
    .A2(net24),
    .ZN(_0183_));
 AND2_X1 _0815_ (.A1(net9),
    .A2(net25),
    .ZN(_0184_));
 AND2_X1 _0816_ (.A1(net8),
    .A2(net26),
    .ZN(_0185_));
 AND2_X1 _0817_ (.A1(net8),
    .A2(net27),
    .ZN(_0186_));
 AND2_X1 _0818_ (.A1(net9),
    .A2(net28),
    .ZN(_0187_));
 AND2_X1 _0819_ (.A1(net9),
    .A2(net29),
    .ZN(_0188_));
 AND2_X1 _0820_ (.A1(net8),
    .A2(net30),
    .ZN(_0189_));
 AND2_X1 _0821_ (.A1(net8),
    .A2(net31),
    .ZN(_0190_));
 AND2_X1 _0822_ (.A1(net8),
    .A2(net33),
    .ZN(_0192_));
 AND2_X1 _0823_ (.A1(net8),
    .A2(net34),
    .ZN(_0193_));
 NAND2_X2 _0824_ (.A1(net9),
    .A2(_0307_),
    .ZN(_0385_));
 OAI21_X1 _0825_ (.A(net9),
    .B1(_0307_),
    .B2(_0382_),
    .ZN(_0386_));
 AOI21_X4 _0826_ (.A(_0372_),
    .B1(_0376_),
    .B2(_0378_),
    .ZN(_0387_));
 AOI22_X1 _0827_ (.A1(init_count[0]),
    .A2(net45),
    .B1(net170),
    .B2(_0387_),
    .ZN(_0388_));
 OAI22_X1 _0828_ (.A1(net171),
    .A2(_0386_),
    .B1(_0388_),
    .B2(_0381_),
    .ZN(_0265_));
 AOI21_X1 _0829_ (.A(net45),
    .B1(_0375_),
    .B2(curr_state[2]),
    .ZN(_0389_));
 INV_X1 _0830_ (.A(_0389_),
    .ZN(_0390_));
 AOI21_X1 _0831_ (.A(init_count[1]),
    .B1(init_count[0]),
    .B2(curr_state[2]),
    .ZN(_0391_));
 OR3_X1 _0832_ (.A1(_0381_),
    .A2(_0389_),
    .A3(_0391_),
    .ZN(_0392_));
 OAI211_X1 _0833_ (.A(_0383_),
    .B(_0392_),
    .C1(_0385_),
    .C2(net188),
    .ZN(_0266_));
 NOR3_X1 _0834_ (.A1(init_count[2]),
    .A2(_0372_),
    .A3(_0375_),
    .ZN(_0393_));
 AOI211_X1 _0835_ (.A(_0382_),
    .B(_0393_),
    .C1(_0390_),
    .C2(init_count[2]),
    .ZN(_0394_));
 OAI22_X1 _0836_ (.A1(net180),
    .A2(_0385_),
    .B1(_0394_),
    .B2(_0381_),
    .ZN(_0267_));
 NOR2_X1 _0837_ (.A1(_0658_),
    .A2(_0375_),
    .ZN(_0395_));
 XOR2_X1 _0838_ (.A(init_count[3]),
    .B(_0395_),
    .Z(_0396_));
 AOI221_X2 _0839_ (.A(_0382_),
    .B1(_0396_),
    .B2(curr_state[2]),
    .C1(net45),
    .C2(init_count[3]),
    .ZN(_0397_));
 OAI22_X1 _0840_ (.A1(net150),
    .A2(_0385_),
    .B1(_0397_),
    .B2(_0381_),
    .ZN(_0268_));
 NAND3_X1 _0841_ (.A1(_0371_),
    .A2(init_count[4]),
    .A3(_0376_),
    .ZN(_0398_));
 OAI21_X1 _0842_ (.A(curr_state[2]),
    .B1(_0376_),
    .B2(init_count[4]),
    .ZN(_0399_));
 INV_X1 _0843_ (.A(_0399_),
    .ZN(_0400_));
 AOI22_X1 _0844_ (.A1(net222),
    .A2(net45),
    .B1(_0398_),
    .B2(_0400_),
    .ZN(_0401_));
 OAI22_X1 _0845_ (.A1(net177),
    .A2(_0385_),
    .B1(_0401_),
    .B2(_0381_),
    .ZN(_0269_));
 OAI21_X1 _0846_ (.A(net182),
    .B1(_0377_),
    .B2(net176),
    .ZN(_0402_));
 AOI22_X1 _0847_ (.A1(net220),
    .A2(net45),
    .B1(_0402_),
    .B2(curr_state[2]),
    .ZN(_0403_));
 OAI22_X1 _0848_ (.A1(net183),
    .A2(_0385_),
    .B1(_0403_),
    .B2(_0381_),
    .ZN(_0270_));
 NOR2_X1 _0849_ (.A1(_0373_),
    .A2(addr_ptr[0]),
    .ZN(_0404_));
 AOI21_X1 _0850_ (.A(_0404_),
    .B1(_0387_),
    .B2(net3),
    .ZN(_0405_));
 OAI22_X1 _0851_ (.A1(net156),
    .A2(_0385_),
    .B1(net4),
    .B2(_0381_),
    .ZN(_0163_));
 NAND2_X1 _0852_ (.A1(addr_ptr[0]),
    .A2(addr_ptr[1]),
    .ZN(_0406_));
 XOR2_X1 _0853_ (.A(addr_ptr[0]),
    .B(net221),
    .Z(_0407_));
 OAI211_X1 _0854_ (.A(_0380_),
    .B(_0407_),
    .C1(_0387_),
    .C2(net45),
    .ZN(_0408_));
 OAI21_X1 _0855_ (.A(_0408_),
    .B1(_0385_),
    .B2(net2),
    .ZN(_0164_));
 AND4_X1 _0856_ (.A1(addr_ptr[0]),
    .A2(addr_ptr[1]),
    .A3(addr_ptr[3]),
    .A4(addr_ptr[2]),
    .ZN(_0409_));
 NAND3_X1 _0857_ (.A1(net197),
    .A2(addr_ptr[4]),
    .A3(_0409_),
    .ZN(_0410_));
 AOI21_X2 _0858_ (.A(_0387_),
    .B1(_0410_),
    .B2(net45),
    .ZN(_0411_));
 AOI21_X1 _0859_ (.A(_0381_),
    .B1(_0406_),
    .B2(net205),
    .ZN(_0412_));
 OAI21_X1 _0860_ (.A(_0412_),
    .B1(_0406_),
    .B2(net205),
    .ZN(_0413_));
 OAI22_X1 _0861_ (.A1(net206),
    .A2(_0385_),
    .B1(_0411_),
    .B2(_0413_),
    .ZN(_0165_));
 NOR3_X1 _0862_ (.A1(_0307_),
    .A2(net205),
    .A3(_0406_),
    .ZN(_0414_));
 OAI21_X1 _0863_ (.A(net9),
    .B1(_0374_),
    .B2(_0414_),
    .ZN(_0415_));
 AOI221_X1 _0864_ (.A(_0415_),
    .B1(_0414_),
    .B2(_0374_),
    .C1(net43),
    .C2(_0411_),
    .ZN(_0166_));
 NAND2_X1 _0865_ (.A1(net43),
    .A2(_0409_),
    .ZN(_0416_));
 OR2_X1 _0866_ (.A1(_0654_),
    .A2(_0416_),
    .ZN(_0417_));
 XNOR2_X1 _0867_ (.A(net189),
    .B(_0416_),
    .ZN(_0418_));
 AOI211_X1 _0868_ (.A(_0370_),
    .B(net190),
    .C1(_0411_),
    .C2(net43),
    .ZN(_0167_));
 XNOR2_X1 _0869_ (.A(net173),
    .B(_0417_),
    .ZN(_0419_));
 AOI211_X1 _0870_ (.A(_0370_),
    .B(net174),
    .C1(_0411_),
    .C2(net43),
    .ZN(_0168_));
 DFF_X1 _0871_ (.D(net153),
    .CK(clknet_4_7__leaf_clk),
    .Q(curr_state[0]),
    .QN(_0518_));
 DFF_X2 _0872_ (.D(_0305_),
    .CK(clknet_4_7__leaf_clk),
    .Q(net45),
    .QN(_0519_));
 DFF_X2 _0873_ (.D(net194),
    .CK(clknet_4_6__leaf_clk),
    .Q(curr_state[2]),
    .QN(_0520_));
 DFF_X2 _0874_ (.D(_0201_),
    .CK(clknet_4_15__leaf_clk),
    .Q(net46),
    .QN(_0521_));
 DFF_X2 _0875_ (.D(_0212_),
    .CK(clknet_4_14__leaf_clk),
    .Q(net57),
    .QN(_0522_));
 DFF_X2 _0876_ (.D(_0223_),
    .CK(clknet_4_15__leaf_clk),
    .Q(net68),
    .QN(_0523_));
 DFF_X2 _0877_ (.D(_0234_),
    .CK(clknet_4_14__leaf_clk),
    .Q(net79),
    .QN(_0524_));
 DFF_X1 _0878_ (.D(_0245_),
    .CK(clknet_4_1__leaf_clk),
    .Q(net90),
    .QN(_0525_));
 DFF_X1 _0879_ (.D(_0256_),
    .CK(clknet_4_1__leaf_clk),
    .Q(net101),
    .QN(_0526_));
 DFF_X2 _0880_ (.D(_0261_),
    .CK(clknet_4_15__leaf_clk),
    .Q(net106),
    .QN(_0527_));
 DFF_X2 _0881_ (.D(_0262_),
    .CK(clknet_4_15__leaf_clk),
    .Q(net107),
    .QN(_0528_));
 DFF_X2 _0882_ (.D(_0263_),
    .CK(clknet_4_4__leaf_clk),
    .Q(net108),
    .QN(_0529_));
 DFF_X2 _0883_ (.D(_0264_),
    .CK(clknet_4_4__leaf_clk),
    .Q(net109),
    .QN(_0530_));
 DFF_X2 _0884_ (.D(_0202_),
    .CK(clknet_4_14__leaf_clk),
    .Q(net47),
    .QN(_0531_));
 DFF_X2 _0885_ (.D(_0203_),
    .CK(clknet_4_3__leaf_clk),
    .Q(net48),
    .QN(_0532_));
 DFF_X2 _0886_ (.D(_0204_),
    .CK(clknet_4_2__leaf_clk),
    .Q(net49),
    .QN(_0533_));
 DFF_X2 _0887_ (.D(_0205_),
    .CK(clknet_4_2__leaf_clk),
    .Q(net50),
    .QN(_0534_));
 DFF_X2 _0888_ (.D(_0206_),
    .CK(clknet_4_11__leaf_clk),
    .Q(net51),
    .QN(_0535_));
 DFF_X2 _0889_ (.D(_0207_),
    .CK(clknet_4_14__leaf_clk),
    .Q(net52),
    .QN(_0536_));
 DFF_X2 _0890_ (.D(_0208_),
    .CK(clknet_4_14__leaf_clk),
    .Q(net53),
    .QN(_0537_));
 DFF_X2 _0891_ (.D(_0209_),
    .CK(clknet_4_13__leaf_clk),
    .Q(net54),
    .QN(_0538_));
 DFF_X2 _0892_ (.D(_0210_),
    .CK(clknet_4_14__leaf_clk),
    .Q(net55),
    .QN(_0539_));
 DFF_X2 _0893_ (.D(_0211_),
    .CK(clknet_4_3__leaf_clk),
    .Q(net56),
    .QN(_0540_));
 DFF_X2 _0894_ (.D(_0213_),
    .CK(clknet_4_15__leaf_clk),
    .Q(net58),
    .QN(_0541_));
 DFF_X2 _0895_ (.D(_0214_),
    .CK(clknet_4_15__leaf_clk),
    .Q(net59),
    .QN(_0542_));
 DFF_X2 _0896_ (.D(_0215_),
    .CK(clknet_4_6__leaf_clk),
    .Q(net60),
    .QN(_0543_));
 DFF_X1 _0897_ (.D(_0216_),
    .CK(clknet_4_6__leaf_clk),
    .Q(net61),
    .QN(_0544_));
 DFF_X2 _0898_ (.D(_0217_),
    .CK(clknet_4_15__leaf_clk),
    .Q(net62),
    .QN(_0545_));
 DFF_X1 _0899_ (.D(_0218_),
    .CK(clknet_4_5__leaf_clk),
    .Q(net63),
    .QN(_0546_));
 DFF_X1 _0900_ (.D(_0219_),
    .CK(clknet_4_4__leaf_clk),
    .Q(net64),
    .QN(_0547_));
 DFF_X2 _0901_ (.D(_0220_),
    .CK(clknet_4_5__leaf_clk),
    .Q(net65),
    .QN(_0548_));
 DFF_X2 _0902_ (.D(_0221_),
    .CK(clknet_4_4__leaf_clk),
    .Q(net66),
    .QN(_0549_));
 DFF_X1 _0903_ (.D(_0222_),
    .CK(clknet_4_14__leaf_clk),
    .Q(net67),
    .QN(_0550_));
 DFF_X1 _0904_ (.D(_0224_),
    .CK(clknet_4_1__leaf_clk),
    .Q(net69),
    .QN(_0551_));
 DFF_X1 _0905_ (.D(_0225_),
    .CK(clknet_4_1__leaf_clk),
    .Q(net70),
    .QN(_0552_));
 DFF_X1 _0906_ (.D(_0226_),
    .CK(clknet_4_2__leaf_clk),
    .Q(net71),
    .QN(_0553_));
 DFF_X2 _0907_ (.D(_0227_),
    .CK(clknet_4_14__leaf_clk),
    .Q(net72),
    .QN(_0554_));
 DFF_X2 _0908_ (.D(_0228_),
    .CK(clknet_4_14__leaf_clk),
    .Q(net73),
    .QN(_0555_));
 DFF_X2 _0909_ (.D(_0229_),
    .CK(clknet_4_13__leaf_clk),
    .Q(net74),
    .QN(_0556_));
 DFF_X1 _0910_ (.D(_0230_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net75),
    .QN(_0557_));
 DFF_X2 _0911_ (.D(_0231_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net76),
    .QN(_0558_));
 DFF_X2 _0912_ (.D(_0232_),
    .CK(clknet_4_12__leaf_clk),
    .Q(net77),
    .QN(_0559_));
 DFF_X2 _0913_ (.D(_0233_),
    .CK(clknet_4_2__leaf_clk),
    .Q(net78),
    .QN(_0560_));
 DFF_X2 _0914_ (.D(_0235_),
    .CK(clknet_4_12__leaf_clk),
    .Q(net80),
    .QN(_0561_));
 DFF_X2 _0915_ (.D(_0236_),
    .CK(clknet_4_8__leaf_clk),
    .Q(net81),
    .QN(_0562_));
 DFF_X2 _0916_ (.D(_0237_),
    .CK(clknet_4_12__leaf_clk),
    .Q(net82),
    .QN(_0563_));
 DFF_X2 _0917_ (.D(_0238_),
    .CK(clknet_4_2__leaf_clk),
    .Q(net83),
    .QN(_0564_));
 DFF_X2 _0918_ (.D(_0239_),
    .CK(clknet_4_3__leaf_clk),
    .Q(net84),
    .QN(_0565_));
 DFF_X2 _0919_ (.D(_0240_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net85),
    .QN(_0566_));
 DFF_X1 _0920_ (.D(_0241_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net86),
    .QN(_0567_));
 DFF_X2 _0921_ (.D(_0242_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net87),
    .QN(_0568_));
 DFF_X2 _0922_ (.D(_0243_),
    .CK(clknet_4_1__leaf_clk),
    .Q(net88),
    .QN(_0569_));
 DFF_X2 _0923_ (.D(_0244_),
    .CK(clknet_4_6__leaf_clk),
    .Q(net89),
    .QN(_0570_));
 DFF_X2 _0924_ (.D(_0246_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net91),
    .QN(_0571_));
 DFF_X1 _0925_ (.D(_0247_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net92),
    .QN(_0572_));
 DFF_X1 _0926_ (.D(_0248_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net93),
    .QN(_0573_));
 DFF_X2 _0927_ (.D(_0249_),
    .CK(clknet_4_12__leaf_clk),
    .Q(net94),
    .QN(_0574_));
 DFF_X2 _0928_ (.D(_0250_),
    .CK(clknet_4_2__leaf_clk),
    .Q(net95),
    .QN(_0575_));
 DFF_X1 _0929_ (.D(_0251_),
    .CK(clknet_4_8__leaf_clk),
    .Q(net96),
    .QN(_0576_));
 DFF_X2 _0930_ (.D(_0252_),
    .CK(clknet_4_13__leaf_clk),
    .Q(net97),
    .QN(_0577_));
 DFF_X2 _0931_ (.D(_0253_),
    .CK(clknet_4_13__leaf_clk),
    .Q(net98),
    .QN(_0578_));
 DFF_X2 _0932_ (.D(_0254_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net99),
    .QN(_0579_));
 DFF_X2 _0933_ (.D(_0255_),
    .CK(clknet_4_13__leaf_clk),
    .Q(net100),
    .QN(_0580_));
 DFF_X2 _0934_ (.D(_0257_),
    .CK(clknet_4_13__leaf_clk),
    .Q(net102),
    .QN(_0581_));
 DFF_X1 _0935_ (.D(_0258_),
    .CK(clknet_4_5__leaf_clk),
    .Q(net103),
    .QN(_0582_));
 DFF_X2 _0936_ (.D(_0259_),
    .CK(clknet_4_14__leaf_clk),
    .Q(net104),
    .QN(_0583_));
 DFF_X2 _0937_ (.D(_0260_),
    .CK(clknet_4_14__leaf_clk),
    .Q(net105),
    .QN(_0584_));
 DFF_X2 _0938_ (.D(_0169_),
    .CK(clknet_4_10__leaf_clk),
    .Q(data_in_reg[0]),
    .QN(_0585_));
 DFF_X2 _0939_ (.D(_0180_),
    .CK(clknet_4_0__leaf_clk),
    .Q(data_in_reg[1]),
    .QN(_0586_));
 DFF_X2 _0940_ (.D(_0191_),
    .CK(clknet_4_13__leaf_clk),
    .Q(data_in_reg[2]),
    .QN(_0587_));
 DFF_X2 _0941_ (.D(_0194_),
    .CK(clknet_4_11__leaf_clk),
    .Q(data_in_reg[3]),
    .QN(_0588_));
 DFF_X2 _0942_ (.D(_0195_),
    .CK(clknet_4_5__leaf_clk),
    .Q(data_in_reg[4]),
    .QN(_0589_));
 DFF_X2 _0943_ (.D(_0196_),
    .CK(clknet_4_15__leaf_clk),
    .Q(data_in_reg[5]),
    .QN(_0590_));
 DFF_X2 _0944_ (.D(_0197_),
    .CK(clknet_4_8__leaf_clk),
    .Q(data_in_reg[6]),
    .QN(_0591_));
 DFF_X2 _0945_ (.D(_0198_),
    .CK(clknet_4_5__leaf_clk),
    .Q(data_in_reg[7]),
    .QN(_0592_));
 DFF_X2 _0946_ (.D(_0199_),
    .CK(clknet_4_13__leaf_clk),
    .Q(data_in_reg[8]),
    .QN(_0593_));
 DFF_X2 _0947_ (.D(_0200_),
    .CK(clknet_4_4__leaf_clk),
    .Q(data_in_reg[9]),
    .QN(_0594_));
 DFF_X2 _0948_ (.D(_0170_),
    .CK(clknet_4_15__leaf_clk),
    .Q(data_in_reg[10]),
    .QN(_0595_));
 DFF_X2 _0949_ (.D(_0171_),
    .CK(clknet_4_5__leaf_clk),
    .Q(data_in_reg[11]),
    .QN(_0596_));
 DFF_X2 _0950_ (.D(_0172_),
    .CK(clknet_4_12__leaf_clk),
    .Q(data_in_reg[12]),
    .QN(_0597_));
 DFF_X2 _0951_ (.D(_0173_),
    .CK(clknet_4_1__leaf_clk),
    .Q(data_in_reg[13]),
    .QN(_0598_));
 DFF_X2 _0952_ (.D(_0174_),
    .CK(clknet_4_14__leaf_clk),
    .Q(data_in_reg[14]),
    .QN(_0599_));
 DFF_X2 _0953_ (.D(_0175_),
    .CK(clknet_4_12__leaf_clk),
    .Q(data_in_reg[15]),
    .QN(_0600_));
 DFF_X2 _0954_ (.D(_0176_),
    .CK(clknet_4_1__leaf_clk),
    .Q(data_in_reg[16]),
    .QN(_0601_));
 DFF_X2 _0955_ (.D(_0177_),
    .CK(clknet_4_4__leaf_clk),
    .Q(data_in_reg[17]),
    .QN(_0602_));
 DFF_X2 _0956_ (.D(_0178_),
    .CK(clknet_4_2__leaf_clk),
    .Q(data_in_reg[18]),
    .QN(_0603_));
 DFF_X2 _0957_ (.D(_0179_),
    .CK(clknet_4_1__leaf_clk),
    .Q(data_in_reg[19]),
    .QN(_0604_));
 DFF_X2 _0958_ (.D(_0181_),
    .CK(clknet_4_5__leaf_clk),
    .Q(data_in_reg[20]),
    .QN(_0605_));
 DFF_X2 _0959_ (.D(_0182_),
    .CK(clknet_4_5__leaf_clk),
    .Q(data_in_reg[21]),
    .QN(_0606_));
 DFF_X2 _0960_ (.D(_0183_),
    .CK(clknet_4_14__leaf_clk),
    .Q(data_in_reg[22]),
    .QN(_0607_));
 DFF_X2 _0961_ (.D(_0184_),
    .CK(clknet_4_9__leaf_clk),
    .Q(data_in_reg[23]),
    .QN(_0608_));
 DFF_X2 _0962_ (.D(_0185_),
    .CK(clknet_4_12__leaf_clk),
    .Q(data_in_reg[24]),
    .QN(_0609_));
 DFF_X2 _0963_ (.D(_0186_),
    .CK(clknet_4_4__leaf_clk),
    .Q(data_in_reg[25]),
    .QN(_0610_));
 DFF_X2 _0964_ (.D(_0187_),
    .CK(clknet_4_1__leaf_clk),
    .Q(data_in_reg[26]),
    .QN(_0611_));
 DFF_X2 _0965_ (.D(_0188_),
    .CK(clknet_4_1__leaf_clk),
    .Q(data_in_reg[27]),
    .QN(_0612_));
 DFF_X2 _0966_ (.D(_0189_),
    .CK(clknet_4_12__leaf_clk),
    .Q(data_in_reg[28]),
    .QN(_0613_));
 DFF_X2 _0967_ (.D(_0190_),
    .CK(clknet_4_8__leaf_clk),
    .Q(data_in_reg[29]),
    .QN(_0614_));
 DFF_X2 _0968_ (.D(_0192_),
    .CK(clknet_4_0__leaf_clk),
    .Q(data_in_reg[30]),
    .QN(_0615_));
 DFF_X2 _0969_ (.D(_0193_),
    .CK(clknet_4_14__leaf_clk),
    .Q(data_in_reg[31]),
    .QN(_0616_));
 DFF_X2 _0970_ (.D(_0271_),
    .CK(clknet_4_3__leaf_clk),
    .Q(sram_rdata_reg[0]),
    .QN(_0617_));
 DFF_X2 _0971_ (.D(_0282_),
    .CK(clknet_4_3__leaf_clk),
    .Q(sram_rdata_reg[1]),
    .QN(_0618_));
 DFF_X2 _0972_ (.D(_0293_),
    .CK(clknet_4_3__leaf_clk),
    .Q(sram_rdata_reg[2]),
    .QN(_0619_));
 DFF_X2 _0973_ (.D(_0296_),
    .CK(clknet_4_3__leaf_clk),
    .Q(sram_rdata_reg[3]),
    .QN(_0620_));
 DFF_X2 _0974_ (.D(_0297_),
    .CK(clknet_4_3__leaf_clk),
    .Q(sram_rdata_reg[4]),
    .QN(_0621_));
 DFF_X2 _0975_ (.D(_0298_),
    .CK(clknet_4_3__leaf_clk),
    .Q(sram_rdata_reg[5]),
    .QN(_0622_));
 DFF_X2 _0976_ (.D(_0299_),
    .CK(clknet_4_11__leaf_clk),
    .Q(sram_rdata_reg[6]),
    .QN(_0623_));
 DFF_X2 _0977_ (.D(_0300_),
    .CK(clknet_4_11__leaf_clk),
    .Q(sram_rdata_reg[7]),
    .QN(_0624_));
 DFF_X2 _0978_ (.D(_0301_),
    .CK(clknet_4_11__leaf_clk),
    .Q(sram_rdata_reg[8]),
    .QN(_0625_));
 DFF_X2 _0979_ (.D(_0302_),
    .CK(clknet_4_11__leaf_clk),
    .Q(sram_rdata_reg[9]),
    .QN(_0626_));
 DFF_X2 _0980_ (.D(_0272_),
    .CK(clknet_4_11__leaf_clk),
    .Q(sram_rdata_reg[10]),
    .QN(_0627_));
 DFF_X2 _0981_ (.D(_0273_),
    .CK(clknet_4_11__leaf_clk),
    .Q(sram_rdata_reg[11]),
    .QN(_0628_));
 DFF_X2 _0982_ (.D(_0274_),
    .CK(clknet_4_9__leaf_clk),
    .Q(sram_rdata_reg[12]),
    .QN(_0629_));
 DFF_X2 _0983_ (.D(_0275_),
    .CK(clknet_4_11__leaf_clk),
    .Q(sram_rdata_reg[13]),
    .QN(_0630_));
 DFF_X2 _0984_ (.D(_0276_),
    .CK(clknet_4_9__leaf_clk),
    .Q(sram_rdata_reg[14]),
    .QN(_0631_));
 DFF_X2 _0985_ (.D(_0277_),
    .CK(clknet_4_9__leaf_clk),
    .Q(sram_rdata_reg[15]),
    .QN(_0632_));
 DFF_X2 _0986_ (.D(_0278_),
    .CK(clknet_4_11__leaf_clk),
    .Q(sram_rdata_reg[16]),
    .QN(_0633_));
 DFF_X2 _0987_ (.D(_0279_),
    .CK(clknet_4_8__leaf_clk),
    .Q(sram_rdata_reg[17]),
    .QN(_0634_));
 DFF_X2 _0988_ (.D(_0280_),
    .CK(clknet_4_10__leaf_clk),
    .Q(sram_rdata_reg[18]),
    .QN(_0635_));
 DFF_X2 _0989_ (.D(_0281_),
    .CK(clknet_4_8__leaf_clk),
    .Q(sram_rdata_reg[19]),
    .QN(_0636_));
 DFF_X2 _0990_ (.D(_0283_),
    .CK(clknet_4_10__leaf_clk),
    .Q(sram_rdata_reg[20]),
    .QN(_0637_));
 DFF_X2 _0991_ (.D(_0284_),
    .CK(clknet_4_9__leaf_clk),
    .Q(sram_rdata_reg[21]),
    .QN(_0638_));
 DFF_X2 _0992_ (.D(_0285_),
    .CK(clknet_4_10__leaf_clk),
    .Q(sram_rdata_reg[22]),
    .QN(_0639_));
 DFF_X2 _0993_ (.D(_0286_),
    .CK(clknet_4_9__leaf_clk),
    .Q(sram_rdata_reg[23]),
    .QN(_0640_));
 DFF_X2 _0994_ (.D(_0287_),
    .CK(clknet_4_10__leaf_clk),
    .Q(sram_rdata_reg[24]),
    .QN(_0641_));
 DFF_X2 _0995_ (.D(_0288_),
    .CK(clknet_4_10__leaf_clk),
    .Q(sram_rdata_reg[25]),
    .QN(_0642_));
 DFF_X2 _0996_ (.D(_0289_),
    .CK(clknet_4_9__leaf_clk),
    .Q(sram_rdata_reg[26]),
    .QN(_0643_));
 DFF_X2 _0997_ (.D(_0290_),
    .CK(clknet_4_11__leaf_clk),
    .Q(sram_rdata_reg[27]),
    .QN(_0644_));
 DFF_X2 _0998_ (.D(_0291_),
    .CK(clknet_4_10__leaf_clk),
    .Q(sram_rdata_reg[28]),
    .QN(_0645_));
 DFF_X2 _0999_ (.D(_0292_),
    .CK(clknet_4_10__leaf_clk),
    .Q(sram_rdata_reg[29]),
    .QN(_0646_));
 DFF_X2 _1000_ (.D(_0294_),
    .CK(clknet_4_9__leaf_clk),
    .Q(sram_rdata_reg[30]),
    .QN(_0647_));
 DFF_X2 _1001_ (.D(_0295_),
    .CK(clknet_4_10__leaf_clk),
    .Q(sram_rdata_reg[31]),
    .QN(_0648_));
 DFF_X2 _1002_ (.D(net7),
    .CK(clknet_4_15__leaf_clk),
    .Q(net110),
    .QN(_0649_));
 DFF_X1 _1003_ (.D(net5),
    .CK(clknet_4_7__leaf_clk),
    .Q(addr_ptr[0]),
    .QN(_0650_));
 DFF_X1 _1004_ (.D(_0164_),
    .CK(clknet_4_7__leaf_clk),
    .Q(addr_ptr[1]),
    .QN(_0651_));
 DFF_X1 _1005_ (.D(_0165_),
    .CK(clknet_4_7__leaf_clk),
    .Q(addr_ptr[2]),
    .QN(_0652_));
 DFF_X1 _1006_ (.D(_0166_),
    .CK(clknet_4_7__leaf_clk),
    .Q(addr_ptr[3]),
    .QN(_0653_));
 DFF_X1 _1007_ (.D(net191),
    .CK(clknet_4_7__leaf_clk),
    .Q(addr_ptr[4]),
    .QN(_0654_));
 DFF_X1 _1008_ (.D(net175),
    .CK(clknet_4_7__leaf_clk),
    .Q(addr_ptr[5]),
    .QN(_0655_));
 DFF_X1 _1009_ (.D(net172),
    .CK(clknet_4_7__leaf_clk),
    .Q(init_count[0]),
    .QN(_0656_));
 DFF_X1 _1010_ (.D(_0266_),
    .CK(clknet_4_7__leaf_clk),
    .Q(init_count[1]),
    .QN(_0657_));
 DFF_X1 _1011_ (.D(net181),
    .CK(clknet_4_6__leaf_clk),
    .Q(init_count[2]),
    .QN(_0658_));
 DFF_X1 _1012_ (.D(net151),
    .CK(clknet_4_6__leaf_clk),
    .Q(init_count[3]),
    .QN(_0659_));
 DFF_X1 _1013_ (.D(net178),
    .CK(clknet_4_6__leaf_clk),
    .Q(init_count[4]),
    .QN(_0660_));
 DFF_X1 _1014_ (.D(net184),
    .CK(clknet_4_6__leaf_clk),
    .Q(init_count[5]),
    .QN(_0661_));
 SRAM_6T_CORE_64x32_MC_TB sram_inst (.ce_in(_0307_),
    .we_in(_0308_),
    .clk(clknet_4_3__leaf_clk),
    .addr_in({net198,
    net196,
    net186,
    net169,
    net200,
    net202}),
    .rd_out({sram_rdata[31],
    sram_rdata[30],
    sram_rdata[29],
    sram_rdata[28],
    sram_rdata[27],
    sram_rdata[26],
    sram_rdata[25],
    sram_rdata[24],
    sram_rdata[23],
    sram_rdata[22],
    sram_rdata[21],
    sram_rdata[20],
    sram_rdata[19],
    sram_rdata[18],
    sram_rdata[17],
    sram_rdata[16],
    sram_rdata[15],
    sram_rdata[14],
    sram_rdata[13],
    sram_rdata[12],
    sram_rdata[11],
    sram_rdata[10],
    sram_rdata[9],
    sram_rdata[8],
    sram_rdata[7],
    sram_rdata[6],
    sram_rdata[5],
    sram_rdata[4],
    sram_rdata[3],
    sram_rdata[2],
    sram_rdata[1],
    sram_rdata[0]}),
    .wd_in({net210,
    data_in_reg[30],
    net219,
    net215,
    data_in_reg[27],
    data_in_reg[26],
    data_in_reg[25],
    net203,
    net204,
    net212,
    data_in_reg[21],
    data_in_reg[20],
    data_in_reg[19],
    data_in_reg[18],
    data_in_reg[17],
    data_in_reg[16],
    net207,
    data_in_reg[14],
    data_in_reg[13],
    net209,
    data_in_reg[11],
    data_in_reg[10],
    data_in_reg[9],
    data_in_reg[8],
    data_in_reg[7],
    net216,
    data_in_reg[5],
    data_in_reg[4],
    net214,
    data_in_reg[2],
    data_in_reg[1],
    net208}));
 AND2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__40_  (.A1(net137),
    .A2(u_multiplier_pp3_0 ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla1__25_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__41_  (.A1(net138),
    .A2(u_multiplier_pp3_0 ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla1__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__42_  (.A(net139),
    .B(u_multiplier_pp3_0 ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla1__27_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__43_  (.A(net142),
    .B(u_multiplier_Final_add_cla1_cla1_cla1_cla1__27_ ),
    .ZN(product[0]));
 AOI21_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__44_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla1__25_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla1_cla1__26_ ),
    .B2(net143),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla1__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__45_  (.A1(u_multiplier_pp3_1 [0]),
    .A2(u_multiplier_pp3_1 [1]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla1__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__46_  (.A1(u_multiplier_pp3_1 [0]),
    .A2(u_multiplier_pp3_1 [1]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla1__30_ ));
 XOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__47_  (.A(u_multiplier_pp3_1 [0]),
    .B(u_multiplier_pp3_1 [1]),
    .Z(u_multiplier_Final_add_cla1_cla1_cla1_cla1__31_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__48_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla1__28_ ),
    .B(u_multiplier_Final_add_cla1_cla1_cla1_cla1__31_ ),
    .ZN(product[1]));
 OAI21_X2 u_multiplier_Final_add_cla1_cla1_cla1_cla1__49_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla1__30_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla1_cla1__29_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla1_cla1__28_ ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla1__32_ ));
 AND2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__50_  (.A1(u_multiplier_pp3_2 [2]),
    .A2(u_multiplier_A [2]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla1__33_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__51_  (.A1(u_multiplier_pp3_2 [2]),
    .A2(u_multiplier_A [2]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla1__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__52_  (.A(u_multiplier_pp3_2 [2]),
    .B(u_multiplier_A [2]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla1__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__53_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla1__32_ ),
    .B(u_multiplier_Final_add_cla1_cla1_cla1_cla1__35_ ),
    .ZN(product[2]));
 AOI21_X2 u_multiplier_Final_add_cla1_cla1_cla1_cla1__54_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla1__33_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla1_cla1__34_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla1_cla1__32_ ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla1__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__55_  (.A1(u_multiplier_B [3]),
    .A2(u_multiplier_A [3]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla1__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__56_  (.A1(u_multiplier_B [3]),
    .A2(u_multiplier_A [3]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla1__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__57_  (.A(u_multiplier_B [3]),
    .B(u_multiplier_A [3]),
    .Z(u_multiplier_Final_add_cla1_cla1_cla1_cla1__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__58_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla1__36_ ),
    .B(u_multiplier_Final_add_cla1_cla1_cla1_cla1__39_ ),
    .ZN(product[3]));
 OAI21_X4 u_multiplier_Final_add_cla1_cla1_cla1_cla1__59_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla1__38_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla1_cla1__37_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla1_cla1__36_ ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_c1 ));
 AND2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__40_  (.A1(u_multiplier_B [4]),
    .A2(u_multiplier_A [4]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla2__25_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__41_  (.A1(u_multiplier_B [4]),
    .A2(u_multiplier_A [4]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla2__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__42_  (.A(u_multiplier_B [4]),
    .B(u_multiplier_A [4]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla2__27_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__43_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_c1 ),
    .B(u_multiplier_Final_add_cla1_cla1_cla1_cla2__27_ ),
    .ZN(product[4]));
 AOI21_X2 u_multiplier_Final_add_cla1_cla1_cla1_cla2__44_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla2__25_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla1_cla2__26_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla1_c1 ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla2__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__45_  (.A1(u_multiplier_B [5]),
    .A2(u_multiplier_A [5]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla2__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__46_  (.A1(u_multiplier_B [5]),
    .A2(u_multiplier_A [5]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla2__30_ ));
 XOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__47_  (.A(u_multiplier_B [5]),
    .B(u_multiplier_A [5]),
    .Z(u_multiplier_Final_add_cla1_cla1_cla1_cla2__31_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__48_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla2__28_ ),
    .B(u_multiplier_Final_add_cla1_cla1_cla1_cla2__31_ ),
    .ZN(product[5]));
 OAI21_X2 u_multiplier_Final_add_cla1_cla1_cla1_cla2__49_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla2__30_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla1_cla2__29_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla1_cla2__28_ ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla2__32_ ));
 AND2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__50_  (.A1(u_multiplier_B [6]),
    .A2(u_multiplier_A [6]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla2__33_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__51_  (.A1(u_multiplier_B [6]),
    .A2(u_multiplier_A [6]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla2__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__52_  (.A(u_multiplier_B [6]),
    .B(u_multiplier_A [6]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla2__35_ ));
 XNOR2_X2 u_multiplier_Final_add_cla1_cla1_cla1_cla2__53_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla2__32_ ),
    .B(u_multiplier_Final_add_cla1_cla1_cla1_cla2__35_ ),
    .ZN(product[6]));
 AOI21_X2 u_multiplier_Final_add_cla1_cla1_cla1_cla2__54_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla2__33_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla1_cla2__34_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla1_cla2__32_ ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla2__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__55_  (.A1(u_multiplier_B [7]),
    .A2(u_multiplier_A [7]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla2__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla2__56_  (.A1(u_multiplier_B [7]),
    .A2(u_multiplier_A [7]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla1_cla2__38_ ));
 XOR2_X2 u_multiplier_Final_add_cla1_cla1_cla1_cla2__57_  (.A(u_multiplier_B [7]),
    .B(u_multiplier_A [7]),
    .Z(u_multiplier_Final_add_cla1_cla1_cla1_cla2__39_ ));
 XNOR2_X2 u_multiplier_Final_add_cla1_cla1_cla1_cla2__58_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla2__36_ ),
    .B(u_multiplier_Final_add_cla1_cla1_cla1_cla2__39_ ),
    .ZN(product[7]));
 OAI21_X2 u_multiplier_Final_add_cla1_cla1_cla1_cla2__59_  (.A(u_multiplier_Final_add_cla1_cla1_cla1_cla2__38_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla1_cla2__37_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla1_cla2__36_ ),
    .ZN(u_multiplier_Final_add_cla1_cla1_c1 ));
 AND2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__40_  (.A1(u_multiplier_B [8]),
    .A2(u_multiplier_A [8]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla1__25_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__41_  (.A1(u_multiplier_B [8]),
    .A2(u_multiplier_A [8]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla1__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__42_  (.A(u_multiplier_B [8]),
    .B(u_multiplier_A [8]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla1__27_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__43_  (.A(u_multiplier_Final_add_cla1_cla1_c1 ),
    .B(u_multiplier_Final_add_cla1_cla1_cla2_cla1__27_ ),
    .ZN(product[8]));
 AOI21_X2 u_multiplier_Final_add_cla1_cla1_cla2_cla1__44_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla1__25_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla2_cla1__26_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_c1 ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla1__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__45_  (.A1(u_multiplier_B [9]),
    .A2(u_multiplier_A [9]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla1__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__46_  (.A1(u_multiplier_B [9]),
    .A2(u_multiplier_A [9]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla1__30_ ));
 XOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__47_  (.A(u_multiplier_B [9]),
    .B(u_multiplier_A [9]),
    .Z(u_multiplier_Final_add_cla1_cla1_cla2_cla1__31_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__48_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla1__28_ ),
    .B(u_multiplier_Final_add_cla1_cla1_cla2_cla1__31_ ),
    .ZN(product[9]));
 OAI21_X2 u_multiplier_Final_add_cla1_cla1_cla2_cla1__49_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla1__30_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla2_cla1__29_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla2_cla1__28_ ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla1__32_ ));
 AND2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__50_  (.A1(u_multiplier_B [10]),
    .A2(u_multiplier_A [10]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla1__33_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__51_  (.A1(u_multiplier_B [10]),
    .A2(u_multiplier_A [10]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla1__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__52_  (.A(u_multiplier_B [10]),
    .B(u_multiplier_A [10]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla1__35_ ));
 XNOR2_X2 u_multiplier_Final_add_cla1_cla1_cla2_cla1__53_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla1__32_ ),
    .B(u_multiplier_Final_add_cla1_cla1_cla2_cla1__35_ ),
    .ZN(product[10]));
 AOI21_X2 u_multiplier_Final_add_cla1_cla1_cla2_cla1__54_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla1__33_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla2_cla1__34_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla2_cla1__32_ ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla1__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__55_  (.A1(u_multiplier_B [11]),
    .A2(u_multiplier_A [11]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla1__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__56_  (.A1(u_multiplier_B [11]),
    .A2(u_multiplier_A [11]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla1__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__57_  (.A(u_multiplier_B [11]),
    .B(u_multiplier_A [11]),
    .Z(u_multiplier_Final_add_cla1_cla1_cla2_cla1__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla1__58_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla1__36_ ),
    .B(u_multiplier_Final_add_cla1_cla1_cla2_cla1__39_ ),
    .ZN(product[11]));
 OAI21_X2 u_multiplier_Final_add_cla1_cla1_cla2_cla1__59_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla1__38_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla2_cla1__37_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla2_cla1__36_ ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_c1 ));
 AND2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__40_  (.A1(u_multiplier_B [12]),
    .A2(u_multiplier_A [12]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla2__25_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__41_  (.A1(u_multiplier_B [12]),
    .A2(u_multiplier_A [12]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla2__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__42_  (.A(u_multiplier_B [12]),
    .B(u_multiplier_A [12]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla2__27_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__43_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_c1 ),
    .B(u_multiplier_Final_add_cla1_cla1_cla2_cla2__27_ ),
    .ZN(product[12]));
 AOI21_X4 u_multiplier_Final_add_cla1_cla1_cla2_cla2__44_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla2__25_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla2_cla2__26_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla2_c1 ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla2__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__45_  (.A1(u_multiplier_B [13]),
    .A2(u_multiplier_A [13]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla2__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__46_  (.A1(u_multiplier_B [13]),
    .A2(u_multiplier_A [13]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla2__30_ ));
 XOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__47_  (.A(u_multiplier_B [13]),
    .B(u_multiplier_A [13]),
    .Z(u_multiplier_Final_add_cla1_cla1_cla2_cla2__31_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__48_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla2__28_ ),
    .B(u_multiplier_Final_add_cla1_cla1_cla2_cla2__31_ ),
    .ZN(product[13]));
 OAI21_X2 u_multiplier_Final_add_cla1_cla1_cla2_cla2__49_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla2__30_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla2_cla2__29_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla2_cla2__28_ ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla2__32_ ));
 AND2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__50_  (.A1(u_multiplier_B [14]),
    .A2(u_multiplier_A [14]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla2__33_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__51_  (.A1(u_multiplier_B [14]),
    .A2(u_multiplier_A [14]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla2__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__52_  (.A(u_multiplier_B [14]),
    .B(u_multiplier_A [14]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla2__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__53_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla2__32_ ),
    .B(u_multiplier_Final_add_cla1_cla1_cla2_cla2__35_ ),
    .ZN(product[14]));
 AOI21_X4 u_multiplier_Final_add_cla1_cla1_cla2_cla2__54_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla2__33_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla2_cla2__34_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla2_cla2__32_ ),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla2__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__55_  (.A1(u_multiplier_B [15]),
    .A2(u_multiplier_A [15]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla2__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla1_cla2_cla2__56_  (.A1(u_multiplier_B [15]),
    .A2(u_multiplier_A [15]),
    .ZN(u_multiplier_Final_add_cla1_cla1_cla2_cla2__38_ ));
 XOR2_X2 u_multiplier_Final_add_cla1_cla1_cla2_cla2__57_  (.A(u_multiplier_B [15]),
    .B(u_multiplier_A [15]),
    .Z(u_multiplier_Final_add_cla1_cla1_cla2_cla2__39_ ));
 XNOR2_X2 u_multiplier_Final_add_cla1_cla1_cla2_cla2__58_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla2__36_ ),
    .B(u_multiplier_Final_add_cla1_cla1_cla2_cla2__39_ ),
    .ZN(product[15]));
 OAI21_X2 u_multiplier_Final_add_cla1_cla1_cla2_cla2__59_  (.A(u_multiplier_Final_add_cla1_cla1_cla2_cla2__38_ ),
    .B1(u_multiplier_Final_add_cla1_cla1_cla2_cla2__37_ ),
    .B2(u_multiplier_Final_add_cla1_cla1_cla2_cla2__36_ ),
    .ZN(u_multiplier_Final_add_cla1_c1 ));
 AND2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__40_  (.A1(u_multiplier_B [16]),
    .A2(u_multiplier_A [16]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla1__25_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__41_  (.A1(u_multiplier_B [16]),
    .A2(u_multiplier_A [16]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla1__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__42_  (.A(u_multiplier_B [16]),
    .B(u_multiplier_A [16]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla1__27_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__43_  (.A(u_multiplier_Final_add_cla1_c1 ),
    .B(u_multiplier_Final_add_cla1_cla2_cla1_cla1__27_ ),
    .ZN(product[16]));
 AOI21_X2 u_multiplier_Final_add_cla1_cla2_cla1_cla1__44_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla1__25_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla1_cla1__26_ ),
    .B2(u_multiplier_Final_add_cla1_c1 ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla1__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__45_  (.A1(u_multiplier_B [17]),
    .A2(u_multiplier_A [17]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla1__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__46_  (.A1(u_multiplier_B [17]),
    .A2(u_multiplier_A [17]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla1__30_ ));
 XOR2_X2 u_multiplier_Final_add_cla1_cla2_cla1_cla1__47_  (.A(u_multiplier_B [17]),
    .B(u_multiplier_A [17]),
    .Z(u_multiplier_Final_add_cla1_cla2_cla1_cla1__31_ ));
 XNOR2_X2 u_multiplier_Final_add_cla1_cla2_cla1_cla1__48_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla1__28_ ),
    .B(u_multiplier_Final_add_cla1_cla2_cla1_cla1__31_ ),
    .ZN(product[17]));
 OAI21_X2 u_multiplier_Final_add_cla1_cla2_cla1_cla1__49_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla1__30_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla1_cla1__29_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla1_cla1__28_ ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla1__32_ ));
 AND2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__50_  (.A1(u_multiplier_B [18]),
    .A2(u_multiplier_A [18]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla1__33_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__51_  (.A1(u_multiplier_B [18]),
    .A2(u_multiplier_A [18]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla1__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__52_  (.A(u_multiplier_B [18]),
    .B(u_multiplier_A [18]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla1__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__53_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla1__32_ ),
    .B(u_multiplier_Final_add_cla1_cla2_cla1_cla1__35_ ),
    .ZN(product[18]));
 AOI21_X4 u_multiplier_Final_add_cla1_cla2_cla1_cla1__54_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla1__33_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla1_cla1__34_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla1_cla1__32_ ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla1__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__55_  (.A1(u_multiplier_B [19]),
    .A2(u_multiplier_A [19]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla1__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__56_  (.A1(u_multiplier_B [19]),
    .A2(u_multiplier_A [19]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla1__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__57_  (.A(u_multiplier_B [19]),
    .B(u_multiplier_A [19]),
    .Z(u_multiplier_Final_add_cla1_cla2_cla1_cla1__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla1__58_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla1__36_ ),
    .B(u_multiplier_Final_add_cla1_cla2_cla1_cla1__39_ ),
    .ZN(product[19]));
 OAI21_X4 u_multiplier_Final_add_cla1_cla2_cla1_cla1__59_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla1__38_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla1_cla1__37_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla1_cla1__36_ ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_c1 ));
 AND2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla2__40_  (.A1(u_multiplier_B [20]),
    .A2(u_multiplier_A [20]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla2__25_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla2__41_  (.A1(u_multiplier_B [20]),
    .A2(u_multiplier_A [20]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla2__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla2__42_  (.A(u_multiplier_B [20]),
    .B(u_multiplier_A [20]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla2__27_ ));
 XNOR2_X2 u_multiplier_Final_add_cla1_cla2_cla1_cla2__43_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_c1 ),
    .B(u_multiplier_Final_add_cla1_cla2_cla1_cla2__27_ ),
    .ZN(product[20]));
 AOI21_X4 u_multiplier_Final_add_cla1_cla2_cla1_cla2__44_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla2__25_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla1_cla2__26_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla1_c1 ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla2__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla2__45_  (.A1(u_multiplier_B [21]),
    .A2(u_multiplier_A [21]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla2__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla2__46_  (.A1(u_multiplier_B [21]),
    .A2(u_multiplier_A [21]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla2__30_ ));
 XOR2_X2 u_multiplier_Final_add_cla1_cla2_cla1_cla2__47_  (.A(u_multiplier_B [21]),
    .B(u_multiplier_A [21]),
    .Z(u_multiplier_Final_add_cla1_cla2_cla1_cla2__31_ ));
 XNOR2_X2 u_multiplier_Final_add_cla1_cla2_cla1_cla2__48_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla2__28_ ),
    .B(u_multiplier_Final_add_cla1_cla2_cla1_cla2__31_ ),
    .ZN(product[21]));
 OAI21_X2 u_multiplier_Final_add_cla1_cla2_cla1_cla2__49_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla2__30_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla1_cla2__29_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla1_cla2__28_ ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla2__32_ ));
 AND2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla2__50_  (.A1(u_multiplier_B [22]),
    .A2(u_multiplier_A [22]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla2__33_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla2__51_  (.A1(u_multiplier_B [22]),
    .A2(u_multiplier_A [22]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla2__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla2__52_  (.A(u_multiplier_B [22]),
    .B(u_multiplier_A [22]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla2__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla2__53_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla2__32_ ),
    .B(u_multiplier_Final_add_cla1_cla2_cla1_cla2__35_ ),
    .ZN(product[22]));
 AOI21_X2 u_multiplier_Final_add_cla1_cla2_cla1_cla2__54_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla2__33_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla1_cla2__34_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla1_cla2__32_ ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla2__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla2__55_  (.A1(u_multiplier_B [23]),
    .A2(u_multiplier_A [23]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla2__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla2__56_  (.A1(u_multiplier_B [23]),
    .A2(u_multiplier_A [23]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla1_cla2__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla2__57_  (.A(u_multiplier_B [23]),
    .B(u_multiplier_A [23]),
    .Z(u_multiplier_Final_add_cla1_cla2_cla1_cla2__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla1_cla2__58_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla2__36_ ),
    .B(u_multiplier_Final_add_cla1_cla2_cla1_cla2__39_ ),
    .ZN(product[23]));
 OAI21_X2 u_multiplier_Final_add_cla1_cla2_cla1_cla2__59_  (.A(u_multiplier_Final_add_cla1_cla2_cla1_cla2__38_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla1_cla2__37_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla1_cla2__36_ ),
    .ZN(u_multiplier_Final_add_cla1_cla2_c1 ));
 AND2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__40_  (.A1(u_multiplier_B [24]),
    .A2(u_multiplier_A [24]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla1__25_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__41_  (.A1(u_multiplier_B [24]),
    .A2(u_multiplier_A [24]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla1__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__42_  (.A(u_multiplier_B [24]),
    .B(u_multiplier_A [24]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla1__27_ ));
 XNOR2_X2 u_multiplier_Final_add_cla1_cla2_cla2_cla1__43_  (.A(u_multiplier_Final_add_cla1_cla2_c1 ),
    .B(u_multiplier_Final_add_cla1_cla2_cla2_cla1__27_ ),
    .ZN(product[24]));
 AOI21_X2 u_multiplier_Final_add_cla1_cla2_cla2_cla1__44_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla1__25_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla2_cla1__26_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_c1 ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla1__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__45_  (.A1(u_multiplier_B [25]),
    .A2(u_multiplier_A [25]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla1__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__46_  (.A1(u_multiplier_B [25]),
    .A2(u_multiplier_A [25]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla1__30_ ));
 XOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__47_  (.A(u_multiplier_B [25]),
    .B(u_multiplier_A [25]),
    .Z(u_multiplier_Final_add_cla1_cla2_cla2_cla1__31_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__48_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla1__28_ ),
    .B(u_multiplier_Final_add_cla1_cla2_cla2_cla1__31_ ),
    .ZN(product[25]));
 OAI21_X2 u_multiplier_Final_add_cla1_cla2_cla2_cla1__49_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla1__30_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla2_cla1__29_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla2_cla1__28_ ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla1__32_ ));
 AND2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__50_  (.A1(u_multiplier_B [26]),
    .A2(u_multiplier_A [26]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla1__33_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__51_  (.A1(u_multiplier_B [26]),
    .A2(u_multiplier_A [26]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla1__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__52_  (.A(u_multiplier_B [26]),
    .B(u_multiplier_A [26]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla1__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__53_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla1__32_ ),
    .B(u_multiplier_Final_add_cla1_cla2_cla2_cla1__35_ ),
    .ZN(product[26]));
 AOI21_X2 u_multiplier_Final_add_cla1_cla2_cla2_cla1__54_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla1__33_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla2_cla1__34_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla2_cla1__32_ ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla1__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__55_  (.A1(u_multiplier_B [27]),
    .A2(u_multiplier_A [27]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla1__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__56_  (.A1(u_multiplier_B [27]),
    .A2(u_multiplier_A [27]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla1__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__57_  (.A(u_multiplier_B [27]),
    .B(u_multiplier_A [27]),
    .Z(u_multiplier_Final_add_cla1_cla2_cla2_cla1__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla1__58_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla1__36_ ),
    .B(u_multiplier_Final_add_cla1_cla2_cla2_cla1__39_ ),
    .ZN(product[27]));
 OAI21_X2 u_multiplier_Final_add_cla1_cla2_cla2_cla1__59_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla1__38_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla2_cla1__37_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla2_cla1__36_ ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_c1 ));
 AND2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__40_  (.A1(u_multiplier_B [28]),
    .A2(u_multiplier_A [28]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla2__25_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__41_  (.A1(u_multiplier_B [28]),
    .A2(u_multiplier_A [28]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla2__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__42_  (.A(u_multiplier_B [28]),
    .B(u_multiplier_A [28]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla2__27_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__43_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_c1 ),
    .B(u_multiplier_Final_add_cla1_cla2_cla2_cla2__27_ ),
    .ZN(product[28]));
 AOI21_X4 u_multiplier_Final_add_cla1_cla2_cla2_cla2__44_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla2__25_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla2_cla2__26_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla2_c1 ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla2__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__45_  (.A1(u_multiplier_B [29]),
    .A2(u_multiplier_A [29]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla2__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__46_  (.A1(u_multiplier_B [29]),
    .A2(u_multiplier_A [29]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla2__30_ ));
 XOR2_X2 u_multiplier_Final_add_cla1_cla2_cla2_cla2__47_  (.A(u_multiplier_B [29]),
    .B(u_multiplier_A [29]),
    .Z(u_multiplier_Final_add_cla1_cla2_cla2_cla2__31_ ));
 XNOR2_X2 u_multiplier_Final_add_cla1_cla2_cla2_cla2__48_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla2__28_ ),
    .B(u_multiplier_Final_add_cla1_cla2_cla2_cla2__31_ ),
    .ZN(product[29]));
 OAI21_X2 u_multiplier_Final_add_cla1_cla2_cla2_cla2__49_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla2__30_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla2_cla2__29_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla2_cla2__28_ ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla2__32_ ));
 AND2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__50_  (.A1(u_multiplier_B [30]),
    .A2(u_multiplier_A [30]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla2__33_ ));
 OR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__51_  (.A1(u_multiplier_B [30]),
    .A2(u_multiplier_A [30]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla2__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__52_  (.A(u_multiplier_B [30]),
    .B(u_multiplier_A [30]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla2__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__53_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla2__32_ ),
    .B(u_multiplier_Final_add_cla1_cla2_cla2_cla2__35_ ),
    .ZN(product[30]));
 AOI21_X4 u_multiplier_Final_add_cla1_cla2_cla2_cla2__54_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla2__33_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla2_cla2__34_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla2_cla2__32_ ),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla2__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__55_  (.A1(u_multiplier_B [31]),
    .A2(u_multiplier_A [31]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla2__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__56_  (.A1(u_multiplier_B [31]),
    .A2(u_multiplier_A [31]),
    .ZN(u_multiplier_Final_add_cla1_cla2_cla2_cla2__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__57_  (.A(u_multiplier_B [31]),
    .B(u_multiplier_A [31]),
    .Z(u_multiplier_Final_add_cla1_cla2_cla2_cla2__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla1_cla2_cla2_cla2__58_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla2__36_ ),
    .B(u_multiplier_Final_add_cla1_cla2_cla2_cla2__39_ ),
    .ZN(product[31]));
 OAI21_X4 u_multiplier_Final_add_cla1_cla2_cla2_cla2__59_  (.A(u_multiplier_Final_add_cla1_cla2_cla2_cla2__38_ ),
    .B1(u_multiplier_Final_add_cla1_cla2_cla2_cla2__37_ ),
    .B2(u_multiplier_Final_add_cla1_cla2_cla2_cla2__36_ ),
    .ZN(u_multiplier_Final_add_c1 ));
 AND2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__40_  (.A1(u_multiplier_B [32]),
    .A2(u_multiplier_A [32]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla1__25_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__41_  (.A1(u_multiplier_B [32]),
    .A2(u_multiplier_A [32]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla1__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__42_  (.A(u_multiplier_B [32]),
    .B(u_multiplier_A [32]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla1__27_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__43_  (.A(u_multiplier_Final_add_c1 ),
    .B(u_multiplier_Final_add_cla2_cla1_cla1_cla1__27_ ),
    .ZN(product[32]));
 AOI21_X4 u_multiplier_Final_add_cla2_cla1_cla1_cla1__44_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla1__25_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla1_cla1__26_ ),
    .B2(u_multiplier_Final_add_c1 ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla1__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__45_  (.A1(u_multiplier_B [33]),
    .A2(u_multiplier_A [33]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla1__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__46_  (.A1(u_multiplier_B [33]),
    .A2(u_multiplier_A [33]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla1__30_ ));
 XOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__47_  (.A(u_multiplier_B [33]),
    .B(u_multiplier_A [33]),
    .Z(u_multiplier_Final_add_cla2_cla1_cla1_cla1__31_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__48_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla1__28_ ),
    .B(u_multiplier_Final_add_cla2_cla1_cla1_cla1__31_ ),
    .ZN(product[33]));
 OAI21_X2 u_multiplier_Final_add_cla2_cla1_cla1_cla1__49_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla1__30_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla1_cla1__29_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla1_cla1__28_ ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla1__32_ ));
 AND2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__50_  (.A1(u_multiplier_B [34]),
    .A2(u_multiplier_A [34]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla1__33_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__51_  (.A1(u_multiplier_B [34]),
    .A2(u_multiplier_A [34]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla1__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__52_  (.A(u_multiplier_B [34]),
    .B(u_multiplier_A [34]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla1__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__53_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla1__32_ ),
    .B(u_multiplier_Final_add_cla2_cla1_cla1_cla1__35_ ),
    .ZN(product[34]));
 AOI21_X4 u_multiplier_Final_add_cla2_cla1_cla1_cla1__54_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla1__33_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla1_cla1__34_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla1_cla1__32_ ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla1__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__55_  (.A1(u_multiplier_B [35]),
    .A2(u_multiplier_A [35]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla1__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__56_  (.A1(u_multiplier_B [35]),
    .A2(u_multiplier_A [35]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla1__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__57_  (.A(u_multiplier_B [35]),
    .B(u_multiplier_A [35]),
    .Z(u_multiplier_Final_add_cla2_cla1_cla1_cla1__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla1__58_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla1__36_ ),
    .B(u_multiplier_Final_add_cla2_cla1_cla1_cla1__39_ ),
    .ZN(product[35]));
 OAI21_X4 u_multiplier_Final_add_cla2_cla1_cla1_cla1__59_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla1__38_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla1_cla1__37_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla1_cla1__36_ ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_c1 ));
 AND2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla2__40_  (.A1(u_multiplier_B [36]),
    .A2(u_multiplier_A [36]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla2__25_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla2__41_  (.A1(u_multiplier_B [36]),
    .A2(u_multiplier_A [36]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla2__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla2__42_  (.A(u_multiplier_B [36]),
    .B(u_multiplier_A [36]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla2__27_ ));
 XNOR2_X2 u_multiplier_Final_add_cla2_cla1_cla1_cla2__43_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_c1 ),
    .B(u_multiplier_Final_add_cla2_cla1_cla1_cla2__27_ ),
    .ZN(product[36]));
 AOI21_X4 u_multiplier_Final_add_cla2_cla1_cla1_cla2__44_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla2__25_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla1_cla2__26_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla1_c1 ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla2__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla2__45_  (.A1(u_multiplier_B [37]),
    .A2(u_multiplier_A [37]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla2__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla2__46_  (.A1(u_multiplier_B [37]),
    .A2(u_multiplier_A [37]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla2__30_ ));
 XOR2_X2 u_multiplier_Final_add_cla2_cla1_cla1_cla2__47_  (.A(u_multiplier_B [37]),
    .B(u_multiplier_A [37]),
    .Z(u_multiplier_Final_add_cla2_cla1_cla1_cla2__31_ ));
 XNOR2_X2 u_multiplier_Final_add_cla2_cla1_cla1_cla2__48_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla2__28_ ),
    .B(u_multiplier_Final_add_cla2_cla1_cla1_cla2__31_ ),
    .ZN(product[37]));
 OAI21_X2 u_multiplier_Final_add_cla2_cla1_cla1_cla2__49_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla2__30_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla1_cla2__29_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla1_cla2__28_ ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla2__32_ ));
 AND2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla2__50_  (.A1(u_multiplier_B [38]),
    .A2(u_multiplier_A [38]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla2__33_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla2__51_  (.A1(u_multiplier_B [38]),
    .A2(u_multiplier_A [38]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla2__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla2__52_  (.A(u_multiplier_B [38]),
    .B(u_multiplier_A [38]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla2__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla2__53_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla2__32_ ),
    .B(u_multiplier_Final_add_cla2_cla1_cla1_cla2__35_ ),
    .ZN(product[38]));
 AOI21_X4 u_multiplier_Final_add_cla2_cla1_cla1_cla2__54_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla2__33_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla1_cla2__34_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla1_cla2__32_ ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla2__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla2__55_  (.A1(u_multiplier_B [39]),
    .A2(u_multiplier_A [39]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla2__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla1_cla1_cla2__56_  (.A1(u_multiplier_B [39]),
    .A2(u_multiplier_A [39]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla1_cla2__38_ ));
 XOR2_X2 u_multiplier_Final_add_cla2_cla1_cla1_cla2__57_  (.A(u_multiplier_B [39]),
    .B(u_multiplier_A [39]),
    .Z(u_multiplier_Final_add_cla2_cla1_cla1_cla2__39_ ));
 XNOR2_X2 u_multiplier_Final_add_cla2_cla1_cla1_cla2__58_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla2__36_ ),
    .B(u_multiplier_Final_add_cla2_cla1_cla1_cla2__39_ ),
    .ZN(product[39]));
 OAI21_X2 u_multiplier_Final_add_cla2_cla1_cla1_cla2__59_  (.A(u_multiplier_Final_add_cla2_cla1_cla1_cla2__38_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla1_cla2__37_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla1_cla2__36_ ),
    .ZN(u_multiplier_Final_add_cla2_cla1_c1 ));
 AND2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__40_  (.A1(u_multiplier_B [40]),
    .A2(u_multiplier_A [40]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla1__25_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__41_  (.A1(u_multiplier_B [40]),
    .A2(u_multiplier_A [40]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla1__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__42_  (.A(u_multiplier_B [40]),
    .B(u_multiplier_A [40]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla1__27_ ));
 XNOR2_X2 u_multiplier_Final_add_cla2_cla1_cla2_cla1__43_  (.A(u_multiplier_Final_add_cla2_cla1_c1 ),
    .B(u_multiplier_Final_add_cla2_cla1_cla2_cla1__27_ ),
    .ZN(product[40]));
 AOI21_X2 u_multiplier_Final_add_cla2_cla1_cla2_cla1__44_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla1__25_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla2_cla1__26_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_c1 ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla1__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__45_  (.A1(u_multiplier_B [41]),
    .A2(u_multiplier_A [41]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla1__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__46_  (.A1(u_multiplier_B [41]),
    .A2(u_multiplier_A [41]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla1__30_ ));
 XOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__47_  (.A(u_multiplier_B [41]),
    .B(u_multiplier_A [41]),
    .Z(u_multiplier_Final_add_cla2_cla1_cla2_cla1__31_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__48_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla1__28_ ),
    .B(u_multiplier_Final_add_cla2_cla1_cla2_cla1__31_ ),
    .ZN(product[41]));
 OAI21_X2 u_multiplier_Final_add_cla2_cla1_cla2_cla1__49_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla1__30_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla2_cla1__29_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla2_cla1__28_ ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla1__32_ ));
 AND2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__50_  (.A1(u_multiplier_B [42]),
    .A2(u_multiplier_A [42]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla1__33_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__51_  (.A1(u_multiplier_B [42]),
    .A2(u_multiplier_A [42]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla1__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__52_  (.A(u_multiplier_B [42]),
    .B(u_multiplier_A [42]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla1__35_ ));
 XNOR2_X2 u_multiplier_Final_add_cla2_cla1_cla2_cla1__53_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla1__32_ ),
    .B(u_multiplier_Final_add_cla2_cla1_cla2_cla1__35_ ),
    .ZN(product[42]));
 AOI21_X4 u_multiplier_Final_add_cla2_cla1_cla2_cla1__54_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla1__33_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla2_cla1__34_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla2_cla1__32_ ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla1__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__55_  (.A1(u_multiplier_B [43]),
    .A2(u_multiplier_A [43]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla1__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__56_  (.A1(u_multiplier_B [43]),
    .A2(u_multiplier_A [43]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla1__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__57_  (.A(u_multiplier_B [43]),
    .B(u_multiplier_A [43]),
    .Z(u_multiplier_Final_add_cla2_cla1_cla2_cla1__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla1__58_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla1__36_ ),
    .B(u_multiplier_Final_add_cla2_cla1_cla2_cla1__39_ ),
    .ZN(product[43]));
 OAI21_X2 u_multiplier_Final_add_cla2_cla1_cla2_cla1__59_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla1__38_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla2_cla1__37_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla2_cla1__36_ ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_c1 ));
 AND2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__40_  (.A1(u_multiplier_B [44]),
    .A2(u_multiplier_A [44]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla2__25_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__41_  (.A1(u_multiplier_B [44]),
    .A2(u_multiplier_A [44]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla2__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__42_  (.A(u_multiplier_B [44]),
    .B(u_multiplier_A [44]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla2__27_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__43_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_c1 ),
    .B(u_multiplier_Final_add_cla2_cla1_cla2_cla2__27_ ),
    .ZN(product[44]));
 AOI21_X2 u_multiplier_Final_add_cla2_cla1_cla2_cla2__44_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla2__25_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla2_cla2__26_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla2_c1 ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla2__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__45_  (.A1(u_multiplier_B [45]),
    .A2(u_multiplier_A [45]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla2__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__46_  (.A1(u_multiplier_B [45]),
    .A2(u_multiplier_A [45]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla2__30_ ));
 XOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__47_  (.A(u_multiplier_B [45]),
    .B(u_multiplier_A [45]),
    .Z(u_multiplier_Final_add_cla2_cla1_cla2_cla2__31_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__48_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla2__28_ ),
    .B(u_multiplier_Final_add_cla2_cla1_cla2_cla2__31_ ),
    .ZN(product[45]));
 OAI21_X2 u_multiplier_Final_add_cla2_cla1_cla2_cla2__49_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla2__30_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla2_cla2__29_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla2_cla2__28_ ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla2__32_ ));
 AND2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__50_  (.A1(u_multiplier_B [46]),
    .A2(u_multiplier_A [46]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla2__33_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__51_  (.A1(u_multiplier_B [46]),
    .A2(u_multiplier_A [46]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla2__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__52_  (.A(u_multiplier_B [46]),
    .B(u_multiplier_A [46]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla2__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__53_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla2__32_ ),
    .B(u_multiplier_Final_add_cla2_cla1_cla2_cla2__35_ ),
    .ZN(product[46]));
 AOI21_X2 u_multiplier_Final_add_cla2_cla1_cla2_cla2__54_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla2__33_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla2_cla2__34_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla2_cla2__32_ ),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla2__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__55_  (.A1(u_multiplier_B [47]),
    .A2(u_multiplier_A [47]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla2__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__56_  (.A1(u_multiplier_B [47]),
    .A2(u_multiplier_A [47]),
    .ZN(u_multiplier_Final_add_cla2_cla1_cla2_cla2__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__57_  (.A(u_multiplier_B [47]),
    .B(u_multiplier_A [47]),
    .Z(u_multiplier_Final_add_cla2_cla1_cla2_cla2__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla1_cla2_cla2__58_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla2__36_ ),
    .B(u_multiplier_Final_add_cla2_cla1_cla2_cla2__39_ ),
    .ZN(product[47]));
 OAI21_X2 u_multiplier_Final_add_cla2_cla1_cla2_cla2__59_  (.A(u_multiplier_Final_add_cla2_cla1_cla2_cla2__38_ ),
    .B1(u_multiplier_Final_add_cla2_cla1_cla2_cla2__37_ ),
    .B2(u_multiplier_Final_add_cla2_cla1_cla2_cla2__36_ ),
    .ZN(u_multiplier_Final_add_cla2_c1 ));
 AND2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__40_  (.A1(u_multiplier_B [48]),
    .A2(u_multiplier_A [48]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla1__25_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__41_  (.A1(u_multiplier_B [48]),
    .A2(u_multiplier_A [48]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla1__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__42_  (.A(u_multiplier_B [48]),
    .B(u_multiplier_A [48]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla1__27_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__43_  (.A(u_multiplier_Final_add_cla2_c1 ),
    .B(u_multiplier_Final_add_cla2_cla2_cla1_cla1__27_ ),
    .ZN(product[48]));
 AOI21_X2 u_multiplier_Final_add_cla2_cla2_cla1_cla1__44_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla1__25_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla1_cla1__26_ ),
    .B2(u_multiplier_Final_add_cla2_c1 ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla1__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__45_  (.A1(u_multiplier_B [49]),
    .A2(u_multiplier_A [49]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla1__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__46_  (.A1(u_multiplier_B [49]),
    .A2(u_multiplier_A [49]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla1__30_ ));
 XOR2_X2 u_multiplier_Final_add_cla2_cla2_cla1_cla1__47_  (.A(u_multiplier_B [49]),
    .B(u_multiplier_A [49]),
    .Z(u_multiplier_Final_add_cla2_cla2_cla1_cla1__31_ ));
 XNOR2_X2 u_multiplier_Final_add_cla2_cla2_cla1_cla1__48_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla1__28_ ),
    .B(u_multiplier_Final_add_cla2_cla2_cla1_cla1__31_ ),
    .ZN(product[49]));
 OAI21_X2 u_multiplier_Final_add_cla2_cla2_cla1_cla1__49_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla1__30_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla1_cla1__29_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla1_cla1__28_ ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla1__32_ ));
 AND2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__50_  (.A1(u_multiplier_B [50]),
    .A2(u_multiplier_A [50]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla1__33_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__51_  (.A1(u_multiplier_B [50]),
    .A2(u_multiplier_A [50]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla1__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__52_  (.A(u_multiplier_B [50]),
    .B(u_multiplier_A [50]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla1__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__53_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla1__32_ ),
    .B(u_multiplier_Final_add_cla2_cla2_cla1_cla1__35_ ),
    .ZN(product[50]));
 AOI21_X2 u_multiplier_Final_add_cla2_cla2_cla1_cla1__54_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla1__33_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla1_cla1__34_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla1_cla1__32_ ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla1__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__55_  (.A1(u_multiplier_B [51]),
    .A2(u_multiplier_A [51]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla1__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__56_  (.A1(u_multiplier_B [51]),
    .A2(u_multiplier_A [51]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla1__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__57_  (.A(u_multiplier_B [51]),
    .B(u_multiplier_A [51]),
    .Z(u_multiplier_Final_add_cla2_cla2_cla1_cla1__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla1__58_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla1__36_ ),
    .B(u_multiplier_Final_add_cla2_cla2_cla1_cla1__39_ ),
    .ZN(product[51]));
 OAI21_X2 u_multiplier_Final_add_cla2_cla2_cla1_cla1__59_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla1__38_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla1_cla1__37_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla1_cla1__36_ ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_c1 ));
 AND2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__40_  (.A1(u_multiplier_B [52]),
    .A2(u_multiplier_A [52]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla2__25_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__41_  (.A1(u_multiplier_B [52]),
    .A2(u_multiplier_A [52]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla2__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__42_  (.A(u_multiplier_B [52]),
    .B(u_multiplier_A [52]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla2__27_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__43_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_c1 ),
    .B(u_multiplier_Final_add_cla2_cla2_cla1_cla2__27_ ),
    .ZN(product[52]));
 AOI21_X4 u_multiplier_Final_add_cla2_cla2_cla1_cla2__44_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla2__25_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla1_cla2__26_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla1_c1 ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla2__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__45_  (.A1(u_multiplier_B [53]),
    .A2(u_multiplier_A [53]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla2__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__46_  (.A1(u_multiplier_B [53]),
    .A2(u_multiplier_A [53]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla2__30_ ));
 XOR2_X2 u_multiplier_Final_add_cla2_cla2_cla1_cla2__47_  (.A(u_multiplier_B [53]),
    .B(u_multiplier_A [53]),
    .Z(u_multiplier_Final_add_cla2_cla2_cla1_cla2__31_ ));
 XNOR2_X2 u_multiplier_Final_add_cla2_cla2_cla1_cla2__48_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla2__28_ ),
    .B(u_multiplier_Final_add_cla2_cla2_cla1_cla2__31_ ),
    .ZN(product[53]));
 OAI21_X2 u_multiplier_Final_add_cla2_cla2_cla1_cla2__49_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla2__30_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla1_cla2__29_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla1_cla2__28_ ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla2__32_ ));
 AND2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__50_  (.A1(u_multiplier_B [54]),
    .A2(u_multiplier_A [54]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla2__33_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__51_  (.A1(u_multiplier_B [54]),
    .A2(u_multiplier_A [54]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla2__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__52_  (.A(u_multiplier_B [54]),
    .B(u_multiplier_A [54]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla2__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__53_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla2__32_ ),
    .B(u_multiplier_Final_add_cla2_cla2_cla1_cla2__35_ ),
    .ZN(product[54]));
 AOI21_X4 u_multiplier_Final_add_cla2_cla2_cla1_cla2__54_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla2__33_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla1_cla2__34_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla1_cla2__32_ ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla2__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__55_  (.A1(u_multiplier_B [55]),
    .A2(u_multiplier_A [55]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla2__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__56_  (.A1(u_multiplier_B [55]),
    .A2(u_multiplier_A [55]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla1_cla2__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__57_  (.A(u_multiplier_B [55]),
    .B(u_multiplier_A [55]),
    .Z(u_multiplier_Final_add_cla2_cla2_cla1_cla2__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla1_cla2__58_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla2__36_ ),
    .B(u_multiplier_Final_add_cla2_cla2_cla1_cla2__39_ ),
    .ZN(product[55]));
 OAI21_X4 u_multiplier_Final_add_cla2_cla2_cla1_cla2__59_  (.A(u_multiplier_Final_add_cla2_cla2_cla1_cla2__38_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla1_cla2__37_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla1_cla2__36_ ),
    .ZN(u_multiplier_Final_add_cla2_cla2_c1 ));
 AND2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__40_  (.A1(u_multiplier_B [56]),
    .A2(u_multiplier_A [56]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla1__25_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__41_  (.A1(u_multiplier_B [56]),
    .A2(u_multiplier_A [56]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla1__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__42_  (.A(u_multiplier_B [56]),
    .B(u_multiplier_A [56]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla1__27_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__43_  (.A(u_multiplier_Final_add_cla2_cla2_c1 ),
    .B(u_multiplier_Final_add_cla2_cla2_cla2_cla1__27_ ),
    .ZN(product[56]));
 AOI21_X2 u_multiplier_Final_add_cla2_cla2_cla2_cla1__44_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla1__25_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla2_cla1__26_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_c1 ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla1__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__45_  (.A1(u_multiplier_B [57]),
    .A2(u_multiplier_A [57]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla1__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__46_  (.A1(u_multiplier_B [57]),
    .A2(u_multiplier_A [57]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla1__30_ ));
 XOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__47_  (.A(u_multiplier_B [57]),
    .B(u_multiplier_A [57]),
    .Z(u_multiplier_Final_add_cla2_cla2_cla2_cla1__31_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__48_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla1__28_ ),
    .B(u_multiplier_Final_add_cla2_cla2_cla2_cla1__31_ ),
    .ZN(product[57]));
 OAI21_X2 u_multiplier_Final_add_cla2_cla2_cla2_cla1__49_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla1__30_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla2_cla1__29_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla2_cla1__28_ ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla1__32_ ));
 AND2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__50_  (.A1(u_multiplier_B [58]),
    .A2(u_multiplier_A [58]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla1__33_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__51_  (.A1(u_multiplier_B [58]),
    .A2(u_multiplier_A [58]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla1__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__52_  (.A(u_multiplier_B [58]),
    .B(u_multiplier_A [58]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla1__35_ ));
 XNOR2_X2 u_multiplier_Final_add_cla2_cla2_cla2_cla1__53_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla1__32_ ),
    .B(u_multiplier_Final_add_cla2_cla2_cla2_cla1__35_ ),
    .ZN(product[58]));
 AOI21_X2 u_multiplier_Final_add_cla2_cla2_cla2_cla1__54_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla1__33_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla2_cla1__34_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla2_cla1__32_ ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla1__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__55_  (.A1(u_multiplier_B [59]),
    .A2(u_multiplier_A [59]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla1__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__56_  (.A1(u_multiplier_B [59]),
    .A2(u_multiplier_A [59]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla1__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__57_  (.A(u_multiplier_B [59]),
    .B(u_multiplier_A [59]),
    .Z(u_multiplier_Final_add_cla2_cla2_cla2_cla1__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla1__58_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla1__36_ ),
    .B(u_multiplier_Final_add_cla2_cla2_cla2_cla1__39_ ),
    .ZN(product[59]));
 OAI21_X2 u_multiplier_Final_add_cla2_cla2_cla2_cla1__59_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla1__38_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla2_cla1__37_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla2_cla1__36_ ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_c1 ));
 AND2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__40_  (.A1(u_multiplier_B [60]),
    .A2(u_multiplier_A [60]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla2__25_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__41_  (.A1(u_multiplier_B [60]),
    .A2(u_multiplier_A [60]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla2__26_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__42_  (.A(u_multiplier_B [60]),
    .B(u_multiplier_A [60]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla2__27_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__43_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_c1 ),
    .B(u_multiplier_Final_add_cla2_cla2_cla2_cla2__27_ ),
    .ZN(product[60]));
 AOI21_X2 u_multiplier_Final_add_cla2_cla2_cla2_cla2__44_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla2__25_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla2_cla2__26_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla2_c1 ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla2__28_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__45_  (.A1(u_multiplier_B [61]),
    .A2(u_multiplier_A [61]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla2__29_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__46_  (.A1(u_multiplier_B [61]),
    .A2(u_multiplier_A [61]),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla2__30_ ));
 XOR2_X2 u_multiplier_Final_add_cla2_cla2_cla2_cla2__47_  (.A(u_multiplier_B [61]),
    .B(u_multiplier_A [61]),
    .Z(u_multiplier_Final_add_cla2_cla2_cla2_cla2__31_ ));
 XNOR2_X2 u_multiplier_Final_add_cla2_cla2_cla2_cla2__48_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla2__28_ ),
    .B(u_multiplier_Final_add_cla2_cla2_cla2_cla2__31_ ),
    .ZN(product[61]));
 OAI21_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__49_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla2__30_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla2_cla2__29_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla2_cla2__28_ ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla2__32_ ));
 AND2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__50_  (.A1(u_multiplier_B [62]),
    .A2(u_multiplier_pp3_62 ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla2__33_ ));
 OR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__51_  (.A1(u_multiplier_B [62]),
    .A2(u_multiplier_pp3_62 ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla2__34_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__52_  (.A(u_multiplier_B [62]),
    .B(u_multiplier_pp3_62 ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla2__35_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__53_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla2__32_ ),
    .B(u_multiplier_Final_add_cla2_cla2_cla2_cla2__35_ ),
    .ZN(product[62]));
 AOI21_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__54_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla2__33_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla2_cla2__34_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla2_cla2__32_ ),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla2__36_ ));
 NOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__55_  (.A1(net144),
    .A2(net145),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla2__37_ ));
 NAND2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__56_  (.A1(net146),
    .A2(net147),
    .ZN(u_multiplier_Final_add_cla2_cla2_cla2_cla2__38_ ));
 XOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__57_  (.A(net148),
    .B(net149),
    .Z(u_multiplier_Final_add_cla2_cla2_cla2_cla2__39_ ));
 XNOR2_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__58_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla2__36_ ),
    .B(u_multiplier_Final_add_cla2_cla2_cla2_cla2__39_ ),
    .ZN(product[63]));
 OAI21_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__59_  (.A(u_multiplier_Final_add_cla2_cla2_cla2_cla2__38_ ),
    .B1(u_multiplier_Final_add_cla2_cla2_cla2_cla2__37_ ),
    .B2(u_multiplier_Final_add_cla2_cla2_cla2_cla2__36_ ),
    .ZN(u_multiplier_Final_add_Cout ));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_32_1__18_  (.A(net111),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_1__19_  (.A1(u_multiplier_STAGE1__0880_ ),
    .A2(u_multiplier_STAGE1__0879_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_1__20_  (.A(u_multiplier_STAGE1__0880_ ),
    .B(u_multiplier_STAGE1__0879_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_1__21_  (.A1(u_multiplier_STAGE1__0881_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_1__22_  (.A(u_multiplier_STAGE1__0881_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_1__23_  (.A1(u_multiplier_STAGE1__0882_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_1__24_  (.A(u_multiplier_STAGE1__0882_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_1__25_  (.A(net112),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_1__16_ ),
    .ZN(u_multiplier_pp1_32 [7]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_32_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_32_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_32_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_32_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_32_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_32_1__17_ ),
    .ZN(u_multiplier_pp1_33 [15]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_32_2__18_  (.A(net113),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_2__19_  (.A1(u_multiplier_STAGE1__0884_ ),
    .A2(u_multiplier_STAGE1__0883_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_2__20_  (.A(u_multiplier_STAGE1__0884_ ),
    .B(u_multiplier_STAGE1__0883_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_2__21_  (.A1(u_multiplier_STAGE1__0885_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_2__22_  (.A(u_multiplier_STAGE1__0885_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_2__23_  (.A1(u_multiplier_STAGE1__0886_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_2__24_  (.A(u_multiplier_STAGE1__0886_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_2__25_  (.A(net114),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_2__16_ ),
    .ZN(u_multiplier_pp1_32 [6]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_32_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_32_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_32_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_32_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_32_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_32_2__17_ ),
    .ZN(u_multiplier_pp1_33 [14]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_32_3__18_  (.A(net115),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_3__19_  (.A1(u_multiplier_STAGE1__0888_ ),
    .A2(u_multiplier_STAGE1__0887_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_3__20_  (.A(u_multiplier_STAGE1__0888_ ),
    .B(u_multiplier_STAGE1__0887_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_3__21_  (.A1(u_multiplier_STAGE1__0889_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_3__22_  (.A(u_multiplier_STAGE1__0889_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_3__23_  (.A1(u_multiplier_STAGE1__0890_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_3__24_  (.A(u_multiplier_STAGE1__0890_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_3__25_  (.A(net116),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_3__16_ ),
    .ZN(u_multiplier_pp1_32 [5]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_32_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_32_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_32_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_32_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_32_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_32_3__17_ ),
    .ZN(u_multiplier_pp1_33 [13]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_32_4__18_  (.A(net117),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_4__19_  (.A1(u_multiplier_STAGE1__0892_ ),
    .A2(u_multiplier_STAGE1__0891_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_4__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_4__20_  (.A(u_multiplier_STAGE1__0892_ ),
    .B(u_multiplier_STAGE1__0891_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_4__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_4__21_  (.A1(u_multiplier_STAGE1__0893_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_4__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_4__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_4__22_  (.A(u_multiplier_STAGE1__0893_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_4__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_4__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_4__23_  (.A1(u_multiplier_STAGE1__0894_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_4__24_  (.A(u_multiplier_STAGE1__0894_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_4__25_  (.A(net118),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_4__16_ ),
    .ZN(u_multiplier_pp1_32 [4]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_4__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_32_4__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_4__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_32_4_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_32_4__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_32_4__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_32_4__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_32_4__17_ ),
    .ZN(u_multiplier_pp1_33 [12]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_32_5__18_  (.A(net119),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_5__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_5__19_  (.A1(u_multiplier_STAGE1__0896_ ),
    .A2(u_multiplier_STAGE1__0895_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_5__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_5__20_  (.A(u_multiplier_STAGE1__0896_ ),
    .B(u_multiplier_STAGE1__0895_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_5__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_5__21_  (.A1(u_multiplier_STAGE1__0897_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_5__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_5__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_5__22_  (.A(u_multiplier_STAGE1__0897_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_5__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_5__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_5__23_  (.A1(u_multiplier_STAGE1__0898_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_5__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_5__24_  (.A(u_multiplier_STAGE1__0898_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_5__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_5__25_  (.A(net120),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_5__16_ ),
    .ZN(u_multiplier_pp1_32 [3]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_5__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_32_5__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_5__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_32_5_cout ));
 OAI21_X1 u_multiplier_STAGE1_E_4_2_pp_32_5__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_32_5__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_32_5__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_32_5__17_ ),
    .ZN(u_multiplier_pp1_33 [11]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_32_6__18_  (.A(net121),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_6__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_6__19_  (.A1(u_multiplier_STAGE1__0900_ ),
    .A2(u_multiplier_STAGE1__0899_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_6__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_6__20_  (.A(u_multiplier_STAGE1__0900_ ),
    .B(u_multiplier_STAGE1__0899_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_6__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_6__21_  (.A1(u_multiplier_STAGE1__0901_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_6__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_6__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_6__22_  (.A(u_multiplier_STAGE1__0901_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_6__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_6__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_6__23_  (.A1(u_multiplier_STAGE1__0902_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_6__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_6__24_  (.A(u_multiplier_STAGE1__0902_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_6__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_6__25_  (.A(net122),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_6__16_ ),
    .ZN(u_multiplier_pp1_32 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_6__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_32_6__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_6__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_32_6_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_32_6__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_32_6__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_32_6__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_32_6__17_ ),
    .ZN(u_multiplier_pp1_33 [10]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_32_7__18_  (.A(net123),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_7__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_7__19_  (.A1(u_multiplier_STAGE1__0904_ ),
    .A2(u_multiplier_STAGE1__0903_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_7__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_7__20_  (.A(u_multiplier_STAGE1__0904_ ),
    .B(u_multiplier_STAGE1__0903_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_7__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_7__21_  (.A1(u_multiplier_STAGE1__0905_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_7__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_7__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_7__22_  (.A(u_multiplier_STAGE1__0905_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_7__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_32_7__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_7__23_  (.A1(u_multiplier_STAGE1__0906_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_7__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_7__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_7__24_  (.A(u_multiplier_STAGE1__0906_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_7__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_32_7__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_32_7__25_  (.A(net124),
    .B(u_multiplier_STAGE1_E_4_2_pp_32_7__16_ ),
    .ZN(u_multiplier_pp1_32 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_32_7__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_32_7__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_32_7__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_32_7_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_32_7__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_32_7__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_32_7__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_32_7__17_ ),
    .ZN(u_multiplier_pp1_33 [9]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_33_1__18_  (.A(u_multiplier_STAGE1_pp1_32_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_1__19_  (.A1(u_multiplier_STAGE1__0911_ ),
    .A2(u_multiplier_STAGE1__0910_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_1__20_  (.A(u_multiplier_STAGE1__0911_ ),
    .B(u_multiplier_STAGE1__0910_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_1__21_  (.A1(u_multiplier_STAGE1__0912_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_1__22_  (.A(u_multiplier_STAGE1__0912_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_1__23_  (.A1(u_multiplier_STAGE1__0913_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_1__24_  (.A(u_multiplier_STAGE1__0913_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_1__25_  (.A(u_multiplier_STAGE1_pp1_32_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_1__16_ ),
    .ZN(u_multiplier_pp1_33 [7]));
 NAND2_X2 u_multiplier_STAGE1_E_4_2_pp_33_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_33_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_33_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_33_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_33_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_33_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_33_1__17_ ),
    .ZN(u_multiplier_pp1_34 [14]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_33_2__18_  (.A(u_multiplier_STAGE1_pp1_32_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_2__19_  (.A1(u_multiplier_STAGE1__0915_ ),
    .A2(u_multiplier_STAGE1__0914_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_2__20_  (.A(u_multiplier_STAGE1__0915_ ),
    .B(u_multiplier_STAGE1__0914_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_2__21_  (.A1(u_multiplier_STAGE1__0916_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_2__22_  (.A(u_multiplier_STAGE1__0916_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_2__23_  (.A1(u_multiplier_STAGE1__0917_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_2__24_  (.A(u_multiplier_STAGE1__0917_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_2__25_  (.A(u_multiplier_STAGE1_pp1_32_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_2__16_ ),
    .ZN(u_multiplier_pp1_33 [6]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_33_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_33_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_33_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_33_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_33_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_33_2__17_ ),
    .ZN(u_multiplier_pp1_34 [13]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_33_3__18_  (.A(u_multiplier_STAGE1_pp1_32_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_3__19_  (.A1(u_multiplier_STAGE1__0919_ ),
    .A2(u_multiplier_STAGE1__0918_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_3__20_  (.A(u_multiplier_STAGE1__0919_ ),
    .B(u_multiplier_STAGE1__0918_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_3__21_  (.A1(u_multiplier_STAGE1__0920_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_3__22_  (.A(u_multiplier_STAGE1__0920_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_3__23_  (.A1(u_multiplier_STAGE1__0921_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_3__24_  (.A(u_multiplier_STAGE1__0921_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_3__25_  (.A(u_multiplier_STAGE1_pp1_32_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_3__16_ ),
    .ZN(u_multiplier_pp1_33 [5]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_33_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_33_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_33_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_33_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_33_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_33_3__17_ ),
    .ZN(u_multiplier_pp1_34 [12]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_33_4__18_  (.A(u_multiplier_STAGE1_pp1_32_4_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_4__19_  (.A1(u_multiplier_STAGE1__0923_ ),
    .A2(u_multiplier_STAGE1__0922_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_4__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_4__20_  (.A(u_multiplier_STAGE1__0923_ ),
    .B(u_multiplier_STAGE1__0922_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_4__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_4__21_  (.A1(u_multiplier_STAGE1__0924_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_4__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_4__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_4__22_  (.A(u_multiplier_STAGE1__0924_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_4__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_4__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_4__23_  (.A1(u_multiplier_STAGE1__0925_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_4__24_  (.A(u_multiplier_STAGE1__0925_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_4__25_  (.A(u_multiplier_STAGE1_pp1_32_4_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_4__16_ ),
    .ZN(u_multiplier_pp1_33 [4]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_4__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_33_4__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_4__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_33_4_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_33_4__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_33_4__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_33_4__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_33_4__17_ ),
    .ZN(u_multiplier_pp1_34 [11]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_33_5__18_  (.A(u_multiplier_STAGE1_pp1_32_5_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_5__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_5__19_  (.A1(u_multiplier_STAGE1__0927_ ),
    .A2(u_multiplier_STAGE1__0926_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_5__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_5__20_  (.A(u_multiplier_STAGE1__0927_ ),
    .B(u_multiplier_STAGE1__0926_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_5__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_5__21_  (.A1(u_multiplier_STAGE1__0928_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_5__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_5__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_5__22_  (.A(u_multiplier_STAGE1__0928_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_5__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_5__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_5__23_  (.A1(u_multiplier_STAGE1__0929_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_5__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_5__24_  (.A(u_multiplier_STAGE1__0929_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_5__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_5__25_  (.A(u_multiplier_STAGE1_pp1_32_5_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_5__16_ ),
    .ZN(u_multiplier_pp1_33 [3]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_5__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_33_5__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_5__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_33_5_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_33_5__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_33_5__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_33_5__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_33_5__17_ ),
    .ZN(u_multiplier_pp1_34 [10]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_33_6__18_  (.A(u_multiplier_STAGE1_pp1_32_6_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_6__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_6__19_  (.A1(u_multiplier_STAGE1__0931_ ),
    .A2(u_multiplier_STAGE1__0930_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_6__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_6__20_  (.A(u_multiplier_STAGE1__0931_ ),
    .B(u_multiplier_STAGE1__0930_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_6__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_6__21_  (.A1(u_multiplier_STAGE1__0932_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_6__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_6__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_6__22_  (.A(u_multiplier_STAGE1__0932_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_6__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_6__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_6__23_  (.A1(u_multiplier_STAGE1__0933_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_6__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_6__24_  (.A(u_multiplier_STAGE1__0933_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_6__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_6__25_  (.A(u_multiplier_STAGE1_pp1_32_6_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_6__16_ ),
    .ZN(u_multiplier_pp1_33 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_6__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_33_6__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_6__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_33_6_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_33_6__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_33_6__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_33_6__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_33_6__17_ ),
    .ZN(u_multiplier_pp1_34 [9]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_33_7__18_  (.A(u_multiplier_STAGE1_pp1_32_7_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_7__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_7__19_  (.A1(u_multiplier_STAGE1__0935_ ),
    .A2(u_multiplier_STAGE1__0934_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_7__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_7__20_  (.A(u_multiplier_STAGE1__0935_ ),
    .B(u_multiplier_STAGE1__0934_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_7__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_7__21_  (.A1(u_multiplier_STAGE1__0936_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_7__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_7__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_7__22_  (.A(u_multiplier_STAGE1__0936_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_7__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_33_7__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_7__23_  (.A1(u_multiplier_STAGE1__0937_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_7__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_7__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_7__24_  (.A(u_multiplier_STAGE1__0937_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_7__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_33_7__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_33_7__25_  (.A(u_multiplier_STAGE1_pp1_32_7_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_33_7__16_ ),
    .ZN(u_multiplier_pp1_33 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_33_7__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_33_7__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_33_7__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_33_7_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_33_7__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_33_7__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_33_7__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_33_7__17_ ),
    .ZN(u_multiplier_pp1_34 [8]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_34_1__18_  (.A(u_multiplier_STAGE1_pp1_33_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_1__19_  (.A1(u_multiplier_STAGE1__0941_ ),
    .A2(u_multiplier_STAGE1__0940_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_1__20_  (.A(u_multiplier_STAGE1__0941_ ),
    .B(u_multiplier_STAGE1__0940_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_1__21_  (.A1(u_multiplier_STAGE1__0942_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_1__22_  (.A(u_multiplier_STAGE1__0942_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_1__23_  (.A1(u_multiplier_STAGE1__0943_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_1__24_  (.A(u_multiplier_STAGE1__0943_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_1__25_  (.A(u_multiplier_STAGE1_pp1_33_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_1__16_ ),
    .ZN(u_multiplier_pp1_34 [6]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_34_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_34_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_34_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_34_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_34_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_34_1__17_ ),
    .ZN(u_multiplier_pp1_35 [13]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_34_2__18_  (.A(u_multiplier_STAGE1_pp1_33_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_2__19_  (.A1(u_multiplier_STAGE1__0945_ ),
    .A2(u_multiplier_STAGE1__0944_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_2__20_  (.A(u_multiplier_STAGE1__0945_ ),
    .B(u_multiplier_STAGE1__0944_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_2__21_  (.A1(u_multiplier_STAGE1__0946_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_2__22_  (.A(u_multiplier_STAGE1__0946_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_2__23_  (.A1(u_multiplier_STAGE1__0947_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_2__24_  (.A(u_multiplier_STAGE1__0947_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_2__25_  (.A(u_multiplier_STAGE1_pp1_33_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_2__16_ ),
    .ZN(u_multiplier_pp1_34 [5]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_34_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_34_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_34_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_34_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_34_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_34_2__17_ ),
    .ZN(u_multiplier_pp1_35 [12]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_34_3__18_  (.A(u_multiplier_STAGE1_pp1_33_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_3__19_  (.A1(u_multiplier_STAGE1__0949_ ),
    .A2(u_multiplier_STAGE1__0948_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_3__20_  (.A(u_multiplier_STAGE1__0949_ ),
    .B(u_multiplier_STAGE1__0948_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_3__21_  (.A1(u_multiplier_STAGE1__0950_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_3__22_  (.A(u_multiplier_STAGE1__0950_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_3__23_  (.A1(u_multiplier_STAGE1__0951_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_3__24_  (.A(u_multiplier_STAGE1__0951_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_3__25_  (.A(u_multiplier_STAGE1_pp1_33_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_3__16_ ),
    .ZN(u_multiplier_pp1_34 [4]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_34_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_34_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_34_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_34_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_34_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_34_3__17_ ),
    .ZN(u_multiplier_pp1_35 [11]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_34_4__18_  (.A(u_multiplier_STAGE1_pp1_33_4_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_4__19_  (.A1(u_multiplier_STAGE1__0953_ ),
    .A2(u_multiplier_STAGE1__0952_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_4__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_4__20_  (.A(u_multiplier_STAGE1__0953_ ),
    .B(u_multiplier_STAGE1__0952_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_4__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_4__21_  (.A1(u_multiplier_STAGE1__0954_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_4__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_4__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_4__22_  (.A(u_multiplier_STAGE1__0954_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_4__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_4__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_4__23_  (.A1(u_multiplier_STAGE1__0955_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_4__24_  (.A(u_multiplier_STAGE1__0955_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_4__25_  (.A(u_multiplier_STAGE1_pp1_33_4_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_4__16_ ),
    .ZN(u_multiplier_pp1_34 [3]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_4__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_34_4__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_4__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_34_4_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_34_4__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_34_4__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_34_4__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_34_4__17_ ),
    .ZN(u_multiplier_pp1_35 [10]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_34_5__18_  (.A(u_multiplier_STAGE1_pp1_33_5_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_5__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_5__19_  (.A1(u_multiplier_STAGE1__0957_ ),
    .A2(u_multiplier_STAGE1__0956_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_5__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_5__20_  (.A(u_multiplier_STAGE1__0957_ ),
    .B(u_multiplier_STAGE1__0956_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_5__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_5__21_  (.A1(u_multiplier_STAGE1__0958_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_5__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_5__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_5__22_  (.A(u_multiplier_STAGE1__0958_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_5__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_5__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_5__23_  (.A1(u_multiplier_STAGE1__0959_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_5__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_5__24_  (.A(u_multiplier_STAGE1__0959_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_5__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_5__25_  (.A(u_multiplier_STAGE1_pp1_33_5_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_5__16_ ),
    .ZN(u_multiplier_pp1_34 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_5__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_34_5__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_5__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_34_5_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_34_5__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_34_5__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_34_5__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_34_5__17_ ),
    .ZN(u_multiplier_pp1_35 [9]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_34_6__18_  (.A(u_multiplier_STAGE1_pp1_33_6_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_6__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_6__19_  (.A1(u_multiplier_STAGE1__0961_ ),
    .A2(u_multiplier_STAGE1__0960_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_6__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_6__20_  (.A(u_multiplier_STAGE1__0961_ ),
    .B(u_multiplier_STAGE1__0960_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_6__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_6__21_  (.A1(u_multiplier_STAGE1__0962_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_6__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_6__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_6__22_  (.A(u_multiplier_STAGE1__0962_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_6__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_6__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_6__23_  (.A1(u_multiplier_STAGE1__0963_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_6__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_6__24_  (.A(u_multiplier_STAGE1__0963_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_6__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_6__25_  (.A(u_multiplier_STAGE1_pp1_33_6_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_6__16_ ),
    .ZN(u_multiplier_pp1_34 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_6__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_34_6__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_6__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_34_6_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_34_6__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_34_6__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_34_6__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_34_6__17_ ),
    .ZN(u_multiplier_pp1_35 [8]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_34_7__18_  (.A(u_multiplier_STAGE1_pp1_33_7_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_7__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_7__19_  (.A1(u_multiplier_STAGE1__0965_ ),
    .A2(u_multiplier_STAGE1__0964_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_7__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_7__20_  (.A(u_multiplier_STAGE1__0965_ ),
    .B(u_multiplier_STAGE1__0964_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_7__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_7__21_  (.A1(u_multiplier_STAGE1__0966_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_7__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_7__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_7__22_  (.A(u_multiplier_STAGE1__0966_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_7__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_34_7__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_34_7__23_  (.A1(u_multiplier_STAGE1__0967_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_7__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_7__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_7__24_  (.A(u_multiplier_STAGE1__0967_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_7__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_34_7__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_34_7__25_  (.A(u_multiplier_STAGE1_pp1_33_7_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_34_7__16_ ),
    .ZN(u_multiplier_pp1_34 [0]));
 NAND2_X2 u_multiplier_STAGE1_E_4_2_pp_34_7__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_34_7__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_34_7__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_34_7_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_34_7__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_34_7__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_34_7__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_34_7__17_ ),
    .ZN(u_multiplier_pp1_35 [7]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_35_1__18_  (.A(u_multiplier_STAGE1_pp1_34_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_1__19_  (.A1(u_multiplier_STAGE1__0969_ ),
    .A2(u_multiplier_STAGE1__0968_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_1__20_  (.A(u_multiplier_STAGE1__0969_ ),
    .B(u_multiplier_STAGE1__0968_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_35_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_1__21_  (.A1(u_multiplier_STAGE1__0970_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_1__22_  (.A(u_multiplier_STAGE1__0970_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_35_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_1__23_  (.A1(u_multiplier_STAGE1__0971_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_1__24_  (.A(u_multiplier_STAGE1__0971_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_1__25_  (.A(u_multiplier_STAGE1_pp1_34_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_1__16_ ),
    .ZN(u_multiplier_pp1_35 [6]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_35_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_35_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_35_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_35_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_35_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_35_1__17_ ),
    .ZN(u_multiplier_pp1_36 [12]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_35_2__18_  (.A(u_multiplier_STAGE1_pp1_34_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_2__19_  (.A1(u_multiplier_STAGE1__0973_ ),
    .A2(u_multiplier_STAGE1__0972_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_2__20_  (.A(u_multiplier_STAGE1__0973_ ),
    .B(u_multiplier_STAGE1__0972_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_35_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_2__21_  (.A1(u_multiplier_STAGE1__0974_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_2__22_  (.A(u_multiplier_STAGE1__0974_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_35_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_2__23_  (.A1(u_multiplier_STAGE1__0975_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_2__24_  (.A(u_multiplier_STAGE1__0975_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_2__25_  (.A(u_multiplier_STAGE1_pp1_34_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_2__16_ ),
    .ZN(u_multiplier_pp1_35 [5]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_35_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_35_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_35_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_35_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_35_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_35_2__17_ ),
    .ZN(u_multiplier_pp1_36 [11]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_35_3__18_  (.A(u_multiplier_STAGE1_pp1_34_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_3__19_  (.A1(u_multiplier_STAGE1__0977_ ),
    .A2(u_multiplier_STAGE1__0976_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_3__20_  (.A(u_multiplier_STAGE1__0977_ ),
    .B(u_multiplier_STAGE1__0976_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_35_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_3__21_  (.A1(u_multiplier_STAGE1__0978_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_3__22_  (.A(u_multiplier_STAGE1__0978_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_35_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_3__23_  (.A1(u_multiplier_STAGE1__0979_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_3__24_  (.A(u_multiplier_STAGE1__0979_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_3__25_  (.A(u_multiplier_STAGE1_pp1_34_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_3__16_ ),
    .ZN(u_multiplier_pp1_35 [4]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_35_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_35_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_35_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_35_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_35_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_35_3__17_ ),
    .ZN(u_multiplier_pp1_36 [10]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_35_4__18_  (.A(u_multiplier_STAGE1_pp1_34_4_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_4__19_  (.A1(u_multiplier_STAGE1__0981_ ),
    .A2(u_multiplier_STAGE1__0980_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_4__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_4__20_  (.A(u_multiplier_STAGE1__0981_ ),
    .B(u_multiplier_STAGE1__0980_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_35_4__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_4__21_  (.A1(u_multiplier_STAGE1__0982_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_4__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_4__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_4__22_  (.A(u_multiplier_STAGE1__0982_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_4__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_35_4__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_4__23_  (.A1(u_multiplier_STAGE1__0983_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_4__24_  (.A(u_multiplier_STAGE1__0983_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_4__25_  (.A(u_multiplier_STAGE1_pp1_34_4_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_4__16_ ),
    .ZN(u_multiplier_pp1_35 [3]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_4__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_35_4__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_4__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_35_4_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_35_4__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_35_4__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_35_4__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_35_4__17_ ),
    .ZN(u_multiplier_pp1_36 [9]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_35_5__18_  (.A(u_multiplier_STAGE1_pp1_34_5_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_5__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_5__19_  (.A1(u_multiplier_STAGE1__0985_ ),
    .A2(u_multiplier_STAGE1__0984_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_5__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_5__20_  (.A(u_multiplier_STAGE1__0985_ ),
    .B(u_multiplier_STAGE1__0984_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_35_5__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_5__21_  (.A1(u_multiplier_STAGE1__0986_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_5__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_5__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_5__22_  (.A(u_multiplier_STAGE1__0986_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_5__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_35_5__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_5__23_  (.A1(u_multiplier_STAGE1__0987_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_5__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_5__24_  (.A(u_multiplier_STAGE1__0987_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_5__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_5__25_  (.A(u_multiplier_STAGE1_pp1_34_5_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_5__16_ ),
    .ZN(u_multiplier_pp1_35 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_5__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_35_5__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_5__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_35_5_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_35_5__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_35_5__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_35_5__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_35_5__17_ ),
    .ZN(u_multiplier_pp1_36 [8]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_35_6__18_  (.A(u_multiplier_STAGE1_pp1_34_6_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_6__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_6__19_  (.A1(u_multiplier_STAGE1__0989_ ),
    .A2(u_multiplier_STAGE1__0988_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_6__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_6__20_  (.A(u_multiplier_STAGE1__0989_ ),
    .B(u_multiplier_STAGE1__0988_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_35_6__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_6__21_  (.A1(u_multiplier_STAGE1__0990_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_6__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_6__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_6__22_  (.A(u_multiplier_STAGE1__0990_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_6__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_35_6__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_6__23_  (.A1(u_multiplier_STAGE1__0991_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_6__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_6__24_  (.A(u_multiplier_STAGE1__0991_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_35_6__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_35_6__25_  (.A(u_multiplier_STAGE1_pp1_34_6_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_35_6__16_ ),
    .ZN(u_multiplier_pp1_35 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_35_6__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_35_6__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_35_6__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_35_6_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_35_6__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_35_6__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_35_6__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_35_6__17_ ),
    .ZN(u_multiplier_pp1_36 [7]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_36_1__18_  (.A(u_multiplier_STAGE1_pp1_35_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_1__19_  (.A1(u_multiplier_STAGE1__0995_ ),
    .A2(u_multiplier_STAGE1__0994_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_1__20_  (.A(u_multiplier_STAGE1__0995_ ),
    .B(u_multiplier_STAGE1__0994_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_36_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_1__21_  (.A1(u_multiplier_STAGE1__0996_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_1__22_  (.A(u_multiplier_STAGE1__0996_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_36_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_1__23_  (.A1(u_multiplier_STAGE1__0997_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_1__24_  (.A(u_multiplier_STAGE1__0997_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_1__25_  (.A(u_multiplier_STAGE1_pp1_35_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_1__16_ ),
    .ZN(u_multiplier_pp1_36 [5]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_36_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_36_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_36_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_36_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_36_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_36_1__17_ ),
    .ZN(u_multiplier_pp1_37 [11]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_36_2__18_  (.A(u_multiplier_STAGE1_pp1_35_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_2__19_  (.A1(u_multiplier_STAGE1__0999_ ),
    .A2(u_multiplier_STAGE1__0998_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_2__20_  (.A(u_multiplier_STAGE1__0999_ ),
    .B(u_multiplier_STAGE1__0998_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_36_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_2__21_  (.A1(u_multiplier_STAGE1__1000_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_2__22_  (.A(u_multiplier_STAGE1__1000_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_36_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_2__23_  (.A1(u_multiplier_STAGE1__1001_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_2__24_  (.A(u_multiplier_STAGE1__1001_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_2__25_  (.A(u_multiplier_STAGE1_pp1_35_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_2__16_ ),
    .ZN(u_multiplier_pp1_36 [4]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_36_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_36_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_36_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_36_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_36_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_36_2__17_ ),
    .ZN(u_multiplier_pp1_37 [10]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_36_3__18_  (.A(u_multiplier_STAGE1_pp1_35_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_3__19_  (.A1(u_multiplier_STAGE1__1003_ ),
    .A2(u_multiplier_STAGE1__1002_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_3__20_  (.A(u_multiplier_STAGE1__1003_ ),
    .B(u_multiplier_STAGE1__1002_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_36_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_3__21_  (.A1(u_multiplier_STAGE1__1004_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_3__22_  (.A(u_multiplier_STAGE1__1004_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_36_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_3__23_  (.A1(u_multiplier_STAGE1__1005_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_3__24_  (.A(u_multiplier_STAGE1__1005_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_3__25_  (.A(u_multiplier_STAGE1_pp1_35_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_3__16_ ),
    .ZN(u_multiplier_pp1_36 [3]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_36_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_36_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_36_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_36_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_36_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_36_3__17_ ),
    .ZN(u_multiplier_pp1_37 [9]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_36_4__18_  (.A(u_multiplier_STAGE1_pp1_35_4_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_4__19_  (.A1(u_multiplier_STAGE1__1007_ ),
    .A2(u_multiplier_STAGE1__1006_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_4__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_4__20_  (.A(u_multiplier_STAGE1__1007_ ),
    .B(u_multiplier_STAGE1__1006_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_36_4__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_4__21_  (.A1(u_multiplier_STAGE1__1008_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_4__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_4__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_4__22_  (.A(u_multiplier_STAGE1__1008_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_4__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_36_4__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_4__23_  (.A1(u_multiplier_STAGE1__1009_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_4__24_  (.A(u_multiplier_STAGE1__1009_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_4__25_  (.A(u_multiplier_STAGE1_pp1_35_4_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_4__16_ ),
    .ZN(u_multiplier_pp1_36 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_4__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_36_4__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_4__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_36_4_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_36_4__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_36_4__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_36_4__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_36_4__17_ ),
    .ZN(u_multiplier_pp1_37 [8]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_36_5__18_  (.A(u_multiplier_STAGE1_pp1_35_5_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_5__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_5__19_  (.A1(u_multiplier_STAGE1__1011_ ),
    .A2(u_multiplier_STAGE1__1010_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_5__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_5__20_  (.A(u_multiplier_STAGE1__1011_ ),
    .B(u_multiplier_STAGE1__1010_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_36_5__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_5__21_  (.A1(u_multiplier_STAGE1__1012_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_5__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_5__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_5__22_  (.A(u_multiplier_STAGE1__1012_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_5__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_36_5__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_5__23_  (.A1(u_multiplier_STAGE1__1013_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_5__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_5__24_  (.A(u_multiplier_STAGE1__1013_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_5__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_5__25_  (.A(u_multiplier_STAGE1_pp1_35_5_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_5__16_ ),
    .ZN(u_multiplier_pp1_36 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_5__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_36_5__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_5__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_36_5_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_36_5__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_36_5__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_36_5__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_36_5__17_ ),
    .ZN(u_multiplier_pp1_37 [7]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_36_6__18_  (.A(u_multiplier_STAGE1_pp1_35_6_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_6__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_6__19_  (.A1(u_multiplier_STAGE1__1015_ ),
    .A2(u_multiplier_STAGE1__1014_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_6__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_6__20_  (.A(u_multiplier_STAGE1__1015_ ),
    .B(u_multiplier_STAGE1__1014_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_36_6__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_6__21_  (.A1(u_multiplier_STAGE1__1016_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_6__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_6__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_6__22_  (.A(u_multiplier_STAGE1__1016_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_6__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_36_6__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_6__23_  (.A1(u_multiplier_STAGE1__1017_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_6__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_6__24_  (.A(u_multiplier_STAGE1__1017_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_6__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_36_6__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_36_6__25_  (.A(u_multiplier_STAGE1_pp1_35_6_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_36_6__16_ ),
    .ZN(u_multiplier_pp1_36 [0]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_36_6__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_36_6__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_36_6__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_36_6_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_36_6__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_36_6__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_36_6__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_36_6__17_ ),
    .ZN(u_multiplier_pp1_37 [6]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_37_1__18_  (.A(u_multiplier_STAGE1_pp1_36_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_1__19_  (.A1(u_multiplier_STAGE1__1019_ ),
    .A2(u_multiplier_STAGE1__1018_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_1__20_  (.A(u_multiplier_STAGE1__1019_ ),
    .B(u_multiplier_STAGE1__1018_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_37_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_1__21_  (.A1(u_multiplier_STAGE1__1020_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_1__22_  (.A(u_multiplier_STAGE1__1020_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_37_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_1__23_  (.A1(u_multiplier_STAGE1__1021_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_1__24_  (.A(u_multiplier_STAGE1__1021_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_1__25_  (.A(u_multiplier_STAGE1_pp1_36_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_1__16_ ),
    .ZN(u_multiplier_pp1_37 [5]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_37_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_37_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_37_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_37_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_37_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_37_1__17_ ),
    .ZN(u_multiplier_pp1_38 [10]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_37_2__18_  (.A(u_multiplier_STAGE1_pp1_36_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_2__19_  (.A1(u_multiplier_STAGE1__1023_ ),
    .A2(u_multiplier_STAGE1__1022_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_2__20_  (.A(u_multiplier_STAGE1__1023_ ),
    .B(u_multiplier_STAGE1__1022_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_37_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_2__21_  (.A1(u_multiplier_STAGE1__1024_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_2__22_  (.A(u_multiplier_STAGE1__1024_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_37_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_2__23_  (.A1(u_multiplier_STAGE1__1025_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_2__24_  (.A(u_multiplier_STAGE1__1025_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_2__25_  (.A(u_multiplier_STAGE1_pp1_36_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_2__16_ ),
    .ZN(u_multiplier_pp1_37 [4]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_37_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_37_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_37_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_37_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_37_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_37_2__17_ ),
    .ZN(u_multiplier_pp1_38 [9]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_37_3__18_  (.A(u_multiplier_STAGE1_pp1_36_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_3__19_  (.A1(u_multiplier_STAGE1__1027_ ),
    .A2(u_multiplier_STAGE1__1026_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_3__20_  (.A(u_multiplier_STAGE1__1027_ ),
    .B(u_multiplier_STAGE1__1026_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_37_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_3__21_  (.A1(u_multiplier_STAGE1__1028_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_3__22_  (.A(u_multiplier_STAGE1__1028_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_37_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_3__23_  (.A1(u_multiplier_STAGE1__1029_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_3__24_  (.A(u_multiplier_STAGE1__1029_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_3__25_  (.A(u_multiplier_STAGE1_pp1_36_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_3__16_ ),
    .ZN(u_multiplier_pp1_37 [3]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_37_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_37_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_37_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_37_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_37_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_37_3__17_ ),
    .ZN(u_multiplier_pp1_38 [8]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_37_4__18_  (.A(u_multiplier_STAGE1_pp1_36_4_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_4__19_  (.A1(u_multiplier_STAGE1__1031_ ),
    .A2(u_multiplier_STAGE1__1030_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_4__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_4__20_  (.A(u_multiplier_STAGE1__1031_ ),
    .B(u_multiplier_STAGE1__1030_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_37_4__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_4__21_  (.A1(u_multiplier_STAGE1__1032_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_4__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_4__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_4__22_  (.A(u_multiplier_STAGE1__1032_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_4__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_37_4__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_4__23_  (.A1(u_multiplier_STAGE1__1033_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_4__24_  (.A(u_multiplier_STAGE1__1033_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_4__25_  (.A(u_multiplier_STAGE1_pp1_36_4_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_4__16_ ),
    .ZN(u_multiplier_pp1_37 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_4__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_37_4__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_4__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_37_4_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_37_4__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_37_4__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_37_4__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_37_4__17_ ),
    .ZN(u_multiplier_pp1_38 [7]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_37_5__18_  (.A(u_multiplier_STAGE1_pp1_36_5_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_5__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_5__19_  (.A1(u_multiplier_STAGE1__1035_ ),
    .A2(u_multiplier_STAGE1__1034_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_5__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_5__20_  (.A(u_multiplier_STAGE1__1035_ ),
    .B(u_multiplier_STAGE1__1034_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_37_5__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_5__21_  (.A1(u_multiplier_STAGE1__1036_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_5__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_5__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_5__22_  (.A(u_multiplier_STAGE1__1036_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_5__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_37_5__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_5__23_  (.A1(u_multiplier_STAGE1__1037_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_5__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_5__24_  (.A(u_multiplier_STAGE1__1037_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_37_5__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_37_5__25_  (.A(u_multiplier_STAGE1_pp1_36_5_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_37_5__16_ ),
    .ZN(u_multiplier_pp1_37 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_37_5__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_37_5__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_37_5__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_37_5_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_37_5__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_37_5__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_37_5__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_37_5__17_ ),
    .ZN(u_multiplier_pp1_38 [6]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_38_1__18_  (.A(u_multiplier_STAGE1_pp1_37_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_1__19_  (.A1(u_multiplier_STAGE1__1041_ ),
    .A2(u_multiplier_STAGE1__1040_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_1__20_  (.A(u_multiplier_STAGE1__1041_ ),
    .B(u_multiplier_STAGE1__1040_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_38_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_1__21_  (.A1(u_multiplier_STAGE1__1042_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_1__22_  (.A(u_multiplier_STAGE1__1042_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_38_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_1__23_  (.A1(u_multiplier_STAGE1__1043_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_1__24_  (.A(u_multiplier_STAGE1__1043_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_1__25_  (.A(u_multiplier_STAGE1_pp1_37_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_1__16_ ),
    .ZN(u_multiplier_pp1_38 [4]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_38_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_38_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_38_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_38_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_38_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_38_1__17_ ),
    .ZN(u_multiplier_pp1_39 [9]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_38_2__18_  (.A(u_multiplier_STAGE1_pp1_37_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_2__19_  (.A1(u_multiplier_STAGE1__1045_ ),
    .A2(u_multiplier_STAGE1__1044_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_2__20_  (.A(u_multiplier_STAGE1__1045_ ),
    .B(u_multiplier_STAGE1__1044_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_38_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_2__21_  (.A1(u_multiplier_STAGE1__1046_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_2__22_  (.A(u_multiplier_STAGE1__1046_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_38_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_2__23_  (.A1(u_multiplier_STAGE1__1047_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_2__24_  (.A(u_multiplier_STAGE1__1047_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_2__25_  (.A(u_multiplier_STAGE1_pp1_37_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_2__16_ ),
    .ZN(u_multiplier_pp1_38 [3]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_38_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_38_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_38_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_38_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_38_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_38_2__17_ ),
    .ZN(u_multiplier_pp1_39 [8]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_38_3__18_  (.A(u_multiplier_STAGE1_pp1_37_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_3__19_  (.A1(u_multiplier_STAGE1__1049_ ),
    .A2(u_multiplier_STAGE1__1048_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_3__20_  (.A(u_multiplier_STAGE1__1049_ ),
    .B(u_multiplier_STAGE1__1048_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_38_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_3__21_  (.A1(u_multiplier_STAGE1__1050_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_3__22_  (.A(u_multiplier_STAGE1__1050_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_38_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_3__23_  (.A1(u_multiplier_STAGE1__1051_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_3__24_  (.A(u_multiplier_STAGE1__1051_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_3__25_  (.A(u_multiplier_STAGE1_pp1_37_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_3__16_ ),
    .ZN(u_multiplier_pp1_38 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_38_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_38_3_cout ));
 OAI21_X1 u_multiplier_STAGE1_E_4_2_pp_38_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_38_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_38_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_38_3__17_ ),
    .ZN(u_multiplier_pp1_39 [7]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_38_4__18_  (.A(u_multiplier_STAGE1_pp1_37_4_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_4__19_  (.A1(u_multiplier_STAGE1__1053_ ),
    .A2(u_multiplier_STAGE1__1052_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_4__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_4__20_  (.A(u_multiplier_STAGE1__1053_ ),
    .B(u_multiplier_STAGE1__1052_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_38_4__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_4__21_  (.A1(u_multiplier_STAGE1__1054_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_4__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_4__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_4__22_  (.A(u_multiplier_STAGE1__1054_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_4__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_38_4__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_4__23_  (.A1(u_multiplier_STAGE1__1055_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_4__24_  (.A(u_multiplier_STAGE1__1055_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_4__25_  (.A(u_multiplier_STAGE1_pp1_37_4_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_4__16_ ),
    .ZN(u_multiplier_pp1_38 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_4__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_38_4__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_4__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_38_4_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_38_4__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_38_4__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_38_4__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_38_4__17_ ),
    .ZN(u_multiplier_pp1_39 [6]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_38_5__18_  (.A(u_multiplier_STAGE1_pp1_37_5_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_5__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_5__19_  (.A1(u_multiplier_STAGE1__1057_ ),
    .A2(u_multiplier_STAGE1__1056_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_5__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_5__20_  (.A(u_multiplier_STAGE1__1057_ ),
    .B(u_multiplier_STAGE1__1056_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_38_5__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_5__21_  (.A1(u_multiplier_STAGE1__1058_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_5__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_5__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_5__22_  (.A(u_multiplier_STAGE1__1058_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_5__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_38_5__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_5__23_  (.A1(u_multiplier_STAGE1__1059_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_5__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_5__24_  (.A(u_multiplier_STAGE1__1059_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_5__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_38_5__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_38_5__25_  (.A(u_multiplier_STAGE1_pp1_37_5_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_38_5__16_ ),
    .ZN(u_multiplier_pp1_38 [0]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_38_5__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_38_5__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_38_5__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_38_5_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_38_5__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_38_5__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_38_5__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_38_5__17_ ),
    .ZN(u_multiplier_pp1_39 [5]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_39_1__18_  (.A(u_multiplier_STAGE1_pp1_38_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_1__19_  (.A1(u_multiplier_STAGE1__1061_ ),
    .A2(u_multiplier_STAGE1__1060_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_1__20_  (.A(u_multiplier_STAGE1__1061_ ),
    .B(u_multiplier_STAGE1__1060_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_39_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_1__21_  (.A1(u_multiplier_STAGE1__1062_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_39_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_1__22_  (.A(u_multiplier_STAGE1__1062_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_39_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_39_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_1__23_  (.A1(u_multiplier_STAGE1__1063_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_39_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_1__24_  (.A(u_multiplier_STAGE1__1063_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_39_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_1__25_  (.A(u_multiplier_STAGE1_pp1_38_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_39_1__16_ ),
    .ZN(u_multiplier_pp1_39 [4]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_39_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_39_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_39_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_39_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_39_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_39_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_39_1__17_ ),
    .ZN(u_multiplier_pp1_40 [8]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_39_2__18_  (.A(u_multiplier_STAGE1_pp1_38_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_2__19_  (.A1(u_multiplier_STAGE1__1065_ ),
    .A2(u_multiplier_STAGE1__1064_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_2__20_  (.A(u_multiplier_STAGE1__1065_ ),
    .B(u_multiplier_STAGE1__1064_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_39_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_2__21_  (.A1(u_multiplier_STAGE1__1066_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_39_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_2__22_  (.A(u_multiplier_STAGE1__1066_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_39_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_39_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_2__23_  (.A1(u_multiplier_STAGE1__1067_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_39_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_2__24_  (.A(u_multiplier_STAGE1__1067_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_39_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_2__25_  (.A(u_multiplier_STAGE1_pp1_38_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_39_2__16_ ),
    .ZN(u_multiplier_pp1_39 [3]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_39_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_39_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_39_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_39_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_39_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_39_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_39_2__17_ ),
    .ZN(u_multiplier_pp1_40 [7]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_39_3__18_  (.A(u_multiplier_STAGE1_pp1_38_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_3__19_  (.A1(u_multiplier_STAGE1__1069_ ),
    .A2(u_multiplier_STAGE1__1068_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_3__20_  (.A(u_multiplier_STAGE1__1069_ ),
    .B(u_multiplier_STAGE1__1068_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_39_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_3__21_  (.A1(u_multiplier_STAGE1__1070_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_39_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_3__22_  (.A(u_multiplier_STAGE1__1070_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_39_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_39_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_3__23_  (.A1(u_multiplier_STAGE1__1071_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_39_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_3__24_  (.A(u_multiplier_STAGE1__1071_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_39_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_3__25_  (.A(u_multiplier_STAGE1_pp1_38_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_39_3__16_ ),
    .ZN(u_multiplier_pp1_39 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_39_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_39_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_39_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_39_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_39_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_39_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_39_3__17_ ),
    .ZN(u_multiplier_pp1_40 [6]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_39_4__18_  (.A(u_multiplier_STAGE1_pp1_38_4_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_4__19_  (.A1(u_multiplier_STAGE1__1073_ ),
    .A2(u_multiplier_STAGE1__1072_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_4__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_4__20_  (.A(u_multiplier_STAGE1__1073_ ),
    .B(u_multiplier_STAGE1__1072_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_39_4__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_4__21_  (.A1(u_multiplier_STAGE1__1074_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_39_4__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_4__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_4__22_  (.A(u_multiplier_STAGE1__1074_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_39_4__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_39_4__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_4__23_  (.A1(u_multiplier_STAGE1__1075_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_39_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_4__24_  (.A(u_multiplier_STAGE1__1075_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_39_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_39_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_39_4__25_  (.A(u_multiplier_STAGE1_pp1_38_4_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_39_4__16_ ),
    .ZN(u_multiplier_pp1_39 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_39_4__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_39_4__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_39_4__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_39_4_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_39_4__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_39_4__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_39_4__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_39_4__17_ ),
    .ZN(u_multiplier_pp1_40 [5]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_40_1__18_  (.A(u_multiplier_STAGE1_pp1_39_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_1__19_  (.A1(u_multiplier_STAGE1__1079_ ),
    .A2(u_multiplier_STAGE1__1078_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_1__20_  (.A(u_multiplier_STAGE1__1079_ ),
    .B(u_multiplier_STAGE1__1078_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_40_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_1__21_  (.A1(u_multiplier_STAGE1__1080_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_40_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_1__22_  (.A(u_multiplier_STAGE1__1080_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_40_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_40_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_1__23_  (.A1(u_multiplier_STAGE1__1081_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_40_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_1__24_  (.A(u_multiplier_STAGE1__1081_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_40_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_1__25_  (.A(u_multiplier_STAGE1_pp1_39_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_40_1__16_ ),
    .ZN(u_multiplier_pp1_40 [3]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_40_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_40_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_40_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_40_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_40_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_40_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_40_1__17_ ),
    .ZN(u_multiplier_pp1_41 [7]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_40_2__18_  (.A(u_multiplier_STAGE1_pp1_39_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_2__19_  (.A1(u_multiplier_STAGE1__1083_ ),
    .A2(u_multiplier_STAGE1__1082_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_2__20_  (.A(u_multiplier_STAGE1__1083_ ),
    .B(u_multiplier_STAGE1__1082_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_40_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_2__21_  (.A1(u_multiplier_STAGE1__1084_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_40_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_2__22_  (.A(u_multiplier_STAGE1__1084_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_40_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_40_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_2__23_  (.A1(u_multiplier_STAGE1__1085_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_40_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_2__24_  (.A(u_multiplier_STAGE1__1085_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_40_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_2__25_  (.A(u_multiplier_STAGE1_pp1_39_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_40_2__16_ ),
    .ZN(u_multiplier_pp1_40 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_40_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_40_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_40_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_40_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_40_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_40_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_40_2__17_ ),
    .ZN(u_multiplier_pp1_41 [6]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_40_3__18_  (.A(u_multiplier_STAGE1_pp1_39_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_3__19_  (.A1(u_multiplier_STAGE1__1087_ ),
    .A2(u_multiplier_STAGE1__1086_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_3__20_  (.A(u_multiplier_STAGE1__1087_ ),
    .B(u_multiplier_STAGE1__1086_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_40_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_3__21_  (.A1(u_multiplier_STAGE1__1088_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_40_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_3__22_  (.A(u_multiplier_STAGE1__1088_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_40_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_40_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_3__23_  (.A1(u_multiplier_STAGE1__1089_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_40_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_3__24_  (.A(u_multiplier_STAGE1__1089_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_40_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_3__25_  (.A(u_multiplier_STAGE1_pp1_39_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_40_3__16_ ),
    .ZN(u_multiplier_pp1_40 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_40_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_40_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_40_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_40_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_40_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_40_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_40_3__17_ ),
    .ZN(u_multiplier_pp1_41 [5]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_40_4__18_  (.A(u_multiplier_STAGE1_pp1_39_4_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_4__19_  (.A1(u_multiplier_STAGE1__1091_ ),
    .A2(u_multiplier_STAGE1__1090_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_4__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_4__20_  (.A(u_multiplier_STAGE1__1091_ ),
    .B(u_multiplier_STAGE1__1090_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_40_4__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_4__21_  (.A1(u_multiplier_STAGE1__1092_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_40_4__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_4__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_4__22_  (.A(u_multiplier_STAGE1__1092_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_40_4__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_40_4__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_4__23_  (.A1(u_multiplier_STAGE1__1093_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_40_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_4__24_  (.A(u_multiplier_STAGE1__1093_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_40_4__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_40_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_40_4__25_  (.A(u_multiplier_STAGE1_pp1_39_4_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_40_4__16_ ),
    .ZN(u_multiplier_pp1_40 [0]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_40_4__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_40_4__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_40_4__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_40_4_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_40_4__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_40_4__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_40_4__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_40_4__17_ ),
    .ZN(u_multiplier_pp1_41 [4]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_41_1__18_  (.A(u_multiplier_STAGE1_pp1_40_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_41_1__19_  (.A1(u_multiplier_STAGE1__1095_ ),
    .A2(u_multiplier_STAGE1__1094_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_41_1__20_  (.A(u_multiplier_STAGE1__1095_ ),
    .B(u_multiplier_STAGE1__1094_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_41_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_41_1__21_  (.A1(u_multiplier_STAGE1__1096_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_41_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_41_1__22_  (.A(u_multiplier_STAGE1__1096_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_41_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_41_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_41_1__23_  (.A1(u_multiplier_STAGE1__1097_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_41_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_41_1__24_  (.A(u_multiplier_STAGE1__1097_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_41_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_41_1__25_  (.A(u_multiplier_STAGE1_pp1_40_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_41_1__16_ ),
    .ZN(u_multiplier_pp1_41 [3]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_41_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_41_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_41_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_41_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_41_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_41_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_41_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_41_1__17_ ),
    .ZN(u_multiplier_pp1_42 [6]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_41_2__18_  (.A(u_multiplier_STAGE1_pp1_40_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_41_2__19_  (.A1(u_multiplier_STAGE1__1099_ ),
    .A2(u_multiplier_STAGE1__1098_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_41_2__20_  (.A(u_multiplier_STAGE1__1099_ ),
    .B(u_multiplier_STAGE1__1098_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_41_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_41_2__21_  (.A1(u_multiplier_STAGE1__1100_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_41_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_41_2__22_  (.A(u_multiplier_STAGE1__1100_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_41_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_41_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_41_2__23_  (.A1(u_multiplier_STAGE1__1101_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_41_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_41_2__24_  (.A(u_multiplier_STAGE1__1101_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_41_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_41_2__25_  (.A(u_multiplier_STAGE1_pp1_40_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_41_2__16_ ),
    .ZN(u_multiplier_pp1_41 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_41_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_41_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_41_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_41_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_41_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_41_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_41_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_41_2__17_ ),
    .ZN(u_multiplier_pp1_42 [5]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_41_3__18_  (.A(u_multiplier_STAGE1_pp1_40_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_41_3__19_  (.A1(u_multiplier_STAGE1__1103_ ),
    .A2(u_multiplier_STAGE1__1102_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_41_3__20_  (.A(u_multiplier_STAGE1__1103_ ),
    .B(u_multiplier_STAGE1__1102_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_41_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_41_3__21_  (.A1(u_multiplier_STAGE1__1104_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_41_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_41_3__22_  (.A(u_multiplier_STAGE1__1104_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_41_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_41_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_41_3__23_  (.A1(u_multiplier_STAGE1__1105_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_41_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_41_3__24_  (.A(u_multiplier_STAGE1__1105_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_41_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_41_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_41_3__25_  (.A(u_multiplier_STAGE1_pp1_40_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_41_3__16_ ),
    .ZN(u_multiplier_pp1_41 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_41_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_41_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_41_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_41_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_41_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_41_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_41_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_41_3__17_ ),
    .ZN(u_multiplier_pp1_42 [4]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_42_1__18_  (.A(u_multiplier_STAGE1_pp1_41_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_42_1__19_  (.A1(u_multiplier_STAGE1__1109_ ),
    .A2(u_multiplier_STAGE1__1108_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_42_1__20_  (.A(u_multiplier_STAGE1__1109_ ),
    .B(u_multiplier_STAGE1__1108_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_42_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_42_1__21_  (.A1(u_multiplier_STAGE1__1110_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_42_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_42_1__22_  (.A(u_multiplier_STAGE1__1110_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_42_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_42_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_42_1__23_  (.A1(u_multiplier_STAGE1__1111_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_42_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_42_1__24_  (.A(u_multiplier_STAGE1__1111_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_42_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_42_1__25_  (.A(u_multiplier_STAGE1_pp1_41_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_42_1__16_ ),
    .ZN(u_multiplier_pp1_42 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_42_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_42_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_42_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_42_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_42_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_42_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_42_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_42_1__17_ ),
    .ZN(u_multiplier_pp1_43 [5]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_42_2__18_  (.A(u_multiplier_STAGE1_pp1_41_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_42_2__19_  (.A1(u_multiplier_STAGE1__1113_ ),
    .A2(u_multiplier_STAGE1__1112_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_42_2__20_  (.A(u_multiplier_STAGE1__1113_ ),
    .B(u_multiplier_STAGE1__1112_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_42_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_42_2__21_  (.A1(u_multiplier_STAGE1__1114_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_42_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_42_2__22_  (.A(u_multiplier_STAGE1__1114_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_42_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_42_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_42_2__23_  (.A1(u_multiplier_STAGE1__1115_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_42_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_42_2__24_  (.A(u_multiplier_STAGE1__1115_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_42_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_42_2__25_  (.A(u_multiplier_STAGE1_pp1_41_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_42_2__16_ ),
    .ZN(u_multiplier_pp1_42 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_42_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_42_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_42_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_42_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_42_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_42_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_42_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_42_2__17_ ),
    .ZN(u_multiplier_pp1_43 [4]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_42_3__18_  (.A(u_multiplier_STAGE1_pp1_41_3_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_42_3__19_  (.A1(u_multiplier_STAGE1__1117_ ),
    .A2(u_multiplier_STAGE1__1116_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_3__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_42_3__20_  (.A(u_multiplier_STAGE1__1117_ ),
    .B(u_multiplier_STAGE1__1116_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_42_3__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_42_3__21_  (.A1(u_multiplier_STAGE1__1118_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_42_3__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_3__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_42_3__22_  (.A(u_multiplier_STAGE1__1118_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_42_3__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_42_3__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_42_3__23_  (.A1(u_multiplier_STAGE1__1119_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_42_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_42_3__24_  (.A(u_multiplier_STAGE1__1119_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_42_3__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_42_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_42_3__25_  (.A(u_multiplier_STAGE1_pp1_41_3_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_42_3__16_ ),
    .ZN(u_multiplier_pp1_42 [0]));
 NAND2_X2 u_multiplier_STAGE1_E_4_2_pp_42_3__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_42_3__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_42_3__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_42_3_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_42_3__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_42_3__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_42_3__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_42_3__17_ ),
    .ZN(u_multiplier_pp1_43 [3]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_43_1__18_  (.A(u_multiplier_STAGE1_pp1_42_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_43_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_43_1__19_  (.A1(u_multiplier_STAGE1__1121_ ),
    .A2(u_multiplier_STAGE1__1120_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_43_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_43_1__20_  (.A(u_multiplier_STAGE1__1121_ ),
    .B(u_multiplier_STAGE1__1120_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_43_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_43_1__21_  (.A1(u_multiplier_STAGE1__1122_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_43_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_43_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_43_1__22_  (.A(u_multiplier_STAGE1__1122_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_43_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_43_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_43_1__23_  (.A1(u_multiplier_STAGE1__1123_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_43_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_43_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_43_1__24_  (.A(u_multiplier_STAGE1__1123_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_43_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_43_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_43_1__25_  (.A(u_multiplier_STAGE1_pp1_42_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_43_1__16_ ),
    .ZN(u_multiplier_pp1_43 [2]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_43_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_43_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_43_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_43_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_43_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_43_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_43_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_43_1__17_ ),
    .ZN(u_multiplier_pp1_44 [4]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_43_2__18_  (.A(u_multiplier_STAGE1_pp1_42_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_43_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_43_2__19_  (.A1(u_multiplier_STAGE1__1125_ ),
    .A2(u_multiplier_STAGE1__1124_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_43_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_43_2__20_  (.A(u_multiplier_STAGE1__1125_ ),
    .B(u_multiplier_STAGE1__1124_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_43_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_43_2__21_  (.A1(u_multiplier_STAGE1__1126_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_43_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_43_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_43_2__22_  (.A(u_multiplier_STAGE1__1126_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_43_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_43_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_43_2__23_  (.A1(u_multiplier_STAGE1__1127_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_43_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_43_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_43_2__24_  (.A(u_multiplier_STAGE1__1127_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_43_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_43_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_43_2__25_  (.A(u_multiplier_STAGE1_pp1_42_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_43_2__16_ ),
    .ZN(u_multiplier_pp1_43 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_43_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_43_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_43_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_43_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_43_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_43_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_43_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_43_2__17_ ),
    .ZN(u_multiplier_pp1_44 [3]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_44_1__18_  (.A(u_multiplier_STAGE1_pp1_43_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_44_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_44_1__19_  (.A1(u_multiplier_STAGE1__1131_ ),
    .A2(u_multiplier_STAGE1__1130_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_44_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_44_1__20_  (.A(u_multiplier_STAGE1__1131_ ),
    .B(u_multiplier_STAGE1__1130_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_44_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_44_1__21_  (.A1(u_multiplier_STAGE1__1132_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_44_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_44_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_44_1__22_  (.A(u_multiplier_STAGE1__1132_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_44_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_44_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_44_1__23_  (.A1(u_multiplier_STAGE1__1133_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_44_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_44_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_44_1__24_  (.A(u_multiplier_STAGE1__1133_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_44_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_44_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_44_1__25_  (.A(u_multiplier_STAGE1_pp1_43_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_44_1__16_ ),
    .ZN(u_multiplier_pp1_44 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_44_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_44_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_44_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_44_1_cout ));
 OAI21_X1 u_multiplier_STAGE1_E_4_2_pp_44_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_44_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_44_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_44_1__17_ ),
    .ZN(u_multiplier_pp1_45 [3]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_44_2__18_  (.A(u_multiplier_STAGE1_pp1_43_2_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_44_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_44_2__19_  (.A1(u_multiplier_STAGE1__1135_ ),
    .A2(u_multiplier_STAGE1__1134_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_44_2__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_44_2__20_  (.A(u_multiplier_STAGE1__1135_ ),
    .B(u_multiplier_STAGE1__1134_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_44_2__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_44_2__21_  (.A1(u_multiplier_STAGE1__1136_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_44_2__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_44_2__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_44_2__22_  (.A(u_multiplier_STAGE1__1136_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_44_2__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_44_2__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_44_2__23_  (.A1(u_multiplier_STAGE1__1137_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_44_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_44_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_44_2__24_  (.A(u_multiplier_STAGE1__1137_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_44_2__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_44_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_44_2__25_  (.A(u_multiplier_STAGE1_pp1_43_2_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_44_2__16_ ),
    .ZN(u_multiplier_pp1_44 [0]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_44_2__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_44_2__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_44_2__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_44_2_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_44_2__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_44_2__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_44_2__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_44_2__17_ ),
    .ZN(u_multiplier_pp1_45 [2]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_45_1__18_  (.A(u_multiplier_STAGE1_pp1_44_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_45_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_45_1__19_  (.A1(u_multiplier_STAGE1__1139_ ),
    .A2(u_multiplier_STAGE1__1138_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_45_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_45_1__20_  (.A(u_multiplier_STAGE1__1139_ ),
    .B(u_multiplier_STAGE1__1138_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_45_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_45_1__21_  (.A1(u_multiplier_STAGE1__1140_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_45_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_45_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_45_1__22_  (.A(u_multiplier_STAGE1__1140_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_45_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_45_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_45_1__23_  (.A1(u_multiplier_STAGE1__1141_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_45_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_45_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_45_1__24_  (.A(u_multiplier_STAGE1__1141_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_45_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_45_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_45_1__25_  (.A(u_multiplier_STAGE1_pp1_44_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_45_1__16_ ),
    .ZN(u_multiplier_pp1_45 [1]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_45_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_45_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_45_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_45_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_45_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_45_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_45_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_45_1__17_ ),
    .ZN(u_multiplier_pp1_46 [2]));
 INV_X1 u_multiplier_STAGE1_E_4_2_pp_46_1__18_  (.A(u_multiplier_STAGE1_pp1_45_1_cout ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_46_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_46_1__19_  (.A1(u_multiplier_STAGE1__1145_ ),
    .A2(u_multiplier_STAGE1__1144_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_46_1__11_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_46_1__20_  (.A(u_multiplier_STAGE1__1145_ ),
    .B(u_multiplier_STAGE1__1144_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_46_1__12_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_46_1__21_  (.A1(u_multiplier_STAGE1__1146_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_46_1__12_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_46_1__13_ ));
 XOR2_X2 u_multiplier_STAGE1_E_4_2_pp_46_1__22_  (.A(u_multiplier_STAGE1__1146_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_46_1__12_ ),
    .Z(u_multiplier_STAGE1_E_4_2_pp_46_1__14_ ));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_46_1__23_  (.A1(u_multiplier_STAGE1__1147_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_46_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_46_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_46_1__24_  (.A(u_multiplier_STAGE1__1147_ ),
    .B(u_multiplier_STAGE1_E_4_2_pp_46_1__14_ ),
    .ZN(u_multiplier_STAGE1_E_4_2_pp_46_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE1_E_4_2_pp_46_1__25_  (.A(u_multiplier_STAGE1_pp1_45_1_cout ),
    .B(u_multiplier_STAGE1_E_4_2_pp_46_1__16_ ),
    .ZN(u_multiplier_pp1_46 [0]));
 NAND2_X1 u_multiplier_STAGE1_E_4_2_pp_46_1__26_  (.A1(u_multiplier_STAGE1_E_4_2_pp_46_1__11_ ),
    .A2(u_multiplier_STAGE1_E_4_2_pp_46_1__13_ ),
    .ZN(u_multiplier_STAGE1_pp1_46_1_cout ));
 OAI21_X2 u_multiplier_STAGE1_E_4_2_pp_46_1__27_  (.A(u_multiplier_STAGE1_E_4_2_pp_46_1__15_ ),
    .B1(u_multiplier_STAGE1_E_4_2_pp_46_1__16_ ),
    .B2(u_multiplier_STAGE1_E_4_2_pp_46_1__17_ ),
    .ZN(u_multiplier_pp1_47 [1]));
 INV_X1 u_multiplier_STAGE1_Full_adder_pp_32_1__12_  (.A(u_multiplier_STAGE1__0909_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_32_1__08_ ));
 NAND3_X1 u_multiplier_STAGE1_Full_adder_pp_32_1__13_  (.A1(u_multiplier_STAGE1__0908_ ),
    .A2(u_multiplier_STAGE1__0907_ ),
    .A3(u_multiplier_STAGE1__0909_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_32_1__09_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_32_1__14_  (.A1(u_multiplier_STAGE1__0908_ ),
    .A2(u_multiplier_STAGE1__0907_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_32_1__10_ ));
 AOI21_X1 u_multiplier_STAGE1_Full_adder_pp_32_1__15_  (.A(u_multiplier_STAGE1__0909_ ),
    .B1(u_multiplier_STAGE1__0907_ ),
    .B2(u_multiplier_STAGE1__0908_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_32_1__11_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_32_1__16_  (.A1(u_multiplier_STAGE1_Full_adder_pp_32_1__10_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_32_1__11_ ),
    .ZN(u_multiplier_pp1_33 [8]));
 AOI22_X2 u_multiplier_STAGE1_Full_adder_pp_32_1__17_  (.A1(u_multiplier_STAGE1_Full_adder_pp_32_1__08_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_32_1__10_ ),
    .B1(u_multiplier_pp1_33 [8]),
    .B2(u_multiplier_STAGE1_Full_adder_pp_32_1__09_ ),
    .ZN(u_multiplier_pp1_32 [0]));
 INV_X1 u_multiplier_STAGE1_Full_adder_pp_35_1__12_  (.A(u_multiplier_STAGE1_pp1_34_7_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_35_1__08_ ));
 NAND3_X2 u_multiplier_STAGE1_Full_adder_pp_35_1__13_  (.A1(u_multiplier_STAGE1__0993_ ),
    .A2(u_multiplier_STAGE1__0992_ ),
    .A3(u_multiplier_STAGE1_pp1_34_7_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_35_1__09_ ));
 NOR2_X4 u_multiplier_STAGE1_Full_adder_pp_35_1__14_  (.A1(u_multiplier_STAGE1__0993_ ),
    .A2(u_multiplier_STAGE1__0992_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_35_1__10_ ));
 AOI21_X2 u_multiplier_STAGE1_Full_adder_pp_35_1__15_  (.A(u_multiplier_STAGE1_pp1_34_7_cout ),
    .B1(u_multiplier_STAGE1__0992_ ),
    .B2(u_multiplier_STAGE1__0993_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_35_1__11_ ));
 NOR2_X4 u_multiplier_STAGE1_Full_adder_pp_35_1__16_  (.A1(u_multiplier_STAGE1_Full_adder_pp_35_1__10_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_35_1__11_ ),
    .ZN(u_multiplier_pp1_36 [6]));
 AOI22_X4 u_multiplier_STAGE1_Full_adder_pp_35_1__17_  (.A1(u_multiplier_STAGE1_Full_adder_pp_35_1__08_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_35_1__10_ ),
    .B1(u_multiplier_pp1_36 [6]),
    .B2(u_multiplier_STAGE1_Full_adder_pp_35_1__09_ ),
    .ZN(u_multiplier_pp1_35 [0]));
 INV_X1 u_multiplier_STAGE1_Full_adder_pp_37_1__12_  (.A(u_multiplier_STAGE1_pp1_36_6_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_37_1__08_ ));
 NAND3_X2 u_multiplier_STAGE1_Full_adder_pp_37_1__13_  (.A1(u_multiplier_STAGE1__1039_ ),
    .A2(u_multiplier_STAGE1__1038_ ),
    .A3(u_multiplier_STAGE1_pp1_36_6_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_37_1__09_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_37_1__14_  (.A1(u_multiplier_STAGE1__1039_ ),
    .A2(u_multiplier_STAGE1__1038_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_37_1__10_ ));
 AOI21_X1 u_multiplier_STAGE1_Full_adder_pp_37_1__15_  (.A(u_multiplier_STAGE1_pp1_36_6_cout ),
    .B1(u_multiplier_STAGE1__1038_ ),
    .B2(u_multiplier_STAGE1__1039_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_37_1__11_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_37_1__16_  (.A1(u_multiplier_STAGE1_Full_adder_pp_37_1__10_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_37_1__11_ ),
    .ZN(u_multiplier_pp1_38 [5]));
 AOI22_X4 u_multiplier_STAGE1_Full_adder_pp_37_1__17_  (.A1(u_multiplier_STAGE1_Full_adder_pp_37_1__08_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_37_1__10_ ),
    .B1(u_multiplier_pp1_38 [5]),
    .B2(u_multiplier_STAGE1_Full_adder_pp_37_1__09_ ),
    .ZN(u_multiplier_pp1_37 [0]));
 INV_X1 u_multiplier_STAGE1_Full_adder_pp_39_1__12_  (.A(u_multiplier_STAGE1_pp1_38_5_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_39_1__08_ ));
 NAND3_X2 u_multiplier_STAGE1_Full_adder_pp_39_1__13_  (.A1(u_multiplier_STAGE1__1077_ ),
    .A2(u_multiplier_STAGE1__1076_ ),
    .A3(u_multiplier_STAGE1_pp1_38_5_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_39_1__09_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_39_1__14_  (.A1(u_multiplier_STAGE1__1077_ ),
    .A2(u_multiplier_STAGE1__1076_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_39_1__10_ ));
 AOI21_X1 u_multiplier_STAGE1_Full_adder_pp_39_1__15_  (.A(u_multiplier_STAGE1_pp1_38_5_cout ),
    .B1(u_multiplier_STAGE1__1076_ ),
    .B2(u_multiplier_STAGE1__1077_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_39_1__11_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_39_1__16_  (.A1(u_multiplier_STAGE1_Full_adder_pp_39_1__10_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_39_1__11_ ),
    .ZN(u_multiplier_pp1_40 [4]));
 AOI22_X4 u_multiplier_STAGE1_Full_adder_pp_39_1__17_  (.A1(u_multiplier_STAGE1_Full_adder_pp_39_1__08_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_39_1__10_ ),
    .B1(u_multiplier_pp1_40 [4]),
    .B2(u_multiplier_STAGE1_Full_adder_pp_39_1__09_ ),
    .ZN(u_multiplier_pp1_39 [0]));
 INV_X1 u_multiplier_STAGE1_Full_adder_pp_41_1__12_  (.A(u_multiplier_STAGE1_pp1_40_4_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_41_1__08_ ));
 NAND3_X2 u_multiplier_STAGE1_Full_adder_pp_41_1__13_  (.A1(u_multiplier_STAGE1__1107_ ),
    .A2(u_multiplier_STAGE1__1106_ ),
    .A3(u_multiplier_STAGE1_pp1_40_4_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_41_1__09_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_41_1__14_  (.A1(u_multiplier_STAGE1__1107_ ),
    .A2(u_multiplier_STAGE1__1106_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_41_1__10_ ));
 AOI21_X1 u_multiplier_STAGE1_Full_adder_pp_41_1__15_  (.A(u_multiplier_STAGE1_pp1_40_4_cout ),
    .B1(u_multiplier_STAGE1__1106_ ),
    .B2(u_multiplier_STAGE1__1107_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_41_1__11_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_41_1__16_  (.A1(u_multiplier_STAGE1_Full_adder_pp_41_1__10_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_41_1__11_ ),
    .ZN(u_multiplier_pp1_42 [3]));
 AOI22_X4 u_multiplier_STAGE1_Full_adder_pp_41_1__17_  (.A1(u_multiplier_STAGE1_Full_adder_pp_41_1__08_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_41_1__10_ ),
    .B1(u_multiplier_pp1_42 [3]),
    .B2(u_multiplier_STAGE1_Full_adder_pp_41_1__09_ ),
    .ZN(u_multiplier_pp1_41 [0]));
 INV_X1 u_multiplier_STAGE1_Full_adder_pp_43_1__12_  (.A(u_multiplier_STAGE1_pp1_42_3_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_43_1__08_ ));
 NAND3_X2 u_multiplier_STAGE1_Full_adder_pp_43_1__13_  (.A1(u_multiplier_STAGE1__1129_ ),
    .A2(u_multiplier_STAGE1__1128_ ),
    .A3(u_multiplier_STAGE1_pp1_42_3_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_43_1__09_ ));
 NOR2_X4 u_multiplier_STAGE1_Full_adder_pp_43_1__14_  (.A1(u_multiplier_STAGE1__1129_ ),
    .A2(u_multiplier_STAGE1__1128_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_43_1__10_ ));
 AOI21_X2 u_multiplier_STAGE1_Full_adder_pp_43_1__15_  (.A(u_multiplier_STAGE1_pp1_42_3_cout ),
    .B1(u_multiplier_STAGE1__1128_ ),
    .B2(u_multiplier_STAGE1__1129_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_43_1__11_ ));
 NOR2_X4 u_multiplier_STAGE1_Full_adder_pp_43_1__16_  (.A1(u_multiplier_STAGE1_Full_adder_pp_43_1__10_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_43_1__11_ ),
    .ZN(u_multiplier_pp1_44 [2]));
 AOI22_X4 u_multiplier_STAGE1_Full_adder_pp_43_1__17_  (.A1(u_multiplier_STAGE1_Full_adder_pp_43_1__08_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_43_1__10_ ),
    .B1(u_multiplier_pp1_44 [2]),
    .B2(u_multiplier_STAGE1_Full_adder_pp_43_1__09_ ),
    .ZN(u_multiplier_pp1_43 [0]));
 INV_X1 u_multiplier_STAGE1_Full_adder_pp_45_1__12_  (.A(u_multiplier_STAGE1_pp1_44_2_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_45_1__08_ ));
 NAND3_X2 u_multiplier_STAGE1_Full_adder_pp_45_1__13_  (.A1(u_multiplier_STAGE1__1143_ ),
    .A2(u_multiplier_STAGE1__1142_ ),
    .A3(u_multiplier_STAGE1_pp1_44_2_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_45_1__09_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_45_1__14_  (.A1(u_multiplier_STAGE1__1143_ ),
    .A2(u_multiplier_STAGE1__1142_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_45_1__10_ ));
 AOI21_X1 u_multiplier_STAGE1_Full_adder_pp_45_1__15_  (.A(u_multiplier_STAGE1_pp1_44_2_cout ),
    .B1(u_multiplier_STAGE1__1142_ ),
    .B2(u_multiplier_STAGE1__1143_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_45_1__11_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_45_1__16_  (.A1(u_multiplier_STAGE1_Full_adder_pp_45_1__10_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_45_1__11_ ),
    .ZN(u_multiplier_pp1_46 [1]));
 AOI22_X4 u_multiplier_STAGE1_Full_adder_pp_45_1__17_  (.A1(u_multiplier_STAGE1_Full_adder_pp_45_1__08_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_45_1__10_ ),
    .B1(u_multiplier_pp1_46 [1]),
    .B2(u_multiplier_STAGE1_Full_adder_pp_45_1__09_ ),
    .ZN(u_multiplier_pp1_45 [0]));
 INV_X1 u_multiplier_STAGE1_Full_adder_pp_47_1__12_  (.A(u_multiplier_STAGE1_pp1_46_1_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_47_1__08_ ));
 NAND3_X2 u_multiplier_STAGE1_Full_adder_pp_47_1__13_  (.A1(u_multiplier_STAGE1__1149_ ),
    .A2(u_multiplier_STAGE1__1148_ ),
    .A3(u_multiplier_STAGE1_pp1_46_1_cout ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_47_1__09_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_47_1__14_  (.A1(u_multiplier_STAGE1__1149_ ),
    .A2(u_multiplier_STAGE1__1148_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_47_1__10_ ));
 AOI21_X1 u_multiplier_STAGE1_Full_adder_pp_47_1__15_  (.A(u_multiplier_STAGE1_pp1_46_1_cout ),
    .B1(u_multiplier_STAGE1__1148_ ),
    .B2(u_multiplier_STAGE1__1149_ ),
    .ZN(u_multiplier_STAGE1_Full_adder_pp_47_1__11_ ));
 NOR2_X2 u_multiplier_STAGE1_Full_adder_pp_47_1__16_  (.A1(u_multiplier_STAGE1_Full_adder_pp_47_1__10_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_47_1__11_ ),
    .ZN(u_multiplier_pp1_48 [0]));
 AOI22_X4 u_multiplier_STAGE1_Full_adder_pp_47_1__17_  (.A1(u_multiplier_STAGE1_Full_adder_pp_47_1__08_ ),
    .A2(u_multiplier_STAGE1_Full_adder_pp_47_1__10_ ),
    .B1(u_multiplier_pp1_48 [0]),
    .B2(u_multiplier_STAGE1_Full_adder_pp_47_1__09_ ),
    .ZN(u_multiplier_pp1_47 [0]));
 AND2_X2 u_multiplier_STAGE1_Half_adder_pp_16__4_  (.A1(u_multiplier_STAGE1__0608_ ),
    .A2(u_multiplier_STAGE1__0607_ ),
    .ZN(u_multiplier_pp1_17 [1]));
 XOR2_X2 u_multiplier_STAGE1_Half_adder_pp_16__5_  (.A(u_multiplier_STAGE1__0608_ ),
    .B(u_multiplier_STAGE1__0607_ ),
    .Z(u_multiplier_pp1_16 [0]));
 AND2_X1 u_multiplier_STAGE1_Half_adder_pp_18__4_  (.A1(u_multiplier_STAGE1__0618_ ),
    .A2(u_multiplier_STAGE1__0617_ ),
    .ZN(u_multiplier_pp1_19 [2]));
 XOR2_X2 u_multiplier_STAGE1_Half_adder_pp_18__5_  (.A(u_multiplier_STAGE1__0618_ ),
    .B(u_multiplier_STAGE1__0617_ ),
    .Z(u_multiplier_pp1_18 [1]));
 AND2_X1 u_multiplier_STAGE1_Half_adder_pp_20__4_  (.A1(u_multiplier_STAGE1__0636_ ),
    .A2(u_multiplier_STAGE1__0635_ ),
    .ZN(u_multiplier_pp1_21 [3]));
 XOR2_X2 u_multiplier_STAGE1_Half_adder_pp_20__5_  (.A(u_multiplier_STAGE1__0636_ ),
    .B(u_multiplier_STAGE1__0635_ ),
    .Z(u_multiplier_pp1_20 [2]));
 AND2_X1 u_multiplier_STAGE1_Half_adder_pp_22__4_  (.A1(u_multiplier_STAGE1__0662_ ),
    .A2(u_multiplier_STAGE1__0661_ ),
    .ZN(u_multiplier_pp1_23 [4]));
 XOR2_X2 u_multiplier_STAGE1_Half_adder_pp_22__5_  (.A(u_multiplier_STAGE1__0662_ ),
    .B(u_multiplier_STAGE1__0661_ ),
    .Z(u_multiplier_pp1_22 [3]));
 AND2_X1 u_multiplier_STAGE1_Half_adder_pp_24__4_  (.A1(u_multiplier_STAGE1__0696_ ),
    .A2(u_multiplier_STAGE1__0695_ ),
    .ZN(u_multiplier_pp1_25 [5]));
 XOR2_X2 u_multiplier_STAGE1_Half_adder_pp_24__5_  (.A(u_multiplier_STAGE1__0696_ ),
    .B(u_multiplier_STAGE1__0695_ ),
    .Z(u_multiplier_pp1_24 [4]));
 AND2_X1 u_multiplier_STAGE1_Half_adder_pp_26__4_  (.A1(u_multiplier_STAGE1__0738_ ),
    .A2(u_multiplier_STAGE1__0737_ ),
    .ZN(u_multiplier_pp1_27 [6]));
 XOR2_X2 u_multiplier_STAGE1_Half_adder_pp_26__5_  (.A(u_multiplier_STAGE1__0738_ ),
    .B(u_multiplier_STAGE1__0737_ ),
    .Z(u_multiplier_pp1_26 [5]));
 AND2_X1 u_multiplier_STAGE1_Half_adder_pp_28__4_  (.A1(u_multiplier_STAGE1__0788_ ),
    .A2(u_multiplier_STAGE1__0787_ ),
    .ZN(u_multiplier_pp1_29 [7]));
 XOR2_X2 u_multiplier_STAGE1_Half_adder_pp_28__5_  (.A(u_multiplier_STAGE1__0788_ ),
    .B(u_multiplier_STAGE1__0787_ ),
    .Z(u_multiplier_pp1_28 [6]));
 AND2_X1 u_multiplier_STAGE1_Half_adder_pp_30__4_  (.A1(u_multiplier_STAGE1__0846_ ),
    .A2(u_multiplier_STAGE1__0845_ ),
    .ZN(u_multiplier_pp1_31 [8]));
 XOR2_X2 u_multiplier_STAGE1_Half_adder_pp_30__5_  (.A(u_multiplier_STAGE1__0846_ ),
    .B(u_multiplier_STAGE1__0845_ ),
    .Z(u_multiplier_pp1_30 [7]));
 AND2_X1 u_multiplier_STAGE1_Half_adder_pp_33_1__4_  (.A1(u_multiplier_STAGE1__0939_ ),
    .A2(u_multiplier_STAGE1__0938_ ),
    .ZN(u_multiplier_pp1_34 [7]));
 XOR2_X2 u_multiplier_STAGE1_Half_adder_pp_33_1__5_  (.A(u_multiplier_STAGE1__0939_ ),
    .B(u_multiplier_STAGE1__0938_ ),
    .Z(u_multiplier_pp1_33 [0]));
 AND2_X1 u_multiplier_STAGE1__1631_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[0]),
    .ZN(u_multiplier_pp3_0 ));
 AND2_X1 u_multiplier_STAGE1__1632_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[1]),
    .ZN(u_multiplier_pp3_1 [0]));
 AND2_X1 u_multiplier_STAGE1__1633_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[1]),
    .ZN(u_multiplier_pp3_1 [1]));
 AND2_X1 u_multiplier_STAGE1__1634_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[2]),
    .ZN(u_multiplier_pp3_2 [0]));
 AND2_X1 u_multiplier_STAGE1__1635_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[1]),
    .ZN(u_multiplier_pp3_2 [1]));
 AND2_X1 u_multiplier_STAGE1__1636_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[2]),
    .ZN(u_multiplier_pp3_2 [2]));
 AND2_X2 u_multiplier_STAGE1__1637_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[3]),
    .ZN(u_multiplier_pp3_3 [0]));
 AND2_X2 u_multiplier_STAGE1__1638_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[2]),
    .ZN(u_multiplier_pp3_3 [1]));
 AND2_X2 u_multiplier_STAGE1__1639_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[2]),
    .ZN(u_multiplier_pp3_3 [2]));
 AND2_X1 u_multiplier_STAGE1__1640_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[3]),
    .ZN(u_multiplier_pp3_3 [3]));
 AND2_X1 u_multiplier_STAGE1__1641_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[4]),
    .ZN(u_multiplier_pp2_4 [4]));
 AND2_X1 u_multiplier_STAGE1__1642_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[3]),
    .ZN(u_multiplier_pp2_4 [3]));
 AND2_X1 u_multiplier_STAGE1__1643_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[2]),
    .ZN(u_multiplier_pp3_4 [1]));
 AND2_X1 u_multiplier_STAGE1__1644_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[3]),
    .ZN(u_multiplier_pp3_4 [2]));
 AND2_X1 u_multiplier_STAGE1__1645_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[4]),
    .ZN(u_multiplier_pp3_4 [3]));
 AND2_X1 u_multiplier_STAGE1__1646_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[5]),
    .ZN(u_multiplier_pp2_5 [5]));
 AND2_X1 u_multiplier_STAGE1__1647_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[4]),
    .ZN(u_multiplier_pp2_5 [4]));
 AND2_X1 u_multiplier_STAGE1__1648_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[3]),
    .ZN(u_multiplier_pp2_5 [3]));
 AND2_X1 u_multiplier_STAGE1__1649_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[3]),
    .ZN(u_multiplier_pp2_5 [2]));
 AND2_X1 u_multiplier_STAGE1__1650_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[4]),
    .ZN(u_multiplier_pp3_5 [2]));
 AND2_X1 u_multiplier_STAGE1__1651_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[5]),
    .ZN(u_multiplier_pp3_5 [3]));
 AND2_X1 u_multiplier_STAGE1__1652_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[6]),
    .ZN(u_multiplier_pp2_6 [6]));
 AND2_X1 u_multiplier_STAGE1__1653_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[5]),
    .ZN(u_multiplier_pp2_6 [5]));
 AND2_X1 u_multiplier_STAGE1__1654_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[4]),
    .ZN(u_multiplier_pp2_6 [4]));
 AND2_X1 u_multiplier_STAGE1__1655_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[3]),
    .ZN(u_multiplier_pp2_6 [3]));
 AND2_X1 u_multiplier_STAGE1__1656_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[4]),
    .ZN(u_multiplier_pp2_6 [2]));
 AND2_X1 u_multiplier_STAGE1__1657_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[5]),
    .ZN(u_multiplier_pp2_6 [1]));
 AND2_X1 u_multiplier_STAGE1__1658_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[6]),
    .ZN(u_multiplier_pp3_6 [3]));
 AND2_X1 u_multiplier_STAGE1__1659_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[7]),
    .ZN(u_multiplier_pp2_7 [7]));
 AND2_X1 u_multiplier_STAGE1__1660_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[6]),
    .ZN(u_multiplier_pp2_7 [6]));
 AND2_X1 u_multiplier_STAGE1__1661_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[5]),
    .ZN(u_multiplier_pp2_7 [5]));
 AND2_X1 u_multiplier_STAGE1__1662_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[4]),
    .ZN(u_multiplier_pp2_7 [4]));
 AND2_X1 u_multiplier_STAGE1__1663_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[4]),
    .ZN(u_multiplier_pp2_7 [3]));
 AND2_X1 u_multiplier_STAGE1__1664_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[5]),
    .ZN(u_multiplier_pp2_7 [2]));
 AND2_X1 u_multiplier_STAGE1__1665_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[6]),
    .ZN(u_multiplier_pp2_7 [1]));
 AND2_X1 u_multiplier_STAGE1__1666_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[7]),
    .ZN(u_multiplier_pp2_7 [0]));
 AND2_X1 u_multiplier_STAGE1__1667_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[8]),
    .ZN(u_multiplier_pp2_8 [7]));
 AND2_X1 u_multiplier_STAGE1__1668_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[7]),
    .ZN(u_multiplier_pp2_8 [6]));
 AND2_X1 u_multiplier_STAGE1__1669_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[6]),
    .ZN(u_multiplier_pp2_8 [5]));
 AND2_X1 u_multiplier_STAGE1__1670_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[5]),
    .ZN(u_multiplier_pp2_8 [4]));
 AND2_X1 u_multiplier_STAGE1__1671_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[4]),
    .ZN(u_multiplier_pp2_8 [3]));
 AND2_X1 u_multiplier_STAGE1__1672_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[5]),
    .ZN(u_multiplier_pp2_8 [2]));
 AND2_X1 u_multiplier_STAGE1__1673_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[6]),
    .ZN(u_multiplier_pp2_8 [1]));
 AND2_X1 u_multiplier_STAGE1__1674_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[7]),
    .ZN(u_multiplier_pp1_8 [7]));
 AND2_X1 u_multiplier_STAGE1__1675_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[8]),
    .ZN(u_multiplier_pp1_8 [8]));
 AND2_X1 u_multiplier_STAGE1__1676_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[9]),
    .ZN(u_multiplier_pp2_9 [7]));
 AND2_X1 u_multiplier_STAGE1__1677_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[8]),
    .ZN(u_multiplier_pp2_9 [6]));
 AND2_X1 u_multiplier_STAGE1__1678_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[7]),
    .ZN(u_multiplier_pp2_9 [5]));
 AND2_X1 u_multiplier_STAGE1__1679_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[6]),
    .ZN(u_multiplier_pp2_9 [4]));
 AND2_X1 u_multiplier_STAGE1__1680_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[5]),
    .ZN(u_multiplier_pp2_9 [3]));
 AND2_X1 u_multiplier_STAGE1__1681_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[5]),
    .ZN(u_multiplier_pp2_9 [2]));
 AND2_X1 u_multiplier_STAGE1__1682_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[6]),
    .ZN(u_multiplier_pp1_9 [6]));
 AND2_X1 u_multiplier_STAGE1__1683_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[7]),
    .ZN(u_multiplier_pp1_9 [7]));
 AND2_X1 u_multiplier_STAGE1__1684_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[8]),
    .ZN(u_multiplier_pp1_9 [8]));
 AND2_X1 u_multiplier_STAGE1__1685_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[9]),
    .ZN(u_multiplier_pp1_9 [9]));
 AND2_X1 u_multiplier_STAGE1__1686_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[10]),
    .ZN(u_multiplier_pp2_10 [7]));
 AND2_X1 u_multiplier_STAGE1__1687_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[9]),
    .ZN(u_multiplier_pp2_10 [6]));
 AND2_X1 u_multiplier_STAGE1__1688_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[8]),
    .ZN(u_multiplier_pp2_10 [5]));
 AND2_X1 u_multiplier_STAGE1__1689_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[7]),
    .ZN(u_multiplier_pp2_10 [4]));
 AND2_X1 u_multiplier_STAGE1__1690_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[6]),
    .ZN(u_multiplier_pp2_10 [3]));
 AND2_X1 u_multiplier_STAGE1__1691_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[5]),
    .ZN(u_multiplier_pp1_10 [5]));
 AND2_X1 u_multiplier_STAGE1__1692_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[6]),
    .ZN(u_multiplier_pp1_10 [6]));
 AND2_X1 u_multiplier_STAGE1__1693_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[7]),
    .ZN(u_multiplier_pp1_10 [7]));
 AND2_X1 u_multiplier_STAGE1__1694_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[8]),
    .ZN(u_multiplier_pp1_10 [8]));
 AND2_X1 u_multiplier_STAGE1__1695_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[9]),
    .ZN(u_multiplier_pp1_10 [9]));
 AND2_X1 u_multiplier_STAGE1__1696_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[10]),
    .ZN(u_multiplier_pp1_10 [10]));
 AND2_X1 u_multiplier_STAGE1__1697_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[11]),
    .ZN(u_multiplier_pp2_11 [7]));
 AND2_X1 u_multiplier_STAGE1__1698_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[10]),
    .ZN(u_multiplier_pp2_11 [6]));
 AND2_X1 u_multiplier_STAGE1__1699_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[9]),
    .ZN(u_multiplier_pp2_11 [5]));
 AND2_X1 u_multiplier_STAGE1__1700_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[8]),
    .ZN(u_multiplier_pp2_11 [4]));
 AND2_X1 u_multiplier_STAGE1__1701_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[7]),
    .ZN(u_multiplier_pp1_11 [4]));
 AND2_X1 u_multiplier_STAGE1__1702_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[6]),
    .ZN(u_multiplier_pp1_11 [5]));
 AND2_X1 u_multiplier_STAGE1__1703_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[6]),
    .ZN(u_multiplier_pp1_11 [6]));
 AND2_X1 u_multiplier_STAGE1__1704_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[7]),
    .ZN(u_multiplier_pp1_11 [7]));
 AND2_X1 u_multiplier_STAGE1__1705_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[8]),
    .ZN(u_multiplier_pp1_11 [8]));
 AND2_X1 u_multiplier_STAGE1__1706_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[9]),
    .ZN(u_multiplier_pp1_11 [9]));
 AND2_X1 u_multiplier_STAGE1__1707_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[10]),
    .ZN(u_multiplier_pp1_11 [10]));
 AND2_X1 u_multiplier_STAGE1__1708_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[11]),
    .ZN(u_multiplier_pp1_11 [11]));
 AND2_X1 u_multiplier_STAGE1__1709_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[12]),
    .ZN(u_multiplier_pp2_12 [7]));
 AND2_X1 u_multiplier_STAGE1__1710_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[11]),
    .ZN(u_multiplier_pp2_12 [6]));
 AND2_X1 u_multiplier_STAGE1__1711_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[10]),
    .ZN(u_multiplier_pp2_12 [5]));
 AND2_X1 u_multiplier_STAGE1__1712_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[9]),
    .ZN(u_multiplier_pp1_12 [3]));
 AND2_X1 u_multiplier_STAGE1__1713_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[8]),
    .ZN(u_multiplier_pp1_12 [4]));
 AND2_X1 u_multiplier_STAGE1__1714_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[7]),
    .ZN(u_multiplier_pp1_12 [5]));
 AND2_X1 u_multiplier_STAGE1__1715_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[6]),
    .ZN(u_multiplier_pp1_12 [6]));
 AND2_X1 u_multiplier_STAGE1__1716_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[7]),
    .ZN(u_multiplier_pp1_12 [7]));
 AND2_X1 u_multiplier_STAGE1__1717_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[8]),
    .ZN(u_multiplier_pp1_12 [8]));
 AND2_X1 u_multiplier_STAGE1__1718_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[9]),
    .ZN(u_multiplier_pp1_12 [9]));
 AND2_X1 u_multiplier_STAGE1__1719_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[10]),
    .ZN(u_multiplier_pp1_12 [10]));
 AND2_X1 u_multiplier_STAGE1__1720_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[11]),
    .ZN(u_multiplier_pp1_12 [11]));
 AND2_X1 u_multiplier_STAGE1__1721_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[12]),
    .ZN(u_multiplier_pp1_12 [12]));
 AND2_X1 u_multiplier_STAGE1__1722_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[13]),
    .ZN(u_multiplier_pp2_13 [7]));
 AND2_X1 u_multiplier_STAGE1__1723_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[12]),
    .ZN(u_multiplier_pp2_13 [6]));
 AND2_X1 u_multiplier_STAGE1__1724_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[11]),
    .ZN(u_multiplier_pp1_13 [2]));
 AND2_X1 u_multiplier_STAGE1__1725_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[10]),
    .ZN(u_multiplier_pp1_13 [3]));
 AND2_X1 u_multiplier_STAGE1__1726_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[9]),
    .ZN(u_multiplier_pp1_13 [4]));
 AND2_X1 u_multiplier_STAGE1__1727_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[8]),
    .ZN(u_multiplier_pp1_13 [5]));
 AND2_X1 u_multiplier_STAGE1__1728_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[7]),
    .ZN(u_multiplier_pp1_13 [6]));
 AND2_X1 u_multiplier_STAGE1__1729_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[7]),
    .ZN(u_multiplier_pp1_13 [7]));
 AND2_X1 u_multiplier_STAGE1__1730_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[8]),
    .ZN(u_multiplier_pp1_13 [8]));
 AND2_X1 u_multiplier_STAGE1__1731_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[9]),
    .ZN(u_multiplier_pp1_13 [9]));
 AND2_X1 u_multiplier_STAGE1__1732_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[10]),
    .ZN(u_multiplier_pp1_13 [10]));
 AND2_X1 u_multiplier_STAGE1__1733_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[11]),
    .ZN(u_multiplier_pp1_13 [11]));
 AND2_X1 u_multiplier_STAGE1__1734_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[12]),
    .ZN(u_multiplier_pp1_13 [12]));
 AND2_X1 u_multiplier_STAGE1__1735_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_pp1_13 [13]));
 AND2_X1 u_multiplier_STAGE1__1736_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_pp2_14 [7]));
 AND2_X1 u_multiplier_STAGE1__1737_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[13]),
    .ZN(u_multiplier_pp1_14 [1]));
 AND2_X1 u_multiplier_STAGE1__1738_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[12]),
    .ZN(u_multiplier_pp1_14 [2]));
 AND2_X1 u_multiplier_STAGE1__1739_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[11]),
    .ZN(u_multiplier_pp1_14 [3]));
 AND2_X1 u_multiplier_STAGE1__1740_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[10]),
    .ZN(u_multiplier_pp1_14 [4]));
 AND2_X1 u_multiplier_STAGE1__1741_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[9]),
    .ZN(u_multiplier_pp1_14 [5]));
 AND2_X1 u_multiplier_STAGE1__1742_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[8]),
    .ZN(u_multiplier_pp1_14 [6]));
 AND2_X1 u_multiplier_STAGE1__1743_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[7]),
    .ZN(u_multiplier_pp1_14 [7]));
 AND2_X1 u_multiplier_STAGE1__1744_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[8]),
    .ZN(u_multiplier_pp1_14 [8]));
 AND2_X1 u_multiplier_STAGE1__1745_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[9]),
    .ZN(u_multiplier_pp1_14 [9]));
 AND2_X1 u_multiplier_STAGE1__1746_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[10]),
    .ZN(u_multiplier_pp1_14 [10]));
 AND2_X1 u_multiplier_STAGE1__1747_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[11]),
    .ZN(u_multiplier_pp1_14 [11]));
 AND2_X1 u_multiplier_STAGE1__1748_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[12]),
    .ZN(u_multiplier_pp1_14 [12]));
 AND2_X1 u_multiplier_STAGE1__1749_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_pp1_14 [13]));
 AND2_X1 u_multiplier_STAGE1__1750_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_pp1_14 [14]));
 AND2_X1 u_multiplier_STAGE1__1751_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_pp1_15 [0]));
 AND2_X1 u_multiplier_STAGE1__1752_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_pp1_15 [1]));
 AND2_X1 u_multiplier_STAGE1__1753_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[13]),
    .ZN(u_multiplier_pp1_15 [2]));
 AND2_X1 u_multiplier_STAGE1__1754_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[12]),
    .ZN(u_multiplier_pp1_15 [3]));
 AND2_X1 u_multiplier_STAGE1__1755_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[11]),
    .ZN(u_multiplier_pp1_15 [4]));
 AND2_X1 u_multiplier_STAGE1__1756_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[10]),
    .ZN(u_multiplier_pp1_15 [5]));
 AND2_X1 u_multiplier_STAGE1__1757_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[9]),
    .ZN(u_multiplier_pp1_15 [6]));
 AND2_X1 u_multiplier_STAGE1__1758_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[8]),
    .ZN(u_multiplier_pp1_15 [7]));
 AND2_X1 u_multiplier_STAGE1__1759_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[8]),
    .ZN(u_multiplier_pp1_15 [8]));
 AND2_X1 u_multiplier_STAGE1__1760_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[9]),
    .ZN(u_multiplier_pp1_15 [9]));
 AND2_X1 u_multiplier_STAGE1__1761_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[10]),
    .ZN(u_multiplier_pp1_15 [10]));
 AND2_X1 u_multiplier_STAGE1__1762_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[11]),
    .ZN(u_multiplier_pp1_15 [11]));
 AND2_X1 u_multiplier_STAGE1__1763_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[12]),
    .ZN(u_multiplier_pp1_15 [12]));
 AND2_X1 u_multiplier_STAGE1__1764_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_pp1_15 [13]));
 AND2_X1 u_multiplier_STAGE1__1765_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_pp1_15 [14]));
 AND2_X1 u_multiplier_STAGE1__1766_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_pp1_15 [15]));
 AND2_X1 u_multiplier_STAGE1__1767_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_STAGE1__0607_ ));
 AND2_X1 u_multiplier_STAGE1__1768_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_STAGE1__0608_ ));
 AND2_X1 u_multiplier_STAGE1__1769_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_pp1_16 [1]));
 AND2_X1 u_multiplier_STAGE1__1770_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[13]),
    .ZN(u_multiplier_pp1_16 [2]));
 AND2_X1 u_multiplier_STAGE1__1771_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[12]),
    .ZN(u_multiplier_pp1_16 [3]));
 AND2_X1 u_multiplier_STAGE1__1772_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[11]),
    .ZN(u_multiplier_pp1_16 [4]));
 AND2_X1 u_multiplier_STAGE1__1773_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[10]),
    .ZN(u_multiplier_pp1_16 [5]));
 AND2_X1 u_multiplier_STAGE1__1774_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[9]),
    .ZN(u_multiplier_pp1_16 [6]));
 AND2_X1 u_multiplier_STAGE1__1775_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[8]),
    .ZN(u_multiplier_pp1_16 [7]));
 AND2_X1 u_multiplier_STAGE1__1776_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[9]),
    .ZN(u_multiplier_pp1_16 [8]));
 AND2_X1 u_multiplier_STAGE1__1777_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[10]),
    .ZN(u_multiplier_pp1_16 [9]));
 AND2_X1 u_multiplier_STAGE1__1778_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[11]),
    .ZN(u_multiplier_pp1_16 [10]));
 AND2_X1 u_multiplier_STAGE1__1779_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[12]),
    .ZN(u_multiplier_pp1_16 [11]));
 AND2_X1 u_multiplier_STAGE1__1780_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_pp1_16 [12]));
 AND2_X1 u_multiplier_STAGE1__1781_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_pp1_16 [13]));
 AND2_X1 u_multiplier_STAGE1__1782_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_pp1_16 [14]));
 AND2_X1 u_multiplier_STAGE1__1783_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_pp1_16 [15]));
 AND2_X1 u_multiplier_STAGE1__1784_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_STAGE1__0609_ ));
 AND2_X1 u_multiplier_STAGE1__1785_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_STAGE1__0610_ ));
 AND2_X1 u_multiplier_STAGE1__1786_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_STAGE1__0611_ ));
 AND2_X1 u_multiplier_STAGE1__1787_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0612_ ));
 AND2_X1 u_multiplier_STAGE1__1788_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[13]),
    .ZN(u_multiplier_pp1_17 [2]));
 AND2_X1 u_multiplier_STAGE1__1789_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[12]),
    .ZN(u_multiplier_pp1_17 [3]));
 AND2_X1 u_multiplier_STAGE1__1790_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[11]),
    .ZN(u_multiplier_pp1_17 [4]));
 AND2_X1 u_multiplier_STAGE1__1791_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[10]),
    .ZN(u_multiplier_pp1_17 [5]));
 AND2_X1 u_multiplier_STAGE1__1792_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[9]),
    .ZN(u_multiplier_pp1_17 [6]));
 AND2_X1 u_multiplier_STAGE1__1793_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[9]),
    .ZN(u_multiplier_pp1_17 [7]));
 AND2_X1 u_multiplier_STAGE1__1794_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[10]),
    .ZN(u_multiplier_pp1_17 [8]));
 AND2_X1 u_multiplier_STAGE1__1795_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[11]),
    .ZN(u_multiplier_pp1_17 [9]));
 AND2_X1 u_multiplier_STAGE1__1796_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[12]),
    .ZN(u_multiplier_pp1_17 [10]));
 AND2_X1 u_multiplier_STAGE1__1797_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_pp1_17 [11]));
 AND2_X1 u_multiplier_STAGE1__1798_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_pp1_17 [12]));
 AND2_X1 u_multiplier_STAGE1__1799_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_pp1_17 [13]));
 AND2_X1 u_multiplier_STAGE1__1800_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_pp1_17 [14]));
 AND2_X1 u_multiplier_STAGE1__1801_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_pp1_17 [15]));
 AND2_X1 u_multiplier_STAGE1__1802_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_STAGE1__0613_ ));
 AND2_X1 u_multiplier_STAGE1__1803_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_STAGE1__0614_ ));
 AND2_X1 u_multiplier_STAGE1__1804_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0615_ ));
 AND2_X1 u_multiplier_STAGE1__1805_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0616_ ));
 AND2_X1 u_multiplier_STAGE1__1806_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[13]),
    .ZN(u_multiplier_STAGE1__0617_ ));
 AND2_X1 u_multiplier_STAGE1__1807_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_STAGE1__0618_ ));
 AND2_X1 u_multiplier_STAGE1__1808_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[12]),
    .ZN(u_multiplier_pp1_18 [3]));
 AND2_X1 u_multiplier_STAGE1__1809_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[11]),
    .ZN(u_multiplier_pp1_18 [4]));
 AND2_X1 u_multiplier_STAGE1__1810_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[10]),
    .ZN(u_multiplier_pp1_18 [5]));
 AND2_X1 u_multiplier_STAGE1__1811_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[9]),
    .ZN(u_multiplier_pp1_18 [6]));
 AND2_X1 u_multiplier_STAGE1__1812_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[10]),
    .ZN(u_multiplier_pp1_18 [7]));
 AND2_X1 u_multiplier_STAGE1__1813_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[11]),
    .ZN(u_multiplier_pp1_18 [8]));
 AND2_X1 u_multiplier_STAGE1__1814_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[12]),
    .ZN(u_multiplier_pp1_18 [9]));
 AND2_X1 u_multiplier_STAGE1__1815_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_pp1_18 [10]));
 AND2_X1 u_multiplier_STAGE1__1816_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_pp1_18 [11]));
 AND2_X1 u_multiplier_STAGE1__1817_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_pp1_18 [12]));
 AND2_X1 u_multiplier_STAGE1__1818_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_pp1_18 [13]));
 AND2_X1 u_multiplier_STAGE1__1819_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_pp1_18 [14]));
 AND2_X1 u_multiplier_STAGE1__1820_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_pp1_18 [15]));
 AND2_X1 u_multiplier_STAGE1__1821_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_STAGE1__0619_ ));
 AND2_X1 u_multiplier_STAGE1__1822_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0620_ ));
 AND2_X1 u_multiplier_STAGE1__1823_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0621_ ));
 AND2_X1 u_multiplier_STAGE1__1824_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0622_ ));
 AND2_X1 u_multiplier_STAGE1__1825_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[12]),
    .ZN(u_multiplier_STAGE1__0623_ ));
 AND2_X1 u_multiplier_STAGE1__1826_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[13]),
    .ZN(u_multiplier_STAGE1__0624_ ));
 AND2_X1 u_multiplier_STAGE1__1827_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_STAGE1__0625_ ));
 AND2_X1 u_multiplier_STAGE1__1828_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_STAGE1__0626_ ));
 AND2_X1 u_multiplier_STAGE1__1829_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[11]),
    .ZN(u_multiplier_pp1_19 [4]));
 AND2_X1 u_multiplier_STAGE1__1830_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[10]),
    .ZN(u_multiplier_pp1_19 [5]));
 AND2_X1 u_multiplier_STAGE1__1831_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[10]),
    .ZN(u_multiplier_pp1_19 [6]));
 AND2_X1 u_multiplier_STAGE1__1832_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[11]),
    .ZN(u_multiplier_pp1_19 [7]));
 AND2_X1 u_multiplier_STAGE1__1833_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[12]),
    .ZN(u_multiplier_pp1_19 [8]));
 AND2_X1 u_multiplier_STAGE1__1834_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_pp1_19 [9]));
 AND2_X1 u_multiplier_STAGE1__1835_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_pp1_19 [10]));
 AND2_X1 u_multiplier_STAGE1__1836_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_pp1_19 [11]));
 AND2_X1 u_multiplier_STAGE1__1837_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_pp1_19 [12]));
 AND2_X1 u_multiplier_STAGE1__1838_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_pp1_19 [13]));
 AND2_X1 u_multiplier_STAGE1__1839_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_pp1_19 [14]));
 AND2_X1 u_multiplier_STAGE1__1840_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_pp1_19 [15]));
 AND2_X1 u_multiplier_STAGE1__1841_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0627_ ));
 AND2_X1 u_multiplier_STAGE1__1842_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0628_ ));
 AND2_X1 u_multiplier_STAGE1__1843_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0629_ ));
 AND2_X1 u_multiplier_STAGE1__1844_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__0630_ ));
 AND2_X1 u_multiplier_STAGE1__1845_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[13]),
    .ZN(u_multiplier_STAGE1__0631_ ));
 AND2_X1 u_multiplier_STAGE1__1846_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_STAGE1__0632_ ));
 AND2_X1 u_multiplier_STAGE1__1847_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_STAGE1__0633_ ));
 AND2_X1 u_multiplier_STAGE1__1848_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_STAGE1__0634_ ));
 AND2_X1 u_multiplier_STAGE1__1849_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[11]),
    .ZN(u_multiplier_STAGE1__0635_ ));
 AND2_X1 u_multiplier_STAGE1__1850_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[12]),
    .ZN(u_multiplier_STAGE1__0636_ ));
 AND2_X1 u_multiplier_STAGE1__1851_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[10]),
    .ZN(u_multiplier_pp1_20 [5]));
 AND2_X1 u_multiplier_STAGE1__1852_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[11]),
    .ZN(u_multiplier_pp1_20 [6]));
 AND2_X1 u_multiplier_STAGE1__1853_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[12]),
    .ZN(u_multiplier_pp1_20 [7]));
 AND2_X1 u_multiplier_STAGE1__1854_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_pp1_20 [8]));
 AND2_X1 u_multiplier_STAGE1__1855_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_pp1_20 [9]));
 AND2_X1 u_multiplier_STAGE1__1856_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_pp1_20 [10]));
 AND2_X1 u_multiplier_STAGE1__1857_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_pp1_20 [11]));
 AND2_X1 u_multiplier_STAGE1__1858_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_pp1_20 [12]));
 AND2_X1 u_multiplier_STAGE1__1859_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_pp1_20 [13]));
 AND2_X1 u_multiplier_STAGE1__1860_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_pp1_20 [14]));
 AND2_X1 u_multiplier_STAGE1__1861_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_pp1_20 [15]));
 AND2_X1 u_multiplier_STAGE1__1862_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0637_ ));
 AND2_X1 u_multiplier_STAGE1__1863_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0638_ ));
 AND2_X1 u_multiplier_STAGE1__1864_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__0639_ ));
 AND2_X1 u_multiplier_STAGE1__1865_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__0640_ ));
 AND2_X1 u_multiplier_STAGE1__1866_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_STAGE1__0641_ ));
 AND2_X1 u_multiplier_STAGE1__1867_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_STAGE1__0642_ ));
 AND2_X1 u_multiplier_STAGE1__1868_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_STAGE1__0643_ ));
 AND2_X1 u_multiplier_STAGE1__1869_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0644_ ));
 AND2_X1 u_multiplier_STAGE1__1870_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[11]),
    .ZN(u_multiplier_STAGE1__0645_ ));
 AND2_X1 u_multiplier_STAGE1__1871_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[11]),
    .ZN(u_multiplier_STAGE1__0646_ ));
 AND2_X1 u_multiplier_STAGE1__1872_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[12]),
    .ZN(u_multiplier_STAGE1__0647_ ));
 AND2_X1 u_multiplier_STAGE1__1873_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[13]),
    .ZN(u_multiplier_STAGE1__0648_ ));
 AND2_X1 u_multiplier_STAGE1__1874_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[12]),
    .ZN(u_multiplier_pp1_21 [6]));
 AND2_X1 u_multiplier_STAGE1__1875_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_pp1_21 [7]));
 AND2_X1 u_multiplier_STAGE1__1876_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_pp1_21 [8]));
 AND2_X1 u_multiplier_STAGE1__1877_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_pp1_21 [9]));
 AND2_X1 u_multiplier_STAGE1__1878_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_pp1_21 [10]));
 AND2_X1 u_multiplier_STAGE1__1879_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_pp1_21 [11]));
 AND2_X1 u_multiplier_STAGE1__1880_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_pp1_21 [12]));
 AND2_X1 u_multiplier_STAGE1__1881_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_pp1_21 [13]));
 AND2_X1 u_multiplier_STAGE1__1882_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_pp1_21 [14]));
 AND2_X1 u_multiplier_STAGE1__1883_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_pp1_21 [15]));
 AND2_X1 u_multiplier_STAGE1__1884_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0649_ ));
 AND2_X1 u_multiplier_STAGE1__1885_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__0650_ ));
 AND2_X1 u_multiplier_STAGE1__1886_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__0651_ ));
 AND2_X1 u_multiplier_STAGE1__1887_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__0652_ ));
 AND2_X1 u_multiplier_STAGE1__1888_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_STAGE1__0653_ ));
 AND2_X1 u_multiplier_STAGE1__1889_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_STAGE1__0654_ ));
 AND2_X1 u_multiplier_STAGE1__1890_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0655_ ));
 AND2_X1 u_multiplier_STAGE1__1891_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0656_ ));
 AND2_X1 u_multiplier_STAGE1__1892_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[11]),
    .ZN(u_multiplier_STAGE1__0657_ ));
 AND2_X1 u_multiplier_STAGE1__1893_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[12]),
    .ZN(u_multiplier_STAGE1__0658_ ));
 AND2_X1 u_multiplier_STAGE1__1894_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[13]),
    .ZN(u_multiplier_STAGE1__0659_ ));
 AND2_X1 u_multiplier_STAGE1__1895_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_STAGE1__0660_ ));
 AND2_X1 u_multiplier_STAGE1__1896_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_STAGE1__0661_ ));
 AND2_X1 u_multiplier_STAGE1__1897_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[12]),
    .ZN(u_multiplier_STAGE1__0662_ ));
 AND2_X1 u_multiplier_STAGE1__1898_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_pp1_22 [7]));
 AND2_X1 u_multiplier_STAGE1__1899_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_pp1_22 [8]));
 AND2_X1 u_multiplier_STAGE1__1900_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_pp1_22 [9]));
 AND2_X1 u_multiplier_STAGE1__1901_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_pp1_22 [10]));
 AND2_X1 u_multiplier_STAGE1__1902_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_pp1_22 [11]));
 AND2_X1 u_multiplier_STAGE1__1903_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_pp1_22 [12]));
 AND2_X1 u_multiplier_STAGE1__1904_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_pp1_22 [13]));
 AND2_X1 u_multiplier_STAGE1__1905_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_pp1_22 [14]));
 AND2_X1 u_multiplier_STAGE1__1906_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_pp1_22 [15]));
 AND2_X1 u_multiplier_STAGE1__1907_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__0663_ ));
 AND2_X1 u_multiplier_STAGE1__1908_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__0664_ ));
 AND2_X1 u_multiplier_STAGE1__1909_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__0665_ ));
 AND2_X1 u_multiplier_STAGE1__1910_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__0666_ ));
 AND2_X1 u_multiplier_STAGE1__1911_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_STAGE1__0667_ ));
 AND2_X1 u_multiplier_STAGE1__1912_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0668_ ));
 AND2_X1 u_multiplier_STAGE1__1913_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0669_ ));
 AND2_X1 u_multiplier_STAGE1__1914_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0670_ ));
 AND2_X1 u_multiplier_STAGE1__1915_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[12]),
    .ZN(u_multiplier_STAGE1__0671_ ));
 AND2_X1 u_multiplier_STAGE1__1916_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[13]),
    .ZN(u_multiplier_STAGE1__0672_ ));
 AND2_X1 u_multiplier_STAGE1__1917_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_STAGE1__0673_ ));
 AND2_X1 u_multiplier_STAGE1__1918_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_STAGE1__0674_ ));
 AND2_X1 u_multiplier_STAGE1__1919_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_STAGE1__0675_ ));
 AND2_X1 u_multiplier_STAGE1__1920_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_STAGE1__0676_ ));
 AND2_X1 u_multiplier_STAGE1__1921_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_STAGE1__0677_ ));
 AND2_X1 u_multiplier_STAGE1__1922_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[12]),
    .ZN(u_multiplier_STAGE1__0678_ ));
 AND2_X1 u_multiplier_STAGE1__1923_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_pp1_23 [8]));
 AND2_X1 u_multiplier_STAGE1__1924_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_pp1_23 [9]));
 AND2_X1 u_multiplier_STAGE1__1925_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_pp1_23 [10]));
 AND2_X1 u_multiplier_STAGE1__1926_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_pp1_23 [11]));
 AND2_X1 u_multiplier_STAGE1__1927_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_pp1_23 [12]));
 AND2_X1 u_multiplier_STAGE1__1928_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_pp1_23 [13]));
 AND2_X1 u_multiplier_STAGE1__1929_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_pp1_23 [14]));
 AND2_X1 u_multiplier_STAGE1__1930_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_pp1_23 [15]));
 AND2_X1 u_multiplier_STAGE1__1931_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__0679_ ));
 AND2_X1 u_multiplier_STAGE1__1932_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__0680_ ));
 AND2_X1 u_multiplier_STAGE1__1933_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__0681_ ));
 AND2_X1 u_multiplier_STAGE1__1934_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__0682_ ));
 AND2_X1 u_multiplier_STAGE1__1935_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0683_ ));
 AND2_X1 u_multiplier_STAGE1__1936_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0684_ ));
 AND2_X1 u_multiplier_STAGE1__1937_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0685_ ));
 AND2_X1 u_multiplier_STAGE1__1938_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__0686_ ));
 AND2_X1 u_multiplier_STAGE1__1939_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[13]),
    .ZN(u_multiplier_STAGE1__0687_ ));
 AND2_X1 u_multiplier_STAGE1__1940_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_STAGE1__0688_ ));
 AND2_X1 u_multiplier_STAGE1__1941_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_STAGE1__0689_ ));
 AND2_X1 u_multiplier_STAGE1__1942_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_STAGE1__0690_ ));
 AND2_X1 u_multiplier_STAGE1__1943_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_STAGE1__0691_ ));
 AND2_X1 u_multiplier_STAGE1__1944_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_STAGE1__0692_ ));
 AND2_X1 u_multiplier_STAGE1__1945_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_STAGE1__0693_ ));
 AND2_X1 u_multiplier_STAGE1__1946_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[12]),
    .ZN(u_multiplier_STAGE1__0694_ ));
 AND2_X1 u_multiplier_STAGE1__1947_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0695_ ));
 AND2_X1 u_multiplier_STAGE1__1948_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_STAGE1__0696_ ));
 AND2_X1 u_multiplier_STAGE1__1949_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_pp1_24 [9]));
 AND2_X1 u_multiplier_STAGE1__1950_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_pp1_24 [10]));
 AND2_X1 u_multiplier_STAGE1__1951_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_pp1_24 [11]));
 AND2_X1 u_multiplier_STAGE1__1952_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_pp1_24 [12]));
 AND2_X1 u_multiplier_STAGE1__1953_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_pp1_24 [13]));
 AND2_X1 u_multiplier_STAGE1__1954_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_pp1_24 [14]));
 AND2_X1 u_multiplier_STAGE1__1955_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_pp1_24 [15]));
 AND2_X1 u_multiplier_STAGE1__1956_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__0697_ ));
 AND2_X1 u_multiplier_STAGE1__1957_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__0698_ ));
 AND2_X1 u_multiplier_STAGE1__1958_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__0699_ ));
 AND2_X1 u_multiplier_STAGE1__1959_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__0700_ ));
 AND2_X1 u_multiplier_STAGE1__1960_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0701_ ));
 AND2_X1 u_multiplier_STAGE1__1961_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0702_ ));
 AND2_X1 u_multiplier_STAGE1__1962_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__0703_ ));
 AND2_X1 u_multiplier_STAGE1__1963_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__0704_ ));
 AND2_X1 u_multiplier_STAGE1__1964_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_STAGE1__0705_ ));
 AND2_X1 u_multiplier_STAGE1__1965_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_STAGE1__0706_ ));
 AND2_X1 u_multiplier_STAGE1__1966_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_STAGE1__0707_ ));
 AND2_X1 u_multiplier_STAGE1__1967_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0708_ ));
 AND2_X1 u_multiplier_STAGE1__1968_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_STAGE1__0709_ ));
 AND2_X1 u_multiplier_STAGE1__1969_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_STAGE1__0710_ ));
 AND2_X1 u_multiplier_STAGE1__1970_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_STAGE1__0711_ ));
 AND2_X1 u_multiplier_STAGE1__1971_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[13]),
    .ZN(u_multiplier_STAGE1__0712_ ));
 AND2_X1 u_multiplier_STAGE1__1972_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0713_ ));
 AND2_X1 u_multiplier_STAGE1__1973_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0714_ ));
 AND2_X1 u_multiplier_STAGE1__1974_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0715_ ));
 AND2_X1 u_multiplier_STAGE1__1975_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_STAGE1__0716_ ));
 AND2_X1 u_multiplier_STAGE1__1976_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_pp1_25 [10]));
 AND2_X1 u_multiplier_STAGE1__1977_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_pp1_25 [11]));
 AND2_X1 u_multiplier_STAGE1__1978_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_pp1_25 [12]));
 AND2_X1 u_multiplier_STAGE1__1979_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_pp1_25 [13]));
 AND2_X1 u_multiplier_STAGE1__1980_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_pp1_25 [14]));
 AND2_X1 u_multiplier_STAGE1__1981_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_pp1_25 [15]));
 AND2_X1 u_multiplier_STAGE1__1982_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__0717_ ));
 AND2_X1 u_multiplier_STAGE1__1983_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__0718_ ));
 AND2_X1 u_multiplier_STAGE1__1984_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__0719_ ));
 AND2_X1 u_multiplier_STAGE1__1985_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__0720_ ));
 AND2_X1 u_multiplier_STAGE1__1986_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0721_ ));
 AND2_X1 u_multiplier_STAGE1__1987_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__0722_ ));
 AND2_X1 u_multiplier_STAGE1__1988_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__0723_ ));
 AND2_X1 u_multiplier_STAGE1__1989_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__0724_ ));
 AND2_X1 u_multiplier_STAGE1__1990_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_STAGE1__0725_ ));
 AND2_X1 u_multiplier_STAGE1__1991_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_STAGE1__0726_ ));
 AND2_X1 u_multiplier_STAGE1__1992_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0727_ ));
 AND2_X1 u_multiplier_STAGE1__1993_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0728_ ));
 AND2_X1 u_multiplier_STAGE1__1994_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_STAGE1__0729_ ));
 AND2_X1 u_multiplier_STAGE1__1995_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_STAGE1__0730_ ));
 AND2_X1 u_multiplier_STAGE1__1996_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[13]),
    .ZN(u_multiplier_STAGE1__0731_ ));
 AND2_X1 u_multiplier_STAGE1__1997_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_STAGE1__0732_ ));
 AND2_X1 u_multiplier_STAGE1__1998_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0733_ ));
 AND2_X1 u_multiplier_STAGE1__1999_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0734_ ));
 AND2_X1 u_multiplier_STAGE1__2000_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0735_ ));
 AND2_X1 u_multiplier_STAGE1__2001_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_STAGE1__0736_ ));
 AND2_X1 u_multiplier_STAGE1__2002_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__0737_ ));
 AND2_X1 u_multiplier_STAGE1__2003_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__0738_ ));
 AND2_X1 u_multiplier_STAGE1__2004_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_pp1_26 [11]));
 AND2_X1 u_multiplier_STAGE1__2005_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_pp1_26 [12]));
 AND2_X1 u_multiplier_STAGE1__2006_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_pp1_26 [13]));
 AND2_X1 u_multiplier_STAGE1__2007_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_pp1_26 [14]));
 AND2_X1 u_multiplier_STAGE1__2008_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_pp1_26 [15]));
 AND2_X1 u_multiplier_STAGE1__2009_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__0739_ ));
 AND2_X1 u_multiplier_STAGE1__2010_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__0740_ ));
 AND2_X1 u_multiplier_STAGE1__2011_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__0741_ ));
 AND2_X1 u_multiplier_STAGE1__2012_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__0742_ ));
 AND2_X1 u_multiplier_STAGE1__2013_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__0743_ ));
 AND2_X1 u_multiplier_STAGE1__2014_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__0744_ ));
 AND2_X1 u_multiplier_STAGE1__2015_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__0745_ ));
 AND2_X1 u_multiplier_STAGE1__2016_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__0746_ ));
 AND2_X1 u_multiplier_STAGE1__2017_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_STAGE1__0747_ ));
 AND2_X1 u_multiplier_STAGE1__2018_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0748_ ));
 AND2_X1 u_multiplier_STAGE1__2019_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0749_ ));
 AND2_X1 u_multiplier_STAGE1__2020_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0750_ ));
 AND2_X1 u_multiplier_STAGE1__2021_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_STAGE1__0751_ ));
 AND2_X1 u_multiplier_STAGE1__2022_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_STAGE1__0752_ ));
 AND2_X1 u_multiplier_STAGE1__2023_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[14]),
    .ZN(u_multiplier_STAGE1__0753_ ));
 AND2_X1 u_multiplier_STAGE1__2024_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_STAGE1__0754_ ));
 AND2_X1 u_multiplier_STAGE1__2025_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0755_ ));
 AND2_X1 u_multiplier_STAGE1__2026_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0756_ ));
 AND2_X1 u_multiplier_STAGE1__2027_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0757_ ));
 AND2_X1 u_multiplier_STAGE1__2028_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_STAGE1__0758_ ));
 AND2_X1 u_multiplier_STAGE1__2029_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__0759_ ));
 AND2_X1 u_multiplier_STAGE1__2030_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__0760_ ));
 AND2_X1 u_multiplier_STAGE1__2031_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__0761_ ));
 AND2_X1 u_multiplier_STAGE1__2032_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__0762_ ));
 AND2_X1 u_multiplier_STAGE1__2033_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_pp1_27 [12]));
 AND2_X1 u_multiplier_STAGE1__2034_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_pp1_27 [13]));
 AND2_X1 u_multiplier_STAGE1__2035_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_pp1_27 [14]));
 AND2_X1 u_multiplier_STAGE1__2036_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_pp1_27 [15]));
 AND2_X1 u_multiplier_STAGE1__2037_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__0763_ ));
 AND2_X1 u_multiplier_STAGE1__2038_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__0764_ ));
 AND2_X1 u_multiplier_STAGE1__2039_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__0765_ ));
 AND2_X1 u_multiplier_STAGE1__2040_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_STAGE1__0766_ ));
 AND2_X1 u_multiplier_STAGE1__2041_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__0767_ ));
 AND2_X1 u_multiplier_STAGE1__2042_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__0768_ ));
 AND2_X1 u_multiplier_STAGE1__2043_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__0769_ ));
 AND2_X1 u_multiplier_STAGE1__2044_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__0770_ ));
 AND2_X1 u_multiplier_STAGE1__2045_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0771_ ));
 AND2_X1 u_multiplier_STAGE1__2046_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0772_ ));
 AND2_X1 u_multiplier_STAGE1__2047_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0773_ ));
 AND2_X1 u_multiplier_STAGE1__2048_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__0774_ ));
 AND2_X1 u_multiplier_STAGE1__2049_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_STAGE1__0775_ ));
 AND2_X1 u_multiplier_STAGE1__2050_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[14]),
    .ZN(u_multiplier_STAGE1__0776_ ));
 AND2_X1 u_multiplier_STAGE1__2051_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_STAGE1__0777_ ));
 AND2_X1 u_multiplier_STAGE1__2052_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_STAGE1__0778_ ));
 AND2_X1 u_multiplier_STAGE1__2053_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0779_ ));
 AND2_X1 u_multiplier_STAGE1__2054_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0780_ ));
 AND2_X1 u_multiplier_STAGE1__2055_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0781_ ));
 AND2_X1 u_multiplier_STAGE1__2056_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_STAGE1__0782_ ));
 AND2_X1 u_multiplier_STAGE1__2057_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__0783_ ));
 AND2_X1 u_multiplier_STAGE1__2058_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__0784_ ));
 AND2_X1 u_multiplier_STAGE1__2059_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__0785_ ));
 AND2_X1 u_multiplier_STAGE1__2060_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__0786_ ));
 AND2_X1 u_multiplier_STAGE1__2061_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__0787_ ));
 AND2_X1 u_multiplier_STAGE1__2062_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__0788_ ));
 AND2_X1 u_multiplier_STAGE1__2063_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_pp1_28 [13]));
 AND2_X1 u_multiplier_STAGE1__2064_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_pp1_28 [14]));
 AND2_X1 u_multiplier_STAGE1__2065_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp1_28 [15]));
 AND2_X1 u_multiplier_STAGE1__2066_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__0789_ ));
 AND2_X1 u_multiplier_STAGE1__2067_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__0790_ ));
 AND2_X1 u_multiplier_STAGE1__2068_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_STAGE1__0791_ ));
 AND2_X1 u_multiplier_STAGE1__2069_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_STAGE1__0792_ ));
 AND2_X1 u_multiplier_STAGE1__2070_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__0793_ ));
 AND2_X1 u_multiplier_STAGE1__2071_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__0794_ ));
 AND2_X1 u_multiplier_STAGE1__2072_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__0795_ ));
 AND2_X1 u_multiplier_STAGE1__2073_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__0796_ ));
 AND2_X1 u_multiplier_STAGE1__2074_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0797_ ));
 AND2_X1 u_multiplier_STAGE1__2075_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0798_ ));
 AND2_X1 u_multiplier_STAGE1__2076_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__0799_ ));
 AND2_X1 u_multiplier_STAGE1__2077_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__0800_ ));
 AND2_X1 u_multiplier_STAGE1__2078_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_STAGE1__0801_ ));
 AND2_X1 u_multiplier_STAGE1__2079_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[15]),
    .ZN(u_multiplier_STAGE1__0802_ ));
 AND2_X1 u_multiplier_STAGE1__2080_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_STAGE1__0803_ ));
 AND2_X1 u_multiplier_STAGE1__2081_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0804_ ));
 AND2_X1 u_multiplier_STAGE1__2082_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0805_ ));
 AND2_X1 u_multiplier_STAGE1__2083_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0806_ ));
 AND2_X1 u_multiplier_STAGE1__2084_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0807_ ));
 AND2_X1 u_multiplier_STAGE1__2085_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_STAGE1__0808_ ));
 AND2_X1 u_multiplier_STAGE1__2086_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__0809_ ));
 AND2_X1 u_multiplier_STAGE1__2087_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__0810_ ));
 AND2_X1 u_multiplier_STAGE1__2088_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__0811_ ));
 AND2_X1 u_multiplier_STAGE1__2089_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__0812_ ));
 AND2_X1 u_multiplier_STAGE1__2090_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__0813_ ));
 AND2_X1 u_multiplier_STAGE1__2091_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__0814_ ));
 AND2_X1 u_multiplier_STAGE1__2092_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__0815_ ));
 AND2_X1 u_multiplier_STAGE1__2093_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__0816_ ));
 AND2_X1 u_multiplier_STAGE1__2094_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp1_29 [14]));
 AND2_X1 u_multiplier_STAGE1__2095_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp1_29 [15]));
 AND2_X1 u_multiplier_STAGE1__2096_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__0817_ ));
 AND2_X1 u_multiplier_STAGE1__2097_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_STAGE1__0818_ ));
 AND2_X1 u_multiplier_STAGE1__2098_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_STAGE1__0819_ ));
 AND2_X1 u_multiplier_STAGE1__2099_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_STAGE1__0820_ ));
 AND2_X1 u_multiplier_STAGE1__2100_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__0821_ ));
 AND2_X1 u_multiplier_STAGE1__2101_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__0822_ ));
 AND2_X1 u_multiplier_STAGE1__2102_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__0823_ ));
 AND2_X1 u_multiplier_STAGE1__2103_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__0824_ ));
 AND2_X1 u_multiplier_STAGE1__2104_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0825_ ));
 AND2_X1 u_multiplier_STAGE1__2105_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__0826_ ));
 AND2_X1 u_multiplier_STAGE1__2106_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__0827_ ));
 AND2_X1 u_multiplier_STAGE1__2107_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__0828_ ));
 AND2_X1 u_multiplier_STAGE1__2108_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[15]),
    .ZN(u_multiplier_STAGE1__0829_ ));
 AND2_X1 u_multiplier_STAGE1__2109_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_STAGE1__0830_ ));
 AND2_X1 u_multiplier_STAGE1__2110_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0831_ ));
 AND2_X1 u_multiplier_STAGE1__2111_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0832_ ));
 AND2_X1 u_multiplier_STAGE1__2112_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0833_ ));
 AND2_X1 u_multiplier_STAGE1__2113_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0834_ ));
 AND2_X1 u_multiplier_STAGE1__2114_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0835_ ));
 AND2_X1 u_multiplier_STAGE1__2115_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_STAGE1__0836_ ));
 AND2_X1 u_multiplier_STAGE1__2116_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__0837_ ));
 AND2_X1 u_multiplier_STAGE1__2117_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__0838_ ));
 AND2_X1 u_multiplier_STAGE1__2118_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__0839_ ));
 AND2_X1 u_multiplier_STAGE1__2119_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__0840_ ));
 AND2_X1 u_multiplier_STAGE1__2120_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__0841_ ));
 AND2_X1 u_multiplier_STAGE1__2121_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__0842_ ));
 AND2_X1 u_multiplier_STAGE1__2122_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__0843_ ));
 AND2_X1 u_multiplier_STAGE1__2123_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__0844_ ));
 AND2_X1 u_multiplier_STAGE1__2124_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_STAGE1__0845_ ));
 AND2_X1 u_multiplier_STAGE1__2125_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_STAGE1__0846_ ));
 AND2_X1 u_multiplier_STAGE1__2126_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp1_30 [15]));
 AND2_X1 u_multiplier_STAGE1__2127_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_STAGE1__0847_ ));
 AND2_X1 u_multiplier_STAGE1__2128_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_STAGE1__0848_ ));
 AND2_X1 u_multiplier_STAGE1__2129_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_STAGE1__0849_ ));
 AND2_X1 u_multiplier_STAGE1__2130_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_STAGE1__0850_ ));
 AND2_X1 u_multiplier_STAGE1__2131_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__0851_ ));
 AND2_X1 u_multiplier_STAGE1__2132_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__0852_ ));
 AND2_X1 u_multiplier_STAGE1__2133_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__0853_ ));
 AND2_X1 u_multiplier_STAGE1__2134_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__0854_ ));
 AND2_X1 u_multiplier_STAGE1__2135_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__0855_ ));
 AND2_X1 u_multiplier_STAGE1__2136_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__0856_ ));
 AND2_X1 u_multiplier_STAGE1__2137_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__0857_ ));
 AND2_X1 u_multiplier_STAGE1__2138_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__0858_ ));
 AND2_X1 u_multiplier_STAGE1__2139_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[16]),
    .ZN(u_multiplier_STAGE1__0859_ ));
 AND2_X1 u_multiplier_STAGE1__2140_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0860_ ));
 AND2_X1 u_multiplier_STAGE1__2141_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0861_ ));
 AND2_X1 u_multiplier_STAGE1__2142_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0862_ ));
 AND2_X1 u_multiplier_STAGE1__2143_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0863_ ));
 AND2_X1 u_multiplier_STAGE1__2144_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0864_ ));
 AND2_X1 u_multiplier_STAGE1__2145_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0865_ ));
 AND2_X1 u_multiplier_STAGE1__2146_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_STAGE1__0866_ ));
 AND2_X1 u_multiplier_STAGE1__2147_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__0867_ ));
 AND2_X1 u_multiplier_STAGE1__2148_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__0868_ ));
 AND2_X1 u_multiplier_STAGE1__2149_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__0869_ ));
 AND2_X1 u_multiplier_STAGE1__2150_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__0870_ ));
 AND2_X1 u_multiplier_STAGE1__2151_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__0871_ ));
 AND2_X1 u_multiplier_STAGE1__2152_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__0872_ ));
 AND2_X1 u_multiplier_STAGE1__2153_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__0873_ ));
 AND2_X1 u_multiplier_STAGE1__2154_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__0874_ ));
 AND2_X1 u_multiplier_STAGE1__2155_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_STAGE1__0875_ ));
 AND2_X1 u_multiplier_STAGE1__2156_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_STAGE1__0876_ ));
 AND2_X1 u_multiplier_STAGE1__2157_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_STAGE1__0877_ ));
 AND2_X1 u_multiplier_STAGE1__2158_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_STAGE1__0878_ ));
 AND2_X1 u_multiplier_STAGE1__2159_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_STAGE1__0879_ ));
 AND2_X1 u_multiplier_STAGE1__2160_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_STAGE1__0880_ ));
 AND2_X1 u_multiplier_STAGE1__2161_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_STAGE1__0881_ ));
 AND2_X1 u_multiplier_STAGE1__2162_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_STAGE1__0882_ ));
 AND2_X1 u_multiplier_STAGE1__2163_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__0883_ ));
 AND2_X1 u_multiplier_STAGE1__2164_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__0884_ ));
 AND2_X1 u_multiplier_STAGE1__2165_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__0885_ ));
 AND2_X1 u_multiplier_STAGE1__2166_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__0886_ ));
 AND2_X1 u_multiplier_STAGE1__2167_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__0887_ ));
 AND2_X1 u_multiplier_STAGE1__2168_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__0888_ ));
 AND2_X1 u_multiplier_STAGE1__2169_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__0889_ ));
 AND2_X1 u_multiplier_STAGE1__2170_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__0890_ ));
 AND2_X1 u_multiplier_STAGE1__2171_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0891_ ));
 AND2_X1 u_multiplier_STAGE1__2172_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0892_ ));
 AND2_X1 u_multiplier_STAGE1__2173_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0893_ ));
 AND2_X1 u_multiplier_STAGE1__2174_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[16]),
    .ZN(u_multiplier_STAGE1__0894_ ));
 AND2_X1 u_multiplier_STAGE1__2175_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0895_ ));
 AND2_X1 u_multiplier_STAGE1__2176_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0896_ ));
 AND2_X1 u_multiplier_STAGE1__2177_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0897_ ));
 AND2_X1 u_multiplier_STAGE1__2178_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__0898_ ));
 AND2_X1 u_multiplier_STAGE1__2179_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__0899_ ));
 AND2_X1 u_multiplier_STAGE1__2180_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__0900_ ));
 AND2_X1 u_multiplier_STAGE1__2181_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__0901_ ));
 AND2_X1 u_multiplier_STAGE1__2182_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__0902_ ));
 AND2_X1 u_multiplier_STAGE1__2183_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__0903_ ));
 AND2_X1 u_multiplier_STAGE1__2184_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__0904_ ));
 AND2_X1 u_multiplier_STAGE1__2185_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__0905_ ));
 AND2_X1 u_multiplier_STAGE1__2186_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_STAGE1__0906_ ));
 AND2_X1 u_multiplier_STAGE1__2187_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_STAGE1__0907_ ));
 AND2_X1 u_multiplier_STAGE1__2188_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_STAGE1__0908_ ));
 AND2_X1 u_multiplier_STAGE1__2189_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_STAGE1__0909_ ));
 AND2_X1 u_multiplier_STAGE1__2190_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_STAGE1__0910_ ));
 AND2_X1 u_multiplier_STAGE1__2191_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_STAGE1__0911_ ));
 AND2_X1 u_multiplier_STAGE1__2192_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_STAGE1__0912_ ));
 AND2_X1 u_multiplier_STAGE1__2193_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_STAGE1__0913_ ));
 AND2_X1 u_multiplier_STAGE1__2194_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__0914_ ));
 AND2_X1 u_multiplier_STAGE1__2195_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__0915_ ));
 AND2_X1 u_multiplier_STAGE1__2196_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__0916_ ));
 AND2_X1 u_multiplier_STAGE1__2197_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__0917_ ));
 AND2_X1 u_multiplier_STAGE1__2198_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__0918_ ));
 AND2_X1 u_multiplier_STAGE1__2199_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__0919_ ));
 AND2_X1 u_multiplier_STAGE1__2200_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__0920_ ));
 AND2_X1 u_multiplier_STAGE1__2201_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__0921_ ));
 AND2_X1 u_multiplier_STAGE1__2202_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0922_ ));
 AND2_X1 u_multiplier_STAGE1__2203_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0923_ ));
 AND2_X1 u_multiplier_STAGE1__2204_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0924_ ));
 AND2_X1 u_multiplier_STAGE1__2205_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[17]),
    .ZN(u_multiplier_STAGE1__0925_ ));
 AND2_X1 u_multiplier_STAGE1__2206_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0926_ ));
 AND2_X1 u_multiplier_STAGE1__2207_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0927_ ));
 AND2_X1 u_multiplier_STAGE1__2208_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__0928_ ));
 AND2_X1 u_multiplier_STAGE1__2209_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__0929_ ));
 AND2_X1 u_multiplier_STAGE1__2210_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__0930_ ));
 AND2_X1 u_multiplier_STAGE1__2211_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__0931_ ));
 AND2_X1 u_multiplier_STAGE1__2212_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__0932_ ));
 AND2_X1 u_multiplier_STAGE1__2213_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__0933_ ));
 AND2_X1 u_multiplier_STAGE1__2214_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__0934_ ));
 AND2_X1 u_multiplier_STAGE1__2215_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__0935_ ));
 AND2_X1 u_multiplier_STAGE1__2216_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_STAGE1__0936_ ));
 AND2_X1 u_multiplier_STAGE1__2217_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_STAGE1__0937_ ));
 AND2_X1 u_multiplier_STAGE1__2218_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_STAGE1__0938_ ));
 AND2_X1 u_multiplier_STAGE1__2219_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_STAGE1__0939_ ));
 AND2_X1 u_multiplier_STAGE1__2220_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_STAGE1__0940_ ));
 AND2_X1 u_multiplier_STAGE1__2221_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_STAGE1__0941_ ));
 AND2_X1 u_multiplier_STAGE1__2222_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_STAGE1__0942_ ));
 AND2_X1 u_multiplier_STAGE1__2223_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__0943_ ));
 AND2_X1 u_multiplier_STAGE1__2224_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__0944_ ));
 AND2_X1 u_multiplier_STAGE1__2225_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__0945_ ));
 AND2_X1 u_multiplier_STAGE1__2226_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__0946_ ));
 AND2_X1 u_multiplier_STAGE1__2227_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__0947_ ));
 AND2_X1 u_multiplier_STAGE1__2228_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__0948_ ));
 AND2_X1 u_multiplier_STAGE1__2229_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__0949_ ));
 AND2_X1 u_multiplier_STAGE1__2230_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__0950_ ));
 AND2_X1 u_multiplier_STAGE1__2231_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0951_ ));
 AND2_X1 u_multiplier_STAGE1__2232_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0952_ ));
 AND2_X1 u_multiplier_STAGE1__2233_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[17]),
    .ZN(u_multiplier_STAGE1__0953_ ));
 AND2_X1 u_multiplier_STAGE1__2234_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0954_ ));
 AND2_X1 u_multiplier_STAGE1__2235_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0955_ ));
 AND2_X1 u_multiplier_STAGE1__2236_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__0956_ ));
 AND2_X1 u_multiplier_STAGE1__2237_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__0957_ ));
 AND2_X1 u_multiplier_STAGE1__2238_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__0958_ ));
 AND2_X1 u_multiplier_STAGE1__2239_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__0959_ ));
 AND2_X1 u_multiplier_STAGE1__2240_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__0960_ ));
 AND2_X1 u_multiplier_STAGE1__2241_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__0961_ ));
 AND2_X1 u_multiplier_STAGE1__2242_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__0962_ ));
 AND2_X1 u_multiplier_STAGE1__2243_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__0963_ ));
 AND2_X1 u_multiplier_STAGE1__2244_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_STAGE1__0964_ ));
 AND2_X1 u_multiplier_STAGE1__2245_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_STAGE1__0965_ ));
 AND2_X1 u_multiplier_STAGE1__2246_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_STAGE1__0966_ ));
 AND2_X1 u_multiplier_STAGE1__2247_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_STAGE1__0967_ ));
 AND2_X1 u_multiplier_STAGE1__2248_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp1_34 [15]));
 AND2_X1 u_multiplier_STAGE1__2249_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_STAGE1__0968_ ));
 AND2_X1 u_multiplier_STAGE1__2250_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_STAGE1__0969_ ));
 AND2_X1 u_multiplier_STAGE1__2251_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__0970_ ));
 AND2_X1 u_multiplier_STAGE1__2252_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__0971_ ));
 AND2_X1 u_multiplier_STAGE1__2253_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__0972_ ));
 AND2_X1 u_multiplier_STAGE1__2254_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__0973_ ));
 AND2_X1 u_multiplier_STAGE1__2255_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__0974_ ));
 AND2_X1 u_multiplier_STAGE1__2256_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__0975_ ));
 AND2_X1 u_multiplier_STAGE1__2257_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__0976_ ));
 AND2_X1 u_multiplier_STAGE1__2258_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__0977_ ));
 AND2_X1 u_multiplier_STAGE1__2259_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__0978_ ));
 AND2_X1 u_multiplier_STAGE1__2260_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__0979_ ));
 AND2_X1 u_multiplier_STAGE1__2261_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[18]),
    .ZN(u_multiplier_STAGE1__0980_ ));
 AND2_X1 u_multiplier_STAGE1__2262_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__0981_ ));
 AND2_X1 u_multiplier_STAGE1__2263_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__0982_ ));
 AND2_X1 u_multiplier_STAGE1__2264_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__0983_ ));
 AND2_X1 u_multiplier_STAGE1__2265_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__0984_ ));
 AND2_X1 u_multiplier_STAGE1__2266_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__0985_ ));
 AND2_X1 u_multiplier_STAGE1__2267_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__0986_ ));
 AND2_X1 u_multiplier_STAGE1__2268_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__0987_ ));
 AND2_X1 u_multiplier_STAGE1__2269_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__0988_ ));
 AND2_X1 u_multiplier_STAGE1__2270_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__0989_ ));
 AND2_X1 u_multiplier_STAGE1__2271_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_STAGE1__0990_ ));
 AND2_X1 u_multiplier_STAGE1__2272_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_STAGE1__0991_ ));
 AND2_X2 u_multiplier_STAGE1__2273_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_STAGE1__0992_ ));
 AND2_X2 u_multiplier_STAGE1__2274_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_STAGE1__0993_ ));
 AND2_X1 u_multiplier_STAGE1__2275_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp1_35 [14]));
 AND2_X1 u_multiplier_STAGE1__2276_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp1_35 [15]));
 AND2_X1 u_multiplier_STAGE1__2277_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_STAGE1__0994_ ));
 AND2_X1 u_multiplier_STAGE1__2278_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__0995_ ));
 AND2_X1 u_multiplier_STAGE1__2279_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__0996_ ));
 AND2_X1 u_multiplier_STAGE1__2280_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__0997_ ));
 AND2_X1 u_multiplier_STAGE1__2281_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__0998_ ));
 AND2_X1 u_multiplier_STAGE1__2282_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__0999_ ));
 AND2_X1 u_multiplier_STAGE1__2283_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__1000_ ));
 AND2_X1 u_multiplier_STAGE1__2284_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__1001_ ));
 AND2_X1 u_multiplier_STAGE1__2285_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__1002_ ));
 AND2_X1 u_multiplier_STAGE1__2286_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__1003_ ));
 AND2_X1 u_multiplier_STAGE1__2287_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[18]),
    .ZN(u_multiplier_STAGE1__1004_ ));
 AND2_X1 u_multiplier_STAGE1__2288_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__1005_ ));
 AND2_X1 u_multiplier_STAGE1__2289_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__1006_ ));
 AND2_X1 u_multiplier_STAGE1__2290_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__1007_ ));
 AND2_X1 u_multiplier_STAGE1__2291_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__1008_ ));
 AND2_X1 u_multiplier_STAGE1__2292_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__1009_ ));
 AND2_X1 u_multiplier_STAGE1__2293_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__1010_ ));
 AND2_X1 u_multiplier_STAGE1__2294_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__1011_ ));
 AND2_X1 u_multiplier_STAGE1__2295_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__1012_ ));
 AND2_X1 u_multiplier_STAGE1__2296_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__1013_ ));
 AND2_X1 u_multiplier_STAGE1__2297_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_STAGE1__1014_ ));
 AND2_X1 u_multiplier_STAGE1__2298_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_STAGE1__1015_ ));
 AND2_X1 u_multiplier_STAGE1__2299_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_STAGE1__1016_ ));
 AND2_X1 u_multiplier_STAGE1__2300_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_STAGE1__1017_ ));
 AND2_X1 u_multiplier_STAGE1__2301_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp1_36 [13]));
 AND2_X1 u_multiplier_STAGE1__2302_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp1_36 [14]));
 AND2_X1 u_multiplier_STAGE1__2303_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp1_36 [15]));
 AND2_X1 u_multiplier_STAGE1__2304_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_STAGE1__1018_ ));
 AND2_X1 u_multiplier_STAGE1__2305_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__1019_ ));
 AND2_X1 u_multiplier_STAGE1__2306_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__1020_ ));
 AND2_X1 u_multiplier_STAGE1__2307_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__1021_ ));
 AND2_X1 u_multiplier_STAGE1__2308_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__1022_ ));
 AND2_X1 u_multiplier_STAGE1__2309_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__1023_ ));
 AND2_X1 u_multiplier_STAGE1__2310_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__1024_ ));
 AND2_X1 u_multiplier_STAGE1__2311_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__1025_ ));
 AND2_X1 u_multiplier_STAGE1__2312_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__1026_ ));
 AND2_X1 u_multiplier_STAGE1__2313_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[19]),
    .ZN(u_multiplier_STAGE1__1027_ ));
 AND2_X1 u_multiplier_STAGE1__2314_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__1028_ ));
 AND2_X1 u_multiplier_STAGE1__2315_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__1029_ ));
 AND2_X1 u_multiplier_STAGE1__2316_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__1030_ ));
 AND2_X1 u_multiplier_STAGE1__2317_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__1031_ ));
 AND2_X1 u_multiplier_STAGE1__2318_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__1032_ ));
 AND2_X1 u_multiplier_STAGE1__2319_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__1033_ ));
 AND2_X1 u_multiplier_STAGE1__2320_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__1034_ ));
 AND2_X1 u_multiplier_STAGE1__2321_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__1035_ ));
 AND2_X1 u_multiplier_STAGE1__2322_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_STAGE1__1036_ ));
 AND2_X1 u_multiplier_STAGE1__2323_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_STAGE1__1037_ ));
 AND2_X1 u_multiplier_STAGE1__2324_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_STAGE1__1038_ ));
 AND2_X1 u_multiplier_STAGE1__2325_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_STAGE1__1039_ ));
 AND2_X1 u_multiplier_STAGE1__2326_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp1_37 [12]));
 AND2_X1 u_multiplier_STAGE1__2327_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp1_37 [13]));
 AND2_X1 u_multiplier_STAGE1__2328_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp1_37 [14]));
 AND2_X1 u_multiplier_STAGE1__2329_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp1_37 [15]));
 AND2_X1 u_multiplier_STAGE1__2330_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_STAGE1__1040_ ));
 AND2_X1 u_multiplier_STAGE1__2331_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__1041_ ));
 AND2_X1 u_multiplier_STAGE1__2332_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__1042_ ));
 AND2_X1 u_multiplier_STAGE1__2333_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__1043_ ));
 AND2_X1 u_multiplier_STAGE1__2334_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__1044_ ));
 AND2_X1 u_multiplier_STAGE1__2335_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__1045_ ));
 AND2_X1 u_multiplier_STAGE1__2336_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__1046_ ));
 AND2_X1 u_multiplier_STAGE1__2337_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[19]),
    .ZN(u_multiplier_STAGE1__1047_ ));
 AND2_X1 u_multiplier_STAGE1__2338_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__1048_ ));
 AND2_X1 u_multiplier_STAGE1__2339_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__1049_ ));
 AND2_X1 u_multiplier_STAGE1__2340_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__1050_ ));
 AND2_X1 u_multiplier_STAGE1__2341_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__1051_ ));
 AND2_X1 u_multiplier_STAGE1__2342_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__1052_ ));
 AND2_X1 u_multiplier_STAGE1__2343_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__1053_ ));
 AND2_X1 u_multiplier_STAGE1__2344_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__1054_ ));
 AND2_X1 u_multiplier_STAGE1__2345_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__1055_ ));
 AND2_X1 u_multiplier_STAGE1__2346_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_STAGE1__1056_ ));
 AND2_X1 u_multiplier_STAGE1__2347_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_STAGE1__1057_ ));
 AND2_X1 u_multiplier_STAGE1__2348_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_STAGE1__1058_ ));
 AND2_X1 u_multiplier_STAGE1__2349_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_STAGE1__1059_ ));
 AND2_X1 u_multiplier_STAGE1__2350_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_pp1_38 [11]));
 AND2_X1 u_multiplier_STAGE1__2351_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp1_38 [12]));
 AND2_X1 u_multiplier_STAGE1__2352_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp1_38 [13]));
 AND2_X1 u_multiplier_STAGE1__2353_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp1_38 [14]));
 AND2_X1 u_multiplier_STAGE1__2354_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp1_38 [15]));
 AND2_X1 u_multiplier_STAGE1__2355_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_STAGE1__1060_ ));
 AND2_X1 u_multiplier_STAGE1__2356_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__1061_ ));
 AND2_X1 u_multiplier_STAGE1__2357_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__1062_ ));
 AND2_X1 u_multiplier_STAGE1__2358_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__1063_ ));
 AND2_X1 u_multiplier_STAGE1__2359_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__1064_ ));
 AND2_X1 u_multiplier_STAGE1__2360_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__1065_ ));
 AND2_X1 u_multiplier_STAGE1__2361_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[20]),
    .ZN(u_multiplier_STAGE1__1066_ ));
 AND2_X1 u_multiplier_STAGE1__2362_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__1067_ ));
 AND2_X1 u_multiplier_STAGE1__2363_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__1068_ ));
 AND2_X1 u_multiplier_STAGE1__2364_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__1069_ ));
 AND2_X1 u_multiplier_STAGE1__2365_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__1070_ ));
 AND2_X1 u_multiplier_STAGE1__2366_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__1071_ ));
 AND2_X1 u_multiplier_STAGE1__2367_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__1072_ ));
 AND2_X1 u_multiplier_STAGE1__2368_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__1073_ ));
 AND2_X1 u_multiplier_STAGE1__2369_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_STAGE1__1074_ ));
 AND2_X1 u_multiplier_STAGE1__2370_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_STAGE1__1075_ ));
 AND2_X1 u_multiplier_STAGE1__2371_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_STAGE1__1076_ ));
 AND2_X1 u_multiplier_STAGE1__2372_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_STAGE1__1077_ ));
 AND2_X1 u_multiplier_STAGE1__2373_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_pp1_39 [10]));
 AND2_X1 u_multiplier_STAGE1__2374_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_pp1_39 [11]));
 AND2_X1 u_multiplier_STAGE1__2375_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp1_39 [12]));
 AND2_X1 u_multiplier_STAGE1__2376_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp1_39 [13]));
 AND2_X1 u_multiplier_STAGE1__2377_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp1_39 [14]));
 AND2_X1 u_multiplier_STAGE1__2378_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp1_39 [15]));
 AND2_X1 u_multiplier_STAGE1__2379_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_STAGE1__1078_ ));
 AND2_X1 u_multiplier_STAGE1__2380_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__1079_ ));
 AND2_X1 u_multiplier_STAGE1__2381_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__1080_ ));
 AND2_X1 u_multiplier_STAGE1__2382_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__1081_ ));
 AND2_X1 u_multiplier_STAGE1__2383_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[20]),
    .ZN(u_multiplier_STAGE1__1082_ ));
 AND2_X1 u_multiplier_STAGE1__2384_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__1083_ ));
 AND2_X1 u_multiplier_STAGE1__2385_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__1084_ ));
 AND2_X1 u_multiplier_STAGE1__2386_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__1085_ ));
 AND2_X1 u_multiplier_STAGE1__2387_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__1086_ ));
 AND2_X1 u_multiplier_STAGE1__2388_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__1087_ ));
 AND2_X1 u_multiplier_STAGE1__2389_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__1088_ ));
 AND2_X1 u_multiplier_STAGE1__2390_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__1089_ ));
 AND2_X1 u_multiplier_STAGE1__2391_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_STAGE1__1090_ ));
 AND2_X1 u_multiplier_STAGE1__2392_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_STAGE1__1091_ ));
 AND2_X1 u_multiplier_STAGE1__2393_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_STAGE1__1092_ ));
 AND2_X1 u_multiplier_STAGE1__2394_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_STAGE1__1093_ ));
 AND2_X1 u_multiplier_STAGE1__2395_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_pp1_40 [9]));
 AND2_X1 u_multiplier_STAGE1__2396_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_pp1_40 [10]));
 AND2_X1 u_multiplier_STAGE1__2397_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_pp1_40 [11]));
 AND2_X1 u_multiplier_STAGE1__2398_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp1_40 [12]));
 AND2_X1 u_multiplier_STAGE1__2399_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp1_40 [13]));
 AND2_X1 u_multiplier_STAGE1__2400_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp1_40 [14]));
 AND2_X1 u_multiplier_STAGE1__2401_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp1_40 [15]));
 AND2_X1 u_multiplier_STAGE1__2402_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_STAGE1__1094_ ));
 AND2_X1 u_multiplier_STAGE1__2403_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__1095_ ));
 AND2_X1 u_multiplier_STAGE1__2404_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__1096_ ));
 AND2_X1 u_multiplier_STAGE1__2405_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[21]),
    .ZN(u_multiplier_STAGE1__1097_ ));
 AND2_X1 u_multiplier_STAGE1__2406_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__1098_ ));
 AND2_X1 u_multiplier_STAGE1__2407_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__1099_ ));
 AND2_X1 u_multiplier_STAGE1__2408_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__1100_ ));
 AND2_X1 u_multiplier_STAGE1__2409_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__1101_ ));
 AND2_X1 u_multiplier_STAGE1__2410_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__1102_ ));
 AND2_X1 u_multiplier_STAGE1__2411_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__1103_ ));
 AND2_X1 u_multiplier_STAGE1__2412_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_STAGE1__1104_ ));
 AND2_X1 u_multiplier_STAGE1__2413_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_STAGE1__1105_ ));
 AND2_X1 u_multiplier_STAGE1__2414_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_STAGE1__1106_ ));
 AND2_X1 u_multiplier_STAGE1__2415_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_STAGE1__1107_ ));
 AND2_X1 u_multiplier_STAGE1__2416_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_pp1_41 [8]));
 AND2_X1 u_multiplier_STAGE1__2417_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_pp1_41 [9]));
 AND2_X1 u_multiplier_STAGE1__2418_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_pp1_41 [10]));
 AND2_X1 u_multiplier_STAGE1__2419_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_pp1_41 [11]));
 AND2_X1 u_multiplier_STAGE1__2420_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp1_41 [12]));
 AND2_X1 u_multiplier_STAGE1__2421_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp1_41 [13]));
 AND2_X1 u_multiplier_STAGE1__2422_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp1_41 [14]));
 AND2_X1 u_multiplier_STAGE1__2423_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp1_41 [15]));
 AND2_X1 u_multiplier_STAGE1__2424_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_STAGE1__1108_ ));
 AND2_X1 u_multiplier_STAGE1__2425_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[21]),
    .ZN(u_multiplier_STAGE1__1109_ ));
 AND2_X1 u_multiplier_STAGE1__2426_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__1110_ ));
 AND2_X1 u_multiplier_STAGE1__2427_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__1111_ ));
 AND2_X1 u_multiplier_STAGE1__2428_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__1112_ ));
 AND2_X1 u_multiplier_STAGE1__2429_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__1113_ ));
 AND2_X1 u_multiplier_STAGE1__2430_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__1114_ ));
 AND2_X1 u_multiplier_STAGE1__2431_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__1115_ ));
 AND2_X1 u_multiplier_STAGE1__2432_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_STAGE1__1116_ ));
 AND2_X1 u_multiplier_STAGE1__2433_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_STAGE1__1117_ ));
 AND2_X1 u_multiplier_STAGE1__2434_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_STAGE1__1118_ ));
 AND2_X1 u_multiplier_STAGE1__2435_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_STAGE1__1119_ ));
 AND2_X1 u_multiplier_STAGE1__2436_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_pp1_42 [7]));
 AND2_X1 u_multiplier_STAGE1__2437_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_pp1_42 [8]));
 AND2_X1 u_multiplier_STAGE1__2438_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_pp1_42 [9]));
 AND2_X1 u_multiplier_STAGE1__2439_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_pp1_42 [10]));
 AND2_X1 u_multiplier_STAGE1__2440_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_pp1_42 [11]));
 AND2_X1 u_multiplier_STAGE1__2441_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp1_42 [12]));
 AND2_X1 u_multiplier_STAGE1__2442_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp1_42 [13]));
 AND2_X1 u_multiplier_STAGE1__2443_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp1_42 [14]));
 AND2_X1 u_multiplier_STAGE1__2444_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp1_42 [15]));
 AND2_X1 u_multiplier_STAGE1__2445_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[22]),
    .ZN(u_multiplier_STAGE1__1120_ ));
 AND2_X1 u_multiplier_STAGE1__2446_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_STAGE1__1121_ ));
 AND2_X1 u_multiplier_STAGE1__2447_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__1122_ ));
 AND2_X1 u_multiplier_STAGE1__2448_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__1123_ ));
 AND2_X1 u_multiplier_STAGE1__2449_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__1124_ ));
 AND2_X1 u_multiplier_STAGE1__2450_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__1125_ ));
 AND2_X1 u_multiplier_STAGE1__2451_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_STAGE1__1126_ ));
 AND2_X1 u_multiplier_STAGE1__2452_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_STAGE1__1127_ ));
 AND2_X2 u_multiplier_STAGE1__2453_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_STAGE1__1128_ ));
 AND2_X2 u_multiplier_STAGE1__2454_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_STAGE1__1129_ ));
 AND2_X1 u_multiplier_STAGE1__2455_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_pp1_43 [6]));
 AND2_X1 u_multiplier_STAGE1__2456_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_pp1_43 [7]));
 AND2_X1 u_multiplier_STAGE1__2457_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_pp1_43 [8]));
 AND2_X1 u_multiplier_STAGE1__2458_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_pp1_43 [9]));
 AND2_X1 u_multiplier_STAGE1__2459_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_pp1_43 [10]));
 AND2_X1 u_multiplier_STAGE1__2460_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_pp1_43 [11]));
 AND2_X1 u_multiplier_STAGE1__2461_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp1_43 [12]));
 AND2_X1 u_multiplier_STAGE1__2462_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp1_43 [13]));
 AND2_X1 u_multiplier_STAGE1__2463_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp1_43 [14]));
 AND2_X1 u_multiplier_STAGE1__2464_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp1_43 [15]));
 AND2_X1 u_multiplier_STAGE1__2465_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_STAGE1__1130_ ));
 AND2_X1 u_multiplier_STAGE1__2466_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_STAGE1__1131_ ));
 AND2_X1 u_multiplier_STAGE1__2467_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__1132_ ));
 AND2_X1 u_multiplier_STAGE1__2468_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__1133_ ));
 AND2_X1 u_multiplier_STAGE1__2469_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_STAGE1__1134_ ));
 AND2_X1 u_multiplier_STAGE1__2470_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_STAGE1__1135_ ));
 AND2_X1 u_multiplier_STAGE1__2471_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_STAGE1__1136_ ));
 AND2_X1 u_multiplier_STAGE1__2472_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_STAGE1__1137_ ));
 AND2_X1 u_multiplier_STAGE1__2473_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_pp1_44 [5]));
 AND2_X1 u_multiplier_STAGE1__2474_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[22]),
    .ZN(u_multiplier_pp1_44 [6]));
 AND2_X1 u_multiplier_STAGE1__2475_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_pp1_44 [7]));
 AND2_X1 u_multiplier_STAGE1__2476_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_pp1_44 [8]));
 AND2_X1 u_multiplier_STAGE1__2477_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_pp1_44 [9]));
 AND2_X1 u_multiplier_STAGE1__2478_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_pp1_44 [10]));
 AND2_X1 u_multiplier_STAGE1__2479_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_pp1_44 [11]));
 AND2_X1 u_multiplier_STAGE1__2480_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp1_44 [12]));
 AND2_X1 u_multiplier_STAGE1__2481_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp1_44 [13]));
 AND2_X1 u_multiplier_STAGE1__2482_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp1_44 [14]));
 AND2_X1 u_multiplier_STAGE1__2483_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp1_44 [15]));
 AND2_X1 u_multiplier_STAGE1__2484_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_STAGE1__1138_ ));
 AND2_X1 u_multiplier_STAGE1__2485_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_STAGE1__1139_ ));
 AND2_X1 u_multiplier_STAGE1__2486_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_STAGE1__1140_ ));
 AND2_X1 u_multiplier_STAGE1__2487_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_STAGE1__1141_ ));
 AND2_X1 u_multiplier_STAGE1__2488_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_STAGE1__1142_ ));
 AND2_X1 u_multiplier_STAGE1__2489_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_STAGE1__1143_ ));
 AND2_X1 u_multiplier_STAGE1__2490_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_pp1_45 [4]));
 AND2_X1 u_multiplier_STAGE1__2491_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_pp1_45 [5]));
 AND2_X1 u_multiplier_STAGE1__2492_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[23]),
    .ZN(u_multiplier_pp1_45 [6]));
 AND2_X1 u_multiplier_STAGE1__2493_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_pp1_45 [7]));
 AND2_X1 u_multiplier_STAGE1__2494_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_pp1_45 [8]));
 AND2_X1 u_multiplier_STAGE1__2495_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_pp1_45 [9]));
 AND2_X1 u_multiplier_STAGE1__2496_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_pp1_45 [10]));
 AND2_X1 u_multiplier_STAGE1__2497_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_pp1_45 [11]));
 AND2_X1 u_multiplier_STAGE1__2498_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp1_45 [12]));
 AND2_X1 u_multiplier_STAGE1__2499_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp1_45 [13]));
 AND2_X1 u_multiplier_STAGE1__2500_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp1_45 [14]));
 AND2_X1 u_multiplier_STAGE1__2501_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp1_45 [15]));
 AND2_X1 u_multiplier_STAGE1__2502_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_STAGE1__1144_ ));
 AND2_X1 u_multiplier_STAGE1__2503_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_STAGE1__1145_ ));
 AND2_X1 u_multiplier_STAGE1__2504_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_STAGE1__1146_ ));
 AND2_X1 u_multiplier_STAGE1__2505_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_STAGE1__1147_ ));
 AND2_X1 u_multiplier_STAGE1__2506_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_pp1_46 [3]));
 AND2_X1 u_multiplier_STAGE1__2507_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_pp1_46 [4]));
 AND2_X1 u_multiplier_STAGE1__2508_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_pp1_46 [5]));
 AND2_X1 u_multiplier_STAGE1__2509_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_pp1_46 [6]));
 AND2_X1 u_multiplier_STAGE1__2510_  (.A1(data_in_reg[23]),
    .A2(sram_rdata_reg[23]),
    .ZN(u_multiplier_pp1_46 [7]));
 AND2_X1 u_multiplier_STAGE1__2511_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_pp1_46 [8]));
 AND2_X1 u_multiplier_STAGE1__2512_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_pp1_46 [9]));
 AND2_X1 u_multiplier_STAGE1__2513_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_pp1_46 [10]));
 AND2_X1 u_multiplier_STAGE1__2514_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_pp1_46 [11]));
 AND2_X1 u_multiplier_STAGE1__2515_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp1_46 [12]));
 AND2_X1 u_multiplier_STAGE1__2516_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp1_46 [13]));
 AND2_X1 u_multiplier_STAGE1__2517_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp1_46 [14]));
 AND2_X1 u_multiplier_STAGE1__2518_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp1_46 [15]));
 AND2_X1 u_multiplier_STAGE1__2519_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_STAGE1__1148_ ));
 AND2_X1 u_multiplier_STAGE1__2520_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_STAGE1__1149_ ));
 AND2_X1 u_multiplier_STAGE1__2521_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_47 [2]));
 AND2_X1 u_multiplier_STAGE1__2522_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_47 [3]));
 AND2_X1 u_multiplier_STAGE1__2523_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_47 [4]));
 AND2_X1 u_multiplier_STAGE1__2524_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_47 [5]));
 AND2_X1 u_multiplier_STAGE1__2525_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_pp1_47 [6]));
 AND2_X1 u_multiplier_STAGE1__2526_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_pp1_47 [7]));
 AND2_X1 u_multiplier_STAGE1__2527_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_pp1_47 [8]));
 AND2_X1 u_multiplier_STAGE1__2528_  (.A1(sram_rdata_reg[23]),
    .A2(data_in_reg[24]),
    .ZN(u_multiplier_pp1_47 [9]));
 AND2_X1 u_multiplier_STAGE1__2529_  (.A1(data_in_reg[23]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_pp1_47 [10]));
 AND2_X1 u_multiplier_STAGE1__2530_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_pp1_47 [11]));
 AND2_X1 u_multiplier_STAGE1__2531_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_pp1_47 [12]));
 AND2_X1 u_multiplier_STAGE1__2532_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_pp1_47 [13]));
 AND2_X1 u_multiplier_STAGE1__2533_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp1_47 [14]));
 AND2_X1 u_multiplier_STAGE1__2534_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp1_47 [15]));
 AND2_X1 u_multiplier_STAGE1__2535_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_48 [1]));
 AND2_X1 u_multiplier_STAGE1__2536_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_48 [2]));
 AND2_X1 u_multiplier_STAGE1__2537_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_48 [3]));
 AND2_X1 u_multiplier_STAGE1__2538_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_48 [4]));
 AND2_X1 u_multiplier_STAGE1__2539_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_pp1_48 [5]));
 AND2_X1 u_multiplier_STAGE1__2540_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_pp1_48 [6]));
 AND2_X1 u_multiplier_STAGE1__2541_  (.A1(sram_rdata_reg[23]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_pp1_48 [7]));
 AND2_X1 u_multiplier_STAGE1__2542_  (.A1(data_in_reg[24]),
    .A2(sram_rdata_reg[24]),
    .ZN(u_multiplier_pp1_48 [8]));
 AND2_X1 u_multiplier_STAGE1__2543_  (.A1(data_in_reg[23]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_pp1_48 [9]));
 AND2_X1 u_multiplier_STAGE1__2544_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_pp1_48 [10]));
 AND2_X1 u_multiplier_STAGE1__2545_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_pp1_48 [11]));
 AND2_X1 u_multiplier_STAGE1__2546_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp1_48 [12]));
 AND2_X1 u_multiplier_STAGE1__2547_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp1_48 [13]));
 AND2_X1 u_multiplier_STAGE1__2548_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp1_48 [14]));
 AND2_X1 u_multiplier_STAGE1__2549_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp1_48 [15]));
 AND2_X1 u_multiplier_STAGE1__2550_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_49 [0]));
 AND2_X1 u_multiplier_STAGE1__2551_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_49 [1]));
 AND2_X1 u_multiplier_STAGE1__2552_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_49 [2]));
 AND2_X1 u_multiplier_STAGE1__2553_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_49 [3]));
 AND2_X1 u_multiplier_STAGE1__2554_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_pp1_49 [4]));
 AND2_X1 u_multiplier_STAGE1__2555_  (.A1(sram_rdata_reg[23]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_pp1_49 [5]));
 AND2_X1 u_multiplier_STAGE1__2556_  (.A1(sram_rdata_reg[24]),
    .A2(data_in_reg[25]),
    .ZN(u_multiplier_pp1_49 [6]));
 AND2_X1 u_multiplier_STAGE1__2557_  (.A1(data_in_reg[24]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_pp1_49 [7]));
 AND2_X1 u_multiplier_STAGE1__2558_  (.A1(data_in_reg[23]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_pp1_49 [8]));
 AND2_X1 u_multiplier_STAGE1__2559_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_pp1_49 [9]));
 AND2_X1 u_multiplier_STAGE1__2560_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp1_49 [10]));
 AND2_X1 u_multiplier_STAGE1__2561_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp1_49 [11]));
 AND2_X1 u_multiplier_STAGE1__2562_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp1_49 [12]));
 AND2_X1 u_multiplier_STAGE1__2563_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp1_49 [13]));
 AND2_X1 u_multiplier_STAGE1__2564_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_50 [0]));
 AND2_X1 u_multiplier_STAGE1__2565_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_50 [1]));
 AND2_X1 u_multiplier_STAGE1__2566_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_50 [2]));
 AND2_X1 u_multiplier_STAGE1__2567_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_50 [3]));
 AND2_X1 u_multiplier_STAGE1__2568_  (.A1(sram_rdata_reg[23]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_pp1_50 [4]));
 AND2_X1 u_multiplier_STAGE1__2569_  (.A1(sram_rdata_reg[24]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_pp1_50 [5]));
 AND2_X1 u_multiplier_STAGE1__2570_  (.A1(data_in_reg[25]),
    .A2(sram_rdata_reg[25]),
    .ZN(u_multiplier_pp1_50 [6]));
 AND2_X1 u_multiplier_STAGE1__2571_  (.A1(data_in_reg[24]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_pp1_50 [7]));
 AND2_X1 u_multiplier_STAGE1__2572_  (.A1(data_in_reg[23]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_pp1_50 [8]));
 AND2_X1 u_multiplier_STAGE1__2573_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp1_50 [9]));
 AND2_X1 u_multiplier_STAGE1__2574_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp1_50 [10]));
 AND2_X1 u_multiplier_STAGE1__2575_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp1_50 [11]));
 AND2_X1 u_multiplier_STAGE1__2576_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp2_50 [7]));
 AND2_X1 u_multiplier_STAGE1__2577_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_51 [0]));
 AND2_X1 u_multiplier_STAGE1__2578_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_51 [1]));
 AND2_X1 u_multiplier_STAGE1__2579_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_51 [2]));
 AND2_X1 u_multiplier_STAGE1__2580_  (.A1(sram_rdata_reg[23]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_51 [3]));
 AND2_X1 u_multiplier_STAGE1__2581_  (.A1(sram_rdata_reg[24]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_pp1_51 [4]));
 AND2_X1 u_multiplier_STAGE1__2582_  (.A1(sram_rdata_reg[25]),
    .A2(data_in_reg[26]),
    .ZN(u_multiplier_pp1_51 [5]));
 AND2_X1 u_multiplier_STAGE1__2583_  (.A1(data_in_reg[25]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_pp1_51 [6]));
 AND2_X1 u_multiplier_STAGE1__2584_  (.A1(data_in_reg[24]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_pp1_51 [7]));
 AND2_X1 u_multiplier_STAGE1__2585_  (.A1(data_in_reg[23]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp1_51 [8]));
 AND2_X1 u_multiplier_STAGE1__2586_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp1_51 [9]));
 AND2_X1 u_multiplier_STAGE1__2587_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp2_51 [7]));
 AND2_X1 u_multiplier_STAGE1__2588_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp2_51 [6]));
 AND2_X1 u_multiplier_STAGE1__2589_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_52 [0]));
 AND2_X1 u_multiplier_STAGE1__2590_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_52 [1]));
 AND2_X1 u_multiplier_STAGE1__2591_  (.A1(sram_rdata_reg[23]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_52 [2]));
 AND2_X1 u_multiplier_STAGE1__2592_  (.A1(sram_rdata_reg[24]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_52 [3]));
 AND2_X1 u_multiplier_STAGE1__2593_  (.A1(sram_rdata_reg[25]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_pp1_52 [4]));
 AND2_X1 u_multiplier_STAGE1__2594_  (.A1(data_in_reg[26]),
    .A2(sram_rdata_reg[26]),
    .ZN(u_multiplier_pp1_52 [5]));
 AND2_X1 u_multiplier_STAGE1__2595_  (.A1(data_in_reg[25]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_pp1_52 [6]));
 AND2_X1 u_multiplier_STAGE1__2596_  (.A1(data_in_reg[24]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp1_52 [7]));
 AND2_X1 u_multiplier_STAGE1__2597_  (.A1(data_in_reg[23]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp2_52 [7]));
 AND2_X1 u_multiplier_STAGE1__2598_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp2_52 [6]));
 AND2_X1 u_multiplier_STAGE1__2599_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp2_52 [5]));
 AND2_X1 u_multiplier_STAGE1__2600_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_53 [0]));
 AND2_X1 u_multiplier_STAGE1__2601_  (.A1(sram_rdata_reg[23]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_53 [1]));
 AND2_X1 u_multiplier_STAGE1__2602_  (.A1(sram_rdata_reg[24]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_53 [2]));
 AND2_X1 u_multiplier_STAGE1__2603_  (.A1(sram_rdata_reg[25]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_53 [3]));
 AND2_X1 u_multiplier_STAGE1__2604_  (.A1(sram_rdata_reg[26]),
    .A2(data_in_reg[27]),
    .ZN(u_multiplier_pp1_53 [4]));
 AND2_X1 u_multiplier_STAGE1__2605_  (.A1(data_in_reg[26]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_pp1_53 [5]));
 AND2_X1 u_multiplier_STAGE1__2606_  (.A1(data_in_reg[25]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp2_53 [7]));
 AND2_X1 u_multiplier_STAGE1__2607_  (.A1(data_in_reg[24]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp2_53 [6]));
 AND2_X1 u_multiplier_STAGE1__2608_  (.A1(data_in_reg[23]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp2_53 [5]));
 AND2_X1 u_multiplier_STAGE1__2609_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp2_53 [4]));
 AND2_X1 u_multiplier_STAGE1__2610_  (.A1(sram_rdata_reg[23]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_54 [0]));
 AND2_X1 u_multiplier_STAGE1__2611_  (.A1(sram_rdata_reg[24]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_54 [1]));
 AND2_X1 u_multiplier_STAGE1__2612_  (.A1(sram_rdata_reg[25]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp1_54 [2]));
 AND2_X1 u_multiplier_STAGE1__2613_  (.A1(sram_rdata_reg[26]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp1_54 [3]));
 AND2_X1 u_multiplier_STAGE1__2614_  (.A1(data_in_reg[27]),
    .A2(sram_rdata_reg[27]),
    .ZN(u_multiplier_pp2_54 [7]));
 AND2_X1 u_multiplier_STAGE1__2615_  (.A1(data_in_reg[26]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp2_54 [6]));
 AND2_X1 u_multiplier_STAGE1__2616_  (.A1(data_in_reg[25]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp2_54 [5]));
 AND2_X1 u_multiplier_STAGE1__2617_  (.A1(data_in_reg[24]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp2_54 [4]));
 AND2_X1 u_multiplier_STAGE1__2618_  (.A1(data_in_reg[23]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp2_54 [3]));
 AND2_X1 u_multiplier_STAGE1__2619_  (.A1(sram_rdata_reg[24]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp1_55 [0]));
 AND2_X1 u_multiplier_STAGE1__2620_  (.A1(sram_rdata_reg[25]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp1_55 [1]));
 AND2_X1 u_multiplier_STAGE1__2621_  (.A1(sram_rdata_reg[26]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp2_55 [7]));
 AND2_X1 u_multiplier_STAGE1__2622_  (.A1(sram_rdata_reg[27]),
    .A2(data_in_reg[28]),
    .ZN(u_multiplier_pp2_55 [6]));
 AND2_X1 u_multiplier_STAGE1__2623_  (.A1(data_in_reg[27]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp2_55 [5]));
 AND2_X1 u_multiplier_STAGE1__2624_  (.A1(data_in_reg[26]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp2_55 [4]));
 AND2_X1 u_multiplier_STAGE1__2625_  (.A1(data_in_reg[25]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp2_55 [3]));
 AND2_X1 u_multiplier_STAGE1__2626_  (.A1(data_in_reg[24]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp2_55 [2]));
 AND2_X1 u_multiplier_STAGE1__2627_  (.A1(sram_rdata_reg[25]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp2_56 [7]));
 AND2_X1 u_multiplier_STAGE1__2628_  (.A1(sram_rdata_reg[26]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp2_56 [6]));
 AND2_X1 u_multiplier_STAGE1__2629_  (.A1(sram_rdata_reg[27]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp2_56 [5]));
 AND2_X1 u_multiplier_STAGE1__2630_  (.A1(data_in_reg[28]),
    .A2(sram_rdata_reg[28]),
    .ZN(u_multiplier_pp2_56 [4]));
 AND2_X1 u_multiplier_STAGE1__2631_  (.A1(data_in_reg[27]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp2_56 [3]));
 AND2_X1 u_multiplier_STAGE1__2632_  (.A1(data_in_reg[26]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp2_56 [2]));
 AND2_X1 u_multiplier_STAGE1__2633_  (.A1(data_in_reg[25]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp2_56 [1]));
 AND2_X1 u_multiplier_STAGE1__2634_  (.A1(sram_rdata_reg[26]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp2_57 [5]));
 AND2_X1 u_multiplier_STAGE1__2635_  (.A1(sram_rdata_reg[27]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp2_57 [4]));
 AND2_X1 u_multiplier_STAGE1__2636_  (.A1(sram_rdata_reg[28]),
    .A2(data_in_reg[29]),
    .ZN(u_multiplier_pp2_57 [3]));
 AND2_X1 u_multiplier_STAGE1__2637_  (.A1(data_in_reg[28]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp2_57 [2]));
 AND2_X1 u_multiplier_STAGE1__2638_  (.A1(data_in_reg[27]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp2_57 [1]));
 AND2_X1 u_multiplier_STAGE1__2639_  (.A1(data_in_reg[26]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp2_57 [0]));
 AND2_X1 u_multiplier_STAGE1__2640_  (.A1(sram_rdata_reg[27]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp3_58 [3]));
 AND2_X1 u_multiplier_STAGE1__2641_  (.A1(sram_rdata_reg[28]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp2_58 [3]));
 AND2_X1 u_multiplier_STAGE1__2642_  (.A1(data_in_reg[29]),
    .A2(sram_rdata_reg[29]),
    .ZN(u_multiplier_pp2_58 [2]));
 AND2_X1 u_multiplier_STAGE1__2643_  (.A1(data_in_reg[28]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp2_58 [1]));
 AND2_X1 u_multiplier_STAGE1__2644_  (.A1(data_in_reg[27]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp2_58 [0]));
 AND2_X1 u_multiplier_STAGE1__2645_  (.A1(sram_rdata_reg[28]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp3_59 [2]));
 AND2_X1 u_multiplier_STAGE1__2646_  (.A1(sram_rdata_reg[29]),
    .A2(data_in_reg[30]),
    .ZN(u_multiplier_pp3_59 [3]));
 AND2_X1 u_multiplier_STAGE1__2647_  (.A1(data_in_reg[29]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp2_59 [1]));
 AND2_X1 u_multiplier_STAGE1__2648_  (.A1(data_in_reg[28]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp2_59 [0]));
 AND2_X1 u_multiplier_STAGE1__2649_  (.A1(sram_rdata_reg[29]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp3_60 [1]));
 AND2_X1 u_multiplier_STAGE1__2650_  (.A1(data_in_reg[30]),
    .A2(sram_rdata_reg[30]),
    .ZN(u_multiplier_pp3_60 [2]));
 AND2_X1 u_multiplier_STAGE1__2651_  (.A1(data_in_reg[29]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp3_60 [3]));
 AND2_X1 u_multiplier_STAGE1__2652_  (.A1(sram_rdata_reg[30]),
    .A2(data_in_reg[31]),
    .ZN(u_multiplier_pp3_61 [0]));
 AND2_X1 u_multiplier_STAGE1__2653_  (.A1(data_in_reg[30]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp3_61 [1]));
 AND2_X1 u_multiplier_STAGE1__2654_  (.A1(data_in_reg[31]),
    .A2(sram_rdata_reg[31]),
    .ZN(u_multiplier_pp3_62 ));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_17_0__21_  (.A1(u_multiplier_STAGE1__0610_ ),
    .A2(u_multiplier_STAGE1__0609_ ),
    .A3(u_multiplier_STAGE1__0611_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_17_0__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_17_0__22_  (.A(u_multiplier_STAGE1__0610_ ),
    .B(u_multiplier_STAGE1__0609_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_17_0__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_17_0__23_  (.A(u_multiplier_STAGE1__0611_ ),
    .B(u_multiplier_STAGE1__0612_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_17_0__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_17_0__24_  (.A1(u_multiplier_STAGE1_acci1_pp_17_0__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_17_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_17_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_17_0__25_  (.A(u_multiplier_STAGE1_acci1_pp_17_0__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_17_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_17_0__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_17_0__26_  (.A1(u_multiplier_STAGE1_acci1_pp_17_0__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_17_0__16_ ),
    .ZN(u_multiplier_pp1_17 [0]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_17_0__27_  (.A1(u_multiplier_STAGE1__0610_ ),
    .A2(u_multiplier_STAGE1__0609_ ),
    .B1(u_multiplier_STAGE1__0611_ ),
    .B2(u_multiplier_STAGE1__0612_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_17_0__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_17_0__28_  (.A1(u_multiplier_STAGE1_acci1_pp_17_0__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_17_0__17_ ),
    .ZN(u_multiplier_pp1_18 [2]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_18_0__21_  (.A1(u_multiplier_STAGE1__0614_ ),
    .A2(u_multiplier_STAGE1__0613_ ),
    .A3(u_multiplier_STAGE1__0615_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_18_0__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_18_0__22_  (.A(u_multiplier_STAGE1__0614_ ),
    .B(u_multiplier_STAGE1__0613_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_18_0__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_18_0__23_  (.A(u_multiplier_STAGE1__0615_ ),
    .B(u_multiplier_STAGE1__0616_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_18_0__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_18_0__24_  (.A1(u_multiplier_STAGE1_acci1_pp_18_0__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_18_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_18_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_18_0__25_  (.A(u_multiplier_STAGE1_acci1_pp_18_0__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_18_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_18_0__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_18_0__26_  (.A1(u_multiplier_STAGE1_acci1_pp_18_0__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_18_0__16_ ),
    .ZN(u_multiplier_pp1_18 [0]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_18_0__27_  (.A1(u_multiplier_STAGE1__0614_ ),
    .A2(u_multiplier_STAGE1__0613_ ),
    .B1(u_multiplier_STAGE1__0615_ ),
    .B2(u_multiplier_STAGE1__0616_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_18_0__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_18_0__28_  (.A1(u_multiplier_STAGE1_acci1_pp_18_0__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_18_0__17_ ),
    .ZN(u_multiplier_pp1_19 [3]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_19_0__21_  (.A1(u_multiplier_STAGE1__0620_ ),
    .A2(u_multiplier_STAGE1__0619_ ),
    .A3(u_multiplier_STAGE1__0621_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_19_0__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_19_0__22_  (.A(u_multiplier_STAGE1__0620_ ),
    .B(u_multiplier_STAGE1__0619_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_19_0__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_19_0__23_  (.A(u_multiplier_STAGE1__0621_ ),
    .B(u_multiplier_STAGE1__0622_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_19_0__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_19_0__24_  (.A1(u_multiplier_STAGE1_acci1_pp_19_0__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_19_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_19_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_19_0__25_  (.A(u_multiplier_STAGE1_acci1_pp_19_0__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_19_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_19_0__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_19_0__26_  (.A1(u_multiplier_STAGE1_acci1_pp_19_0__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_19_0__16_ ),
    .ZN(u_multiplier_pp1_19 [0]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_19_0__27_  (.A1(u_multiplier_STAGE1__0620_ ),
    .A2(u_multiplier_STAGE1__0619_ ),
    .B1(u_multiplier_STAGE1__0621_ ),
    .B2(u_multiplier_STAGE1__0622_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_19_0__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_19_0__28_  (.A1(u_multiplier_STAGE1_acci1_pp_19_0__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_19_0__17_ ),
    .ZN(u_multiplier_pp1_20 [4]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_19_1__21_  (.A1(u_multiplier_STAGE1__0624_ ),
    .A2(u_multiplier_STAGE1__0623_ ),
    .A3(u_multiplier_STAGE1__0625_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_19_1__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_19_1__22_  (.A(u_multiplier_STAGE1__0624_ ),
    .B(u_multiplier_STAGE1__0623_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_19_1__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_19_1__23_  (.A(u_multiplier_STAGE1__0625_ ),
    .B(u_multiplier_STAGE1__0626_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_19_1__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_19_1__24_  (.A1(u_multiplier_STAGE1_acci1_pp_19_1__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_19_1__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_19_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_19_1__25_  (.A(u_multiplier_STAGE1_acci1_pp_19_1__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_19_1__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_19_1__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_19_1__26_  (.A1(u_multiplier_STAGE1_acci1_pp_19_1__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_19_1__16_ ),
    .ZN(u_multiplier_pp1_19 [1]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_19_1__27_  (.A1(u_multiplier_STAGE1__0624_ ),
    .A2(u_multiplier_STAGE1__0623_ ),
    .B1(u_multiplier_STAGE1__0625_ ),
    .B2(u_multiplier_STAGE1__0626_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_19_1__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_19_1__28_  (.A1(u_multiplier_STAGE1_acci1_pp_19_1__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_19_1__17_ ),
    .ZN(u_multiplier_pp1_20 [3]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_20_0__21_  (.A1(u_multiplier_STAGE1__0628_ ),
    .A2(u_multiplier_STAGE1__0627_ ),
    .A3(u_multiplier_STAGE1__0629_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_20_0__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_20_0__22_  (.A(u_multiplier_STAGE1__0628_ ),
    .B(u_multiplier_STAGE1__0627_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_20_0__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_20_0__23_  (.A(u_multiplier_STAGE1__0629_ ),
    .B(u_multiplier_STAGE1__0630_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_20_0__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_20_0__24_  (.A1(u_multiplier_STAGE1_acci1_pp_20_0__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_20_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_20_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_20_0__25_  (.A(u_multiplier_STAGE1_acci1_pp_20_0__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_20_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_20_0__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_20_0__26_  (.A1(u_multiplier_STAGE1_acci1_pp_20_0__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_20_0__16_ ),
    .ZN(u_multiplier_pp1_20 [0]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_20_0__27_  (.A1(u_multiplier_STAGE1__0628_ ),
    .A2(u_multiplier_STAGE1__0627_ ),
    .B1(u_multiplier_STAGE1__0629_ ),
    .B2(u_multiplier_STAGE1__0630_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_20_0__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_20_0__28_  (.A1(u_multiplier_STAGE1_acci1_pp_20_0__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_20_0__17_ ),
    .ZN(u_multiplier_pp1_21 [5]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_20_1__21_  (.A1(u_multiplier_STAGE1__0632_ ),
    .A2(u_multiplier_STAGE1__0631_ ),
    .A3(u_multiplier_STAGE1__0633_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_20_1__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_20_1__22_  (.A(u_multiplier_STAGE1__0632_ ),
    .B(u_multiplier_STAGE1__0631_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_20_1__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_20_1__23_  (.A(u_multiplier_STAGE1__0633_ ),
    .B(u_multiplier_STAGE1__0634_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_20_1__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_20_1__24_  (.A1(u_multiplier_STAGE1_acci1_pp_20_1__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_20_1__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_20_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_20_1__25_  (.A(u_multiplier_STAGE1_acci1_pp_20_1__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_20_1__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_20_1__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_20_1__26_  (.A1(u_multiplier_STAGE1_acci1_pp_20_1__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_20_1__16_ ),
    .ZN(u_multiplier_pp1_20 [1]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_20_1__27_  (.A1(u_multiplier_STAGE1__0632_ ),
    .A2(u_multiplier_STAGE1__0631_ ),
    .B1(u_multiplier_STAGE1__0633_ ),
    .B2(u_multiplier_STAGE1__0634_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_20_1__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_20_1__28_  (.A1(u_multiplier_STAGE1_acci1_pp_20_1__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_20_1__17_ ),
    .ZN(u_multiplier_pp1_21 [4]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_21_0__21_  (.A1(u_multiplier_STAGE1__0638_ ),
    .A2(u_multiplier_STAGE1__0637_ ),
    .A3(u_multiplier_STAGE1__0639_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_21_0__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_21_0__22_  (.A(u_multiplier_STAGE1__0638_ ),
    .B(u_multiplier_STAGE1__0637_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_21_0__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_21_0__23_  (.A(u_multiplier_STAGE1__0639_ ),
    .B(u_multiplier_STAGE1__0640_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_21_0__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_21_0__24_  (.A1(u_multiplier_STAGE1_acci1_pp_21_0__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_21_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_21_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_21_0__25_  (.A(u_multiplier_STAGE1_acci1_pp_21_0__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_21_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_21_0__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_21_0__26_  (.A1(u_multiplier_STAGE1_acci1_pp_21_0__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_21_0__16_ ),
    .ZN(u_multiplier_pp1_21 [0]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_21_0__27_  (.A1(u_multiplier_STAGE1__0638_ ),
    .A2(u_multiplier_STAGE1__0637_ ),
    .B1(u_multiplier_STAGE1__0639_ ),
    .B2(u_multiplier_STAGE1__0640_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_21_0__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_21_0__28_  (.A1(u_multiplier_STAGE1_acci1_pp_21_0__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_21_0__17_ ),
    .ZN(u_multiplier_pp1_22 [6]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_21_1__21_  (.A1(u_multiplier_STAGE1__0642_ ),
    .A2(u_multiplier_STAGE1__0641_ ),
    .A3(u_multiplier_STAGE1__0643_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_21_1__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_21_1__22_  (.A(u_multiplier_STAGE1__0642_ ),
    .B(u_multiplier_STAGE1__0641_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_21_1__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_21_1__23_  (.A(u_multiplier_STAGE1__0643_ ),
    .B(u_multiplier_STAGE1__0644_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_21_1__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_21_1__24_  (.A1(u_multiplier_STAGE1_acci1_pp_21_1__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_21_1__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_21_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_21_1__25_  (.A(u_multiplier_STAGE1_acci1_pp_21_1__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_21_1__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_21_1__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_21_1__26_  (.A1(u_multiplier_STAGE1_acci1_pp_21_1__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_21_1__16_ ),
    .ZN(u_multiplier_pp1_21 [1]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_21_1__27_  (.A1(u_multiplier_STAGE1__0642_ ),
    .A2(u_multiplier_STAGE1__0641_ ),
    .B1(u_multiplier_STAGE1__0643_ ),
    .B2(u_multiplier_STAGE1__0644_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_21_1__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_21_1__28_  (.A1(u_multiplier_STAGE1_acci1_pp_21_1__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_21_1__17_ ),
    .ZN(u_multiplier_pp1_22 [5]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_21_2__21_  (.A1(u_multiplier_STAGE1__0646_ ),
    .A2(u_multiplier_STAGE1__0645_ ),
    .A3(u_multiplier_STAGE1__0647_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_21_2__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_21_2__22_  (.A(u_multiplier_STAGE1__0646_ ),
    .B(u_multiplier_STAGE1__0645_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_21_2__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_21_2__23_  (.A(u_multiplier_STAGE1__0647_ ),
    .B(u_multiplier_STAGE1__0648_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_21_2__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_21_2__24_  (.A1(u_multiplier_STAGE1_acci1_pp_21_2__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_21_2__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_21_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_21_2__25_  (.A(u_multiplier_STAGE1_acci1_pp_21_2__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_21_2__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_21_2__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_21_2__26_  (.A1(u_multiplier_STAGE1_acci1_pp_21_2__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_21_2__16_ ),
    .ZN(u_multiplier_pp1_21 [2]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_21_2__27_  (.A1(u_multiplier_STAGE1__0646_ ),
    .A2(u_multiplier_STAGE1__0645_ ),
    .B1(u_multiplier_STAGE1__0647_ ),
    .B2(u_multiplier_STAGE1__0648_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_21_2__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_21_2__28_  (.A1(u_multiplier_STAGE1_acci1_pp_21_2__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_21_2__17_ ),
    .ZN(u_multiplier_pp1_22 [4]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_22_0__21_  (.A1(u_multiplier_STAGE1__0650_ ),
    .A2(u_multiplier_STAGE1__0649_ ),
    .A3(u_multiplier_STAGE1__0651_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_22_0__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_22_0__22_  (.A(u_multiplier_STAGE1__0650_ ),
    .B(u_multiplier_STAGE1__0649_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_22_0__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_22_0__23_  (.A(u_multiplier_STAGE1__0651_ ),
    .B(u_multiplier_STAGE1__0652_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_22_0__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_22_0__24_  (.A1(u_multiplier_STAGE1_acci1_pp_22_0__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_22_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_22_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_22_0__25_  (.A(u_multiplier_STAGE1_acci1_pp_22_0__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_22_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_22_0__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_22_0__26_  (.A1(u_multiplier_STAGE1_acci1_pp_22_0__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_22_0__16_ ),
    .ZN(u_multiplier_pp1_22 [0]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_22_0__27_  (.A1(u_multiplier_STAGE1__0650_ ),
    .A2(u_multiplier_STAGE1__0649_ ),
    .B1(u_multiplier_STAGE1__0651_ ),
    .B2(u_multiplier_STAGE1__0652_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_22_0__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_22_0__28_  (.A1(u_multiplier_STAGE1_acci1_pp_22_0__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_22_0__17_ ),
    .ZN(u_multiplier_pp1_23 [7]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_22_1__21_  (.A1(u_multiplier_STAGE1__0654_ ),
    .A2(u_multiplier_STAGE1__0653_ ),
    .A3(u_multiplier_STAGE1__0655_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_22_1__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_22_1__22_  (.A(u_multiplier_STAGE1__0654_ ),
    .B(u_multiplier_STAGE1__0653_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_22_1__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_22_1__23_  (.A(u_multiplier_STAGE1__0655_ ),
    .B(u_multiplier_STAGE1__0656_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_22_1__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_22_1__24_  (.A1(u_multiplier_STAGE1_acci1_pp_22_1__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_22_1__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_22_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_22_1__25_  (.A(u_multiplier_STAGE1_acci1_pp_22_1__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_22_1__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_22_1__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_22_1__26_  (.A1(u_multiplier_STAGE1_acci1_pp_22_1__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_22_1__16_ ),
    .ZN(u_multiplier_pp1_22 [1]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_22_1__27_  (.A1(u_multiplier_STAGE1__0654_ ),
    .A2(u_multiplier_STAGE1__0653_ ),
    .B1(u_multiplier_STAGE1__0655_ ),
    .B2(u_multiplier_STAGE1__0656_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_22_1__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_22_1__28_  (.A1(u_multiplier_STAGE1_acci1_pp_22_1__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_22_1__17_ ),
    .ZN(u_multiplier_pp1_23 [6]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_22_2__21_  (.A1(u_multiplier_STAGE1__0658_ ),
    .A2(u_multiplier_STAGE1__0657_ ),
    .A3(u_multiplier_STAGE1__0659_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_22_2__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_22_2__22_  (.A(u_multiplier_STAGE1__0658_ ),
    .B(u_multiplier_STAGE1__0657_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_22_2__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_22_2__23_  (.A(u_multiplier_STAGE1__0659_ ),
    .B(u_multiplier_STAGE1__0660_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_22_2__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_22_2__24_  (.A1(u_multiplier_STAGE1_acci1_pp_22_2__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_22_2__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_22_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_22_2__25_  (.A(u_multiplier_STAGE1_acci1_pp_22_2__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_22_2__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_22_2__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_22_2__26_  (.A1(u_multiplier_STAGE1_acci1_pp_22_2__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_22_2__16_ ),
    .ZN(u_multiplier_pp1_22 [2]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_22_2__27_  (.A1(u_multiplier_STAGE1__0658_ ),
    .A2(u_multiplier_STAGE1__0657_ ),
    .B1(u_multiplier_STAGE1__0659_ ),
    .B2(u_multiplier_STAGE1__0660_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_22_2__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_22_2__28_  (.A1(u_multiplier_STAGE1_acci1_pp_22_2__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_22_2__17_ ),
    .ZN(u_multiplier_pp1_23 [5]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_23_0__21_  (.A1(u_multiplier_STAGE1__0664_ ),
    .A2(u_multiplier_STAGE1__0663_ ),
    .A3(u_multiplier_STAGE1__0665_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_23_0__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_23_0__22_  (.A(u_multiplier_STAGE1__0664_ ),
    .B(u_multiplier_STAGE1__0663_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_23_0__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_23_0__23_  (.A(u_multiplier_STAGE1__0665_ ),
    .B(u_multiplier_STAGE1__0666_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_23_0__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_23_0__24_  (.A1(u_multiplier_STAGE1_acci1_pp_23_0__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_23_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_23_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_23_0__25_  (.A(u_multiplier_STAGE1_acci1_pp_23_0__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_23_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_23_0__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_23_0__26_  (.A1(u_multiplier_STAGE1_acci1_pp_23_0__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_23_0__16_ ),
    .ZN(u_multiplier_pp1_23 [0]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_23_0__27_  (.A1(u_multiplier_STAGE1__0664_ ),
    .A2(u_multiplier_STAGE1__0663_ ),
    .B1(u_multiplier_STAGE1__0665_ ),
    .B2(u_multiplier_STAGE1__0666_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_23_0__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_23_0__28_  (.A1(u_multiplier_STAGE1_acci1_pp_23_0__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_23_0__17_ ),
    .ZN(u_multiplier_pp1_24 [8]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_23_1__21_  (.A1(u_multiplier_STAGE1__0668_ ),
    .A2(u_multiplier_STAGE1__0667_ ),
    .A3(u_multiplier_STAGE1__0669_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_23_1__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_23_1__22_  (.A(u_multiplier_STAGE1__0668_ ),
    .B(u_multiplier_STAGE1__0667_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_23_1__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_23_1__23_  (.A(u_multiplier_STAGE1__0669_ ),
    .B(u_multiplier_STAGE1__0670_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_23_1__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_23_1__24_  (.A1(u_multiplier_STAGE1_acci1_pp_23_1__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_23_1__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_23_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_23_1__25_  (.A(u_multiplier_STAGE1_acci1_pp_23_1__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_23_1__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_23_1__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_23_1__26_  (.A1(u_multiplier_STAGE1_acci1_pp_23_1__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_23_1__16_ ),
    .ZN(u_multiplier_pp1_23 [1]));
 AOI22_X1 u_multiplier_STAGE1_acci1_pp_23_1__27_  (.A1(u_multiplier_STAGE1__0668_ ),
    .A2(u_multiplier_STAGE1__0667_ ),
    .B1(u_multiplier_STAGE1__0669_ ),
    .B2(u_multiplier_STAGE1__0670_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_23_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_23_1__28_  (.A1(u_multiplier_STAGE1_acci1_pp_23_1__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_23_1__17_ ),
    .ZN(u_multiplier_pp1_24 [7]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_23_2__21_  (.A1(u_multiplier_STAGE1__0672_ ),
    .A2(u_multiplier_STAGE1__0671_ ),
    .A3(u_multiplier_STAGE1__0673_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_23_2__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_23_2__22_  (.A(u_multiplier_STAGE1__0672_ ),
    .B(u_multiplier_STAGE1__0671_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_23_2__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_23_2__23_  (.A(u_multiplier_STAGE1__0673_ ),
    .B(u_multiplier_STAGE1__0674_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_23_2__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_23_2__24_  (.A1(u_multiplier_STAGE1_acci1_pp_23_2__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_23_2__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_23_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_23_2__25_  (.A(u_multiplier_STAGE1_acci1_pp_23_2__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_23_2__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_23_2__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_23_2__26_  (.A1(u_multiplier_STAGE1_acci1_pp_23_2__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_23_2__16_ ),
    .ZN(u_multiplier_pp1_23 [2]));
 AOI22_X1 u_multiplier_STAGE1_acci1_pp_23_2__27_  (.A1(u_multiplier_STAGE1__0672_ ),
    .A2(u_multiplier_STAGE1__0671_ ),
    .B1(u_multiplier_STAGE1__0673_ ),
    .B2(u_multiplier_STAGE1__0674_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_23_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_23_2__28_  (.A1(u_multiplier_STAGE1_acci1_pp_23_2__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_23_2__17_ ),
    .ZN(u_multiplier_pp1_24 [6]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_23_3__21_  (.A1(u_multiplier_STAGE1__0676_ ),
    .A2(u_multiplier_STAGE1__0675_ ),
    .A3(u_multiplier_STAGE1__0677_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_23_3__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_23_3__22_  (.A(u_multiplier_STAGE1__0676_ ),
    .B(u_multiplier_STAGE1__0675_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_23_3__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_23_3__23_  (.A(u_multiplier_STAGE1__0677_ ),
    .B(u_multiplier_STAGE1__0678_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_23_3__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_23_3__24_  (.A1(u_multiplier_STAGE1_acci1_pp_23_3__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_23_3__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_23_3__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_23_3__25_  (.A(u_multiplier_STAGE1_acci1_pp_23_3__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_23_3__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_23_3__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_23_3__26_  (.A1(u_multiplier_STAGE1_acci1_pp_23_3__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_23_3__16_ ),
    .ZN(u_multiplier_pp1_23 [3]));
 AOI22_X1 u_multiplier_STAGE1_acci1_pp_23_3__27_  (.A1(u_multiplier_STAGE1__0676_ ),
    .A2(u_multiplier_STAGE1__0675_ ),
    .B1(u_multiplier_STAGE1__0677_ ),
    .B2(u_multiplier_STAGE1__0678_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_23_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_23_3__28_  (.A1(u_multiplier_STAGE1_acci1_pp_23_3__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_23_3__17_ ),
    .ZN(u_multiplier_pp1_24 [5]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_24_0__21_  (.A1(u_multiplier_STAGE1__0680_ ),
    .A2(u_multiplier_STAGE1__0679_ ),
    .A3(u_multiplier_STAGE1__0681_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_24_0__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_24_0__22_  (.A(u_multiplier_STAGE1__0680_ ),
    .B(u_multiplier_STAGE1__0679_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_24_0__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_24_0__23_  (.A(u_multiplier_STAGE1__0681_ ),
    .B(u_multiplier_STAGE1__0682_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_24_0__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_24_0__24_  (.A1(u_multiplier_STAGE1_acci1_pp_24_0__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_24_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_24_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_24_0__25_  (.A(u_multiplier_STAGE1_acci1_pp_24_0__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_24_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_24_0__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_24_0__26_  (.A1(u_multiplier_STAGE1_acci1_pp_24_0__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_24_0__16_ ),
    .ZN(u_multiplier_pp1_24 [0]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_24_0__27_  (.A1(u_multiplier_STAGE1__0680_ ),
    .A2(u_multiplier_STAGE1__0679_ ),
    .B1(u_multiplier_STAGE1__0681_ ),
    .B2(u_multiplier_STAGE1__0682_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_24_0__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_24_0__28_  (.A1(u_multiplier_STAGE1_acci1_pp_24_0__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_24_0__17_ ),
    .ZN(u_multiplier_pp1_25 [9]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_24_1__21_  (.A1(u_multiplier_STAGE1__0684_ ),
    .A2(u_multiplier_STAGE1__0683_ ),
    .A3(u_multiplier_STAGE1__0685_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_24_1__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_24_1__22_  (.A(u_multiplier_STAGE1__0684_ ),
    .B(u_multiplier_STAGE1__0683_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_24_1__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_24_1__23_  (.A(u_multiplier_STAGE1__0685_ ),
    .B(u_multiplier_STAGE1__0686_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_24_1__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_24_1__24_  (.A1(u_multiplier_STAGE1_acci1_pp_24_1__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_24_1__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_24_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_24_1__25_  (.A(u_multiplier_STAGE1_acci1_pp_24_1__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_24_1__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_24_1__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_24_1__26_  (.A1(u_multiplier_STAGE1_acci1_pp_24_1__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_24_1__16_ ),
    .ZN(u_multiplier_pp1_24 [1]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_24_1__27_  (.A1(u_multiplier_STAGE1__0684_ ),
    .A2(u_multiplier_STAGE1__0683_ ),
    .B1(u_multiplier_STAGE1__0685_ ),
    .B2(u_multiplier_STAGE1__0686_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_24_1__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_24_1__28_  (.A1(u_multiplier_STAGE1_acci1_pp_24_1__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_24_1__17_ ),
    .ZN(u_multiplier_pp1_25 [8]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_24_2__21_  (.A1(u_multiplier_STAGE1__0688_ ),
    .A2(u_multiplier_STAGE1__0687_ ),
    .A3(u_multiplier_STAGE1__0689_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_24_2__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_24_2__22_  (.A(u_multiplier_STAGE1__0688_ ),
    .B(u_multiplier_STAGE1__0687_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_24_2__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_24_2__23_  (.A(u_multiplier_STAGE1__0689_ ),
    .B(u_multiplier_STAGE1__0690_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_24_2__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_24_2__24_  (.A1(u_multiplier_STAGE1_acci1_pp_24_2__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_24_2__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_24_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_24_2__25_  (.A(u_multiplier_STAGE1_acci1_pp_24_2__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_24_2__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_24_2__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_24_2__26_  (.A1(u_multiplier_STAGE1_acci1_pp_24_2__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_24_2__16_ ),
    .ZN(u_multiplier_pp1_24 [2]));
 AOI22_X1 u_multiplier_STAGE1_acci1_pp_24_2__27_  (.A1(u_multiplier_STAGE1__0688_ ),
    .A2(u_multiplier_STAGE1__0687_ ),
    .B1(u_multiplier_STAGE1__0689_ ),
    .B2(u_multiplier_STAGE1__0690_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_24_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_24_2__28_  (.A1(u_multiplier_STAGE1_acci1_pp_24_2__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_24_2__17_ ),
    .ZN(u_multiplier_pp1_25 [7]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_24_3__21_  (.A1(u_multiplier_STAGE1__0692_ ),
    .A2(u_multiplier_STAGE1__0691_ ),
    .A3(u_multiplier_STAGE1__0693_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_24_3__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_24_3__22_  (.A(u_multiplier_STAGE1__0692_ ),
    .B(u_multiplier_STAGE1__0691_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_24_3__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_24_3__23_  (.A(u_multiplier_STAGE1__0693_ ),
    .B(u_multiplier_STAGE1__0694_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_24_3__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_24_3__24_  (.A1(u_multiplier_STAGE1_acci1_pp_24_3__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_24_3__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_24_3__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_24_3__25_  (.A(u_multiplier_STAGE1_acci1_pp_24_3__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_24_3__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_24_3__16_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_24_3__26_  (.A1(u_multiplier_STAGE1_acci1_pp_24_3__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_24_3__16_ ),
    .ZN(u_multiplier_pp1_24 [3]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_24_3__27_  (.A1(u_multiplier_STAGE1__0692_ ),
    .A2(u_multiplier_STAGE1__0691_ ),
    .B1(u_multiplier_STAGE1__0693_ ),
    .B2(u_multiplier_STAGE1__0694_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_24_3__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_24_3__28_  (.A1(u_multiplier_STAGE1_acci1_pp_24_3__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_24_3__17_ ),
    .ZN(u_multiplier_pp1_25 [6]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_25_0__21_  (.A1(u_multiplier_STAGE1__0698_ ),
    .A2(u_multiplier_STAGE1__0697_ ),
    .A3(u_multiplier_STAGE1__0699_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_25_0__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_25_0__22_  (.A(u_multiplier_STAGE1__0698_ ),
    .B(u_multiplier_STAGE1__0697_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_25_0__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_25_0__23_  (.A(u_multiplier_STAGE1__0699_ ),
    .B(u_multiplier_STAGE1__0700_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_25_0__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_25_0__24_  (.A1(u_multiplier_STAGE1_acci1_pp_25_0__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_25_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_25_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_25_0__25_  (.A(u_multiplier_STAGE1_acci1_pp_25_0__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_25_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_25_0__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_25_0__26_  (.A1(u_multiplier_STAGE1_acci1_pp_25_0__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_25_0__16_ ),
    .ZN(u_multiplier_pp1_25 [0]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_25_0__27_  (.A1(u_multiplier_STAGE1__0698_ ),
    .A2(u_multiplier_STAGE1__0697_ ),
    .B1(u_multiplier_STAGE1__0699_ ),
    .B2(u_multiplier_STAGE1__0700_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_25_0__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_25_0__28_  (.A1(u_multiplier_STAGE1_acci1_pp_25_0__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_25_0__17_ ),
    .ZN(u_multiplier_pp1_26 [10]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_25_1__21_  (.A1(u_multiplier_STAGE1__0702_ ),
    .A2(u_multiplier_STAGE1__0701_ ),
    .A3(u_multiplier_STAGE1__0703_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_25_1__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_25_1__22_  (.A(u_multiplier_STAGE1__0702_ ),
    .B(u_multiplier_STAGE1__0701_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_25_1__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_25_1__23_  (.A(u_multiplier_STAGE1__0703_ ),
    .B(u_multiplier_STAGE1__0704_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_25_1__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_25_1__24_  (.A1(u_multiplier_STAGE1_acci1_pp_25_1__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_25_1__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_25_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_25_1__25_  (.A(u_multiplier_STAGE1_acci1_pp_25_1__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_25_1__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_25_1__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_25_1__26_  (.A1(u_multiplier_STAGE1_acci1_pp_25_1__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_25_1__16_ ),
    .ZN(u_multiplier_pp1_25 [1]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_25_1__27_  (.A1(u_multiplier_STAGE1__0702_ ),
    .A2(u_multiplier_STAGE1__0701_ ),
    .B1(u_multiplier_STAGE1__0703_ ),
    .B2(u_multiplier_STAGE1__0704_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_25_1__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_25_1__28_  (.A1(u_multiplier_STAGE1_acci1_pp_25_1__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_25_1__17_ ),
    .ZN(u_multiplier_pp1_26 [9]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_25_2__21_  (.A1(u_multiplier_STAGE1__0706_ ),
    .A2(u_multiplier_STAGE1__0705_ ),
    .A3(u_multiplier_STAGE1__0707_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_25_2__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_25_2__22_  (.A(u_multiplier_STAGE1__0706_ ),
    .B(u_multiplier_STAGE1__0705_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_25_2__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_25_2__23_  (.A(u_multiplier_STAGE1__0707_ ),
    .B(u_multiplier_STAGE1__0708_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_25_2__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_25_2__24_  (.A1(u_multiplier_STAGE1_acci1_pp_25_2__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_25_2__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_25_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_25_2__25_  (.A(u_multiplier_STAGE1_acci1_pp_25_2__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_25_2__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_25_2__16_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_25_2__26_  (.A1(u_multiplier_STAGE1_acci1_pp_25_2__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_25_2__16_ ),
    .ZN(u_multiplier_pp1_25 [2]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_25_2__27_  (.A1(u_multiplier_STAGE1__0706_ ),
    .A2(u_multiplier_STAGE1__0705_ ),
    .B1(u_multiplier_STAGE1__0707_ ),
    .B2(u_multiplier_STAGE1__0708_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_25_2__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_25_2__28_  (.A1(u_multiplier_STAGE1_acci1_pp_25_2__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_25_2__17_ ),
    .ZN(u_multiplier_pp1_26 [8]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_25_3__21_  (.A1(u_multiplier_STAGE1__0710_ ),
    .A2(u_multiplier_STAGE1__0709_ ),
    .A3(u_multiplier_STAGE1__0711_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_25_3__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_25_3__22_  (.A(u_multiplier_STAGE1__0710_ ),
    .B(u_multiplier_STAGE1__0709_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_25_3__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_25_3__23_  (.A(u_multiplier_STAGE1__0711_ ),
    .B(u_multiplier_STAGE1__0712_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_25_3__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_25_3__24_  (.A1(u_multiplier_STAGE1_acci1_pp_25_3__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_25_3__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_25_3__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_25_3__25_  (.A(u_multiplier_STAGE1_acci1_pp_25_3__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_25_3__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_25_3__16_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_25_3__26_  (.A1(u_multiplier_STAGE1_acci1_pp_25_3__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_25_3__16_ ),
    .ZN(u_multiplier_pp1_25 [3]));
 AOI22_X1 u_multiplier_STAGE1_acci1_pp_25_3__27_  (.A1(u_multiplier_STAGE1__0710_ ),
    .A2(u_multiplier_STAGE1__0709_ ),
    .B1(u_multiplier_STAGE1__0711_ ),
    .B2(u_multiplier_STAGE1__0712_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_25_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_25_3__28_  (.A1(u_multiplier_STAGE1_acci1_pp_25_3__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_25_3__17_ ),
    .ZN(u_multiplier_pp1_26 [7]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_25_4__21_  (.A1(u_multiplier_STAGE1__0714_ ),
    .A2(u_multiplier_STAGE1__0713_ ),
    .A3(u_multiplier_STAGE1__0715_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_25_4__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_25_4__22_  (.A(u_multiplier_STAGE1__0714_ ),
    .B(u_multiplier_STAGE1__0713_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_25_4__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_25_4__23_  (.A(u_multiplier_STAGE1__0715_ ),
    .B(u_multiplier_STAGE1__0716_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_25_4__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_25_4__24_  (.A1(u_multiplier_STAGE1_acci1_pp_25_4__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_25_4__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_25_4__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_25_4__25_  (.A(u_multiplier_STAGE1_acci1_pp_25_4__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_25_4__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_25_4__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_25_4__26_  (.A1(u_multiplier_STAGE1_acci1_pp_25_4__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_25_4__16_ ),
    .ZN(u_multiplier_pp1_25 [4]));
 AOI22_X1 u_multiplier_STAGE1_acci1_pp_25_4__27_  (.A1(u_multiplier_STAGE1__0714_ ),
    .A2(u_multiplier_STAGE1__0713_ ),
    .B1(u_multiplier_STAGE1__0715_ ),
    .B2(u_multiplier_STAGE1__0716_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_25_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_25_4__28_  (.A1(u_multiplier_STAGE1_acci1_pp_25_4__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_25_4__17_ ),
    .ZN(u_multiplier_pp1_26 [6]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_26_0__21_  (.A1(u_multiplier_STAGE1__0718_ ),
    .A2(u_multiplier_STAGE1__0717_ ),
    .A3(u_multiplier_STAGE1__0719_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_26_0__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_26_0__22_  (.A(u_multiplier_STAGE1__0718_ ),
    .B(u_multiplier_STAGE1__0717_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_26_0__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_26_0__23_  (.A(u_multiplier_STAGE1__0719_ ),
    .B(u_multiplier_STAGE1__0720_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_26_0__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_26_0__24_  (.A1(u_multiplier_STAGE1_acci1_pp_26_0__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_26_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_26_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_26_0__25_  (.A(u_multiplier_STAGE1_acci1_pp_26_0__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_26_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_26_0__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_26_0__26_  (.A1(u_multiplier_STAGE1_acci1_pp_26_0__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_26_0__16_ ),
    .ZN(u_multiplier_pp1_26 [0]));
 AOI22_X1 u_multiplier_STAGE1_acci1_pp_26_0__27_  (.A1(u_multiplier_STAGE1__0718_ ),
    .A2(u_multiplier_STAGE1__0717_ ),
    .B1(u_multiplier_STAGE1__0719_ ),
    .B2(u_multiplier_STAGE1__0720_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_26_0__17_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_26_0__28_  (.A1(u_multiplier_STAGE1_acci1_pp_26_0__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_26_0__17_ ),
    .ZN(u_multiplier_pp1_27 [11]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_26_1__21_  (.A1(u_multiplier_STAGE1__0722_ ),
    .A2(u_multiplier_STAGE1__0721_ ),
    .A3(u_multiplier_STAGE1__0723_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_26_1__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_26_1__22_  (.A(u_multiplier_STAGE1__0722_ ),
    .B(u_multiplier_STAGE1__0721_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_26_1__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_26_1__23_  (.A(u_multiplier_STAGE1__0723_ ),
    .B(u_multiplier_STAGE1__0724_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_26_1__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_26_1__24_  (.A1(u_multiplier_STAGE1_acci1_pp_26_1__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_26_1__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_26_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_26_1__25_  (.A(u_multiplier_STAGE1_acci1_pp_26_1__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_26_1__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_26_1__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_26_1__26_  (.A1(u_multiplier_STAGE1_acci1_pp_26_1__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_26_1__16_ ),
    .ZN(u_multiplier_pp1_26 [1]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_26_1__27_  (.A1(u_multiplier_STAGE1__0722_ ),
    .A2(u_multiplier_STAGE1__0721_ ),
    .B1(u_multiplier_STAGE1__0723_ ),
    .B2(u_multiplier_STAGE1__0724_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_26_1__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_26_1__28_  (.A1(u_multiplier_STAGE1_acci1_pp_26_1__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_26_1__17_ ),
    .ZN(u_multiplier_pp1_27 [10]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_26_2__21_  (.A1(u_multiplier_STAGE1__0726_ ),
    .A2(u_multiplier_STAGE1__0725_ ),
    .A3(u_multiplier_STAGE1__0727_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_26_2__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_26_2__22_  (.A(u_multiplier_STAGE1__0726_ ),
    .B(u_multiplier_STAGE1__0725_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_26_2__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_26_2__23_  (.A(u_multiplier_STAGE1__0727_ ),
    .B(u_multiplier_STAGE1__0728_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_26_2__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_26_2__24_  (.A1(u_multiplier_STAGE1_acci1_pp_26_2__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_26_2__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_26_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_26_2__25_  (.A(u_multiplier_STAGE1_acci1_pp_26_2__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_26_2__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_26_2__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_26_2__26_  (.A1(u_multiplier_STAGE1_acci1_pp_26_2__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_26_2__16_ ),
    .ZN(u_multiplier_pp1_26 [2]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_26_2__27_  (.A1(u_multiplier_STAGE1__0726_ ),
    .A2(u_multiplier_STAGE1__0725_ ),
    .B1(u_multiplier_STAGE1__0727_ ),
    .B2(u_multiplier_STAGE1__0728_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_26_2__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_26_2__28_  (.A1(u_multiplier_STAGE1_acci1_pp_26_2__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_26_2__17_ ),
    .ZN(u_multiplier_pp1_27 [9]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_26_3__21_  (.A1(u_multiplier_STAGE1__0730_ ),
    .A2(u_multiplier_STAGE1__0729_ ),
    .A3(u_multiplier_STAGE1__0731_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_26_3__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_26_3__22_  (.A(u_multiplier_STAGE1__0730_ ),
    .B(u_multiplier_STAGE1__0729_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_26_3__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_26_3__23_  (.A(u_multiplier_STAGE1__0731_ ),
    .B(u_multiplier_STAGE1__0732_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_26_3__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_26_3__24_  (.A1(u_multiplier_STAGE1_acci1_pp_26_3__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_26_3__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_26_3__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_26_3__25_  (.A(u_multiplier_STAGE1_acci1_pp_26_3__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_26_3__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_26_3__16_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_26_3__26_  (.A1(u_multiplier_STAGE1_acci1_pp_26_3__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_26_3__16_ ),
    .ZN(u_multiplier_pp1_26 [3]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_26_3__27_  (.A1(u_multiplier_STAGE1__0730_ ),
    .A2(u_multiplier_STAGE1__0729_ ),
    .B1(u_multiplier_STAGE1__0731_ ),
    .B2(u_multiplier_STAGE1__0732_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_26_3__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_26_3__28_  (.A1(u_multiplier_STAGE1_acci1_pp_26_3__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_26_3__17_ ),
    .ZN(u_multiplier_pp1_27 [8]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_26_4__21_  (.A1(u_multiplier_STAGE1__0734_ ),
    .A2(u_multiplier_STAGE1__0733_ ),
    .A3(u_multiplier_STAGE1__0735_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_26_4__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_26_4__22_  (.A(u_multiplier_STAGE1__0734_ ),
    .B(u_multiplier_STAGE1__0733_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_26_4__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_26_4__23_  (.A(u_multiplier_STAGE1__0735_ ),
    .B(u_multiplier_STAGE1__0736_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_26_4__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_26_4__24_  (.A1(u_multiplier_STAGE1_acci1_pp_26_4__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_26_4__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_26_4__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_26_4__25_  (.A(u_multiplier_STAGE1_acci1_pp_26_4__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_26_4__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_26_4__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_26_4__26_  (.A1(u_multiplier_STAGE1_acci1_pp_26_4__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_26_4__16_ ),
    .ZN(u_multiplier_pp1_26 [4]));
 AOI22_X1 u_multiplier_STAGE1_acci1_pp_26_4__27_  (.A1(u_multiplier_STAGE1__0734_ ),
    .A2(u_multiplier_STAGE1__0733_ ),
    .B1(u_multiplier_STAGE1__0735_ ),
    .B2(u_multiplier_STAGE1__0736_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_26_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_26_4__28_  (.A1(u_multiplier_STAGE1_acci1_pp_26_4__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_26_4__17_ ),
    .ZN(u_multiplier_pp1_27 [7]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_27_0__21_  (.A1(u_multiplier_STAGE1__0740_ ),
    .A2(u_multiplier_STAGE1__0739_ ),
    .A3(u_multiplier_STAGE1__0741_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_27_0__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_27_0__22_  (.A(u_multiplier_STAGE1__0740_ ),
    .B(u_multiplier_STAGE1__0739_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_27_0__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_27_0__23_  (.A(u_multiplier_STAGE1__0741_ ),
    .B(u_multiplier_STAGE1__0742_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_27_0__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_27_0__24_  (.A1(u_multiplier_STAGE1_acci1_pp_27_0__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_27_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_27_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_27_0__25_  (.A(u_multiplier_STAGE1_acci1_pp_27_0__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_27_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_27_0__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_27_0__26_  (.A1(u_multiplier_STAGE1_acci1_pp_27_0__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_27_0__16_ ),
    .ZN(u_multiplier_pp1_27 [0]));
 AOI22_X1 u_multiplier_STAGE1_acci1_pp_27_0__27_  (.A1(u_multiplier_STAGE1__0740_ ),
    .A2(u_multiplier_STAGE1__0739_ ),
    .B1(u_multiplier_STAGE1__0741_ ),
    .B2(u_multiplier_STAGE1__0742_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_27_0__17_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_27_0__28_  (.A1(u_multiplier_STAGE1_acci1_pp_27_0__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_27_0__17_ ),
    .ZN(u_multiplier_pp1_28 [12]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_27_1__21_  (.A1(u_multiplier_STAGE1__0744_ ),
    .A2(u_multiplier_STAGE1__0743_ ),
    .A3(u_multiplier_STAGE1__0745_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_27_1__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_27_1__22_  (.A(u_multiplier_STAGE1__0744_ ),
    .B(u_multiplier_STAGE1__0743_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_27_1__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_27_1__23_  (.A(u_multiplier_STAGE1__0745_ ),
    .B(u_multiplier_STAGE1__0746_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_27_1__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_27_1__24_  (.A1(u_multiplier_STAGE1_acci1_pp_27_1__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_27_1__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_27_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_27_1__25_  (.A(u_multiplier_STAGE1_acci1_pp_27_1__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_27_1__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_27_1__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_27_1__26_  (.A1(u_multiplier_STAGE1_acci1_pp_27_1__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_27_1__16_ ),
    .ZN(u_multiplier_pp1_27 [1]));
 AOI22_X1 u_multiplier_STAGE1_acci1_pp_27_1__27_  (.A1(u_multiplier_STAGE1__0744_ ),
    .A2(u_multiplier_STAGE1__0743_ ),
    .B1(u_multiplier_STAGE1__0745_ ),
    .B2(u_multiplier_STAGE1__0746_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_27_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_27_1__28_  (.A1(u_multiplier_STAGE1_acci1_pp_27_1__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_27_1__17_ ),
    .ZN(u_multiplier_pp1_28 [11]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_27_2__21_  (.A1(u_multiplier_STAGE1__0748_ ),
    .A2(u_multiplier_STAGE1__0747_ ),
    .A3(u_multiplier_STAGE1__0749_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_27_2__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_27_2__22_  (.A(u_multiplier_STAGE1__0748_ ),
    .B(u_multiplier_STAGE1__0747_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_27_2__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_27_2__23_  (.A(u_multiplier_STAGE1__0749_ ),
    .B(u_multiplier_STAGE1__0750_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_27_2__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_27_2__24_  (.A1(u_multiplier_STAGE1_acci1_pp_27_2__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_27_2__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_27_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_27_2__25_  (.A(u_multiplier_STAGE1_acci1_pp_27_2__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_27_2__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_27_2__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_27_2__26_  (.A1(u_multiplier_STAGE1_acci1_pp_27_2__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_27_2__16_ ),
    .ZN(u_multiplier_pp1_27 [2]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_27_2__27_  (.A1(u_multiplier_STAGE1__0748_ ),
    .A2(u_multiplier_STAGE1__0747_ ),
    .B1(u_multiplier_STAGE1__0749_ ),
    .B2(u_multiplier_STAGE1__0750_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_27_2__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_27_2__28_  (.A1(u_multiplier_STAGE1_acci1_pp_27_2__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_27_2__17_ ),
    .ZN(u_multiplier_pp1_28 [10]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_27_3__21_  (.A1(u_multiplier_STAGE1__0752_ ),
    .A2(u_multiplier_STAGE1__0751_ ),
    .A3(u_multiplier_STAGE1__0753_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_27_3__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_27_3__22_  (.A(u_multiplier_STAGE1__0752_ ),
    .B(u_multiplier_STAGE1__0751_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_27_3__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_27_3__23_  (.A(u_multiplier_STAGE1__0753_ ),
    .B(u_multiplier_STAGE1__0754_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_27_3__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_27_3__24_  (.A1(u_multiplier_STAGE1_acci1_pp_27_3__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_27_3__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_27_3__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_27_3__25_  (.A(u_multiplier_STAGE1_acci1_pp_27_3__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_27_3__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_27_3__16_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_27_3__26_  (.A1(u_multiplier_STAGE1_acci1_pp_27_3__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_27_3__16_ ),
    .ZN(u_multiplier_pp1_27 [3]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_27_3__27_  (.A1(u_multiplier_STAGE1__0752_ ),
    .A2(u_multiplier_STAGE1__0751_ ),
    .B1(u_multiplier_STAGE1__0753_ ),
    .B2(u_multiplier_STAGE1__0754_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_27_3__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_27_3__28_  (.A1(u_multiplier_STAGE1_acci1_pp_27_3__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_27_3__17_ ),
    .ZN(u_multiplier_pp1_28 [9]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_27_4__21_  (.A1(u_multiplier_STAGE1__0756_ ),
    .A2(u_multiplier_STAGE1__0755_ ),
    .A3(u_multiplier_STAGE1__0757_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_27_4__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_27_4__22_  (.A(u_multiplier_STAGE1__0756_ ),
    .B(u_multiplier_STAGE1__0755_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_27_4__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_27_4__23_  (.A(u_multiplier_STAGE1__0757_ ),
    .B(u_multiplier_STAGE1__0758_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_27_4__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_27_4__24_  (.A1(u_multiplier_STAGE1_acci1_pp_27_4__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_27_4__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_27_4__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_27_4__25_  (.A(u_multiplier_STAGE1_acci1_pp_27_4__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_27_4__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_27_4__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_27_4__26_  (.A1(u_multiplier_STAGE1_acci1_pp_27_4__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_27_4__16_ ),
    .ZN(u_multiplier_pp1_27 [4]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_27_4__27_  (.A1(u_multiplier_STAGE1__0756_ ),
    .A2(u_multiplier_STAGE1__0755_ ),
    .B1(u_multiplier_STAGE1__0757_ ),
    .B2(u_multiplier_STAGE1__0758_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_27_4__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_27_4__28_  (.A1(u_multiplier_STAGE1_acci1_pp_27_4__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_27_4__17_ ),
    .ZN(u_multiplier_pp1_28 [8]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_27_5__21_  (.A1(u_multiplier_STAGE1__0760_ ),
    .A2(u_multiplier_STAGE1__0759_ ),
    .A3(u_multiplier_STAGE1__0761_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_27_5__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_27_5__22_  (.A(u_multiplier_STAGE1__0760_ ),
    .B(u_multiplier_STAGE1__0759_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_27_5__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_27_5__23_  (.A(u_multiplier_STAGE1__0761_ ),
    .B(u_multiplier_STAGE1__0762_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_27_5__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_27_5__24_  (.A1(u_multiplier_STAGE1_acci1_pp_27_5__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_27_5__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_27_5__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_27_5__25_  (.A(u_multiplier_STAGE1_acci1_pp_27_5__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_27_5__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_27_5__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_27_5__26_  (.A1(u_multiplier_STAGE1_acci1_pp_27_5__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_27_5__16_ ),
    .ZN(u_multiplier_pp1_27 [5]));
 AOI22_X1 u_multiplier_STAGE1_acci1_pp_27_5__27_  (.A1(u_multiplier_STAGE1__0760_ ),
    .A2(u_multiplier_STAGE1__0759_ ),
    .B1(u_multiplier_STAGE1__0761_ ),
    .B2(u_multiplier_STAGE1__0762_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_27_5__17_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_27_5__28_  (.A1(u_multiplier_STAGE1_acci1_pp_27_5__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_27_5__17_ ),
    .ZN(u_multiplier_pp1_28 [7]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_28_0__21_  (.A1(u_multiplier_STAGE1__0764_ ),
    .A2(u_multiplier_STAGE1__0763_ ),
    .A3(u_multiplier_STAGE1__0765_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_28_0__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_28_0__22_  (.A(u_multiplier_STAGE1__0764_ ),
    .B(u_multiplier_STAGE1__0763_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_28_0__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_28_0__23_  (.A(u_multiplier_STAGE1__0765_ ),
    .B(u_multiplier_STAGE1__0766_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_28_0__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_28_0__24_  (.A1(u_multiplier_STAGE1_acci1_pp_28_0__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_28_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_28_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_28_0__25_  (.A(u_multiplier_STAGE1_acci1_pp_28_0__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_28_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_28_0__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_28_0__26_  (.A1(u_multiplier_STAGE1_acci1_pp_28_0__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_28_0__16_ ),
    .ZN(u_multiplier_pp1_28 [0]));
 AOI22_X1 u_multiplier_STAGE1_acci1_pp_28_0__27_  (.A1(u_multiplier_STAGE1__0764_ ),
    .A2(u_multiplier_STAGE1__0763_ ),
    .B1(u_multiplier_STAGE1__0765_ ),
    .B2(u_multiplier_STAGE1__0766_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_28_0__17_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_28_0__28_  (.A1(u_multiplier_STAGE1_acci1_pp_28_0__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_28_0__17_ ),
    .ZN(u_multiplier_pp1_29 [13]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_28_1__21_  (.A1(u_multiplier_STAGE1__0768_ ),
    .A2(u_multiplier_STAGE1__0767_ ),
    .A3(u_multiplier_STAGE1__0769_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_28_1__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_28_1__22_  (.A(u_multiplier_STAGE1__0768_ ),
    .B(u_multiplier_STAGE1__0767_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_28_1__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_28_1__23_  (.A(u_multiplier_STAGE1__0769_ ),
    .B(u_multiplier_STAGE1__0770_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_28_1__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_28_1__24_  (.A1(u_multiplier_STAGE1_acci1_pp_28_1__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_28_1__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_28_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_28_1__25_  (.A(u_multiplier_STAGE1_acci1_pp_28_1__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_28_1__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_28_1__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_28_1__26_  (.A1(u_multiplier_STAGE1_acci1_pp_28_1__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_28_1__16_ ),
    .ZN(u_multiplier_pp1_28 [1]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_28_1__27_  (.A1(u_multiplier_STAGE1__0768_ ),
    .A2(u_multiplier_STAGE1__0767_ ),
    .B1(u_multiplier_STAGE1__0769_ ),
    .B2(u_multiplier_STAGE1__0770_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_28_1__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_28_1__28_  (.A1(u_multiplier_STAGE1_acci1_pp_28_1__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_28_1__17_ ),
    .ZN(u_multiplier_pp1_29 [12]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_28_2__21_  (.A1(u_multiplier_STAGE1__0772_ ),
    .A2(u_multiplier_STAGE1__0771_ ),
    .A3(u_multiplier_STAGE1__0773_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_28_2__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_28_2__22_  (.A(u_multiplier_STAGE1__0772_ ),
    .B(u_multiplier_STAGE1__0771_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_28_2__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_28_2__23_  (.A(u_multiplier_STAGE1__0773_ ),
    .B(u_multiplier_STAGE1__0774_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_28_2__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_28_2__24_  (.A1(u_multiplier_STAGE1_acci1_pp_28_2__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_28_2__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_28_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_28_2__25_  (.A(u_multiplier_STAGE1_acci1_pp_28_2__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_28_2__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_28_2__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_28_2__26_  (.A1(u_multiplier_STAGE1_acci1_pp_28_2__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_28_2__16_ ),
    .ZN(u_multiplier_pp1_28 [2]));
 AOI22_X1 u_multiplier_STAGE1_acci1_pp_28_2__27_  (.A1(u_multiplier_STAGE1__0772_ ),
    .A2(u_multiplier_STAGE1__0771_ ),
    .B1(u_multiplier_STAGE1__0773_ ),
    .B2(u_multiplier_STAGE1__0774_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_28_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_28_2__28_  (.A1(u_multiplier_STAGE1_acci1_pp_28_2__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_28_2__17_ ),
    .ZN(u_multiplier_pp1_29 [11]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_28_3__21_  (.A1(u_multiplier_STAGE1__0776_ ),
    .A2(u_multiplier_STAGE1__0775_ ),
    .A3(u_multiplier_STAGE1__0777_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_28_3__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_28_3__22_  (.A(u_multiplier_STAGE1__0776_ ),
    .B(u_multiplier_STAGE1__0775_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_28_3__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_28_3__23_  (.A(u_multiplier_STAGE1__0777_ ),
    .B(u_multiplier_STAGE1__0778_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_28_3__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_28_3__24_  (.A1(u_multiplier_STAGE1_acci1_pp_28_3__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_28_3__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_28_3__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_28_3__25_  (.A(u_multiplier_STAGE1_acci1_pp_28_3__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_28_3__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_28_3__16_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_28_3__26_  (.A1(u_multiplier_STAGE1_acci1_pp_28_3__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_28_3__16_ ),
    .ZN(u_multiplier_pp1_28 [3]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_28_3__27_  (.A1(u_multiplier_STAGE1__0776_ ),
    .A2(u_multiplier_STAGE1__0775_ ),
    .B1(u_multiplier_STAGE1__0777_ ),
    .B2(u_multiplier_STAGE1__0778_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_28_3__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_28_3__28_  (.A1(u_multiplier_STAGE1_acci1_pp_28_3__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_28_3__17_ ),
    .ZN(u_multiplier_pp1_29 [10]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_28_4__21_  (.A1(u_multiplier_STAGE1__0780_ ),
    .A2(u_multiplier_STAGE1__0779_ ),
    .A3(u_multiplier_STAGE1__0781_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_28_4__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_28_4__22_  (.A(u_multiplier_STAGE1__0780_ ),
    .B(u_multiplier_STAGE1__0779_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_28_4__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_28_4__23_  (.A(u_multiplier_STAGE1__0781_ ),
    .B(u_multiplier_STAGE1__0782_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_28_4__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_28_4__24_  (.A1(u_multiplier_STAGE1_acci1_pp_28_4__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_28_4__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_28_4__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_28_4__25_  (.A(u_multiplier_STAGE1_acci1_pp_28_4__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_28_4__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_28_4__16_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_28_4__26_  (.A1(u_multiplier_STAGE1_acci1_pp_28_4__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_28_4__16_ ),
    .ZN(u_multiplier_pp1_28 [4]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_28_4__27_  (.A1(u_multiplier_STAGE1__0780_ ),
    .A2(u_multiplier_STAGE1__0779_ ),
    .B1(u_multiplier_STAGE1__0781_ ),
    .B2(u_multiplier_STAGE1__0782_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_28_4__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_28_4__28_  (.A1(u_multiplier_STAGE1_acci1_pp_28_4__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_28_4__17_ ),
    .ZN(u_multiplier_pp1_29 [9]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_28_5__21_  (.A1(u_multiplier_STAGE1__0784_ ),
    .A2(u_multiplier_STAGE1__0783_ ),
    .A3(u_multiplier_STAGE1__0785_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_28_5__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_28_5__22_  (.A(u_multiplier_STAGE1__0784_ ),
    .B(u_multiplier_STAGE1__0783_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_28_5__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_28_5__23_  (.A(u_multiplier_STAGE1__0785_ ),
    .B(u_multiplier_STAGE1__0786_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_28_5__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_28_5__24_  (.A1(u_multiplier_STAGE1_acci1_pp_28_5__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_28_5__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_28_5__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_28_5__25_  (.A(u_multiplier_STAGE1_acci1_pp_28_5__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_28_5__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_28_5__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_28_5__26_  (.A1(u_multiplier_STAGE1_acci1_pp_28_5__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_28_5__16_ ),
    .ZN(u_multiplier_pp1_28 [5]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_28_5__27_  (.A1(u_multiplier_STAGE1__0784_ ),
    .A2(u_multiplier_STAGE1__0783_ ),
    .B1(u_multiplier_STAGE1__0785_ ),
    .B2(u_multiplier_STAGE1__0786_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_28_5__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_28_5__28_  (.A1(u_multiplier_STAGE1_acci1_pp_28_5__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_28_5__17_ ),
    .ZN(u_multiplier_pp1_29 [8]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_29_0__21_  (.A1(u_multiplier_STAGE1__0790_ ),
    .A2(u_multiplier_STAGE1__0789_ ),
    .A3(u_multiplier_STAGE1__0791_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_0__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_29_0__22_  (.A(u_multiplier_STAGE1__0790_ ),
    .B(u_multiplier_STAGE1__0789_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_29_0__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_29_0__23_  (.A(u_multiplier_STAGE1__0791_ ),
    .B(u_multiplier_STAGE1__0792_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_29_0__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_29_0__24_  (.A1(u_multiplier_STAGE1_acci1_pp_29_0__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_29_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_29_0__25_  (.A(u_multiplier_STAGE1_acci1_pp_29_0__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_29_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_0__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_29_0__26_  (.A1(u_multiplier_STAGE1_acci1_pp_29_0__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_29_0__16_ ),
    .ZN(u_multiplier_pp1_29 [0]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_29_0__27_  (.A1(u_multiplier_STAGE1__0790_ ),
    .A2(u_multiplier_STAGE1__0789_ ),
    .B1(u_multiplier_STAGE1__0791_ ),
    .B2(u_multiplier_STAGE1__0792_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_0__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_29_0__28_  (.A1(u_multiplier_STAGE1_acci1_pp_29_0__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_29_0__17_ ),
    .ZN(u_multiplier_pp1_30 [14]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_29_1__21_  (.A1(u_multiplier_STAGE1__0794_ ),
    .A2(u_multiplier_STAGE1__0793_ ),
    .A3(u_multiplier_STAGE1__0795_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_1__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_29_1__22_  (.A(u_multiplier_STAGE1__0794_ ),
    .B(u_multiplier_STAGE1__0793_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_29_1__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_29_1__23_  (.A(u_multiplier_STAGE1__0795_ ),
    .B(u_multiplier_STAGE1__0796_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_29_1__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_29_1__24_  (.A1(u_multiplier_STAGE1_acci1_pp_29_1__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_29_1__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_29_1__25_  (.A(u_multiplier_STAGE1_acci1_pp_29_1__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_29_1__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_1__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_29_1__26_  (.A1(u_multiplier_STAGE1_acci1_pp_29_1__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_29_1__16_ ),
    .ZN(u_multiplier_pp1_29 [1]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_29_1__27_  (.A1(u_multiplier_STAGE1__0794_ ),
    .A2(u_multiplier_STAGE1__0793_ ),
    .B1(u_multiplier_STAGE1__0795_ ),
    .B2(u_multiplier_STAGE1__0796_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_1__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_29_1__28_  (.A1(u_multiplier_STAGE1_acci1_pp_29_1__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_29_1__17_ ),
    .ZN(u_multiplier_pp1_30 [13]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_29_2__21_  (.A1(u_multiplier_STAGE1__0798_ ),
    .A2(u_multiplier_STAGE1__0797_ ),
    .A3(u_multiplier_STAGE1__0799_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_2__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_29_2__22_  (.A(u_multiplier_STAGE1__0798_ ),
    .B(u_multiplier_STAGE1__0797_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_29_2__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_29_2__23_  (.A(u_multiplier_STAGE1__0799_ ),
    .B(u_multiplier_STAGE1__0800_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_29_2__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_29_2__24_  (.A1(u_multiplier_STAGE1_acci1_pp_29_2__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_29_2__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_29_2__25_  (.A(u_multiplier_STAGE1_acci1_pp_29_2__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_29_2__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_2__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_29_2__26_  (.A1(u_multiplier_STAGE1_acci1_pp_29_2__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_29_2__16_ ),
    .ZN(u_multiplier_pp1_29 [2]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_29_2__27_  (.A1(u_multiplier_STAGE1__0798_ ),
    .A2(u_multiplier_STAGE1__0797_ ),
    .B1(u_multiplier_STAGE1__0799_ ),
    .B2(u_multiplier_STAGE1__0800_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_2__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_29_2__28_  (.A1(u_multiplier_STAGE1_acci1_pp_29_2__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_29_2__17_ ),
    .ZN(u_multiplier_pp1_30 [12]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_29_3__21_  (.A1(u_multiplier_STAGE1__0802_ ),
    .A2(u_multiplier_STAGE1__0801_ ),
    .A3(u_multiplier_STAGE1__0803_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_3__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_29_3__22_  (.A(u_multiplier_STAGE1__0802_ ),
    .B(u_multiplier_STAGE1__0801_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_29_3__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_29_3__23_  (.A(u_multiplier_STAGE1__0803_ ),
    .B(u_multiplier_STAGE1__0804_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_29_3__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_29_3__24_  (.A1(u_multiplier_STAGE1_acci1_pp_29_3__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_29_3__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_3__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_29_3__25_  (.A(u_multiplier_STAGE1_acci1_pp_29_3__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_29_3__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_3__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_29_3__26_  (.A1(u_multiplier_STAGE1_acci1_pp_29_3__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_29_3__16_ ),
    .ZN(u_multiplier_pp1_29 [3]));
 AOI22_X1 u_multiplier_STAGE1_acci1_pp_29_3__27_  (.A1(u_multiplier_STAGE1__0802_ ),
    .A2(u_multiplier_STAGE1__0801_ ),
    .B1(u_multiplier_STAGE1__0803_ ),
    .B2(u_multiplier_STAGE1__0804_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_29_3__28_  (.A1(u_multiplier_STAGE1_acci1_pp_29_3__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_29_3__17_ ),
    .ZN(u_multiplier_pp1_30 [11]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_29_4__21_  (.A1(u_multiplier_STAGE1__0806_ ),
    .A2(u_multiplier_STAGE1__0805_ ),
    .A3(u_multiplier_STAGE1__0807_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_4__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_29_4__22_  (.A(u_multiplier_STAGE1__0806_ ),
    .B(u_multiplier_STAGE1__0805_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_29_4__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_29_4__23_  (.A(u_multiplier_STAGE1__0807_ ),
    .B(u_multiplier_STAGE1__0808_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_29_4__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_29_4__24_  (.A1(u_multiplier_STAGE1_acci1_pp_29_4__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_29_4__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_4__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_29_4__25_  (.A(u_multiplier_STAGE1_acci1_pp_29_4__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_29_4__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_4__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_29_4__26_  (.A1(u_multiplier_STAGE1_acci1_pp_29_4__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_29_4__16_ ),
    .ZN(u_multiplier_pp1_29 [4]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_29_4__27_  (.A1(u_multiplier_STAGE1__0806_ ),
    .A2(u_multiplier_STAGE1__0805_ ),
    .B1(u_multiplier_STAGE1__0807_ ),
    .B2(u_multiplier_STAGE1__0808_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_4__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_29_4__28_  (.A1(u_multiplier_STAGE1_acci1_pp_29_4__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_29_4__17_ ),
    .ZN(u_multiplier_pp1_30 [10]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_29_5__21_  (.A1(u_multiplier_STAGE1__0810_ ),
    .A2(u_multiplier_STAGE1__0809_ ),
    .A3(u_multiplier_STAGE1__0811_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_5__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_29_5__22_  (.A(u_multiplier_STAGE1__0810_ ),
    .B(u_multiplier_STAGE1__0809_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_29_5__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_29_5__23_  (.A(u_multiplier_STAGE1__0811_ ),
    .B(u_multiplier_STAGE1__0812_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_29_5__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_29_5__24_  (.A1(u_multiplier_STAGE1_acci1_pp_29_5__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_29_5__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_5__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_29_5__25_  (.A(u_multiplier_STAGE1_acci1_pp_29_5__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_29_5__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_5__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_29_5__26_  (.A1(u_multiplier_STAGE1_acci1_pp_29_5__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_29_5__16_ ),
    .ZN(u_multiplier_pp1_29 [5]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_29_5__27_  (.A1(u_multiplier_STAGE1__0810_ ),
    .A2(u_multiplier_STAGE1__0809_ ),
    .B1(u_multiplier_STAGE1__0811_ ),
    .B2(u_multiplier_STAGE1__0812_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_5__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_29_5__28_  (.A1(u_multiplier_STAGE1_acci1_pp_29_5__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_29_5__17_ ),
    .ZN(u_multiplier_pp1_30 [9]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_29_6__21_  (.A1(u_multiplier_STAGE1__0814_ ),
    .A2(u_multiplier_STAGE1__0813_ ),
    .A3(u_multiplier_STAGE1__0815_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_6__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_29_6__22_  (.A(u_multiplier_STAGE1__0814_ ),
    .B(u_multiplier_STAGE1__0813_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_29_6__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_29_6__23_  (.A(u_multiplier_STAGE1__0815_ ),
    .B(u_multiplier_STAGE1__0816_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_29_6__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_29_6__24_  (.A1(u_multiplier_STAGE1_acci1_pp_29_6__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_29_6__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_6__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_29_6__25_  (.A(u_multiplier_STAGE1_acci1_pp_29_6__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_29_6__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_6__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_29_6__26_  (.A1(u_multiplier_STAGE1_acci1_pp_29_6__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_29_6__16_ ),
    .ZN(u_multiplier_pp1_29 [6]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_29_6__27_  (.A1(u_multiplier_STAGE1__0814_ ),
    .A2(u_multiplier_STAGE1__0813_ ),
    .B1(u_multiplier_STAGE1__0815_ ),
    .B2(u_multiplier_STAGE1__0816_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_29_6__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_29_6__28_  (.A1(u_multiplier_STAGE1_acci1_pp_29_6__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_29_6__17_ ),
    .ZN(u_multiplier_pp1_30 [8]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_30_0__21_  (.A1(u_multiplier_STAGE1__0818_ ),
    .A2(u_multiplier_STAGE1__0817_ ),
    .A3(u_multiplier_STAGE1__0819_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_0__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_30_0__22_  (.A(u_multiplier_STAGE1__0818_ ),
    .B(u_multiplier_STAGE1__0817_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_30_0__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_30_0__23_  (.A(u_multiplier_STAGE1__0819_ ),
    .B(u_multiplier_STAGE1__0820_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_30_0__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_30_0__24_  (.A1(u_multiplier_STAGE1_acci1_pp_30_0__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_30_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_30_0__25_  (.A(u_multiplier_STAGE1_acci1_pp_30_0__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_30_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_0__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_30_0__26_  (.A1(u_multiplier_STAGE1_acci1_pp_30_0__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_30_0__16_ ),
    .ZN(u_multiplier_pp1_30 [0]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_30_0__27_  (.A1(u_multiplier_STAGE1__0818_ ),
    .A2(u_multiplier_STAGE1__0817_ ),
    .B1(u_multiplier_STAGE1__0819_ ),
    .B2(u_multiplier_STAGE1__0820_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_0__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_30_0__28_  (.A1(u_multiplier_STAGE1_acci1_pp_30_0__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_30_0__17_ ),
    .ZN(u_multiplier_pp1_31 [15]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_30_1__21_  (.A1(u_multiplier_STAGE1__0822_ ),
    .A2(u_multiplier_STAGE1__0821_ ),
    .A3(u_multiplier_STAGE1__0823_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_1__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_30_1__22_  (.A(u_multiplier_STAGE1__0822_ ),
    .B(u_multiplier_STAGE1__0821_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_30_1__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_30_1__23_  (.A(u_multiplier_STAGE1__0823_ ),
    .B(u_multiplier_STAGE1__0824_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_30_1__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_30_1__24_  (.A1(u_multiplier_STAGE1_acci1_pp_30_1__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_30_1__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_30_1__25_  (.A(u_multiplier_STAGE1_acci1_pp_30_1__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_30_1__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_1__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_30_1__26_  (.A1(u_multiplier_STAGE1_acci1_pp_30_1__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_30_1__16_ ),
    .ZN(u_multiplier_pp1_30 [1]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_30_1__27_  (.A1(u_multiplier_STAGE1__0822_ ),
    .A2(u_multiplier_STAGE1__0821_ ),
    .B1(u_multiplier_STAGE1__0823_ ),
    .B2(u_multiplier_STAGE1__0824_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_1__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_30_1__28_  (.A1(u_multiplier_STAGE1_acci1_pp_30_1__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_30_1__17_ ),
    .ZN(u_multiplier_pp1_31 [14]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_30_2__21_  (.A1(u_multiplier_STAGE1__0826_ ),
    .A2(u_multiplier_STAGE1__0825_ ),
    .A3(u_multiplier_STAGE1__0827_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_2__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_30_2__22_  (.A(u_multiplier_STAGE1__0826_ ),
    .B(u_multiplier_STAGE1__0825_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_30_2__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_30_2__23_  (.A(u_multiplier_STAGE1__0827_ ),
    .B(u_multiplier_STAGE1__0828_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_30_2__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_30_2__24_  (.A1(u_multiplier_STAGE1_acci1_pp_30_2__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_30_2__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_30_2__25_  (.A(u_multiplier_STAGE1_acci1_pp_30_2__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_30_2__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_2__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_30_2__26_  (.A1(u_multiplier_STAGE1_acci1_pp_30_2__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_30_2__16_ ),
    .ZN(u_multiplier_pp1_30 [2]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_30_2__27_  (.A1(u_multiplier_STAGE1__0826_ ),
    .A2(u_multiplier_STAGE1__0825_ ),
    .B1(u_multiplier_STAGE1__0827_ ),
    .B2(u_multiplier_STAGE1__0828_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_2__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_30_2__28_  (.A1(u_multiplier_STAGE1_acci1_pp_30_2__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_30_2__17_ ),
    .ZN(u_multiplier_pp1_31 [13]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_30_3__21_  (.A1(u_multiplier_STAGE1__0830_ ),
    .A2(u_multiplier_STAGE1__0829_ ),
    .A3(u_multiplier_STAGE1__0831_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_3__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_30_3__22_  (.A(u_multiplier_STAGE1__0830_ ),
    .B(u_multiplier_STAGE1__0829_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_30_3__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_30_3__23_  (.A(u_multiplier_STAGE1__0831_ ),
    .B(u_multiplier_STAGE1__0832_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_30_3__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_30_3__24_  (.A1(u_multiplier_STAGE1_acci1_pp_30_3__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_30_3__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_3__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_30_3__25_  (.A(u_multiplier_STAGE1_acci1_pp_30_3__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_30_3__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_3__16_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_30_3__26_  (.A1(u_multiplier_STAGE1_acci1_pp_30_3__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_30_3__16_ ),
    .ZN(u_multiplier_pp1_30 [3]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_30_3__27_  (.A1(u_multiplier_STAGE1__0830_ ),
    .A2(u_multiplier_STAGE1__0829_ ),
    .B1(u_multiplier_STAGE1__0831_ ),
    .B2(u_multiplier_STAGE1__0832_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_3__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_30_3__28_  (.A1(u_multiplier_STAGE1_acci1_pp_30_3__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_30_3__17_ ),
    .ZN(u_multiplier_pp1_31 [12]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_30_4__21_  (.A1(u_multiplier_STAGE1__0834_ ),
    .A2(u_multiplier_STAGE1__0833_ ),
    .A3(u_multiplier_STAGE1__0835_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_4__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_30_4__22_  (.A(u_multiplier_STAGE1__0834_ ),
    .B(u_multiplier_STAGE1__0833_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_30_4__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_30_4__23_  (.A(u_multiplier_STAGE1__0835_ ),
    .B(u_multiplier_STAGE1__0836_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_30_4__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_30_4__24_  (.A1(u_multiplier_STAGE1_acci1_pp_30_4__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_30_4__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_4__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_30_4__25_  (.A(u_multiplier_STAGE1_acci1_pp_30_4__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_30_4__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_4__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_30_4__26_  (.A1(u_multiplier_STAGE1_acci1_pp_30_4__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_30_4__16_ ),
    .ZN(u_multiplier_pp1_30 [4]));
 AOI22_X1 u_multiplier_STAGE1_acci1_pp_30_4__27_  (.A1(u_multiplier_STAGE1__0834_ ),
    .A2(u_multiplier_STAGE1__0833_ ),
    .B1(u_multiplier_STAGE1__0835_ ),
    .B2(u_multiplier_STAGE1__0836_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_30_4__28_  (.A1(u_multiplier_STAGE1_acci1_pp_30_4__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_30_4__17_ ),
    .ZN(u_multiplier_pp1_31 [11]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_30_5__21_  (.A1(u_multiplier_STAGE1__0838_ ),
    .A2(u_multiplier_STAGE1__0837_ ),
    .A3(u_multiplier_STAGE1__0839_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_5__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_30_5__22_  (.A(u_multiplier_STAGE1__0838_ ),
    .B(u_multiplier_STAGE1__0837_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_30_5__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_30_5__23_  (.A(u_multiplier_STAGE1__0839_ ),
    .B(u_multiplier_STAGE1__0840_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_30_5__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_30_5__24_  (.A1(u_multiplier_STAGE1_acci1_pp_30_5__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_30_5__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_5__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_30_5__25_  (.A(u_multiplier_STAGE1_acci1_pp_30_5__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_30_5__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_5__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_30_5__26_  (.A1(u_multiplier_STAGE1_acci1_pp_30_5__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_30_5__16_ ),
    .ZN(u_multiplier_pp1_30 [5]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_30_5__27_  (.A1(u_multiplier_STAGE1__0838_ ),
    .A2(u_multiplier_STAGE1__0837_ ),
    .B1(u_multiplier_STAGE1__0839_ ),
    .B2(u_multiplier_STAGE1__0840_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_5__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_30_5__28_  (.A1(u_multiplier_STAGE1_acci1_pp_30_5__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_30_5__17_ ),
    .ZN(u_multiplier_pp1_31 [10]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_30_6__21_  (.A1(u_multiplier_STAGE1__0842_ ),
    .A2(u_multiplier_STAGE1__0841_ ),
    .A3(u_multiplier_STAGE1__0843_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_6__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_30_6__22_  (.A(u_multiplier_STAGE1__0842_ ),
    .B(u_multiplier_STAGE1__0841_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_30_6__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_30_6__23_  (.A(u_multiplier_STAGE1__0843_ ),
    .B(u_multiplier_STAGE1__0844_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_30_6__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_30_6__24_  (.A1(u_multiplier_STAGE1_acci1_pp_30_6__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_30_6__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_6__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_30_6__25_  (.A(u_multiplier_STAGE1_acci1_pp_30_6__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_30_6__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_6__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_30_6__26_  (.A1(u_multiplier_STAGE1_acci1_pp_30_6__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_30_6__16_ ),
    .ZN(u_multiplier_pp1_30 [6]));
 AOI22_X2 u_multiplier_STAGE1_acci1_pp_30_6__27_  (.A1(u_multiplier_STAGE1__0842_ ),
    .A2(u_multiplier_STAGE1__0841_ ),
    .B1(u_multiplier_STAGE1__0843_ ),
    .B2(u_multiplier_STAGE1__0844_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_30_6__17_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_30_6__28_  (.A1(u_multiplier_STAGE1_acci1_pp_30_6__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_30_6__17_ ),
    .ZN(u_multiplier_pp1_31 [9]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_31_0__21_  (.A1(u_multiplier_STAGE1__0848_ ),
    .A2(u_multiplier_STAGE1__0847_ ),
    .A3(u_multiplier_STAGE1__0849_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_0__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_31_0__22_  (.A(u_multiplier_STAGE1__0848_ ),
    .B(u_multiplier_STAGE1__0847_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_31_0__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_31_0__23_  (.A(u_multiplier_STAGE1__0849_ ),
    .B(u_multiplier_STAGE1__0850_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_31_0__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_31_0__24_  (.A1(u_multiplier_STAGE1_acci1_pp_31_0__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_31_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_31_0__25_  (.A(u_multiplier_STAGE1_acci1_pp_31_0__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_31_0__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_0__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_31_0__26_  (.A1(u_multiplier_STAGE1_acci1_pp_31_0__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_31_0__16_ ),
    .ZN(u_multiplier_pp1_31 [0]));
 AOI22_X1 u_multiplier_STAGE1_acci1_pp_31_0__27_  (.A1(u_multiplier_STAGE1__0848_ ),
    .A2(u_multiplier_STAGE1__0847_ ),
    .B1(u_multiplier_STAGE1__0849_ ),
    .B2(u_multiplier_STAGE1__0850_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_0__17_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_31_0__28_  (.A1(u_multiplier_STAGE1_acci1_pp_31_0__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_31_0__17_ ),
    .ZN(u_multiplier_pp1_32 [15]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_31_1__21_  (.A1(u_multiplier_STAGE1__0852_ ),
    .A2(u_multiplier_STAGE1__0851_ ),
    .A3(u_multiplier_STAGE1__0853_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_1__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_31_1__22_  (.A(u_multiplier_STAGE1__0852_ ),
    .B(u_multiplier_STAGE1__0851_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_31_1__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_31_1__23_  (.A(u_multiplier_STAGE1__0853_ ),
    .B(u_multiplier_STAGE1__0854_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_31_1__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_31_1__24_  (.A1(u_multiplier_STAGE1_acci1_pp_31_1__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_31_1__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_31_1__25_  (.A(u_multiplier_STAGE1_acci1_pp_31_1__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_31_1__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_1__16_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_31_1__26_  (.A1(u_multiplier_STAGE1_acci1_pp_31_1__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_31_1__16_ ),
    .ZN(u_multiplier_pp1_31 [1]));
 AOI22_X1 u_multiplier_STAGE1_acci1_pp_31_1__27_  (.A1(u_multiplier_STAGE1__0852_ ),
    .A2(u_multiplier_STAGE1__0851_ ),
    .B1(u_multiplier_STAGE1__0853_ ),
    .B2(u_multiplier_STAGE1__0854_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_1__17_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_31_1__28_  (.A1(u_multiplier_STAGE1_acci1_pp_31_1__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_31_1__17_ ),
    .ZN(u_multiplier_pp1_32 [14]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_31_2__21_  (.A1(u_multiplier_STAGE1__0856_ ),
    .A2(u_multiplier_STAGE1__0855_ ),
    .A3(u_multiplier_STAGE1__0857_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_2__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_31_2__22_  (.A(u_multiplier_STAGE1__0856_ ),
    .B(u_multiplier_STAGE1__0855_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_31_2__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_31_2__23_  (.A(u_multiplier_STAGE1__0857_ ),
    .B(u_multiplier_STAGE1__0858_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_31_2__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_31_2__24_  (.A1(u_multiplier_STAGE1_acci1_pp_31_2__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_31_2__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_31_2__25_  (.A(u_multiplier_STAGE1_acci1_pp_31_2__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_31_2__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_2__16_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_31_2__26_  (.A1(u_multiplier_STAGE1_acci1_pp_31_2__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_31_2__16_ ),
    .ZN(u_multiplier_pp1_31 [2]));
 AOI22_X1 u_multiplier_STAGE1_acci1_pp_31_2__27_  (.A1(u_multiplier_STAGE1__0856_ ),
    .A2(u_multiplier_STAGE1__0855_ ),
    .B1(u_multiplier_STAGE1__0857_ ),
    .B2(u_multiplier_STAGE1__0858_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_2__17_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_31_2__28_  (.A1(u_multiplier_STAGE1_acci1_pp_31_2__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_31_2__17_ ),
    .ZN(u_multiplier_pp1_32 [13]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_31_3__21_  (.A1(u_multiplier_STAGE1__0860_ ),
    .A2(u_multiplier_STAGE1__0859_ ),
    .A3(u_multiplier_STAGE1__0861_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_3__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_31_3__22_  (.A(u_multiplier_STAGE1__0860_ ),
    .B(u_multiplier_STAGE1__0859_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_31_3__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_31_3__23_  (.A(u_multiplier_STAGE1__0861_ ),
    .B(u_multiplier_STAGE1__0862_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_31_3__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_31_3__24_  (.A1(u_multiplier_STAGE1_acci1_pp_31_3__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_31_3__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_3__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_31_3__25_  (.A(u_multiplier_STAGE1_acci1_pp_31_3__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_31_3__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_3__16_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_31_3__26_  (.A1(u_multiplier_STAGE1_acci1_pp_31_3__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_31_3__16_ ),
    .ZN(u_multiplier_pp1_31 [3]));
 AOI22_X1 u_multiplier_STAGE1_acci1_pp_31_3__27_  (.A1(u_multiplier_STAGE1__0860_ ),
    .A2(u_multiplier_STAGE1__0859_ ),
    .B1(u_multiplier_STAGE1__0861_ ),
    .B2(u_multiplier_STAGE1__0862_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_3__17_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_31_3__28_  (.A1(u_multiplier_STAGE1_acci1_pp_31_3__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_31_3__17_ ),
    .ZN(u_multiplier_pp1_32 [12]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_31_4__21_  (.A1(u_multiplier_STAGE1__0864_ ),
    .A2(u_multiplier_STAGE1__0863_ ),
    .A3(u_multiplier_STAGE1__0865_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_4__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_31_4__22_  (.A(u_multiplier_STAGE1__0864_ ),
    .B(u_multiplier_STAGE1__0863_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_31_4__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_31_4__23_  (.A(u_multiplier_STAGE1__0865_ ),
    .B(u_multiplier_STAGE1__0866_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_31_4__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_31_4__24_  (.A1(u_multiplier_STAGE1_acci1_pp_31_4__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_31_4__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_4__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_31_4__25_  (.A(u_multiplier_STAGE1_acci1_pp_31_4__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_31_4__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_4__16_ ));
 NAND2_X2 u_multiplier_STAGE1_acci1_pp_31_4__26_  (.A1(u_multiplier_STAGE1_acci1_pp_31_4__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_31_4__16_ ),
    .ZN(u_multiplier_pp1_31 [4]));
 AOI22_X1 u_multiplier_STAGE1_acci1_pp_31_4__27_  (.A1(u_multiplier_STAGE1__0864_ ),
    .A2(u_multiplier_STAGE1__0863_ ),
    .B1(u_multiplier_STAGE1__0865_ ),
    .B2(u_multiplier_STAGE1__0866_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_4__17_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_31_4__28_  (.A1(u_multiplier_STAGE1_acci1_pp_31_4__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_31_4__17_ ),
    .ZN(u_multiplier_pp1_32 [11]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_31_5__21_  (.A1(u_multiplier_STAGE1__0868_ ),
    .A2(u_multiplier_STAGE1__0867_ ),
    .A3(u_multiplier_STAGE1__0869_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_5__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_31_5__22_  (.A(u_multiplier_STAGE1__0868_ ),
    .B(u_multiplier_STAGE1__0867_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_31_5__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_31_5__23_  (.A(u_multiplier_STAGE1__0869_ ),
    .B(u_multiplier_STAGE1__0870_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_31_5__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_31_5__24_  (.A1(u_multiplier_STAGE1_acci1_pp_31_5__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_31_5__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_5__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_31_5__25_  (.A(u_multiplier_STAGE1_acci1_pp_31_5__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_31_5__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_5__16_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_31_5__26_  (.A1(u_multiplier_STAGE1_acci1_pp_31_5__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_31_5__16_ ),
    .ZN(u_multiplier_pp1_31 [5]));
 AOI22_X1 u_multiplier_STAGE1_acci1_pp_31_5__27_  (.A1(u_multiplier_STAGE1__0868_ ),
    .A2(u_multiplier_STAGE1__0867_ ),
    .B1(u_multiplier_STAGE1__0869_ ),
    .B2(u_multiplier_STAGE1__0870_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_5__17_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_31_5__28_  (.A1(u_multiplier_STAGE1_acci1_pp_31_5__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_31_5__17_ ),
    .ZN(u_multiplier_pp1_32 [10]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_31_6__21_  (.A1(u_multiplier_STAGE1__0872_ ),
    .A2(u_multiplier_STAGE1__0871_ ),
    .A3(u_multiplier_STAGE1__0873_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_6__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_31_6__22_  (.A(u_multiplier_STAGE1__0872_ ),
    .B(u_multiplier_STAGE1__0871_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_31_6__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_31_6__23_  (.A(u_multiplier_STAGE1__0873_ ),
    .B(u_multiplier_STAGE1__0874_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_31_6__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_31_6__24_  (.A1(u_multiplier_STAGE1_acci1_pp_31_6__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_31_6__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_6__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_31_6__25_  (.A(u_multiplier_STAGE1_acci1_pp_31_6__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_31_6__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_6__16_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_31_6__26_  (.A1(u_multiplier_STAGE1_acci1_pp_31_6__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_31_6__16_ ),
    .ZN(u_multiplier_pp1_31 [6]));
 AOI22_X1 u_multiplier_STAGE1_acci1_pp_31_6__27_  (.A1(u_multiplier_STAGE1__0872_ ),
    .A2(u_multiplier_STAGE1__0871_ ),
    .B1(u_multiplier_STAGE1__0873_ ),
    .B2(u_multiplier_STAGE1__0874_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_6__17_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_31_6__28_  (.A1(u_multiplier_STAGE1_acci1_pp_31_6__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_31_6__17_ ),
    .ZN(u_multiplier_pp1_32 [9]));
 NAND3_X1 u_multiplier_STAGE1_acci1_pp_31_7__21_  (.A1(u_multiplier_STAGE1__0876_ ),
    .A2(u_multiplier_STAGE1__0875_ ),
    .A3(u_multiplier_STAGE1__0877_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_7__18_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_31_7__22_  (.A(u_multiplier_STAGE1__0876_ ),
    .B(u_multiplier_STAGE1__0875_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_31_7__19_ ));
 XOR2_X2 u_multiplier_STAGE1_acci1_pp_31_7__23_  (.A(u_multiplier_STAGE1__0877_ ),
    .B(u_multiplier_STAGE1__0878_ ),
    .Z(u_multiplier_STAGE1_acci1_pp_31_7__20_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_31_7__24_  (.A1(u_multiplier_STAGE1_acci1_pp_31_7__19_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_31_7__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_7__15_ ));
 XNOR2_X1 u_multiplier_STAGE1_acci1_pp_31_7__25_  (.A(u_multiplier_STAGE1_acci1_pp_31_7__19_ ),
    .B(u_multiplier_STAGE1_acci1_pp_31_7__20_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_7__16_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_31_7__26_  (.A1(u_multiplier_STAGE1_acci1_pp_31_7__18_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_31_7__16_ ),
    .ZN(u_multiplier_pp1_31 [7]));
 AOI22_X1 u_multiplier_STAGE1_acci1_pp_31_7__27_  (.A1(u_multiplier_STAGE1__0876_ ),
    .A2(u_multiplier_STAGE1__0875_ ),
    .B1(u_multiplier_STAGE1__0877_ ),
    .B2(u_multiplier_STAGE1__0878_ ),
    .ZN(u_multiplier_STAGE1_acci1_pp_31_7__17_ ));
 NAND2_X1 u_multiplier_STAGE1_acci1_pp_31_7__28_  (.A1(u_multiplier_STAGE1_acci1_pp_31_7__15_ ),
    .A2(u_multiplier_STAGE1_acci1_pp_31_7__17_ ),
    .ZN(u_multiplier_pp1_32 [8]));
 LOGIC0_X1 u_multiplier_STAGE2_E_4_2_pp2_32_1__18__125  (.Z(net125));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_32_1__18_  (.A(net125),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_1__19_  (.A1(u_multiplier_pp1_32 [1]),
    .A2(u_multiplier_pp1_32 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_1__20_  (.A(u_multiplier_pp1_32 [1]),
    .B(u_multiplier_pp1_32 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_32_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_1__21_  (.A1(u_multiplier_pp1_32 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_32_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_1__22_  (.A(u_multiplier_pp1_32 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_32_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_32_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_1__23_  (.A1(u_multiplier_pp1_32 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_32_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_1__24_  (.A(u_multiplier_pp1_32 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_32_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_1__25_  (.A(net126),
    .B(u_multiplier_STAGE2_E_4_2_pp2_32_1__16_ ),
    .ZN(u_multiplier_pp2_32 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_32_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_32_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_32_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_32_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_32_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_32_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_32_1__17_ ),
    .ZN(u_multiplier_pp2_33 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_32_2__18_  (.A(net127),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_2__19_  (.A1(u_multiplier_pp1_32 [5]),
    .A2(u_multiplier_pp1_32 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_2__20_  (.A(u_multiplier_pp1_32 [5]),
    .B(u_multiplier_pp1_32 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_32_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_2__21_  (.A1(u_multiplier_pp1_32 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_32_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_2__22_  (.A(u_multiplier_pp1_32 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_32_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_32_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_2__23_  (.A1(u_multiplier_pp1_32 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_32_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_2__24_  (.A(u_multiplier_pp1_32 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_32_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_2__25_  (.A(net128),
    .B(u_multiplier_STAGE2_E_4_2_pp2_32_2__16_ ),
    .ZN(u_multiplier_pp2_32 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_32_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_32_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_32_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_32_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_32_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_32_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_32_2__17_ ),
    .ZN(u_multiplier_pp2_33 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_32_3__18_  (.A(net129),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_3__19_  (.A1(u_multiplier_pp1_32 [9]),
    .A2(u_multiplier_pp1_32 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_3__20_  (.A(u_multiplier_pp1_32 [9]),
    .B(u_multiplier_pp1_32 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_32_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_3__21_  (.A1(u_multiplier_pp1_32 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_32_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_3__22_  (.A(u_multiplier_pp1_32 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_32_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_32_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_3__23_  (.A1(u_multiplier_pp1_32 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_32_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_3__24_  (.A(u_multiplier_pp1_32 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_32_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_3__25_  (.A(net130),
    .B(u_multiplier_STAGE2_E_4_2_pp2_32_3__16_ ),
    .ZN(u_multiplier_pp2_32 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_32_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_32_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_32_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_32_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_32_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_32_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_32_3__17_ ),
    .ZN(u_multiplier_pp2_33 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_32_4__18_  (.A(net131),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_4__19_  (.A1(u_multiplier_pp1_32 [13]),
    .A2(u_multiplier_pp1_32 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_4__20_  (.A(u_multiplier_pp1_32 [13]),
    .B(u_multiplier_pp1_32 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_32_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_4__21_  (.A1(u_multiplier_pp1_32 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_32_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_4__22_  (.A(u_multiplier_pp1_32 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_32_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_32_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_32_4__23_  (.A1(u_multiplier_pp1_32 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_32_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_4__24_  (.A(u_multiplier_pp1_32 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_32_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_32_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_4__25_  (.A(net132),
    .B(u_multiplier_STAGE2_E_4_2_pp2_32_4__16_ ),
    .ZN(u_multiplier_pp2_32 [0]));
 NAND2_X2 u_multiplier_STAGE2_E_4_2_pp2_32_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_32_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_32_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_32_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_32_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_32_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_32_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_32_4__17_ ),
    .ZN(u_multiplier_pp2_33 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_33_1__18_  (.A(u_multiplier_STAGE2_pp2_32_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_1__19_  (.A1(u_multiplier_pp1_33 [1]),
    .A2(u_multiplier_pp1_33 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_1__20_  (.A(u_multiplier_pp1_33 [1]),
    .B(u_multiplier_pp1_33 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_33_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_1__21_  (.A1(u_multiplier_pp1_33 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_33_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_1__22_  (.A(u_multiplier_pp1_33 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_33_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_33_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_1__23_  (.A1(u_multiplier_pp1_33 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_33_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_1__24_  (.A(u_multiplier_pp1_33 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_33_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_1__25_  (.A(u_multiplier_STAGE2_pp2_32_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_33_1__16_ ),
    .ZN(u_multiplier_pp2_33 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_33_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_33_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_33_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE2_E_4_2_pp2_33_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_33_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_33_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_33_1__17_ ),
    .ZN(u_multiplier_pp2_34 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_33_2__18_  (.A(u_multiplier_STAGE2_pp2_32_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_2__19_  (.A1(u_multiplier_pp1_33 [5]),
    .A2(u_multiplier_pp1_33 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_2__20_  (.A(u_multiplier_pp1_33 [5]),
    .B(u_multiplier_pp1_33 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_33_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_2__21_  (.A1(u_multiplier_pp1_33 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_33_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_2__22_  (.A(u_multiplier_pp1_33 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_33_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_33_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_2__23_  (.A1(u_multiplier_pp1_33 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_33_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_2__24_  (.A(u_multiplier_pp1_33 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_33_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_2__25_  (.A(u_multiplier_STAGE2_pp2_32_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_33_2__16_ ),
    .ZN(u_multiplier_pp2_33 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_33_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_33_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_33_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_33_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_33_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_33_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_33_2__17_ ),
    .ZN(u_multiplier_pp2_34 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_33_3__18_  (.A(u_multiplier_STAGE2_pp2_32_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_3__19_  (.A1(u_multiplier_pp1_33 [9]),
    .A2(u_multiplier_pp1_33 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_3__20_  (.A(u_multiplier_pp1_33 [9]),
    .B(u_multiplier_pp1_33 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_33_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_3__21_  (.A1(u_multiplier_pp1_33 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_33_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_3__22_  (.A(u_multiplier_pp1_33 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_33_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_33_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_3__23_  (.A1(u_multiplier_pp1_33 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_33_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_3__24_  (.A(u_multiplier_pp1_33 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_33_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_3__25_  (.A(u_multiplier_STAGE2_pp2_32_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_33_3__16_ ),
    .ZN(u_multiplier_pp2_33 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_33_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_33_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_33_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_33_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_33_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_33_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_33_3__17_ ),
    .ZN(u_multiplier_pp2_34 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_33_4__18_  (.A(u_multiplier_STAGE2_pp2_32_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_4__19_  (.A1(u_multiplier_pp1_33 [13]),
    .A2(u_multiplier_pp1_33 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_4__20_  (.A(u_multiplier_pp1_33 [13]),
    .B(u_multiplier_pp1_33 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_33_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_4__21_  (.A1(u_multiplier_pp1_33 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_33_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_4__22_  (.A(u_multiplier_pp1_33 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_33_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_33_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_4__23_  (.A1(u_multiplier_pp1_33 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_33_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_4__24_  (.A(u_multiplier_pp1_33 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_33_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_33_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_33_4__25_  (.A(u_multiplier_STAGE2_pp2_32_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_33_4__16_ ),
    .ZN(u_multiplier_pp2_33 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_33_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_33_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_33_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_33_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_33_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_33_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_33_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_33_4__17_ ),
    .ZN(u_multiplier_pp2_34 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_34_1__18_  (.A(u_multiplier_STAGE2_pp2_33_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_1__19_  (.A1(u_multiplier_pp1_34 [1]),
    .A2(u_multiplier_pp1_34 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_1__20_  (.A(u_multiplier_pp1_34 [1]),
    .B(u_multiplier_pp1_34 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_34_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_1__21_  (.A1(u_multiplier_pp1_34 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_34_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_1__22_  (.A(u_multiplier_pp1_34 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_34_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_34_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_1__23_  (.A1(u_multiplier_pp1_34 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_34_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_1__24_  (.A(u_multiplier_pp1_34 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_34_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_1__25_  (.A(u_multiplier_STAGE2_pp2_33_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_34_1__16_ ),
    .ZN(u_multiplier_pp2_34 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_34_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_34_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_34_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_34_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_34_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_34_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_34_1__17_ ),
    .ZN(u_multiplier_pp2_35 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_34_2__18_  (.A(u_multiplier_STAGE2_pp2_33_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_2__19_  (.A1(u_multiplier_pp1_34 [5]),
    .A2(u_multiplier_pp1_34 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_2__20_  (.A(u_multiplier_pp1_34 [5]),
    .B(u_multiplier_pp1_34 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_34_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_2__21_  (.A1(u_multiplier_pp1_34 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_34_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_2__22_  (.A(u_multiplier_pp1_34 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_34_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_34_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_2__23_  (.A1(u_multiplier_pp1_34 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_34_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_2__24_  (.A(u_multiplier_pp1_34 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_34_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_2__25_  (.A(u_multiplier_STAGE2_pp2_33_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_34_2__16_ ),
    .ZN(u_multiplier_pp2_34 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_34_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_34_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_34_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_34_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_34_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_34_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_34_2__17_ ),
    .ZN(u_multiplier_pp2_35 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_34_3__18_  (.A(u_multiplier_STAGE2_pp2_33_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_3__19_  (.A1(u_multiplier_pp1_34 [9]),
    .A2(u_multiplier_pp1_34 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_3__20_  (.A(u_multiplier_pp1_34 [9]),
    .B(u_multiplier_pp1_34 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_34_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_3__21_  (.A1(u_multiplier_pp1_34 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_34_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_3__22_  (.A(u_multiplier_pp1_34 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_34_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_34_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_3__23_  (.A1(u_multiplier_pp1_34 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_34_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_3__24_  (.A(u_multiplier_pp1_34 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_34_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_3__25_  (.A(u_multiplier_STAGE2_pp2_33_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_34_3__16_ ),
    .ZN(u_multiplier_pp2_34 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_34_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_34_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_34_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_34_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_34_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_34_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_34_3__17_ ),
    .ZN(u_multiplier_pp2_35 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_34_4__18_  (.A(u_multiplier_STAGE2_pp2_33_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_4__19_  (.A1(u_multiplier_pp1_34 [13]),
    .A2(u_multiplier_pp1_34 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_4__20_  (.A(u_multiplier_pp1_34 [13]),
    .B(u_multiplier_pp1_34 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_34_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_4__21_  (.A1(u_multiplier_pp1_34 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_34_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_4__22_  (.A(u_multiplier_pp1_34 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_34_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_34_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_4__23_  (.A1(u_multiplier_pp1_34 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_34_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_4__24_  (.A(u_multiplier_pp1_34 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_34_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_34_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_34_4__25_  (.A(u_multiplier_STAGE2_pp2_33_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_34_4__16_ ),
    .ZN(u_multiplier_pp2_34 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_34_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_34_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_34_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_34_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_34_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_34_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_34_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_34_4__17_ ),
    .ZN(u_multiplier_pp2_35 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_35_1__18_  (.A(u_multiplier_STAGE2_pp2_34_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_1__19_  (.A1(u_multiplier_pp1_35 [1]),
    .A2(u_multiplier_pp1_35 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_1__20_  (.A(u_multiplier_pp1_35 [1]),
    .B(u_multiplier_pp1_35 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_35_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_1__21_  (.A1(u_multiplier_pp1_35 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_35_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_1__22_  (.A(u_multiplier_pp1_35 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_35_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_35_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_1__23_  (.A1(u_multiplier_pp1_35 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_35_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_1__24_  (.A(u_multiplier_pp1_35 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_35_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_1__25_  (.A(u_multiplier_STAGE2_pp2_34_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_35_1__16_ ),
    .ZN(u_multiplier_pp2_35 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_35_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_35_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_35_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_35_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_35_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_35_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_35_1__17_ ),
    .ZN(u_multiplier_pp2_36 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_35_2__18_  (.A(u_multiplier_STAGE2_pp2_34_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_2__19_  (.A1(u_multiplier_pp1_35 [5]),
    .A2(u_multiplier_pp1_35 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_2__20_  (.A(u_multiplier_pp1_35 [5]),
    .B(u_multiplier_pp1_35 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_35_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_2__21_  (.A1(u_multiplier_pp1_35 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_35_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_2__22_  (.A(u_multiplier_pp1_35 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_35_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_35_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_2__23_  (.A1(u_multiplier_pp1_35 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_35_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_2__24_  (.A(u_multiplier_pp1_35 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_35_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_2__25_  (.A(u_multiplier_STAGE2_pp2_34_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_35_2__16_ ),
    .ZN(u_multiplier_pp2_35 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_35_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_35_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_35_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_35_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_35_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_35_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_35_2__17_ ),
    .ZN(u_multiplier_pp2_36 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_35_3__18_  (.A(u_multiplier_STAGE2_pp2_34_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_3__19_  (.A1(u_multiplier_pp1_35 [9]),
    .A2(u_multiplier_pp1_35 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_3__20_  (.A(u_multiplier_pp1_35 [9]),
    .B(u_multiplier_pp1_35 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_35_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_3__21_  (.A1(u_multiplier_pp1_35 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_35_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_3__22_  (.A(u_multiplier_pp1_35 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_35_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_35_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_3__23_  (.A1(u_multiplier_pp1_35 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_35_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_3__24_  (.A(u_multiplier_pp1_35 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_35_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_3__25_  (.A(u_multiplier_STAGE2_pp2_34_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_35_3__16_ ),
    .ZN(u_multiplier_pp2_35 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_35_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_35_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_35_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_35_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_35_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_35_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_35_3__17_ ),
    .ZN(u_multiplier_pp2_36 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_35_4__18_  (.A(u_multiplier_STAGE2_pp2_34_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_4__19_  (.A1(u_multiplier_pp1_35 [13]),
    .A2(u_multiplier_pp1_35 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_4__20_  (.A(u_multiplier_pp1_35 [13]),
    .B(u_multiplier_pp1_35 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_35_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_4__21_  (.A1(u_multiplier_pp1_35 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_35_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_4__22_  (.A(u_multiplier_pp1_35 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_35_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_35_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_4__23_  (.A1(u_multiplier_pp1_35 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_35_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_4__24_  (.A(u_multiplier_pp1_35 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_35_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_35_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_35_4__25_  (.A(u_multiplier_STAGE2_pp2_34_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_35_4__16_ ),
    .ZN(u_multiplier_pp2_35 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_35_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_35_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_35_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_35_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_35_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_35_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_35_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_35_4__17_ ),
    .ZN(u_multiplier_pp2_36 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_36_1__18_  (.A(u_multiplier_STAGE2_pp2_35_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_1__19_  (.A1(u_multiplier_pp1_36 [1]),
    .A2(u_multiplier_pp1_36 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_1__20_  (.A(u_multiplier_pp1_36 [1]),
    .B(u_multiplier_pp1_36 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_36_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_1__21_  (.A1(u_multiplier_pp1_36 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_36_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_1__22_  (.A(u_multiplier_pp1_36 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_36_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_36_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_1__23_  (.A1(u_multiplier_pp1_36 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_36_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_1__24_  (.A(u_multiplier_pp1_36 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_36_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_1__25_  (.A(u_multiplier_STAGE2_pp2_35_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_36_1__16_ ),
    .ZN(u_multiplier_pp2_36 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_36_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_36_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_36_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_36_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_36_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_36_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_36_1__17_ ),
    .ZN(u_multiplier_pp2_37 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_36_2__18_  (.A(u_multiplier_STAGE2_pp2_35_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_2__19_  (.A1(u_multiplier_pp1_36 [5]),
    .A2(u_multiplier_pp1_36 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_2__20_  (.A(u_multiplier_pp1_36 [5]),
    .B(u_multiplier_pp1_36 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_36_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_2__21_  (.A1(u_multiplier_pp1_36 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_36_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_2__22_  (.A(u_multiplier_pp1_36 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_36_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_36_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_2__23_  (.A1(u_multiplier_pp1_36 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_36_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_2__24_  (.A(u_multiplier_pp1_36 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_36_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_2__25_  (.A(u_multiplier_STAGE2_pp2_35_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_36_2__16_ ),
    .ZN(u_multiplier_pp2_36 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_36_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_36_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_36_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_36_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_36_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_36_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_36_2__17_ ),
    .ZN(u_multiplier_pp2_37 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_36_3__18_  (.A(u_multiplier_STAGE2_pp2_35_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_3__19_  (.A1(u_multiplier_pp1_36 [9]),
    .A2(u_multiplier_pp1_36 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_3__20_  (.A(u_multiplier_pp1_36 [9]),
    .B(u_multiplier_pp1_36 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_36_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_3__21_  (.A1(u_multiplier_pp1_36 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_36_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_3__22_  (.A(u_multiplier_pp1_36 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_36_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_36_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_3__23_  (.A1(u_multiplier_pp1_36 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_36_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_3__24_  (.A(u_multiplier_pp1_36 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_36_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_3__25_  (.A(u_multiplier_STAGE2_pp2_35_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_36_3__16_ ),
    .ZN(u_multiplier_pp2_36 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_36_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_36_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_36_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_36_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_36_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_36_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_36_3__17_ ),
    .ZN(u_multiplier_pp2_37 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_36_4__18_  (.A(u_multiplier_STAGE2_pp2_35_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_4__19_  (.A1(u_multiplier_pp1_36 [13]),
    .A2(u_multiplier_pp1_36 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_4__20_  (.A(u_multiplier_pp1_36 [13]),
    .B(u_multiplier_pp1_36 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_36_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_4__21_  (.A1(u_multiplier_pp1_36 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_36_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_4__22_  (.A(u_multiplier_pp1_36 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_36_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_36_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_4__23_  (.A1(u_multiplier_pp1_36 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_36_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_4__24_  (.A(u_multiplier_pp1_36 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_36_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_36_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_36_4__25_  (.A(u_multiplier_STAGE2_pp2_35_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_36_4__16_ ),
    .ZN(u_multiplier_pp2_36 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_36_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_36_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_36_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_36_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_36_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_36_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_36_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_36_4__17_ ),
    .ZN(u_multiplier_pp2_37 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_37_1__18_  (.A(u_multiplier_STAGE2_pp2_36_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_1__19_  (.A1(u_multiplier_pp1_37 [1]),
    .A2(u_multiplier_pp1_37 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_1__20_  (.A(u_multiplier_pp1_37 [1]),
    .B(u_multiplier_pp1_37 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_37_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_1__21_  (.A1(u_multiplier_pp1_37 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_37_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_1__22_  (.A(u_multiplier_pp1_37 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_37_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_37_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_1__23_  (.A1(u_multiplier_pp1_37 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_37_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_1__24_  (.A(u_multiplier_pp1_37 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_37_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_1__25_  (.A(u_multiplier_STAGE2_pp2_36_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_37_1__16_ ),
    .ZN(u_multiplier_pp2_37 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_37_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_37_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_37_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_37_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_37_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_37_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_37_1__17_ ),
    .ZN(u_multiplier_pp2_38 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_37_2__18_  (.A(u_multiplier_STAGE2_pp2_36_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_2__19_  (.A1(u_multiplier_pp1_37 [5]),
    .A2(u_multiplier_pp1_37 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_2__20_  (.A(u_multiplier_pp1_37 [5]),
    .B(u_multiplier_pp1_37 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_37_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_2__21_  (.A1(u_multiplier_pp1_37 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_37_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_2__22_  (.A(u_multiplier_pp1_37 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_37_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_37_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_2__23_  (.A1(u_multiplier_pp1_37 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_37_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_2__24_  (.A(u_multiplier_pp1_37 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_37_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_2__25_  (.A(u_multiplier_STAGE2_pp2_36_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_37_2__16_ ),
    .ZN(u_multiplier_pp2_37 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_37_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_37_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_37_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_37_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_37_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_37_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_37_2__17_ ),
    .ZN(u_multiplier_pp2_38 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_37_3__18_  (.A(u_multiplier_STAGE2_pp2_36_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_3__19_  (.A1(u_multiplier_pp1_37 [9]),
    .A2(u_multiplier_pp1_37 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_3__20_  (.A(u_multiplier_pp1_37 [9]),
    .B(u_multiplier_pp1_37 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_37_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_3__21_  (.A1(u_multiplier_pp1_37 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_37_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_3__22_  (.A(u_multiplier_pp1_37 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_37_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_37_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_3__23_  (.A1(u_multiplier_pp1_37 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_37_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_3__24_  (.A(u_multiplier_pp1_37 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_37_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_3__25_  (.A(u_multiplier_STAGE2_pp2_36_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_37_3__16_ ),
    .ZN(u_multiplier_pp2_37 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_37_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_37_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_37_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_37_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_37_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_37_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_37_3__17_ ),
    .ZN(u_multiplier_pp2_38 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_37_4__18_  (.A(u_multiplier_STAGE2_pp2_36_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_4__19_  (.A1(u_multiplier_pp1_37 [13]),
    .A2(u_multiplier_pp1_37 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_4__20_  (.A(u_multiplier_pp1_37 [13]),
    .B(u_multiplier_pp1_37 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_37_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_4__21_  (.A1(u_multiplier_pp1_37 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_37_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_4__22_  (.A(u_multiplier_pp1_37 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_37_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_37_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_4__23_  (.A1(u_multiplier_pp1_37 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_37_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_4__24_  (.A(u_multiplier_pp1_37 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_37_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_37_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_37_4__25_  (.A(u_multiplier_STAGE2_pp2_36_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_37_4__16_ ),
    .ZN(u_multiplier_pp2_37 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_37_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_37_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_37_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_37_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_37_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_37_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_37_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_37_4__17_ ),
    .ZN(u_multiplier_pp2_38 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_38_1__18_  (.A(u_multiplier_STAGE2_pp2_37_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_1__19_  (.A1(u_multiplier_pp1_38 [1]),
    .A2(u_multiplier_pp1_38 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_1__20_  (.A(u_multiplier_pp1_38 [1]),
    .B(u_multiplier_pp1_38 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_38_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_1__21_  (.A1(u_multiplier_pp1_38 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_38_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_1__22_  (.A(u_multiplier_pp1_38 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_38_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_38_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_1__23_  (.A1(u_multiplier_pp1_38 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_38_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_1__24_  (.A(u_multiplier_pp1_38 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_38_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_1__25_  (.A(u_multiplier_STAGE2_pp2_37_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_38_1__16_ ),
    .ZN(u_multiplier_pp2_38 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_38_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_38_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_38_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_38_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_38_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_38_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_38_1__17_ ),
    .ZN(u_multiplier_pp2_39 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_38_2__18_  (.A(u_multiplier_STAGE2_pp2_37_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_2__19_  (.A1(u_multiplier_pp1_38 [5]),
    .A2(u_multiplier_pp1_38 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_2__20_  (.A(u_multiplier_pp1_38 [5]),
    .B(u_multiplier_pp1_38 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_38_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_2__21_  (.A1(u_multiplier_pp1_38 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_38_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_2__22_  (.A(u_multiplier_pp1_38 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_38_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_38_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_2__23_  (.A1(u_multiplier_pp1_38 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_38_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_2__24_  (.A(u_multiplier_pp1_38 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_38_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_2__25_  (.A(u_multiplier_STAGE2_pp2_37_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_38_2__16_ ),
    .ZN(u_multiplier_pp2_38 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_38_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_38_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_38_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_38_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_38_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_38_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_38_2__17_ ),
    .ZN(u_multiplier_pp2_39 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_38_3__18_  (.A(u_multiplier_STAGE2_pp2_37_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_3__19_  (.A1(u_multiplier_pp1_38 [9]),
    .A2(u_multiplier_pp1_38 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_3__20_  (.A(u_multiplier_pp1_38 [9]),
    .B(u_multiplier_pp1_38 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_38_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_3__21_  (.A1(u_multiplier_pp1_38 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_38_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_3__22_  (.A(u_multiplier_pp1_38 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_38_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_38_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_3__23_  (.A1(u_multiplier_pp1_38 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_38_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_3__24_  (.A(u_multiplier_pp1_38 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_38_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_3__25_  (.A(u_multiplier_STAGE2_pp2_37_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_38_3__16_ ),
    .ZN(u_multiplier_pp2_38 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_38_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_38_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_38_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_38_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_38_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_38_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_38_3__17_ ),
    .ZN(u_multiplier_pp2_39 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_38_4__18_  (.A(u_multiplier_STAGE2_pp2_37_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_4__19_  (.A1(u_multiplier_pp1_38 [13]),
    .A2(u_multiplier_pp1_38 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_4__20_  (.A(u_multiplier_pp1_38 [13]),
    .B(u_multiplier_pp1_38 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_38_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_4__21_  (.A1(u_multiplier_pp1_38 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_38_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_4__22_  (.A(u_multiplier_pp1_38 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_38_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_38_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_4__23_  (.A1(u_multiplier_pp1_38 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_38_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_4__24_  (.A(u_multiplier_pp1_38 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_38_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_38_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_38_4__25_  (.A(u_multiplier_STAGE2_pp2_37_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_38_4__16_ ),
    .ZN(u_multiplier_pp2_38 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_38_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_38_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_38_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_38_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_38_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_38_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_38_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_38_4__17_ ),
    .ZN(u_multiplier_pp2_39 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_39_1__18_  (.A(u_multiplier_STAGE2_pp2_38_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_1__19_  (.A1(u_multiplier_pp1_39 [1]),
    .A2(u_multiplier_pp1_39 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_1__20_  (.A(u_multiplier_pp1_39 [1]),
    .B(u_multiplier_pp1_39 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_39_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_1__21_  (.A1(u_multiplier_pp1_39 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_39_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_1__22_  (.A(u_multiplier_pp1_39 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_39_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_39_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_1__23_  (.A1(u_multiplier_pp1_39 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_39_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_1__24_  (.A(u_multiplier_pp1_39 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_39_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_1__25_  (.A(u_multiplier_STAGE2_pp2_38_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_39_1__16_ ),
    .ZN(u_multiplier_pp2_39 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_39_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_39_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_39_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_39_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_39_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_39_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_39_1__17_ ),
    .ZN(u_multiplier_pp2_40 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_39_2__18_  (.A(u_multiplier_STAGE2_pp2_38_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_2__19_  (.A1(u_multiplier_pp1_39 [5]),
    .A2(u_multiplier_pp1_39 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_2__20_  (.A(u_multiplier_pp1_39 [5]),
    .B(u_multiplier_pp1_39 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_39_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_2__21_  (.A1(u_multiplier_pp1_39 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_39_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_2__22_  (.A(u_multiplier_pp1_39 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_39_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_39_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_2__23_  (.A1(u_multiplier_pp1_39 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_39_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_2__24_  (.A(u_multiplier_pp1_39 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_39_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_2__25_  (.A(u_multiplier_STAGE2_pp2_38_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_39_2__16_ ),
    .ZN(u_multiplier_pp2_39 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_39_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_39_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_39_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_39_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_39_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_39_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_39_2__17_ ),
    .ZN(u_multiplier_pp2_40 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_39_3__18_  (.A(u_multiplier_STAGE2_pp2_38_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_3__19_  (.A1(u_multiplier_pp1_39 [9]),
    .A2(u_multiplier_pp1_39 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_3__20_  (.A(u_multiplier_pp1_39 [9]),
    .B(u_multiplier_pp1_39 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_39_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_3__21_  (.A1(u_multiplier_pp1_39 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_39_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_3__22_  (.A(u_multiplier_pp1_39 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_39_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_39_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_3__23_  (.A1(u_multiplier_pp1_39 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_39_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_3__24_  (.A(u_multiplier_pp1_39 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_39_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_3__25_  (.A(u_multiplier_STAGE2_pp2_38_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_39_3__16_ ),
    .ZN(u_multiplier_pp2_39 [1]));
 NAND2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_39_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_39_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_39_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_39_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_39_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_39_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_39_3__17_ ),
    .ZN(u_multiplier_pp2_40 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_39_4__18_  (.A(u_multiplier_STAGE2_pp2_38_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_4__19_  (.A1(u_multiplier_pp1_39 [13]),
    .A2(u_multiplier_pp1_39 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_4__20_  (.A(u_multiplier_pp1_39 [13]),
    .B(u_multiplier_pp1_39 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_39_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_4__21_  (.A1(u_multiplier_pp1_39 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_39_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_4__22_  (.A(u_multiplier_pp1_39 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_39_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_39_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_4__23_  (.A1(u_multiplier_pp1_39 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_39_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_4__24_  (.A(u_multiplier_pp1_39 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_39_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_39_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_39_4__25_  (.A(u_multiplier_STAGE2_pp2_38_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_39_4__16_ ),
    .ZN(u_multiplier_pp2_39 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_39_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_39_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_39_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_39_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_39_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_39_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_39_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_39_4__17_ ),
    .ZN(u_multiplier_pp2_40 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_40_1__18_  (.A(u_multiplier_STAGE2_pp2_39_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_1__19_  (.A1(u_multiplier_pp1_40 [1]),
    .A2(u_multiplier_pp1_40 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_1__20_  (.A(u_multiplier_pp1_40 [1]),
    .B(u_multiplier_pp1_40 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_40_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_1__21_  (.A1(u_multiplier_pp1_40 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_40_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_1__22_  (.A(u_multiplier_pp1_40 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_40_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_40_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_1__23_  (.A1(u_multiplier_pp1_40 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_40_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_1__24_  (.A(u_multiplier_pp1_40 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_40_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_1__25_  (.A(u_multiplier_STAGE2_pp2_39_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_40_1__16_ ),
    .ZN(u_multiplier_pp2_40 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_40_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_40_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_40_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE2_E_4_2_pp2_40_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_40_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_40_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_40_1__17_ ),
    .ZN(u_multiplier_pp2_41 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_40_2__18_  (.A(u_multiplier_STAGE2_pp2_39_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_2__19_  (.A1(u_multiplier_pp1_40 [5]),
    .A2(u_multiplier_pp1_40 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_2__20_  (.A(u_multiplier_pp1_40 [5]),
    .B(u_multiplier_pp1_40 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_40_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_2__21_  (.A1(u_multiplier_pp1_40 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_40_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_2__22_  (.A(u_multiplier_pp1_40 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_40_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_40_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_2__23_  (.A1(u_multiplier_pp1_40 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_40_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_2__24_  (.A(u_multiplier_pp1_40 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_40_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_2__25_  (.A(u_multiplier_STAGE2_pp2_39_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_40_2__16_ ),
    .ZN(u_multiplier_pp2_40 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_40_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_40_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_40_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_40_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_40_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_40_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_40_2__17_ ),
    .ZN(u_multiplier_pp2_41 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_40_3__18_  (.A(u_multiplier_STAGE2_pp2_39_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_3__19_  (.A1(u_multiplier_pp1_40 [9]),
    .A2(u_multiplier_pp1_40 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_3__20_  (.A(u_multiplier_pp1_40 [9]),
    .B(u_multiplier_pp1_40 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_40_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_3__21_  (.A1(u_multiplier_pp1_40 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_40_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_3__22_  (.A(u_multiplier_pp1_40 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_40_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_40_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_3__23_  (.A1(u_multiplier_pp1_40 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_40_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_3__24_  (.A(u_multiplier_pp1_40 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_40_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_3__25_  (.A(u_multiplier_STAGE2_pp2_39_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_40_3__16_ ),
    .ZN(u_multiplier_pp2_40 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_40_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_40_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_40_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_40_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_40_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_40_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_40_3__17_ ),
    .ZN(u_multiplier_pp2_41 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_40_4__18_  (.A(u_multiplier_STAGE2_pp2_39_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_4__19_  (.A1(u_multiplier_pp1_40 [13]),
    .A2(u_multiplier_pp1_40 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_4__20_  (.A(u_multiplier_pp1_40 [13]),
    .B(u_multiplier_pp1_40 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_40_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_4__21_  (.A1(u_multiplier_pp1_40 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_40_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_4__22_  (.A(u_multiplier_pp1_40 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_40_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_40_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_4__23_  (.A1(u_multiplier_pp1_40 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_40_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_4__24_  (.A(u_multiplier_pp1_40 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_40_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_40_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_40_4__25_  (.A(u_multiplier_STAGE2_pp2_39_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_40_4__16_ ),
    .ZN(u_multiplier_pp2_40 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_40_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_40_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_40_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_40_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_40_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_40_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_40_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_40_4__17_ ),
    .ZN(u_multiplier_pp2_41 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_41_1__18_  (.A(u_multiplier_STAGE2_pp2_40_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_1__19_  (.A1(u_multiplier_pp1_41 [1]),
    .A2(u_multiplier_pp1_41 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_1__20_  (.A(u_multiplier_pp1_41 [1]),
    .B(u_multiplier_pp1_41 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_41_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_1__21_  (.A1(u_multiplier_pp1_41 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_41_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_1__22_  (.A(u_multiplier_pp1_41 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_41_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_41_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_1__23_  (.A1(u_multiplier_pp1_41 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_41_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_1__24_  (.A(u_multiplier_pp1_41 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_41_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_1__25_  (.A(u_multiplier_STAGE2_pp2_40_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_41_1__16_ ),
    .ZN(u_multiplier_pp2_41 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_41_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_41_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_41_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_41_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_41_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_41_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_41_1__17_ ),
    .ZN(u_multiplier_pp2_42 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_41_2__18_  (.A(u_multiplier_STAGE2_pp2_40_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_2__19_  (.A1(u_multiplier_pp1_41 [5]),
    .A2(u_multiplier_pp1_41 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_2__20_  (.A(u_multiplier_pp1_41 [5]),
    .B(u_multiplier_pp1_41 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_41_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_2__21_  (.A1(u_multiplier_pp1_41 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_41_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_2__22_  (.A(u_multiplier_pp1_41 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_41_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_41_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_2__23_  (.A1(u_multiplier_pp1_41 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_41_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_2__24_  (.A(u_multiplier_pp1_41 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_41_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_2__25_  (.A(u_multiplier_STAGE2_pp2_40_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_41_2__16_ ),
    .ZN(u_multiplier_pp2_41 [2]));
 NAND2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_41_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_41_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_41_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_41_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_41_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_41_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_41_2__17_ ),
    .ZN(u_multiplier_pp2_42 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_41_3__18_  (.A(u_multiplier_STAGE2_pp2_40_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_3__19_  (.A1(u_multiplier_pp1_41 [9]),
    .A2(u_multiplier_pp1_41 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_3__20_  (.A(u_multiplier_pp1_41 [9]),
    .B(u_multiplier_pp1_41 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_41_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_3__21_  (.A1(u_multiplier_pp1_41 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_41_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_3__22_  (.A(u_multiplier_pp1_41 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_41_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_41_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_3__23_  (.A1(u_multiplier_pp1_41 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_41_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_3__24_  (.A(u_multiplier_pp1_41 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_41_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_3__25_  (.A(u_multiplier_STAGE2_pp2_40_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_41_3__16_ ),
    .ZN(u_multiplier_pp2_41 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_41_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_41_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_41_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_41_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_41_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_41_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_41_3__17_ ),
    .ZN(u_multiplier_pp2_42 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_41_4__18_  (.A(u_multiplier_STAGE2_pp2_40_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_4__19_  (.A1(u_multiplier_pp1_41 [13]),
    .A2(u_multiplier_pp1_41 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_4__20_  (.A(u_multiplier_pp1_41 [13]),
    .B(u_multiplier_pp1_41 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_41_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_4__21_  (.A1(u_multiplier_pp1_41 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_41_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_4__22_  (.A(u_multiplier_pp1_41 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_41_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_41_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_4__23_  (.A1(u_multiplier_pp1_41 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_41_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_4__24_  (.A(u_multiplier_pp1_41 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_41_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_41_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_41_4__25_  (.A(u_multiplier_STAGE2_pp2_40_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_41_4__16_ ),
    .ZN(u_multiplier_pp2_41 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_41_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_41_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_41_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_41_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_41_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_41_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_41_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_41_4__17_ ),
    .ZN(u_multiplier_pp2_42 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_42_1__18_  (.A(u_multiplier_STAGE2_pp2_41_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_1__19_  (.A1(u_multiplier_pp1_42 [1]),
    .A2(u_multiplier_pp1_42 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_1__20_  (.A(u_multiplier_pp1_42 [1]),
    .B(u_multiplier_pp1_42 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_42_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_1__21_  (.A1(u_multiplier_pp1_42 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_42_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_1__22_  (.A(u_multiplier_pp1_42 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_42_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_42_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_1__23_  (.A1(u_multiplier_pp1_42 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_42_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_1__24_  (.A(u_multiplier_pp1_42 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_42_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_1__25_  (.A(u_multiplier_STAGE2_pp2_41_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_42_1__16_ ),
    .ZN(u_multiplier_pp2_42 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_42_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_42_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_42_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_42_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_42_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_42_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_42_1__17_ ),
    .ZN(u_multiplier_pp2_43 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_42_2__18_  (.A(u_multiplier_STAGE2_pp2_41_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_2__19_  (.A1(u_multiplier_pp1_42 [5]),
    .A2(u_multiplier_pp1_42 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_2__20_  (.A(u_multiplier_pp1_42 [5]),
    .B(u_multiplier_pp1_42 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_42_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_2__21_  (.A1(u_multiplier_pp1_42 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_42_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_2__22_  (.A(u_multiplier_pp1_42 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_42_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_42_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_2__23_  (.A1(u_multiplier_pp1_42 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_42_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_2__24_  (.A(u_multiplier_pp1_42 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_42_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_2__25_  (.A(u_multiplier_STAGE2_pp2_41_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_42_2__16_ ),
    .ZN(u_multiplier_pp2_42 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_42_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_42_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_42_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_42_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_42_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_42_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_42_2__17_ ),
    .ZN(u_multiplier_pp2_43 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_42_3__18_  (.A(u_multiplier_STAGE2_pp2_41_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_3__19_  (.A1(u_multiplier_pp1_42 [9]),
    .A2(u_multiplier_pp1_42 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_3__20_  (.A(u_multiplier_pp1_42 [9]),
    .B(u_multiplier_pp1_42 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_42_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_3__21_  (.A1(u_multiplier_pp1_42 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_42_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_3__22_  (.A(u_multiplier_pp1_42 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_42_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_42_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_3__23_  (.A1(u_multiplier_pp1_42 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_42_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_3__24_  (.A(u_multiplier_pp1_42 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_42_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_3__25_  (.A(u_multiplier_STAGE2_pp2_41_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_42_3__16_ ),
    .ZN(u_multiplier_pp2_42 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_42_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_42_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_42_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_42_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_42_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_42_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_42_3__17_ ),
    .ZN(u_multiplier_pp2_43 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_42_4__18_  (.A(u_multiplier_STAGE2_pp2_41_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_4__19_  (.A1(u_multiplier_pp1_42 [13]),
    .A2(u_multiplier_pp1_42 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_4__20_  (.A(u_multiplier_pp1_42 [13]),
    .B(u_multiplier_pp1_42 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_42_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_4__21_  (.A1(u_multiplier_pp1_42 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_42_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_4__22_  (.A(u_multiplier_pp1_42 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_42_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_42_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_4__23_  (.A1(u_multiplier_pp1_42 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_42_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_4__24_  (.A(u_multiplier_pp1_42 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_42_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_42_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_42_4__25_  (.A(u_multiplier_STAGE2_pp2_41_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_42_4__16_ ),
    .ZN(u_multiplier_pp2_42 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_42_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_42_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_42_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_42_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_42_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_42_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_42_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_42_4__17_ ),
    .ZN(u_multiplier_pp2_43 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_43_1__18_  (.A(u_multiplier_STAGE2_pp2_42_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_1__19_  (.A1(u_multiplier_pp1_43 [1]),
    .A2(u_multiplier_pp1_43 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_1__20_  (.A(u_multiplier_pp1_43 [1]),
    .B(u_multiplier_pp1_43 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_43_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_1__21_  (.A1(u_multiplier_pp1_43 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_43_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_1__22_  (.A(u_multiplier_pp1_43 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_43_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_43_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_1__23_  (.A1(u_multiplier_pp1_43 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_43_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_1__24_  (.A(u_multiplier_pp1_43 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_43_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_1__25_  (.A(u_multiplier_STAGE2_pp2_42_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_43_1__16_ ),
    .ZN(u_multiplier_pp2_43 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_43_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_43_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_43_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_43_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_43_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_43_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_43_1__17_ ),
    .ZN(u_multiplier_pp2_44 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_43_2__18_  (.A(u_multiplier_STAGE2_pp2_42_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_2__19_  (.A1(u_multiplier_pp1_43 [5]),
    .A2(u_multiplier_pp1_43 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_2__20_  (.A(u_multiplier_pp1_43 [5]),
    .B(u_multiplier_pp1_43 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_43_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_2__21_  (.A1(u_multiplier_pp1_43 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_43_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_2__22_  (.A(u_multiplier_pp1_43 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_43_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_43_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_2__23_  (.A1(u_multiplier_pp1_43 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_43_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_2__24_  (.A(u_multiplier_pp1_43 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_43_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_2__25_  (.A(u_multiplier_STAGE2_pp2_42_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_43_2__16_ ),
    .ZN(u_multiplier_pp2_43 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_43_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_43_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_43_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_43_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_43_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_43_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_43_2__17_ ),
    .ZN(u_multiplier_pp2_44 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_43_3__18_  (.A(u_multiplier_STAGE2_pp2_42_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_3__19_  (.A1(u_multiplier_pp1_43 [9]),
    .A2(u_multiplier_pp1_43 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_3__20_  (.A(u_multiplier_pp1_43 [9]),
    .B(u_multiplier_pp1_43 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_43_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_3__21_  (.A1(u_multiplier_pp1_43 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_43_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_3__22_  (.A(u_multiplier_pp1_43 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_43_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_43_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_3__23_  (.A1(u_multiplier_pp1_43 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_43_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_3__24_  (.A(u_multiplier_pp1_43 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_43_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_3__25_  (.A(u_multiplier_STAGE2_pp2_42_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_43_3__16_ ),
    .ZN(u_multiplier_pp2_43 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_43_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_43_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_43_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_43_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_43_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_43_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_43_3__17_ ),
    .ZN(u_multiplier_pp2_44 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_43_4__18_  (.A(u_multiplier_STAGE2_pp2_42_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_4__19_  (.A1(u_multiplier_pp1_43 [13]),
    .A2(u_multiplier_pp1_43 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_4__20_  (.A(u_multiplier_pp1_43 [13]),
    .B(u_multiplier_pp1_43 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_43_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_4__21_  (.A1(u_multiplier_pp1_43 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_43_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_4__22_  (.A(u_multiplier_pp1_43 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_43_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_43_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_4__23_  (.A1(u_multiplier_pp1_43 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_43_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_4__24_  (.A(u_multiplier_pp1_43 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_43_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_43_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_43_4__25_  (.A(u_multiplier_STAGE2_pp2_42_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_43_4__16_ ),
    .ZN(u_multiplier_pp2_43 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_43_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_43_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_43_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_43_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_43_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_43_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_43_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_43_4__17_ ),
    .ZN(u_multiplier_pp2_44 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_44_1__18_  (.A(u_multiplier_STAGE2_pp2_43_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_1__19_  (.A1(u_multiplier_pp1_44 [1]),
    .A2(u_multiplier_pp1_44 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_1__20_  (.A(u_multiplier_pp1_44 [1]),
    .B(u_multiplier_pp1_44 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_44_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_1__21_  (.A1(u_multiplier_pp1_44 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_44_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_1__22_  (.A(u_multiplier_pp1_44 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_44_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_44_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_1__23_  (.A1(u_multiplier_pp1_44 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_44_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_1__24_  (.A(u_multiplier_pp1_44 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_44_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_1__25_  (.A(u_multiplier_STAGE2_pp2_43_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_44_1__16_ ),
    .ZN(u_multiplier_pp2_44 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_44_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_44_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_44_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_44_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_44_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_44_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_44_1__17_ ),
    .ZN(u_multiplier_pp2_45 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_44_2__18_  (.A(u_multiplier_STAGE2_pp2_43_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_2__19_  (.A1(u_multiplier_pp1_44 [5]),
    .A2(u_multiplier_pp1_44 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_2__20_  (.A(u_multiplier_pp1_44 [5]),
    .B(u_multiplier_pp1_44 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_44_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_2__21_  (.A1(u_multiplier_pp1_44 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_44_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_2__22_  (.A(u_multiplier_pp1_44 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_44_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_44_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_2__23_  (.A1(u_multiplier_pp1_44 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_44_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_2__24_  (.A(u_multiplier_pp1_44 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_44_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_2__25_  (.A(u_multiplier_STAGE2_pp2_43_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_44_2__16_ ),
    .ZN(u_multiplier_pp2_44 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_44_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_44_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_44_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_44_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_44_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_44_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_44_2__17_ ),
    .ZN(u_multiplier_pp2_45 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_44_3__18_  (.A(u_multiplier_STAGE2_pp2_43_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_3__19_  (.A1(u_multiplier_pp1_44 [9]),
    .A2(u_multiplier_pp1_44 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_3__20_  (.A(u_multiplier_pp1_44 [9]),
    .B(u_multiplier_pp1_44 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_44_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_3__21_  (.A1(u_multiplier_pp1_44 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_44_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_3__22_  (.A(u_multiplier_pp1_44 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_44_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_44_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_3__23_  (.A1(u_multiplier_pp1_44 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_44_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_3__24_  (.A(u_multiplier_pp1_44 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_44_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_3__25_  (.A(u_multiplier_STAGE2_pp2_43_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_44_3__16_ ),
    .ZN(u_multiplier_pp2_44 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_44_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_44_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_44_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_44_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_44_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_44_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_44_3__17_ ),
    .ZN(u_multiplier_pp2_45 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_44_4__18_  (.A(u_multiplier_STAGE2_pp2_43_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_4__19_  (.A1(u_multiplier_pp1_44 [13]),
    .A2(u_multiplier_pp1_44 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_4__20_  (.A(u_multiplier_pp1_44 [13]),
    .B(u_multiplier_pp1_44 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_44_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_4__21_  (.A1(u_multiplier_pp1_44 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_44_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_4__22_  (.A(u_multiplier_pp1_44 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_44_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_44_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_4__23_  (.A1(u_multiplier_pp1_44 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_44_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_4__24_  (.A(u_multiplier_pp1_44 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_44_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_44_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_44_4__25_  (.A(u_multiplier_STAGE2_pp2_43_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_44_4__16_ ),
    .ZN(u_multiplier_pp2_44 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_44_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_44_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_44_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_44_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_44_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_44_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_44_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_44_4__17_ ),
    .ZN(u_multiplier_pp2_45 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_45_1__18_  (.A(u_multiplier_STAGE2_pp2_44_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_1__19_  (.A1(u_multiplier_pp1_45 [1]),
    .A2(u_multiplier_pp1_45 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_1__20_  (.A(u_multiplier_pp1_45 [1]),
    .B(u_multiplier_pp1_45 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_45_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_1__21_  (.A1(u_multiplier_pp1_45 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_45_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_1__22_  (.A(u_multiplier_pp1_45 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_45_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_45_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_1__23_  (.A1(u_multiplier_pp1_45 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_45_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_1__24_  (.A(u_multiplier_pp1_45 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_45_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_1__25_  (.A(u_multiplier_STAGE2_pp2_44_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_45_1__16_ ),
    .ZN(u_multiplier_pp2_45 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_45_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_45_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_45_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_45_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_45_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_45_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_45_1__17_ ),
    .ZN(u_multiplier_pp2_46 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_45_2__18_  (.A(u_multiplier_STAGE2_pp2_44_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_2__19_  (.A1(u_multiplier_pp1_45 [5]),
    .A2(u_multiplier_pp1_45 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_2__20_  (.A(u_multiplier_pp1_45 [5]),
    .B(u_multiplier_pp1_45 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_45_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_2__21_  (.A1(u_multiplier_pp1_45 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_45_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_2__22_  (.A(u_multiplier_pp1_45 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_45_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_45_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_2__23_  (.A1(u_multiplier_pp1_45 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_45_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_2__24_  (.A(u_multiplier_pp1_45 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_45_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_2__25_  (.A(u_multiplier_STAGE2_pp2_44_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_45_2__16_ ),
    .ZN(u_multiplier_pp2_45 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_45_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_45_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_45_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_45_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_45_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_45_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_45_2__17_ ),
    .ZN(u_multiplier_pp2_46 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_45_3__18_  (.A(u_multiplier_STAGE2_pp2_44_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_3__19_  (.A1(u_multiplier_pp1_45 [9]),
    .A2(u_multiplier_pp1_45 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_3__20_  (.A(u_multiplier_pp1_45 [9]),
    .B(u_multiplier_pp1_45 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_45_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_3__21_  (.A1(u_multiplier_pp1_45 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_45_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_3__22_  (.A(u_multiplier_pp1_45 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_45_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_45_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_3__23_  (.A1(u_multiplier_pp1_45 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_45_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_3__24_  (.A(u_multiplier_pp1_45 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_45_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_3__25_  (.A(u_multiplier_STAGE2_pp2_44_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_45_3__16_ ),
    .ZN(u_multiplier_pp2_45 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_45_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_45_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_45_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_45_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_45_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_45_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_45_3__17_ ),
    .ZN(u_multiplier_pp2_46 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_45_4__18_  (.A(u_multiplier_STAGE2_pp2_44_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_4__19_  (.A1(u_multiplier_pp1_45 [13]),
    .A2(u_multiplier_pp1_45 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_4__20_  (.A(u_multiplier_pp1_45 [13]),
    .B(u_multiplier_pp1_45 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_45_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_4__21_  (.A1(u_multiplier_pp1_45 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_45_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_4__22_  (.A(u_multiplier_pp1_45 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_45_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_45_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_4__23_  (.A1(u_multiplier_pp1_45 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_45_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_4__24_  (.A(u_multiplier_pp1_45 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_45_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_45_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_45_4__25_  (.A(u_multiplier_STAGE2_pp2_44_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_45_4__16_ ),
    .ZN(u_multiplier_pp2_45 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_45_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_45_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_45_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_45_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_45_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_45_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_45_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_45_4__17_ ),
    .ZN(u_multiplier_pp2_46 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_46_1__18_  (.A(u_multiplier_STAGE2_pp2_45_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_1__19_  (.A1(u_multiplier_pp1_46 [1]),
    .A2(u_multiplier_pp1_46 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_1__20_  (.A(u_multiplier_pp1_46 [1]),
    .B(u_multiplier_pp1_46 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_46_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_1__21_  (.A1(u_multiplier_pp1_46 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_46_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_1__22_  (.A(u_multiplier_pp1_46 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_46_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_46_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_1__23_  (.A1(u_multiplier_pp1_46 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_46_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_1__24_  (.A(u_multiplier_pp1_46 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_46_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_1__25_  (.A(u_multiplier_STAGE2_pp2_45_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_46_1__16_ ),
    .ZN(u_multiplier_pp2_46 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_46_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_46_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_46_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_46_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_46_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_46_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_46_1__17_ ),
    .ZN(u_multiplier_pp2_47 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_46_2__18_  (.A(u_multiplier_STAGE2_pp2_45_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_2__19_  (.A1(u_multiplier_pp1_46 [5]),
    .A2(u_multiplier_pp1_46 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_2__20_  (.A(u_multiplier_pp1_46 [5]),
    .B(u_multiplier_pp1_46 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_46_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_2__21_  (.A1(u_multiplier_pp1_46 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_46_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_2__22_  (.A(u_multiplier_pp1_46 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_46_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_46_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_2__23_  (.A1(u_multiplier_pp1_46 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_46_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_2__24_  (.A(u_multiplier_pp1_46 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_46_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_2__25_  (.A(u_multiplier_STAGE2_pp2_45_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_46_2__16_ ),
    .ZN(u_multiplier_pp2_46 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_46_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_46_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_46_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_46_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_46_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_46_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_46_2__17_ ),
    .ZN(u_multiplier_pp2_47 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_46_3__18_  (.A(u_multiplier_STAGE2_pp2_45_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_3__19_  (.A1(u_multiplier_pp1_46 [9]),
    .A2(u_multiplier_pp1_46 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_3__20_  (.A(u_multiplier_pp1_46 [9]),
    .B(u_multiplier_pp1_46 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_46_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_3__21_  (.A1(u_multiplier_pp1_46 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_46_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_3__22_  (.A(u_multiplier_pp1_46 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_46_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_46_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_3__23_  (.A1(u_multiplier_pp1_46 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_46_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_3__24_  (.A(u_multiplier_pp1_46 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_46_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_3__25_  (.A(u_multiplier_STAGE2_pp2_45_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_46_3__16_ ),
    .ZN(u_multiplier_pp2_46 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_46_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_46_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_46_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_46_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_46_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_46_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_46_3__17_ ),
    .ZN(u_multiplier_pp2_47 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_46_4__18_  (.A(u_multiplier_STAGE2_pp2_45_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_4__19_  (.A1(u_multiplier_pp1_46 [13]),
    .A2(u_multiplier_pp1_46 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_4__20_  (.A(u_multiplier_pp1_46 [13]),
    .B(u_multiplier_pp1_46 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_46_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_4__21_  (.A1(u_multiplier_pp1_46 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_46_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_4__22_  (.A(u_multiplier_pp1_46 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_46_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_46_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_4__23_  (.A1(u_multiplier_pp1_46 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_46_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_4__24_  (.A(u_multiplier_pp1_46 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_46_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_46_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_46_4__25_  (.A(u_multiplier_STAGE2_pp2_45_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_46_4__16_ ),
    .ZN(u_multiplier_pp2_46 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_46_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_46_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_46_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_46_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_46_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_46_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_46_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_46_4__17_ ),
    .ZN(u_multiplier_pp2_47 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_47_1__18_  (.A(u_multiplier_STAGE2_pp2_46_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_1__19_  (.A1(u_multiplier_pp1_47 [1]),
    .A2(u_multiplier_pp1_47 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_1__20_  (.A(u_multiplier_pp1_47 [1]),
    .B(u_multiplier_pp1_47 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_47_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_1__21_  (.A1(u_multiplier_pp1_47 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_47_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_1__22_  (.A(u_multiplier_pp1_47 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_47_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_47_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_1__23_  (.A1(u_multiplier_pp1_47 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_47_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_1__24_  (.A(u_multiplier_pp1_47 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_47_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_1__25_  (.A(u_multiplier_STAGE2_pp2_46_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_47_1__16_ ),
    .ZN(u_multiplier_pp2_47 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_47_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_47_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_47_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_47_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_47_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_47_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_47_1__17_ ),
    .ZN(u_multiplier_pp2_48 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_47_2__18_  (.A(u_multiplier_STAGE2_pp2_46_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_2__19_  (.A1(u_multiplier_pp1_47 [5]),
    .A2(u_multiplier_pp1_47 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_2__20_  (.A(u_multiplier_pp1_47 [5]),
    .B(u_multiplier_pp1_47 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_47_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_2__21_  (.A1(u_multiplier_pp1_47 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_47_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_2__22_  (.A(u_multiplier_pp1_47 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_47_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_47_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_2__23_  (.A1(u_multiplier_pp1_47 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_47_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_2__24_  (.A(u_multiplier_pp1_47 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_47_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_2__25_  (.A(u_multiplier_STAGE2_pp2_46_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_47_2__16_ ),
    .ZN(u_multiplier_pp2_47 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_47_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_47_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_47_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_47_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_47_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_47_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_47_2__17_ ),
    .ZN(u_multiplier_pp2_48 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_47_3__18_  (.A(u_multiplier_STAGE2_pp2_46_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_3__19_  (.A1(u_multiplier_pp1_47 [9]),
    .A2(u_multiplier_pp1_47 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_3__20_  (.A(u_multiplier_pp1_47 [9]),
    .B(u_multiplier_pp1_47 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_47_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_3__21_  (.A1(u_multiplier_pp1_47 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_47_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_3__22_  (.A(u_multiplier_pp1_47 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_47_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_47_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_3__23_  (.A1(u_multiplier_pp1_47 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_47_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_3__24_  (.A(u_multiplier_pp1_47 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_47_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_3__25_  (.A(u_multiplier_STAGE2_pp2_46_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_47_3__16_ ),
    .ZN(u_multiplier_pp2_47 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_47_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_47_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_47_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_47_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_47_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_47_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_47_3__17_ ),
    .ZN(u_multiplier_pp2_48 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_47_4__18_  (.A(u_multiplier_STAGE2_pp2_46_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_4__19_  (.A1(u_multiplier_pp1_47 [13]),
    .A2(u_multiplier_pp1_47 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_4__20_  (.A(u_multiplier_pp1_47 [13]),
    .B(u_multiplier_pp1_47 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_47_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_4__21_  (.A1(u_multiplier_pp1_47 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_47_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_4__22_  (.A(u_multiplier_pp1_47 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_47_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_47_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_4__23_  (.A1(u_multiplier_pp1_47 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_47_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_4__24_  (.A(u_multiplier_pp1_47 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_47_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_47_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_47_4__25_  (.A(u_multiplier_STAGE2_pp2_46_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_47_4__16_ ),
    .ZN(u_multiplier_pp2_47 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_47_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_47_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_47_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_47_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_47_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_47_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_47_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_47_4__17_ ),
    .ZN(u_multiplier_pp2_48 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_48_1__18_  (.A(u_multiplier_STAGE2_pp2_47_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_1__19_  (.A1(u_multiplier_pp1_48 [1]),
    .A2(u_multiplier_pp1_48 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_1__20_  (.A(u_multiplier_pp1_48 [1]),
    .B(u_multiplier_pp1_48 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_48_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_1__21_  (.A1(u_multiplier_pp1_48 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_48_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_1__22_  (.A(u_multiplier_pp1_48 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_48_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_48_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_1__23_  (.A1(u_multiplier_pp1_48 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_48_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_1__24_  (.A(u_multiplier_pp1_48 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_48_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_1__25_  (.A(u_multiplier_STAGE2_pp2_47_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_48_1__16_ ),
    .ZN(u_multiplier_pp2_48 [3]));
 NAND2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_48_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_48_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_48_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_48_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_48_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_48_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_48_1__17_ ),
    .ZN(u_multiplier_pp2_49 [7]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_48_2__18_  (.A(u_multiplier_STAGE2_pp2_47_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_2__19_  (.A1(u_multiplier_pp1_48 [5]),
    .A2(u_multiplier_pp1_48 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_2__20_  (.A(u_multiplier_pp1_48 [5]),
    .B(u_multiplier_pp1_48 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_48_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_2__21_  (.A1(u_multiplier_pp1_48 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_48_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_2__22_  (.A(u_multiplier_pp1_48 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_48_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_48_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_2__23_  (.A1(u_multiplier_pp1_48 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_48_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_2__24_  (.A(u_multiplier_pp1_48 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_48_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_2__25_  (.A(u_multiplier_STAGE2_pp2_47_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_48_2__16_ ),
    .ZN(u_multiplier_pp2_48 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_48_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_48_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_48_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_48_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_48_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_48_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_48_2__17_ ),
    .ZN(u_multiplier_pp2_49 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_48_3__18_  (.A(u_multiplier_STAGE2_pp2_47_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_3__19_  (.A1(u_multiplier_pp1_48 [9]),
    .A2(u_multiplier_pp1_48 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_3__20_  (.A(u_multiplier_pp1_48 [9]),
    .B(u_multiplier_pp1_48 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_48_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_3__21_  (.A1(u_multiplier_pp1_48 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_48_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_3__22_  (.A(u_multiplier_pp1_48 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_48_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_48_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_3__23_  (.A1(u_multiplier_pp1_48 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_48_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_3__24_  (.A(u_multiplier_pp1_48 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_48_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_3__25_  (.A(u_multiplier_STAGE2_pp2_47_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_48_3__16_ ),
    .ZN(u_multiplier_pp2_48 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_48_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_48_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_48_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_48_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_48_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_48_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_48_3__17_ ),
    .ZN(u_multiplier_pp2_49 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_48_4__18_  (.A(u_multiplier_STAGE2_pp2_47_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_4__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_4__19_  (.A1(u_multiplier_pp1_48 [13]),
    .A2(u_multiplier_pp1_48 [12]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_4__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_4__20_  (.A(u_multiplier_pp1_48 [13]),
    .B(u_multiplier_pp1_48 [12]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_48_4__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_4__21_  (.A1(u_multiplier_pp1_48 [14]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_48_4__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_4__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_4__22_  (.A(u_multiplier_pp1_48 [14]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_48_4__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_48_4__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_4__23_  (.A1(u_multiplier_pp1_48 [15]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_48_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_4__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_4__24_  (.A(u_multiplier_pp1_48 [15]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_48_4__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_48_4__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_48_4__25_  (.A(u_multiplier_STAGE2_pp2_47_e42_4_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_48_4__16_ ),
    .ZN(u_multiplier_pp2_48 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_48_4__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_48_4__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_48_4__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_48_e42_4_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_48_4__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_48_4__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_48_4__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_48_4__17_ ),
    .ZN(u_multiplier_pp2_49 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_49_1__18_  (.A(u_multiplier_STAGE2_pp2_48_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_49_1__19_  (.A1(u_multiplier_pp1_49 [1]),
    .A2(u_multiplier_pp1_49 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_49_1__20_  (.A(u_multiplier_pp1_49 [1]),
    .B(u_multiplier_pp1_49 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_49_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_49_1__21_  (.A1(u_multiplier_pp1_49 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_49_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_49_1__22_  (.A(u_multiplier_pp1_49 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_49_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_49_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_49_1__23_  (.A1(u_multiplier_pp1_49 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_49_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_49_1__24_  (.A(u_multiplier_pp1_49 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_49_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_49_1__25_  (.A(u_multiplier_STAGE2_pp2_48_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_49_1__16_ ),
    .ZN(u_multiplier_pp2_49 [3]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_49_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_49_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_49_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_49_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_49_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_49_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_49_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_49_1__17_ ),
    .ZN(u_multiplier_pp2_50 [6]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_49_2__18_  (.A(u_multiplier_STAGE2_pp2_48_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_49_2__19_  (.A1(u_multiplier_pp1_49 [5]),
    .A2(u_multiplier_pp1_49 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_49_2__20_  (.A(u_multiplier_pp1_49 [5]),
    .B(u_multiplier_pp1_49 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_49_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_49_2__21_  (.A1(u_multiplier_pp1_49 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_49_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_49_2__22_  (.A(u_multiplier_pp1_49 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_49_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_49_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_49_2__23_  (.A1(u_multiplier_pp1_49 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_49_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_49_2__24_  (.A(u_multiplier_pp1_49 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_49_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_49_2__25_  (.A(u_multiplier_STAGE2_pp2_48_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_49_2__16_ ),
    .ZN(u_multiplier_pp2_49 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_49_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_49_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_49_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_49_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_49_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_49_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_49_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_49_2__17_ ),
    .ZN(u_multiplier_pp2_50 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_49_3__18_  (.A(u_multiplier_STAGE2_pp2_48_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_49_3__19_  (.A1(u_multiplier_pp1_49 [9]),
    .A2(u_multiplier_pp1_49 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_49_3__20_  (.A(u_multiplier_pp1_49 [9]),
    .B(u_multiplier_pp1_49 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_49_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_49_3__21_  (.A1(u_multiplier_pp1_49 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_49_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_49_3__22_  (.A(u_multiplier_pp1_49 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_49_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_49_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_49_3__23_  (.A1(u_multiplier_pp1_49 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_49_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_49_3__24_  (.A(u_multiplier_pp1_49 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_49_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_49_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_49_3__25_  (.A(u_multiplier_STAGE2_pp2_48_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_49_3__16_ ),
    .ZN(u_multiplier_pp2_49 [1]));
 NAND2_X2 u_multiplier_STAGE2_E_4_2_pp2_49_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_49_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_49_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_49_e42_3_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_49_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_49_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_49_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_49_3__17_ ),
    .ZN(u_multiplier_pp2_50 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_50_1__18_  (.A(u_multiplier_STAGE2_pp2_49_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_50_1__19_  (.A1(u_multiplier_pp1_50 [1]),
    .A2(u_multiplier_pp1_50 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_50_1__20_  (.A(u_multiplier_pp1_50 [1]),
    .B(u_multiplier_pp1_50 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_50_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_50_1__21_  (.A1(u_multiplier_pp1_50 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_50_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_50_1__22_  (.A(u_multiplier_pp1_50 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_50_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_50_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_50_1__23_  (.A1(u_multiplier_pp1_50 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_50_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_50_1__24_  (.A(u_multiplier_pp1_50 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_50_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_50_1__25_  (.A(u_multiplier_STAGE2_pp2_49_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_50_1__16_ ),
    .ZN(u_multiplier_pp2_50 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_50_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_50_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_50_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_50_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_50_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_50_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_50_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_50_1__17_ ),
    .ZN(u_multiplier_pp2_51 [5]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_50_2__18_  (.A(u_multiplier_STAGE2_pp2_49_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_50_2__19_  (.A1(u_multiplier_pp1_50 [5]),
    .A2(u_multiplier_pp1_50 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_50_2__20_  (.A(u_multiplier_pp1_50 [5]),
    .B(u_multiplier_pp1_50 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_50_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_50_2__21_  (.A1(u_multiplier_pp1_50 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_50_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_50_2__22_  (.A(u_multiplier_pp1_50 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_50_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_50_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_50_2__23_  (.A1(u_multiplier_pp1_50 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_50_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_50_2__24_  (.A(u_multiplier_pp1_50 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_50_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_50_2__25_  (.A(u_multiplier_STAGE2_pp2_49_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_50_2__16_ ),
    .ZN(u_multiplier_pp2_50 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_50_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_50_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_50_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_50_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_50_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_50_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_50_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_50_2__17_ ),
    .ZN(u_multiplier_pp2_51 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_50_3__18_  (.A(u_multiplier_STAGE2_pp2_49_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_50_3__19_  (.A1(u_multiplier_pp1_50 [9]),
    .A2(u_multiplier_pp1_50 [8]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_3__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_50_3__20_  (.A(u_multiplier_pp1_50 [9]),
    .B(u_multiplier_pp1_50 [8]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_50_3__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_50_3__21_  (.A1(u_multiplier_pp1_50 [10]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_50_3__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_3__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_50_3__22_  (.A(u_multiplier_pp1_50 [10]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_50_3__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_50_3__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_50_3__23_  (.A1(u_multiplier_pp1_50 [11]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_50_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_3__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_50_3__24_  (.A(u_multiplier_pp1_50 [11]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_50_3__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_50_3__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_50_3__25_  (.A(u_multiplier_STAGE2_pp2_49_e42_3_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_50_3__16_ ),
    .ZN(u_multiplier_pp2_50 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_50_3__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_50_3__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_50_3__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_50_e42_3_cout ));
 OAI21_X1 u_multiplier_STAGE2_E_4_2_pp2_50_3__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_50_3__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_50_3__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_50_3__17_ ),
    .ZN(u_multiplier_pp2_51 [3]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_51_1__18_  (.A(u_multiplier_STAGE2_pp2_50_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_51_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_51_1__19_  (.A1(u_multiplier_pp1_51 [1]),
    .A2(u_multiplier_pp1_51 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_51_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_51_1__20_  (.A(u_multiplier_pp1_51 [1]),
    .B(u_multiplier_pp1_51 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_51_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_51_1__21_  (.A1(u_multiplier_pp1_51 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_51_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_51_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_51_1__22_  (.A(u_multiplier_pp1_51 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_51_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_51_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_51_1__23_  (.A1(u_multiplier_pp1_51 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_51_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_51_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_51_1__24_  (.A(u_multiplier_pp1_51 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_51_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_51_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_51_1__25_  (.A(u_multiplier_STAGE2_pp2_50_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_51_1__16_ ),
    .ZN(u_multiplier_pp2_51 [2]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_51_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_51_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_51_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_51_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_51_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_51_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_51_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_51_1__17_ ),
    .ZN(u_multiplier_pp2_52 [4]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_51_2__18_  (.A(u_multiplier_STAGE2_pp2_50_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_51_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_51_2__19_  (.A1(u_multiplier_pp1_51 [5]),
    .A2(u_multiplier_pp1_51 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_51_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_51_2__20_  (.A(u_multiplier_pp1_51 [5]),
    .B(u_multiplier_pp1_51 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_51_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_51_2__21_  (.A1(u_multiplier_pp1_51 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_51_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_51_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_51_2__22_  (.A(u_multiplier_pp1_51 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_51_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_51_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_51_2__23_  (.A1(u_multiplier_pp1_51 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_51_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_51_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_51_2__24_  (.A(u_multiplier_pp1_51 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_51_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_51_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_51_2__25_  (.A(u_multiplier_STAGE2_pp2_50_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_51_2__16_ ),
    .ZN(u_multiplier_pp2_51 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_51_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_51_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_51_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_51_e42_2_cout ));
 OAI21_X1 u_multiplier_STAGE2_E_4_2_pp2_51_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_51_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_51_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_51_2__17_ ),
    .ZN(u_multiplier_pp2_52 [3]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_52_1__18_  (.A(u_multiplier_STAGE2_pp2_51_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_52_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_52_1__19_  (.A1(u_multiplier_pp1_52 [1]),
    .A2(u_multiplier_pp1_52 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_52_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_52_1__20_  (.A(u_multiplier_pp1_52 [1]),
    .B(u_multiplier_pp1_52 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_52_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_52_1__21_  (.A1(u_multiplier_pp1_52 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_52_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_52_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_52_1__22_  (.A(u_multiplier_pp1_52 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_52_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_52_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_52_1__23_  (.A1(u_multiplier_pp1_52 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_52_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_52_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_52_1__24_  (.A(u_multiplier_pp1_52 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_52_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_52_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_52_1__25_  (.A(u_multiplier_STAGE2_pp2_51_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_52_1__16_ ),
    .ZN(u_multiplier_pp2_52 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_52_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_52_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_52_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_52_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE2_E_4_2_pp2_52_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_52_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_52_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_52_1__17_ ),
    .ZN(u_multiplier_pp2_53 [3]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_52_2__18_  (.A(u_multiplier_STAGE2_pp2_51_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_52_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_52_2__19_  (.A1(u_multiplier_pp1_52 [5]),
    .A2(u_multiplier_pp1_52 [4]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_52_2__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_52_2__20_  (.A(u_multiplier_pp1_52 [5]),
    .B(u_multiplier_pp1_52 [4]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_52_2__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_52_2__21_  (.A1(u_multiplier_pp1_52 [6]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_52_2__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_52_2__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_52_2__22_  (.A(u_multiplier_pp1_52 [6]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_52_2__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_52_2__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_52_2__23_  (.A1(u_multiplier_pp1_52 [7]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_52_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_52_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_52_2__24_  (.A(u_multiplier_pp1_52 [7]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_52_2__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_52_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_52_2__25_  (.A(u_multiplier_STAGE2_pp2_51_e42_2_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_52_2__16_ ),
    .ZN(u_multiplier_pp2_52 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_52_2__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_52_2__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_52_2__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_52_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_52_2__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_52_2__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_52_2__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_52_2__17_ ),
    .ZN(u_multiplier_pp2_53 [2]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_53_1__18_  (.A(u_multiplier_STAGE2_pp2_52_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_53_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_53_1__19_  (.A1(u_multiplier_pp1_53 [1]),
    .A2(u_multiplier_pp1_53 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_53_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_53_1__20_  (.A(u_multiplier_pp1_53 [1]),
    .B(u_multiplier_pp1_53 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_53_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_53_1__21_  (.A1(u_multiplier_pp1_53 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_53_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_53_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_53_1__22_  (.A(u_multiplier_pp1_53 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_53_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_53_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_53_1__23_  (.A1(u_multiplier_pp1_53 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_53_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_53_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_53_1__24_  (.A(u_multiplier_pp1_53 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_53_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_53_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_53_1__25_  (.A(u_multiplier_STAGE2_pp2_52_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_53_1__16_ ),
    .ZN(u_multiplier_pp2_53 [1]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_53_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_53_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_53_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_53_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_53_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_53_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_53_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_53_1__17_ ),
    .ZN(u_multiplier_pp2_54 [2]));
 INV_X1 u_multiplier_STAGE2_E_4_2_pp2_54_1__18_  (.A(u_multiplier_STAGE2_pp2_53_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_54_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_54_1__19_  (.A1(u_multiplier_pp1_54 [1]),
    .A2(u_multiplier_pp1_54 [0]),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_54_1__11_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_54_1__20_  (.A(u_multiplier_pp1_54 [1]),
    .B(u_multiplier_pp1_54 [0]),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_54_1__12_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_54_1__21_  (.A1(u_multiplier_pp1_54 [2]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_54_1__12_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_54_1__13_ ));
 XOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_54_1__22_  (.A(u_multiplier_pp1_54 [2]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_54_1__12_ ),
    .Z(u_multiplier_STAGE2_E_4_2_pp2_54_1__14_ ));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_54_1__23_  (.A1(u_multiplier_pp1_54 [3]),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_54_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_54_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_54_1__24_  (.A(u_multiplier_pp1_54 [3]),
    .B(u_multiplier_STAGE2_E_4_2_pp2_54_1__14_ ),
    .ZN(u_multiplier_STAGE2_E_4_2_pp2_54_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE2_E_4_2_pp2_54_1__25_  (.A(u_multiplier_STAGE2_pp2_53_e42_1_cout ),
    .B(u_multiplier_STAGE2_E_4_2_pp2_54_1__16_ ),
    .ZN(u_multiplier_pp2_54 [0]));
 NAND2_X1 u_multiplier_STAGE2_E_4_2_pp2_54_1__26_  (.A1(u_multiplier_STAGE2_E_4_2_pp2_54_1__11_ ),
    .A2(u_multiplier_STAGE2_E_4_2_pp2_54_1__13_ ),
    .ZN(u_multiplier_STAGE2_pp2_54_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE2_E_4_2_pp2_54_1__27_  (.A(u_multiplier_STAGE2_E_4_2_pp2_54_1__15_ ),
    .B1(u_multiplier_STAGE2_E_4_2_pp2_54_1__16_ ),
    .B2(u_multiplier_STAGE2_E_4_2_pp2_54_1__17_ ),
    .ZN(u_multiplier_pp2_55 [1]));
 INV_X1 u_multiplier_STAGE2_Full_adder_pp2_49_1__12_  (.A(u_multiplier_STAGE2_pp2_48_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_49_1__08_ ));
 NAND3_X1 u_multiplier_STAGE2_Full_adder_pp2_49_1__13_  (.A1(u_multiplier_pp1_49 [13]),
    .A2(u_multiplier_pp1_49 [12]),
    .A3(u_multiplier_STAGE2_pp2_48_e42_4_cout ),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_49_1__09_ ));
 NOR2_X2 u_multiplier_STAGE2_Full_adder_pp2_49_1__14_  (.A1(u_multiplier_pp1_49 [13]),
    .A2(u_multiplier_pp1_49 [12]),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_49_1__10_ ));
 AOI21_X1 u_multiplier_STAGE2_Full_adder_pp2_49_1__15_  (.A(u_multiplier_STAGE2_pp2_48_e42_4_cout ),
    .B1(u_multiplier_pp1_49 [12]),
    .B2(u_multiplier_pp1_49 [13]),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_49_1__11_ ));
 NOR2_X2 u_multiplier_STAGE2_Full_adder_pp2_49_1__16_  (.A1(u_multiplier_STAGE2_Full_adder_pp2_49_1__10_ ),
    .A2(u_multiplier_STAGE2_Full_adder_pp2_49_1__11_ ),
    .ZN(u_multiplier_pp2_50 [3]));
 AOI22_X2 u_multiplier_STAGE2_Full_adder_pp2_49_1__17_  (.A1(u_multiplier_STAGE2_Full_adder_pp2_49_1__08_ ),
    .A2(u_multiplier_STAGE2_Full_adder_pp2_49_1__10_ ),
    .B1(u_multiplier_pp2_50 [3]),
    .B2(u_multiplier_STAGE2_Full_adder_pp2_49_1__09_ ),
    .ZN(u_multiplier_pp2_49 [0]));
 INV_X1 u_multiplier_STAGE2_Full_adder_pp2_51_1__12_  (.A(u_multiplier_STAGE2_pp2_50_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_51_1__08_ ));
 NAND3_X1 u_multiplier_STAGE2_Full_adder_pp2_51_1__13_  (.A1(u_multiplier_pp1_51 [9]),
    .A2(u_multiplier_pp1_51 [8]),
    .A3(u_multiplier_STAGE2_pp2_50_e42_3_cout ),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_51_1__09_ ));
 NOR2_X2 u_multiplier_STAGE2_Full_adder_pp2_51_1__14_  (.A1(u_multiplier_pp1_51 [9]),
    .A2(u_multiplier_pp1_51 [8]),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_51_1__10_ ));
 AOI21_X1 u_multiplier_STAGE2_Full_adder_pp2_51_1__15_  (.A(u_multiplier_STAGE2_pp2_50_e42_3_cout ),
    .B1(u_multiplier_pp1_51 [8]),
    .B2(u_multiplier_pp1_51 [9]),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_51_1__11_ ));
 NOR2_X2 u_multiplier_STAGE2_Full_adder_pp2_51_1__16_  (.A1(u_multiplier_STAGE2_Full_adder_pp2_51_1__10_ ),
    .A2(u_multiplier_STAGE2_Full_adder_pp2_51_1__11_ ),
    .ZN(u_multiplier_pp2_52 [2]));
 AOI22_X2 u_multiplier_STAGE2_Full_adder_pp2_51_1__17_  (.A1(u_multiplier_STAGE2_Full_adder_pp2_51_1__08_ ),
    .A2(u_multiplier_STAGE2_Full_adder_pp2_51_1__10_ ),
    .B1(u_multiplier_pp2_52 [2]),
    .B2(u_multiplier_STAGE2_Full_adder_pp2_51_1__09_ ),
    .ZN(u_multiplier_pp2_51 [0]));
 INV_X1 u_multiplier_STAGE2_Full_adder_pp2_53_1__12_  (.A(u_multiplier_STAGE2_pp2_52_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_53_1__08_ ));
 NAND3_X1 u_multiplier_STAGE2_Full_adder_pp2_53_1__13_  (.A1(u_multiplier_pp1_53 [5]),
    .A2(u_multiplier_pp1_53 [4]),
    .A3(u_multiplier_STAGE2_pp2_52_e42_2_cout ),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_53_1__09_ ));
 NOR2_X2 u_multiplier_STAGE2_Full_adder_pp2_53_1__14_  (.A1(u_multiplier_pp1_53 [5]),
    .A2(u_multiplier_pp1_53 [4]),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_53_1__10_ ));
 AOI21_X1 u_multiplier_STAGE2_Full_adder_pp2_53_1__15_  (.A(u_multiplier_STAGE2_pp2_52_e42_2_cout ),
    .B1(u_multiplier_pp1_53 [4]),
    .B2(u_multiplier_pp1_53 [5]),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_53_1__11_ ));
 NOR2_X2 u_multiplier_STAGE2_Full_adder_pp2_53_1__16_  (.A1(u_multiplier_STAGE2_Full_adder_pp2_53_1__10_ ),
    .A2(u_multiplier_STAGE2_Full_adder_pp2_53_1__11_ ),
    .ZN(u_multiplier_pp2_54 [1]));
 AOI22_X2 u_multiplier_STAGE2_Full_adder_pp2_53_1__17_  (.A1(u_multiplier_STAGE2_Full_adder_pp2_53_1__08_ ),
    .A2(u_multiplier_STAGE2_Full_adder_pp2_53_1__10_ ),
    .B1(u_multiplier_pp2_54 [1]),
    .B2(u_multiplier_STAGE2_Full_adder_pp2_53_1__09_ ),
    .ZN(u_multiplier_pp2_53 [0]));
 INV_X1 u_multiplier_STAGE2_Full_adder_pp2_55_1__12_  (.A(u_multiplier_STAGE2_pp2_54_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_55_1__08_ ));
 NAND3_X2 u_multiplier_STAGE2_Full_adder_pp2_55_1__13_  (.A1(u_multiplier_pp1_55 [1]),
    .A2(u_multiplier_pp1_55 [0]),
    .A3(u_multiplier_STAGE2_pp2_54_e42_1_cout ),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_55_1__09_ ));
 NOR2_X2 u_multiplier_STAGE2_Full_adder_pp2_55_1__14_  (.A1(u_multiplier_pp1_55 [1]),
    .A2(u_multiplier_pp1_55 [0]),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_55_1__10_ ));
 AOI21_X1 u_multiplier_STAGE2_Full_adder_pp2_55_1__15_  (.A(u_multiplier_STAGE2_pp2_54_e42_1_cout ),
    .B1(u_multiplier_pp1_55 [0]),
    .B2(u_multiplier_pp1_55 [1]),
    .ZN(u_multiplier_STAGE2_Full_adder_pp2_55_1__11_ ));
 NOR2_X2 u_multiplier_STAGE2_Full_adder_pp2_55_1__16_  (.A1(u_multiplier_STAGE2_Full_adder_pp2_55_1__10_ ),
    .A2(u_multiplier_STAGE2_Full_adder_pp2_55_1__11_ ),
    .ZN(u_multiplier_pp2_56 [0]));
 AOI22_X4 u_multiplier_STAGE2_Full_adder_pp2_55_1__17_  (.A1(u_multiplier_STAGE2_Full_adder_pp2_55_1__08_ ),
    .A2(u_multiplier_STAGE2_Full_adder_pp2_55_1__10_ ),
    .B1(u_multiplier_pp2_56 [0]),
    .B2(u_multiplier_STAGE2_Full_adder_pp2_55_1__09_ ),
    .ZN(u_multiplier_pp2_55 [0]));
 AND2_X1 u_multiplier_STAGE2_Half_adder_pp2_10__4_  (.A1(u_multiplier_pp1_10 [6]),
    .A2(u_multiplier_pp1_10 [5]),
    .ZN(u_multiplier_pp2_11 [2]));
 XOR2_X2 u_multiplier_STAGE2_Half_adder_pp2_10__5_  (.A(u_multiplier_pp1_10 [6]),
    .B(u_multiplier_pp1_10 [5]),
    .Z(u_multiplier_pp2_10 [1]));
 AND2_X1 u_multiplier_STAGE2_Half_adder_pp2_12__4_  (.A1(u_multiplier_pp1_12 [4]),
    .A2(u_multiplier_pp1_12 [3]),
    .ZN(u_multiplier_pp2_13 [3]));
 XOR2_X2 u_multiplier_STAGE2_Half_adder_pp2_12__5_  (.A(u_multiplier_pp1_12 [4]),
    .B(u_multiplier_pp1_12 [3]),
    .Z(u_multiplier_pp2_12 [2]));
 AND2_X1 u_multiplier_STAGE2_Half_adder_pp2_14__4_  (.A1(u_multiplier_pp1_14 [2]),
    .A2(u_multiplier_pp1_14 [1]),
    .ZN(u_multiplier_pp2_15 [4]));
 XOR2_X2 u_multiplier_STAGE2_Half_adder_pp2_14__5_  (.A(u_multiplier_pp1_14 [2]),
    .B(u_multiplier_pp1_14 [1]),
    .Z(u_multiplier_pp2_14 [3]));
 AND2_X1 u_multiplier_STAGE2_Half_adder_pp2_8__4_  (.A1(u_multiplier_pp1_8 [8]),
    .A2(u_multiplier_pp1_8 [7]),
    .ZN(u_multiplier_pp2_9 [1]));
 XOR2_X2 u_multiplier_STAGE2_Half_adder_pp2_8__5_  (.A(u_multiplier_pp1_8 [8]),
    .B(u_multiplier_pp1_8 [7]),
    .Z(u_multiplier_pp2_8 [0]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_10_0__21_  (.A1(u_multiplier_pp1_10 [8]),
    .A2(u_multiplier_pp1_10 [7]),
    .A3(u_multiplier_pp1_10 [9]),
    .ZN(u_multiplier_STAGE2_acci_pp2_10_0__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_10_0__22_  (.A(u_multiplier_pp1_10 [8]),
    .B(u_multiplier_pp1_10 [7]),
    .Z(u_multiplier_STAGE2_acci_pp2_10_0__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_10_0__23_  (.A(u_multiplier_pp1_10 [9]),
    .B(u_multiplier_pp1_10 [10]),
    .Z(u_multiplier_STAGE2_acci_pp2_10_0__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_10_0__24_  (.A1(u_multiplier_STAGE2_acci_pp2_10_0__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_10_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_10_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_10_0__25_  (.A(u_multiplier_STAGE2_acci_pp2_10_0__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_10_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_10_0__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_10_0__26_  (.A1(u_multiplier_STAGE2_acci_pp2_10_0__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_10_0__16_ ),
    .ZN(u_multiplier_pp2_10 [0]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_10_0__27_  (.A1(u_multiplier_pp1_10 [8]),
    .A2(u_multiplier_pp1_10 [7]),
    .B1(u_multiplier_pp1_10 [9]),
    .B2(u_multiplier_pp1_10 [10]),
    .ZN(u_multiplier_STAGE2_acci_pp2_10_0__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_10_0__28_  (.A1(u_multiplier_STAGE2_acci_pp2_10_0__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_10_0__17_ ),
    .ZN(u_multiplier_pp2_11 [3]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_11_0__21_  (.A1(u_multiplier_pp1_11 [9]),
    .A2(u_multiplier_pp1_11 [8]),
    .A3(u_multiplier_pp1_11 [10]),
    .ZN(u_multiplier_STAGE2_acci_pp2_11_0__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_11_0__22_  (.A(u_multiplier_pp1_11 [9]),
    .B(u_multiplier_pp1_11 [8]),
    .Z(u_multiplier_STAGE2_acci_pp2_11_0__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_11_0__23_  (.A(u_multiplier_pp1_11 [10]),
    .B(u_multiplier_pp1_11 [11]),
    .Z(u_multiplier_STAGE2_acci_pp2_11_0__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_11_0__24_  (.A1(u_multiplier_STAGE2_acci_pp2_11_0__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_11_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_11_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_11_0__25_  (.A(u_multiplier_STAGE2_acci_pp2_11_0__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_11_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_11_0__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_11_0__26_  (.A1(u_multiplier_STAGE2_acci_pp2_11_0__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_11_0__16_ ),
    .ZN(u_multiplier_pp2_11 [0]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_11_0__27_  (.A1(u_multiplier_pp1_11 [9]),
    .A2(u_multiplier_pp1_11 [8]),
    .B1(u_multiplier_pp1_11 [10]),
    .B2(u_multiplier_pp1_11 [11]),
    .ZN(u_multiplier_STAGE2_acci_pp2_11_0__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_11_0__28_  (.A1(u_multiplier_STAGE2_acci_pp2_11_0__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_11_0__17_ ),
    .ZN(u_multiplier_pp2_12 [4]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_11_1__21_  (.A1(u_multiplier_pp1_11 [5]),
    .A2(u_multiplier_pp1_11 [4]),
    .A3(u_multiplier_pp1_11 [6]),
    .ZN(u_multiplier_STAGE2_acci_pp2_11_1__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_11_1__22_  (.A(u_multiplier_pp1_11 [5]),
    .B(u_multiplier_pp1_11 [4]),
    .Z(u_multiplier_STAGE2_acci_pp2_11_1__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_11_1__23_  (.A(u_multiplier_pp1_11 [6]),
    .B(u_multiplier_pp1_11 [7]),
    .Z(u_multiplier_STAGE2_acci_pp2_11_1__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_11_1__24_  (.A1(u_multiplier_STAGE2_acci_pp2_11_1__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_11_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_11_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_11_1__25_  (.A(u_multiplier_STAGE2_acci_pp2_11_1__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_11_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_11_1__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_11_1__26_  (.A1(u_multiplier_STAGE2_acci_pp2_11_1__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_11_1__16_ ),
    .ZN(u_multiplier_pp2_11 [1]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_11_1__27_  (.A1(u_multiplier_pp1_11 [5]),
    .A2(u_multiplier_pp1_11 [4]),
    .B1(u_multiplier_pp1_11 [6]),
    .B2(u_multiplier_pp1_11 [7]),
    .ZN(u_multiplier_STAGE2_acci_pp2_11_1__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_11_1__28_  (.A1(u_multiplier_STAGE2_acci_pp2_11_1__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_11_1__17_ ),
    .ZN(u_multiplier_pp2_12 [3]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_12_0__21_  (.A1(u_multiplier_pp1_12 [10]),
    .A2(u_multiplier_pp1_12 [9]),
    .A3(u_multiplier_pp1_12 [11]),
    .ZN(u_multiplier_STAGE2_acci_pp2_12_0__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_12_0__22_  (.A(u_multiplier_pp1_12 [10]),
    .B(u_multiplier_pp1_12 [9]),
    .Z(u_multiplier_STAGE2_acci_pp2_12_0__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_12_0__23_  (.A(u_multiplier_pp1_12 [11]),
    .B(u_multiplier_pp1_12 [12]),
    .Z(u_multiplier_STAGE2_acci_pp2_12_0__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_12_0__24_  (.A1(u_multiplier_STAGE2_acci_pp2_12_0__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_12_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_12_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_12_0__25_  (.A(u_multiplier_STAGE2_acci_pp2_12_0__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_12_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_12_0__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_12_0__26_  (.A1(u_multiplier_STAGE2_acci_pp2_12_0__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_12_0__16_ ),
    .ZN(u_multiplier_pp2_12 [0]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_12_0__27_  (.A1(u_multiplier_pp1_12 [10]),
    .A2(u_multiplier_pp1_12 [9]),
    .B1(u_multiplier_pp1_12 [11]),
    .B2(u_multiplier_pp1_12 [12]),
    .ZN(u_multiplier_STAGE2_acci_pp2_12_0__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_12_0__28_  (.A1(u_multiplier_STAGE2_acci_pp2_12_0__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_12_0__17_ ),
    .ZN(u_multiplier_pp2_13 [5]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_12_1__21_  (.A1(u_multiplier_pp1_12 [6]),
    .A2(u_multiplier_pp1_12 [5]),
    .A3(u_multiplier_pp1_12 [7]),
    .ZN(u_multiplier_STAGE2_acci_pp2_12_1__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_12_1__22_  (.A(u_multiplier_pp1_12 [6]),
    .B(u_multiplier_pp1_12 [5]),
    .Z(u_multiplier_STAGE2_acci_pp2_12_1__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_12_1__23_  (.A(u_multiplier_pp1_12 [7]),
    .B(u_multiplier_pp1_12 [8]),
    .Z(u_multiplier_STAGE2_acci_pp2_12_1__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_12_1__24_  (.A1(u_multiplier_STAGE2_acci_pp2_12_1__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_12_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_12_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_12_1__25_  (.A(u_multiplier_STAGE2_acci_pp2_12_1__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_12_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_12_1__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_12_1__26_  (.A1(u_multiplier_STAGE2_acci_pp2_12_1__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_12_1__16_ ),
    .ZN(u_multiplier_pp2_12 [1]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_12_1__27_  (.A1(u_multiplier_pp1_12 [6]),
    .A2(u_multiplier_pp1_12 [5]),
    .B1(u_multiplier_pp1_12 [7]),
    .B2(u_multiplier_pp1_12 [8]),
    .ZN(u_multiplier_STAGE2_acci_pp2_12_1__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_12_1__28_  (.A1(u_multiplier_STAGE2_acci_pp2_12_1__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_12_1__17_ ),
    .ZN(u_multiplier_pp2_13 [4]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_13_0__21_  (.A1(u_multiplier_pp1_13 [11]),
    .A2(u_multiplier_pp1_13 [10]),
    .A3(u_multiplier_pp1_13 [12]),
    .ZN(u_multiplier_STAGE2_acci_pp2_13_0__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_13_0__22_  (.A(u_multiplier_pp1_13 [11]),
    .B(u_multiplier_pp1_13 [10]),
    .Z(u_multiplier_STAGE2_acci_pp2_13_0__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_13_0__23_  (.A(u_multiplier_pp1_13 [12]),
    .B(u_multiplier_pp1_13 [13]),
    .Z(u_multiplier_STAGE2_acci_pp2_13_0__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_13_0__24_  (.A1(u_multiplier_STAGE2_acci_pp2_13_0__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_13_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_13_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_13_0__25_  (.A(u_multiplier_STAGE2_acci_pp2_13_0__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_13_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_13_0__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_13_0__26_  (.A1(u_multiplier_STAGE2_acci_pp2_13_0__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_13_0__16_ ),
    .ZN(u_multiplier_pp2_13 [0]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_13_0__27_  (.A1(u_multiplier_pp1_13 [11]),
    .A2(u_multiplier_pp1_13 [10]),
    .B1(u_multiplier_pp1_13 [12]),
    .B2(u_multiplier_pp1_13 [13]),
    .ZN(u_multiplier_STAGE2_acci_pp2_13_0__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_13_0__28_  (.A1(u_multiplier_STAGE2_acci_pp2_13_0__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_13_0__17_ ),
    .ZN(u_multiplier_pp2_14 [6]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_13_1__21_  (.A1(u_multiplier_pp1_13 [7]),
    .A2(u_multiplier_pp1_13 [6]),
    .A3(u_multiplier_pp1_13 [8]),
    .ZN(u_multiplier_STAGE2_acci_pp2_13_1__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_13_1__22_  (.A(u_multiplier_pp1_13 [7]),
    .B(u_multiplier_pp1_13 [6]),
    .Z(u_multiplier_STAGE2_acci_pp2_13_1__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_13_1__23_  (.A(u_multiplier_pp1_13 [8]),
    .B(u_multiplier_pp1_13 [9]),
    .Z(u_multiplier_STAGE2_acci_pp2_13_1__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_13_1__24_  (.A1(u_multiplier_STAGE2_acci_pp2_13_1__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_13_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_13_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_13_1__25_  (.A(u_multiplier_STAGE2_acci_pp2_13_1__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_13_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_13_1__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_13_1__26_  (.A1(u_multiplier_STAGE2_acci_pp2_13_1__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_13_1__16_ ),
    .ZN(u_multiplier_pp2_13 [1]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_13_1__27_  (.A1(u_multiplier_pp1_13 [7]),
    .A2(u_multiplier_pp1_13 [6]),
    .B1(u_multiplier_pp1_13 [8]),
    .B2(u_multiplier_pp1_13 [9]),
    .ZN(u_multiplier_STAGE2_acci_pp2_13_1__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_13_1__28_  (.A1(u_multiplier_STAGE2_acci_pp2_13_1__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_13_1__17_ ),
    .ZN(u_multiplier_pp2_14 [5]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_13_2__21_  (.A1(u_multiplier_pp1_13 [3]),
    .A2(u_multiplier_pp1_13 [2]),
    .A3(u_multiplier_pp1_13 [4]),
    .ZN(u_multiplier_STAGE2_acci_pp2_13_2__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_13_2__22_  (.A(u_multiplier_pp1_13 [3]),
    .B(u_multiplier_pp1_13 [2]),
    .Z(u_multiplier_STAGE2_acci_pp2_13_2__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_13_2__23_  (.A(u_multiplier_pp1_13 [4]),
    .B(u_multiplier_pp1_13 [5]),
    .Z(u_multiplier_STAGE2_acci_pp2_13_2__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_13_2__24_  (.A1(u_multiplier_STAGE2_acci_pp2_13_2__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_13_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_13_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_13_2__25_  (.A(u_multiplier_STAGE2_acci_pp2_13_2__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_13_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_13_2__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_13_2__26_  (.A1(u_multiplier_STAGE2_acci_pp2_13_2__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_13_2__16_ ),
    .ZN(u_multiplier_pp2_13 [2]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_13_2__27_  (.A1(u_multiplier_pp1_13 [3]),
    .A2(u_multiplier_pp1_13 [2]),
    .B1(u_multiplier_pp1_13 [4]),
    .B2(u_multiplier_pp1_13 [5]),
    .ZN(u_multiplier_STAGE2_acci_pp2_13_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_13_2__28_  (.A1(u_multiplier_STAGE2_acci_pp2_13_2__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_13_2__17_ ),
    .ZN(u_multiplier_pp2_14 [4]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_14_0__21_  (.A1(u_multiplier_pp1_14 [12]),
    .A2(u_multiplier_pp1_14 [11]),
    .A3(u_multiplier_pp1_14 [13]),
    .ZN(u_multiplier_STAGE2_acci_pp2_14_0__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_14_0__22_  (.A(u_multiplier_pp1_14 [12]),
    .B(u_multiplier_pp1_14 [11]),
    .Z(u_multiplier_STAGE2_acci_pp2_14_0__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_14_0__23_  (.A(u_multiplier_pp1_14 [13]),
    .B(u_multiplier_pp1_14 [14]),
    .Z(u_multiplier_STAGE2_acci_pp2_14_0__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_14_0__24_  (.A1(u_multiplier_STAGE2_acci_pp2_14_0__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_14_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_14_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_14_0__25_  (.A(u_multiplier_STAGE2_acci_pp2_14_0__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_14_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_14_0__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_14_0__26_  (.A1(u_multiplier_STAGE2_acci_pp2_14_0__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_14_0__16_ ),
    .ZN(u_multiplier_pp2_14 [0]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_14_0__27_  (.A1(u_multiplier_pp1_14 [12]),
    .A2(u_multiplier_pp1_14 [11]),
    .B1(u_multiplier_pp1_14 [13]),
    .B2(u_multiplier_pp1_14 [14]),
    .ZN(u_multiplier_STAGE2_acci_pp2_14_0__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_14_0__28_  (.A1(u_multiplier_STAGE2_acci_pp2_14_0__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_14_0__17_ ),
    .ZN(u_multiplier_pp2_15 [7]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_14_1__21_  (.A1(u_multiplier_pp1_14 [8]),
    .A2(u_multiplier_pp1_14 [7]),
    .A3(u_multiplier_pp1_14 [9]),
    .ZN(u_multiplier_STAGE2_acci_pp2_14_1__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_14_1__22_  (.A(u_multiplier_pp1_14 [8]),
    .B(u_multiplier_pp1_14 [7]),
    .Z(u_multiplier_STAGE2_acci_pp2_14_1__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_14_1__23_  (.A(u_multiplier_pp1_14 [9]),
    .B(u_multiplier_pp1_14 [10]),
    .Z(u_multiplier_STAGE2_acci_pp2_14_1__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_14_1__24_  (.A1(u_multiplier_STAGE2_acci_pp2_14_1__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_14_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_14_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_14_1__25_  (.A(u_multiplier_STAGE2_acci_pp2_14_1__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_14_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_14_1__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_14_1__26_  (.A1(u_multiplier_STAGE2_acci_pp2_14_1__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_14_1__16_ ),
    .ZN(u_multiplier_pp2_14 [1]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_14_1__27_  (.A1(u_multiplier_pp1_14 [8]),
    .A2(u_multiplier_pp1_14 [7]),
    .B1(u_multiplier_pp1_14 [9]),
    .B2(u_multiplier_pp1_14 [10]),
    .ZN(u_multiplier_STAGE2_acci_pp2_14_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_14_1__28_  (.A1(u_multiplier_STAGE2_acci_pp2_14_1__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_14_1__17_ ),
    .ZN(u_multiplier_pp2_15 [6]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_14_2__21_  (.A1(u_multiplier_pp1_14 [4]),
    .A2(u_multiplier_pp1_14 [3]),
    .A3(u_multiplier_pp1_14 [5]),
    .ZN(u_multiplier_STAGE2_acci_pp2_14_2__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_14_2__22_  (.A(u_multiplier_pp1_14 [4]),
    .B(u_multiplier_pp1_14 [3]),
    .Z(u_multiplier_STAGE2_acci_pp2_14_2__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_14_2__23_  (.A(u_multiplier_pp1_14 [5]),
    .B(u_multiplier_pp1_14 [6]),
    .Z(u_multiplier_STAGE2_acci_pp2_14_2__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_14_2__24_  (.A1(u_multiplier_STAGE2_acci_pp2_14_2__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_14_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_14_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_14_2__25_  (.A(u_multiplier_STAGE2_acci_pp2_14_2__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_14_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_14_2__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_14_2__26_  (.A1(u_multiplier_STAGE2_acci_pp2_14_2__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_14_2__16_ ),
    .ZN(u_multiplier_pp2_14 [2]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_14_2__27_  (.A1(u_multiplier_pp1_14 [4]),
    .A2(u_multiplier_pp1_14 [3]),
    .B1(u_multiplier_pp1_14 [5]),
    .B2(u_multiplier_pp1_14 [6]),
    .ZN(u_multiplier_STAGE2_acci_pp2_14_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_14_2__28_  (.A1(u_multiplier_STAGE2_acci_pp2_14_2__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_14_2__17_ ),
    .ZN(u_multiplier_pp2_15 [5]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_15_0__21_  (.A1(u_multiplier_pp1_15 [13]),
    .A2(u_multiplier_pp1_15 [12]),
    .A3(u_multiplier_pp1_15 [14]),
    .ZN(u_multiplier_STAGE2_acci_pp2_15_0__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_15_0__22_  (.A(u_multiplier_pp1_15 [13]),
    .B(u_multiplier_pp1_15 [12]),
    .Z(u_multiplier_STAGE2_acci_pp2_15_0__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_15_0__23_  (.A(u_multiplier_pp1_15 [14]),
    .B(u_multiplier_pp1_15 [15]),
    .Z(u_multiplier_STAGE2_acci_pp2_15_0__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_15_0__24_  (.A1(u_multiplier_STAGE2_acci_pp2_15_0__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_15_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_15_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_15_0__25_  (.A(u_multiplier_STAGE2_acci_pp2_15_0__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_15_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_15_0__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_15_0__26_  (.A1(u_multiplier_STAGE2_acci_pp2_15_0__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_15_0__16_ ),
    .ZN(u_multiplier_pp2_15 [0]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_15_0__27_  (.A1(u_multiplier_pp1_15 [13]),
    .A2(u_multiplier_pp1_15 [12]),
    .B1(u_multiplier_pp1_15 [14]),
    .B2(u_multiplier_pp1_15 [15]),
    .ZN(u_multiplier_STAGE2_acci_pp2_15_0__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_15_0__28_  (.A1(u_multiplier_STAGE2_acci_pp2_15_0__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_15_0__17_ ),
    .ZN(u_multiplier_pp2_16 [7]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_15_1__21_  (.A1(u_multiplier_pp1_15 [9]),
    .A2(u_multiplier_pp1_15 [8]),
    .A3(u_multiplier_pp1_15 [10]),
    .ZN(u_multiplier_STAGE2_acci_pp2_15_1__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_15_1__22_  (.A(u_multiplier_pp1_15 [9]),
    .B(u_multiplier_pp1_15 [8]),
    .Z(u_multiplier_STAGE2_acci_pp2_15_1__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_15_1__23_  (.A(u_multiplier_pp1_15 [10]),
    .B(u_multiplier_pp1_15 [11]),
    .Z(u_multiplier_STAGE2_acci_pp2_15_1__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_15_1__24_  (.A1(u_multiplier_STAGE2_acci_pp2_15_1__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_15_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_15_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_15_1__25_  (.A(u_multiplier_STAGE2_acci_pp2_15_1__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_15_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_15_1__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_15_1__26_  (.A1(u_multiplier_STAGE2_acci_pp2_15_1__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_15_1__16_ ),
    .ZN(u_multiplier_pp2_15 [1]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_15_1__27_  (.A1(u_multiplier_pp1_15 [9]),
    .A2(u_multiplier_pp1_15 [8]),
    .B1(u_multiplier_pp1_15 [10]),
    .B2(u_multiplier_pp1_15 [11]),
    .ZN(u_multiplier_STAGE2_acci_pp2_15_1__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_15_1__28_  (.A1(u_multiplier_STAGE2_acci_pp2_15_1__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_15_1__17_ ),
    .ZN(u_multiplier_pp2_16 [6]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_15_2__21_  (.A1(u_multiplier_pp1_15 [5]),
    .A2(u_multiplier_pp1_15 [4]),
    .A3(u_multiplier_pp1_15 [6]),
    .ZN(u_multiplier_STAGE2_acci_pp2_15_2__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_15_2__22_  (.A(u_multiplier_pp1_15 [5]),
    .B(u_multiplier_pp1_15 [4]),
    .Z(u_multiplier_STAGE2_acci_pp2_15_2__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_15_2__23_  (.A(u_multiplier_pp1_15 [6]),
    .B(u_multiplier_pp1_15 [7]),
    .Z(u_multiplier_STAGE2_acci_pp2_15_2__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_15_2__24_  (.A1(u_multiplier_STAGE2_acci_pp2_15_2__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_15_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_15_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_15_2__25_  (.A(u_multiplier_STAGE2_acci_pp2_15_2__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_15_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_15_2__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_15_2__26_  (.A1(u_multiplier_STAGE2_acci_pp2_15_2__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_15_2__16_ ),
    .ZN(u_multiplier_pp2_15 [2]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_15_2__27_  (.A1(u_multiplier_pp1_15 [5]),
    .A2(u_multiplier_pp1_15 [4]),
    .B1(u_multiplier_pp1_15 [6]),
    .B2(u_multiplier_pp1_15 [7]),
    .ZN(u_multiplier_STAGE2_acci_pp2_15_2__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_15_2__28_  (.A1(u_multiplier_STAGE2_acci_pp2_15_2__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_15_2__17_ ),
    .ZN(u_multiplier_pp2_16 [5]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_15_3__21_  (.A1(u_multiplier_pp1_15 [1]),
    .A2(u_multiplier_pp1_15 [0]),
    .A3(u_multiplier_pp1_15 [2]),
    .ZN(u_multiplier_STAGE2_acci_pp2_15_3__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_15_3__22_  (.A(u_multiplier_pp1_15 [1]),
    .B(u_multiplier_pp1_15 [0]),
    .Z(u_multiplier_STAGE2_acci_pp2_15_3__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_15_3__23_  (.A(u_multiplier_pp1_15 [2]),
    .B(u_multiplier_pp1_15 [3]),
    .Z(u_multiplier_STAGE2_acci_pp2_15_3__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_15_3__24_  (.A1(u_multiplier_STAGE2_acci_pp2_15_3__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_15_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_15_3__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_15_3__25_  (.A(u_multiplier_STAGE2_acci_pp2_15_3__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_15_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_15_3__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_15_3__26_  (.A1(u_multiplier_STAGE2_acci_pp2_15_3__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_15_3__16_ ),
    .ZN(u_multiplier_pp2_15 [3]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_15_3__27_  (.A1(u_multiplier_pp1_15 [1]),
    .A2(u_multiplier_pp1_15 [0]),
    .B1(u_multiplier_pp1_15 [2]),
    .B2(u_multiplier_pp1_15 [3]),
    .ZN(u_multiplier_STAGE2_acci_pp2_15_3__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_15_3__28_  (.A1(u_multiplier_STAGE2_acci_pp2_15_3__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_15_3__17_ ),
    .ZN(u_multiplier_pp2_16 [4]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_16_0__21_  (.A1(u_multiplier_pp1_16 [13]),
    .A2(u_multiplier_pp1_16 [12]),
    .A3(u_multiplier_pp1_16 [14]),
    .ZN(u_multiplier_STAGE2_acci_pp2_16_0__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_16_0__22_  (.A(u_multiplier_pp1_16 [13]),
    .B(u_multiplier_pp1_16 [12]),
    .Z(u_multiplier_STAGE2_acci_pp2_16_0__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_16_0__23_  (.A(u_multiplier_pp1_16 [14]),
    .B(u_multiplier_pp1_16 [15]),
    .Z(u_multiplier_STAGE2_acci_pp2_16_0__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_16_0__24_  (.A1(u_multiplier_STAGE2_acci_pp2_16_0__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_16_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_16_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_16_0__25_  (.A(u_multiplier_STAGE2_acci_pp2_16_0__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_16_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_16_0__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_16_0__26_  (.A1(u_multiplier_STAGE2_acci_pp2_16_0__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_16_0__16_ ),
    .ZN(u_multiplier_pp2_16 [0]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_16_0__27_  (.A1(u_multiplier_pp1_16 [13]),
    .A2(u_multiplier_pp1_16 [12]),
    .B1(u_multiplier_pp1_16 [14]),
    .B2(u_multiplier_pp1_16 [15]),
    .ZN(u_multiplier_STAGE2_acci_pp2_16_0__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_16_0__28_  (.A1(u_multiplier_STAGE2_acci_pp2_16_0__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_16_0__17_ ),
    .ZN(u_multiplier_pp2_17 [7]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_16_1__21_  (.A1(u_multiplier_pp1_16 [9]),
    .A2(u_multiplier_pp1_16 [8]),
    .A3(u_multiplier_pp1_16 [10]),
    .ZN(u_multiplier_STAGE2_acci_pp2_16_1__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_16_1__22_  (.A(u_multiplier_pp1_16 [9]),
    .B(u_multiplier_pp1_16 [8]),
    .Z(u_multiplier_STAGE2_acci_pp2_16_1__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_16_1__23_  (.A(u_multiplier_pp1_16 [10]),
    .B(u_multiplier_pp1_16 [11]),
    .Z(u_multiplier_STAGE2_acci_pp2_16_1__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_16_1__24_  (.A1(u_multiplier_STAGE2_acci_pp2_16_1__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_16_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_16_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_16_1__25_  (.A(u_multiplier_STAGE2_acci_pp2_16_1__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_16_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_16_1__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_16_1__26_  (.A1(u_multiplier_STAGE2_acci_pp2_16_1__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_16_1__16_ ),
    .ZN(u_multiplier_pp2_16 [1]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_16_1__27_  (.A1(u_multiplier_pp1_16 [9]),
    .A2(u_multiplier_pp1_16 [8]),
    .B1(u_multiplier_pp1_16 [10]),
    .B2(u_multiplier_pp1_16 [11]),
    .ZN(u_multiplier_STAGE2_acci_pp2_16_1__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_16_1__28_  (.A1(u_multiplier_STAGE2_acci_pp2_16_1__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_16_1__17_ ),
    .ZN(u_multiplier_pp2_17 [6]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_16_2__21_  (.A1(u_multiplier_pp1_16 [5]),
    .A2(u_multiplier_pp1_16 [4]),
    .A3(u_multiplier_pp1_16 [6]),
    .ZN(u_multiplier_STAGE2_acci_pp2_16_2__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_16_2__22_  (.A(u_multiplier_pp1_16 [5]),
    .B(u_multiplier_pp1_16 [4]),
    .Z(u_multiplier_STAGE2_acci_pp2_16_2__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_16_2__23_  (.A(u_multiplier_pp1_16 [6]),
    .B(u_multiplier_pp1_16 [7]),
    .Z(u_multiplier_STAGE2_acci_pp2_16_2__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_16_2__24_  (.A1(u_multiplier_STAGE2_acci_pp2_16_2__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_16_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_16_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_16_2__25_  (.A(u_multiplier_STAGE2_acci_pp2_16_2__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_16_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_16_2__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_16_2__26_  (.A1(u_multiplier_STAGE2_acci_pp2_16_2__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_16_2__16_ ),
    .ZN(u_multiplier_pp2_16 [2]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_16_2__27_  (.A1(u_multiplier_pp1_16 [5]),
    .A2(u_multiplier_pp1_16 [4]),
    .B1(u_multiplier_pp1_16 [6]),
    .B2(u_multiplier_pp1_16 [7]),
    .ZN(u_multiplier_STAGE2_acci_pp2_16_2__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_16_2__28_  (.A1(u_multiplier_STAGE2_acci_pp2_16_2__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_16_2__17_ ),
    .ZN(u_multiplier_pp2_17 [5]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_16_3__21_  (.A1(u_multiplier_pp1_16 [1]),
    .A2(u_multiplier_pp1_16 [0]),
    .A3(u_multiplier_pp1_16 [2]),
    .ZN(u_multiplier_STAGE2_acci_pp2_16_3__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_16_3__22_  (.A(u_multiplier_pp1_16 [1]),
    .B(u_multiplier_pp1_16 [0]),
    .Z(u_multiplier_STAGE2_acci_pp2_16_3__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_16_3__23_  (.A(u_multiplier_pp1_16 [2]),
    .B(u_multiplier_pp1_16 [3]),
    .Z(u_multiplier_STAGE2_acci_pp2_16_3__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_16_3__24_  (.A1(u_multiplier_STAGE2_acci_pp2_16_3__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_16_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_16_3__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_16_3__25_  (.A(u_multiplier_STAGE2_acci_pp2_16_3__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_16_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_16_3__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_16_3__26_  (.A1(u_multiplier_STAGE2_acci_pp2_16_3__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_16_3__16_ ),
    .ZN(u_multiplier_pp2_16 [3]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_16_3__27_  (.A1(u_multiplier_pp1_16 [1]),
    .A2(u_multiplier_pp1_16 [0]),
    .B1(u_multiplier_pp1_16 [2]),
    .B2(u_multiplier_pp1_16 [3]),
    .ZN(u_multiplier_STAGE2_acci_pp2_16_3__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_16_3__28_  (.A1(u_multiplier_STAGE2_acci_pp2_16_3__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_16_3__17_ ),
    .ZN(u_multiplier_pp2_17 [4]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_17_0__21_  (.A1(u_multiplier_pp1_17 [13]),
    .A2(u_multiplier_pp1_17 [12]),
    .A3(u_multiplier_pp1_17 [14]),
    .ZN(u_multiplier_STAGE2_acci_pp2_17_0__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_17_0__22_  (.A(u_multiplier_pp1_17 [13]),
    .B(u_multiplier_pp1_17 [12]),
    .Z(u_multiplier_STAGE2_acci_pp2_17_0__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_17_0__23_  (.A(u_multiplier_pp1_17 [14]),
    .B(u_multiplier_pp1_17 [15]),
    .Z(u_multiplier_STAGE2_acci_pp2_17_0__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_17_0__24_  (.A1(u_multiplier_STAGE2_acci_pp2_17_0__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_17_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_17_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_17_0__25_  (.A(u_multiplier_STAGE2_acci_pp2_17_0__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_17_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_17_0__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_17_0__26_  (.A1(u_multiplier_STAGE2_acci_pp2_17_0__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_17_0__16_ ),
    .ZN(u_multiplier_pp2_17 [0]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_17_0__27_  (.A1(u_multiplier_pp1_17 [13]),
    .A2(u_multiplier_pp1_17 [12]),
    .B1(u_multiplier_pp1_17 [14]),
    .B2(u_multiplier_pp1_17 [15]),
    .ZN(u_multiplier_STAGE2_acci_pp2_17_0__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_17_0__28_  (.A1(u_multiplier_STAGE2_acci_pp2_17_0__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_17_0__17_ ),
    .ZN(u_multiplier_pp2_18 [7]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_17_1__21_  (.A1(u_multiplier_pp1_17 [9]),
    .A2(u_multiplier_pp1_17 [8]),
    .A3(u_multiplier_pp1_17 [10]),
    .ZN(u_multiplier_STAGE2_acci_pp2_17_1__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_17_1__22_  (.A(u_multiplier_pp1_17 [9]),
    .B(u_multiplier_pp1_17 [8]),
    .Z(u_multiplier_STAGE2_acci_pp2_17_1__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_17_1__23_  (.A(u_multiplier_pp1_17 [10]),
    .B(u_multiplier_pp1_17 [11]),
    .Z(u_multiplier_STAGE2_acci_pp2_17_1__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_17_1__24_  (.A1(u_multiplier_STAGE2_acci_pp2_17_1__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_17_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_17_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_17_1__25_  (.A(u_multiplier_STAGE2_acci_pp2_17_1__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_17_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_17_1__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_17_1__26_  (.A1(u_multiplier_STAGE2_acci_pp2_17_1__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_17_1__16_ ),
    .ZN(u_multiplier_pp2_17 [1]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_17_1__27_  (.A1(u_multiplier_pp1_17 [9]),
    .A2(u_multiplier_pp1_17 [8]),
    .B1(u_multiplier_pp1_17 [10]),
    .B2(u_multiplier_pp1_17 [11]),
    .ZN(u_multiplier_STAGE2_acci_pp2_17_1__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_17_1__28_  (.A1(u_multiplier_STAGE2_acci_pp2_17_1__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_17_1__17_ ),
    .ZN(u_multiplier_pp2_18 [6]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_17_2__21_  (.A1(u_multiplier_pp1_17 [5]),
    .A2(u_multiplier_pp1_17 [4]),
    .A3(u_multiplier_pp1_17 [6]),
    .ZN(u_multiplier_STAGE2_acci_pp2_17_2__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_17_2__22_  (.A(u_multiplier_pp1_17 [5]),
    .B(u_multiplier_pp1_17 [4]),
    .Z(u_multiplier_STAGE2_acci_pp2_17_2__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_17_2__23_  (.A(u_multiplier_pp1_17 [6]),
    .B(u_multiplier_pp1_17 [7]),
    .Z(u_multiplier_STAGE2_acci_pp2_17_2__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_17_2__24_  (.A1(u_multiplier_STAGE2_acci_pp2_17_2__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_17_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_17_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_17_2__25_  (.A(u_multiplier_STAGE2_acci_pp2_17_2__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_17_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_17_2__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_17_2__26_  (.A1(u_multiplier_STAGE2_acci_pp2_17_2__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_17_2__16_ ),
    .ZN(u_multiplier_pp2_17 [2]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_17_2__27_  (.A1(u_multiplier_pp1_17 [5]),
    .A2(u_multiplier_pp1_17 [4]),
    .B1(u_multiplier_pp1_17 [6]),
    .B2(u_multiplier_pp1_17 [7]),
    .ZN(u_multiplier_STAGE2_acci_pp2_17_2__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_17_2__28_  (.A1(u_multiplier_STAGE2_acci_pp2_17_2__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_17_2__17_ ),
    .ZN(u_multiplier_pp2_18 [5]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_17_3__21_  (.A1(u_multiplier_pp1_17 [1]),
    .A2(u_multiplier_pp1_17 [0]),
    .A3(u_multiplier_pp1_17 [2]),
    .ZN(u_multiplier_STAGE2_acci_pp2_17_3__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_17_3__22_  (.A(u_multiplier_pp1_17 [1]),
    .B(u_multiplier_pp1_17 [0]),
    .Z(u_multiplier_STAGE2_acci_pp2_17_3__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_17_3__23_  (.A(u_multiplier_pp1_17 [2]),
    .B(u_multiplier_pp1_17 [3]),
    .Z(u_multiplier_STAGE2_acci_pp2_17_3__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_17_3__24_  (.A1(u_multiplier_STAGE2_acci_pp2_17_3__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_17_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_17_3__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_17_3__25_  (.A(u_multiplier_STAGE2_acci_pp2_17_3__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_17_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_17_3__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_17_3__26_  (.A1(u_multiplier_STAGE2_acci_pp2_17_3__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_17_3__16_ ),
    .ZN(u_multiplier_pp2_17 [3]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_17_3__27_  (.A1(u_multiplier_pp1_17 [1]),
    .A2(u_multiplier_pp1_17 [0]),
    .B1(u_multiplier_pp1_17 [2]),
    .B2(u_multiplier_pp1_17 [3]),
    .ZN(u_multiplier_STAGE2_acci_pp2_17_3__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_17_3__28_  (.A1(u_multiplier_STAGE2_acci_pp2_17_3__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_17_3__17_ ),
    .ZN(u_multiplier_pp2_18 [4]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_18_0__21_  (.A1(u_multiplier_pp1_18 [13]),
    .A2(u_multiplier_pp1_18 [12]),
    .A3(u_multiplier_pp1_18 [14]),
    .ZN(u_multiplier_STAGE2_acci_pp2_18_0__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_18_0__22_  (.A(u_multiplier_pp1_18 [13]),
    .B(u_multiplier_pp1_18 [12]),
    .Z(u_multiplier_STAGE2_acci_pp2_18_0__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_18_0__23_  (.A(u_multiplier_pp1_18 [14]),
    .B(u_multiplier_pp1_18 [15]),
    .Z(u_multiplier_STAGE2_acci_pp2_18_0__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_18_0__24_  (.A1(u_multiplier_STAGE2_acci_pp2_18_0__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_18_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_18_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_18_0__25_  (.A(u_multiplier_STAGE2_acci_pp2_18_0__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_18_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_18_0__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_18_0__26_  (.A1(u_multiplier_STAGE2_acci_pp2_18_0__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_18_0__16_ ),
    .ZN(u_multiplier_pp2_18 [0]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_18_0__27_  (.A1(u_multiplier_pp1_18 [13]),
    .A2(u_multiplier_pp1_18 [12]),
    .B1(u_multiplier_pp1_18 [14]),
    .B2(u_multiplier_pp1_18 [15]),
    .ZN(u_multiplier_STAGE2_acci_pp2_18_0__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_18_0__28_  (.A1(u_multiplier_STAGE2_acci_pp2_18_0__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_18_0__17_ ),
    .ZN(u_multiplier_pp2_19 [7]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_18_1__21_  (.A1(u_multiplier_pp1_18 [9]),
    .A2(u_multiplier_pp1_18 [8]),
    .A3(u_multiplier_pp1_18 [10]),
    .ZN(u_multiplier_STAGE2_acci_pp2_18_1__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_18_1__22_  (.A(u_multiplier_pp1_18 [9]),
    .B(u_multiplier_pp1_18 [8]),
    .Z(u_multiplier_STAGE2_acci_pp2_18_1__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_18_1__23_  (.A(u_multiplier_pp1_18 [10]),
    .B(u_multiplier_pp1_18 [11]),
    .Z(u_multiplier_STAGE2_acci_pp2_18_1__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_18_1__24_  (.A1(u_multiplier_STAGE2_acci_pp2_18_1__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_18_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_18_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_18_1__25_  (.A(u_multiplier_STAGE2_acci_pp2_18_1__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_18_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_18_1__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_18_1__26_  (.A1(u_multiplier_STAGE2_acci_pp2_18_1__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_18_1__16_ ),
    .ZN(u_multiplier_pp2_18 [1]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_18_1__27_  (.A1(u_multiplier_pp1_18 [9]),
    .A2(u_multiplier_pp1_18 [8]),
    .B1(u_multiplier_pp1_18 [10]),
    .B2(u_multiplier_pp1_18 [11]),
    .ZN(u_multiplier_STAGE2_acci_pp2_18_1__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_18_1__28_  (.A1(u_multiplier_STAGE2_acci_pp2_18_1__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_18_1__17_ ),
    .ZN(u_multiplier_pp2_19 [6]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_18_2__21_  (.A1(u_multiplier_pp1_18 [5]),
    .A2(u_multiplier_pp1_18 [4]),
    .A3(u_multiplier_pp1_18 [6]),
    .ZN(u_multiplier_STAGE2_acci_pp2_18_2__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_18_2__22_  (.A(u_multiplier_pp1_18 [5]),
    .B(u_multiplier_pp1_18 [4]),
    .Z(u_multiplier_STAGE2_acci_pp2_18_2__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_18_2__23_  (.A(u_multiplier_pp1_18 [6]),
    .B(u_multiplier_pp1_18 [7]),
    .Z(u_multiplier_STAGE2_acci_pp2_18_2__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_18_2__24_  (.A1(u_multiplier_STAGE2_acci_pp2_18_2__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_18_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_18_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_18_2__25_  (.A(u_multiplier_STAGE2_acci_pp2_18_2__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_18_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_18_2__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_18_2__26_  (.A1(u_multiplier_STAGE2_acci_pp2_18_2__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_18_2__16_ ),
    .ZN(u_multiplier_pp2_18 [2]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_18_2__27_  (.A1(u_multiplier_pp1_18 [5]),
    .A2(u_multiplier_pp1_18 [4]),
    .B1(u_multiplier_pp1_18 [6]),
    .B2(u_multiplier_pp1_18 [7]),
    .ZN(u_multiplier_STAGE2_acci_pp2_18_2__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_18_2__28_  (.A1(u_multiplier_STAGE2_acci_pp2_18_2__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_18_2__17_ ),
    .ZN(u_multiplier_pp2_19 [5]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_18_3__21_  (.A1(u_multiplier_pp1_18 [1]),
    .A2(u_multiplier_pp1_18 [0]),
    .A3(u_multiplier_pp1_18 [2]),
    .ZN(u_multiplier_STAGE2_acci_pp2_18_3__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_18_3__22_  (.A(u_multiplier_pp1_18 [1]),
    .B(u_multiplier_pp1_18 [0]),
    .Z(u_multiplier_STAGE2_acci_pp2_18_3__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_18_3__23_  (.A(u_multiplier_pp1_18 [2]),
    .B(u_multiplier_pp1_18 [3]),
    .Z(u_multiplier_STAGE2_acci_pp2_18_3__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_18_3__24_  (.A1(u_multiplier_STAGE2_acci_pp2_18_3__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_18_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_18_3__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_18_3__25_  (.A(u_multiplier_STAGE2_acci_pp2_18_3__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_18_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_18_3__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_18_3__26_  (.A1(u_multiplier_STAGE2_acci_pp2_18_3__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_18_3__16_ ),
    .ZN(u_multiplier_pp2_18 [3]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_18_3__27_  (.A1(u_multiplier_pp1_18 [1]),
    .A2(u_multiplier_pp1_18 [0]),
    .B1(u_multiplier_pp1_18 [2]),
    .B2(u_multiplier_pp1_18 [3]),
    .ZN(u_multiplier_STAGE2_acci_pp2_18_3__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_18_3__28_  (.A1(u_multiplier_STAGE2_acci_pp2_18_3__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_18_3__17_ ),
    .ZN(u_multiplier_pp2_19 [4]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_19_0__21_  (.A1(u_multiplier_pp1_19 [13]),
    .A2(u_multiplier_pp1_19 [12]),
    .A3(u_multiplier_pp1_19 [14]),
    .ZN(u_multiplier_STAGE2_acci_pp2_19_0__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_19_0__22_  (.A(u_multiplier_pp1_19 [13]),
    .B(u_multiplier_pp1_19 [12]),
    .Z(u_multiplier_STAGE2_acci_pp2_19_0__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_19_0__23_  (.A(u_multiplier_pp1_19 [14]),
    .B(u_multiplier_pp1_19 [15]),
    .Z(u_multiplier_STAGE2_acci_pp2_19_0__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_19_0__24_  (.A1(u_multiplier_STAGE2_acci_pp2_19_0__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_19_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_19_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_19_0__25_  (.A(u_multiplier_STAGE2_acci_pp2_19_0__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_19_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_19_0__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_19_0__26_  (.A1(u_multiplier_STAGE2_acci_pp2_19_0__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_19_0__16_ ),
    .ZN(u_multiplier_pp2_19 [0]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_19_0__27_  (.A1(u_multiplier_pp1_19 [13]),
    .A2(u_multiplier_pp1_19 [12]),
    .B1(u_multiplier_pp1_19 [14]),
    .B2(u_multiplier_pp1_19 [15]),
    .ZN(u_multiplier_STAGE2_acci_pp2_19_0__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_19_0__28_  (.A1(u_multiplier_STAGE2_acci_pp2_19_0__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_19_0__17_ ),
    .ZN(u_multiplier_pp2_20 [7]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_19_1__21_  (.A1(u_multiplier_pp1_19 [9]),
    .A2(u_multiplier_pp1_19 [8]),
    .A3(u_multiplier_pp1_19 [10]),
    .ZN(u_multiplier_STAGE2_acci_pp2_19_1__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_19_1__22_  (.A(u_multiplier_pp1_19 [9]),
    .B(u_multiplier_pp1_19 [8]),
    .Z(u_multiplier_STAGE2_acci_pp2_19_1__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_19_1__23_  (.A(u_multiplier_pp1_19 [10]),
    .B(u_multiplier_pp1_19 [11]),
    .Z(u_multiplier_STAGE2_acci_pp2_19_1__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_19_1__24_  (.A1(u_multiplier_STAGE2_acci_pp2_19_1__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_19_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_19_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_19_1__25_  (.A(u_multiplier_STAGE2_acci_pp2_19_1__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_19_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_19_1__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_19_1__26_  (.A1(u_multiplier_STAGE2_acci_pp2_19_1__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_19_1__16_ ),
    .ZN(u_multiplier_pp2_19 [1]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_19_1__27_  (.A1(u_multiplier_pp1_19 [9]),
    .A2(u_multiplier_pp1_19 [8]),
    .B1(u_multiplier_pp1_19 [10]),
    .B2(u_multiplier_pp1_19 [11]),
    .ZN(u_multiplier_STAGE2_acci_pp2_19_1__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_19_1__28_  (.A1(u_multiplier_STAGE2_acci_pp2_19_1__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_19_1__17_ ),
    .ZN(u_multiplier_pp2_20 [6]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_19_2__21_  (.A1(u_multiplier_pp1_19 [5]),
    .A2(u_multiplier_pp1_19 [4]),
    .A3(u_multiplier_pp1_19 [6]),
    .ZN(u_multiplier_STAGE2_acci_pp2_19_2__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_19_2__22_  (.A(u_multiplier_pp1_19 [5]),
    .B(u_multiplier_pp1_19 [4]),
    .Z(u_multiplier_STAGE2_acci_pp2_19_2__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_19_2__23_  (.A(u_multiplier_pp1_19 [6]),
    .B(u_multiplier_pp1_19 [7]),
    .Z(u_multiplier_STAGE2_acci_pp2_19_2__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_19_2__24_  (.A1(u_multiplier_STAGE2_acci_pp2_19_2__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_19_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_19_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_19_2__25_  (.A(u_multiplier_STAGE2_acci_pp2_19_2__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_19_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_19_2__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_19_2__26_  (.A1(u_multiplier_STAGE2_acci_pp2_19_2__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_19_2__16_ ),
    .ZN(u_multiplier_pp2_19 [2]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_19_2__27_  (.A1(u_multiplier_pp1_19 [5]),
    .A2(u_multiplier_pp1_19 [4]),
    .B1(u_multiplier_pp1_19 [6]),
    .B2(u_multiplier_pp1_19 [7]),
    .ZN(u_multiplier_STAGE2_acci_pp2_19_2__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_19_2__28_  (.A1(u_multiplier_STAGE2_acci_pp2_19_2__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_19_2__17_ ),
    .ZN(u_multiplier_pp2_20 [5]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_19_3__21_  (.A1(u_multiplier_pp1_19 [1]),
    .A2(u_multiplier_pp1_19 [0]),
    .A3(u_multiplier_pp1_19 [2]),
    .ZN(u_multiplier_STAGE2_acci_pp2_19_3__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_19_3__22_  (.A(u_multiplier_pp1_19 [1]),
    .B(u_multiplier_pp1_19 [0]),
    .Z(u_multiplier_STAGE2_acci_pp2_19_3__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_19_3__23_  (.A(u_multiplier_pp1_19 [2]),
    .B(u_multiplier_pp1_19 [3]),
    .Z(u_multiplier_STAGE2_acci_pp2_19_3__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_19_3__24_  (.A1(u_multiplier_STAGE2_acci_pp2_19_3__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_19_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_19_3__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_19_3__25_  (.A(u_multiplier_STAGE2_acci_pp2_19_3__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_19_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_19_3__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_19_3__26_  (.A1(u_multiplier_STAGE2_acci_pp2_19_3__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_19_3__16_ ),
    .ZN(u_multiplier_pp2_19 [3]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_19_3__27_  (.A1(u_multiplier_pp1_19 [1]),
    .A2(u_multiplier_pp1_19 [0]),
    .B1(u_multiplier_pp1_19 [2]),
    .B2(u_multiplier_pp1_19 [3]),
    .ZN(u_multiplier_STAGE2_acci_pp2_19_3__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_19_3__28_  (.A1(u_multiplier_STAGE2_acci_pp2_19_3__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_19_3__17_ ),
    .ZN(u_multiplier_pp2_20 [4]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_20_0__21_  (.A1(u_multiplier_pp1_20 [13]),
    .A2(u_multiplier_pp1_20 [12]),
    .A3(u_multiplier_pp1_20 [14]),
    .ZN(u_multiplier_STAGE2_acci_pp2_20_0__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_20_0__22_  (.A(u_multiplier_pp1_20 [13]),
    .B(u_multiplier_pp1_20 [12]),
    .Z(u_multiplier_STAGE2_acci_pp2_20_0__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_20_0__23_  (.A(u_multiplier_pp1_20 [14]),
    .B(u_multiplier_pp1_20 [15]),
    .Z(u_multiplier_STAGE2_acci_pp2_20_0__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_20_0__24_  (.A1(u_multiplier_STAGE2_acci_pp2_20_0__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_20_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_20_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_20_0__25_  (.A(u_multiplier_STAGE2_acci_pp2_20_0__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_20_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_20_0__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_20_0__26_  (.A1(u_multiplier_STAGE2_acci_pp2_20_0__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_20_0__16_ ),
    .ZN(u_multiplier_pp2_20 [0]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_20_0__27_  (.A1(u_multiplier_pp1_20 [13]),
    .A2(u_multiplier_pp1_20 [12]),
    .B1(u_multiplier_pp1_20 [14]),
    .B2(u_multiplier_pp1_20 [15]),
    .ZN(u_multiplier_STAGE2_acci_pp2_20_0__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_20_0__28_  (.A1(u_multiplier_STAGE2_acci_pp2_20_0__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_20_0__17_ ),
    .ZN(u_multiplier_pp2_21 [7]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_20_1__21_  (.A1(u_multiplier_pp1_20 [9]),
    .A2(u_multiplier_pp1_20 [8]),
    .A3(u_multiplier_pp1_20 [10]),
    .ZN(u_multiplier_STAGE2_acci_pp2_20_1__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_20_1__22_  (.A(u_multiplier_pp1_20 [9]),
    .B(u_multiplier_pp1_20 [8]),
    .Z(u_multiplier_STAGE2_acci_pp2_20_1__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_20_1__23_  (.A(u_multiplier_pp1_20 [10]),
    .B(u_multiplier_pp1_20 [11]),
    .Z(u_multiplier_STAGE2_acci_pp2_20_1__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_20_1__24_  (.A1(u_multiplier_STAGE2_acci_pp2_20_1__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_20_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_20_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_20_1__25_  (.A(u_multiplier_STAGE2_acci_pp2_20_1__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_20_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_20_1__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_20_1__26_  (.A1(u_multiplier_STAGE2_acci_pp2_20_1__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_20_1__16_ ),
    .ZN(u_multiplier_pp2_20 [1]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_20_1__27_  (.A1(u_multiplier_pp1_20 [9]),
    .A2(u_multiplier_pp1_20 [8]),
    .B1(u_multiplier_pp1_20 [10]),
    .B2(u_multiplier_pp1_20 [11]),
    .ZN(u_multiplier_STAGE2_acci_pp2_20_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_20_1__28_  (.A1(u_multiplier_STAGE2_acci_pp2_20_1__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_20_1__17_ ),
    .ZN(u_multiplier_pp2_21 [6]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_20_2__21_  (.A1(u_multiplier_pp1_20 [5]),
    .A2(u_multiplier_pp1_20 [4]),
    .A3(u_multiplier_pp1_20 [6]),
    .ZN(u_multiplier_STAGE2_acci_pp2_20_2__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_20_2__22_  (.A(u_multiplier_pp1_20 [5]),
    .B(u_multiplier_pp1_20 [4]),
    .Z(u_multiplier_STAGE2_acci_pp2_20_2__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_20_2__23_  (.A(u_multiplier_pp1_20 [6]),
    .B(u_multiplier_pp1_20 [7]),
    .Z(u_multiplier_STAGE2_acci_pp2_20_2__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_20_2__24_  (.A1(u_multiplier_STAGE2_acci_pp2_20_2__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_20_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_20_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_20_2__25_  (.A(u_multiplier_STAGE2_acci_pp2_20_2__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_20_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_20_2__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_20_2__26_  (.A1(u_multiplier_STAGE2_acci_pp2_20_2__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_20_2__16_ ),
    .ZN(u_multiplier_pp2_20 [2]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_20_2__27_  (.A1(u_multiplier_pp1_20 [5]),
    .A2(u_multiplier_pp1_20 [4]),
    .B1(u_multiplier_pp1_20 [6]),
    .B2(u_multiplier_pp1_20 [7]),
    .ZN(u_multiplier_STAGE2_acci_pp2_20_2__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_20_2__28_  (.A1(u_multiplier_STAGE2_acci_pp2_20_2__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_20_2__17_ ),
    .ZN(u_multiplier_pp2_21 [5]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_20_3__21_  (.A1(u_multiplier_pp1_20 [1]),
    .A2(u_multiplier_pp1_20 [0]),
    .A3(u_multiplier_pp1_20 [2]),
    .ZN(u_multiplier_STAGE2_acci_pp2_20_3__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_20_3__22_  (.A(u_multiplier_pp1_20 [1]),
    .B(u_multiplier_pp1_20 [0]),
    .Z(u_multiplier_STAGE2_acci_pp2_20_3__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_20_3__23_  (.A(u_multiplier_pp1_20 [2]),
    .B(u_multiplier_pp1_20 [3]),
    .Z(u_multiplier_STAGE2_acci_pp2_20_3__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_20_3__24_  (.A1(u_multiplier_STAGE2_acci_pp2_20_3__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_20_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_20_3__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_20_3__25_  (.A(u_multiplier_STAGE2_acci_pp2_20_3__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_20_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_20_3__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_20_3__26_  (.A1(u_multiplier_STAGE2_acci_pp2_20_3__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_20_3__16_ ),
    .ZN(u_multiplier_pp2_20 [3]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_20_3__27_  (.A1(u_multiplier_pp1_20 [1]),
    .A2(u_multiplier_pp1_20 [0]),
    .B1(u_multiplier_pp1_20 [2]),
    .B2(u_multiplier_pp1_20 [3]),
    .ZN(u_multiplier_STAGE2_acci_pp2_20_3__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_20_3__28_  (.A1(u_multiplier_STAGE2_acci_pp2_20_3__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_20_3__17_ ),
    .ZN(u_multiplier_pp2_21 [4]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_21_0__21_  (.A1(u_multiplier_pp1_21 [13]),
    .A2(u_multiplier_pp1_21 [12]),
    .A3(u_multiplier_pp1_21 [14]),
    .ZN(u_multiplier_STAGE2_acci_pp2_21_0__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_21_0__22_  (.A(u_multiplier_pp1_21 [13]),
    .B(u_multiplier_pp1_21 [12]),
    .Z(u_multiplier_STAGE2_acci_pp2_21_0__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_21_0__23_  (.A(u_multiplier_pp1_21 [14]),
    .B(u_multiplier_pp1_21 [15]),
    .Z(u_multiplier_STAGE2_acci_pp2_21_0__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_21_0__24_  (.A1(u_multiplier_STAGE2_acci_pp2_21_0__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_21_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_21_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_21_0__25_  (.A(u_multiplier_STAGE2_acci_pp2_21_0__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_21_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_21_0__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_21_0__26_  (.A1(u_multiplier_STAGE2_acci_pp2_21_0__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_21_0__16_ ),
    .ZN(u_multiplier_pp2_21 [0]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_21_0__27_  (.A1(u_multiplier_pp1_21 [13]),
    .A2(u_multiplier_pp1_21 [12]),
    .B1(u_multiplier_pp1_21 [14]),
    .B2(u_multiplier_pp1_21 [15]),
    .ZN(u_multiplier_STAGE2_acci_pp2_21_0__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_21_0__28_  (.A1(u_multiplier_STAGE2_acci_pp2_21_0__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_21_0__17_ ),
    .ZN(u_multiplier_pp2_22 [7]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_21_1__21_  (.A1(u_multiplier_pp1_21 [9]),
    .A2(u_multiplier_pp1_21 [8]),
    .A3(u_multiplier_pp1_21 [10]),
    .ZN(u_multiplier_STAGE2_acci_pp2_21_1__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_21_1__22_  (.A(u_multiplier_pp1_21 [9]),
    .B(u_multiplier_pp1_21 [8]),
    .Z(u_multiplier_STAGE2_acci_pp2_21_1__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_21_1__23_  (.A(u_multiplier_pp1_21 [10]),
    .B(u_multiplier_pp1_21 [11]),
    .Z(u_multiplier_STAGE2_acci_pp2_21_1__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_21_1__24_  (.A1(u_multiplier_STAGE2_acci_pp2_21_1__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_21_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_21_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_21_1__25_  (.A(u_multiplier_STAGE2_acci_pp2_21_1__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_21_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_21_1__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_21_1__26_  (.A1(u_multiplier_STAGE2_acci_pp2_21_1__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_21_1__16_ ),
    .ZN(u_multiplier_pp2_21 [1]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_21_1__27_  (.A1(u_multiplier_pp1_21 [9]),
    .A2(u_multiplier_pp1_21 [8]),
    .B1(u_multiplier_pp1_21 [10]),
    .B2(u_multiplier_pp1_21 [11]),
    .ZN(u_multiplier_STAGE2_acci_pp2_21_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_21_1__28_  (.A1(u_multiplier_STAGE2_acci_pp2_21_1__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_21_1__17_ ),
    .ZN(u_multiplier_pp2_22 [6]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_21_2__21_  (.A1(u_multiplier_pp1_21 [5]),
    .A2(u_multiplier_pp1_21 [4]),
    .A3(u_multiplier_pp1_21 [6]),
    .ZN(u_multiplier_STAGE2_acci_pp2_21_2__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_21_2__22_  (.A(u_multiplier_pp1_21 [5]),
    .B(u_multiplier_pp1_21 [4]),
    .Z(u_multiplier_STAGE2_acci_pp2_21_2__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_21_2__23_  (.A(u_multiplier_pp1_21 [6]),
    .B(u_multiplier_pp1_21 [7]),
    .Z(u_multiplier_STAGE2_acci_pp2_21_2__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_21_2__24_  (.A1(u_multiplier_STAGE2_acci_pp2_21_2__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_21_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_21_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_21_2__25_  (.A(u_multiplier_STAGE2_acci_pp2_21_2__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_21_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_21_2__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_21_2__26_  (.A1(u_multiplier_STAGE2_acci_pp2_21_2__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_21_2__16_ ),
    .ZN(u_multiplier_pp2_21 [2]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_21_2__27_  (.A1(u_multiplier_pp1_21 [5]),
    .A2(u_multiplier_pp1_21 [4]),
    .B1(u_multiplier_pp1_21 [6]),
    .B2(u_multiplier_pp1_21 [7]),
    .ZN(u_multiplier_STAGE2_acci_pp2_21_2__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_21_2__28_  (.A1(u_multiplier_STAGE2_acci_pp2_21_2__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_21_2__17_ ),
    .ZN(u_multiplier_pp2_22 [5]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_21_3__21_  (.A1(u_multiplier_pp1_21 [1]),
    .A2(u_multiplier_pp1_21 [0]),
    .A3(u_multiplier_pp1_21 [2]),
    .ZN(u_multiplier_STAGE2_acci_pp2_21_3__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_21_3__22_  (.A(u_multiplier_pp1_21 [1]),
    .B(u_multiplier_pp1_21 [0]),
    .Z(u_multiplier_STAGE2_acci_pp2_21_3__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_21_3__23_  (.A(u_multiplier_pp1_21 [2]),
    .B(u_multiplier_pp1_21 [3]),
    .Z(u_multiplier_STAGE2_acci_pp2_21_3__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_21_3__24_  (.A1(u_multiplier_STAGE2_acci_pp2_21_3__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_21_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_21_3__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_21_3__25_  (.A(u_multiplier_STAGE2_acci_pp2_21_3__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_21_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_21_3__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_21_3__26_  (.A1(u_multiplier_STAGE2_acci_pp2_21_3__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_21_3__16_ ),
    .ZN(u_multiplier_pp2_21 [3]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_21_3__27_  (.A1(u_multiplier_pp1_21 [1]),
    .A2(u_multiplier_pp1_21 [0]),
    .B1(u_multiplier_pp1_21 [2]),
    .B2(u_multiplier_pp1_21 [3]),
    .ZN(u_multiplier_STAGE2_acci_pp2_21_3__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_21_3__28_  (.A1(u_multiplier_STAGE2_acci_pp2_21_3__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_21_3__17_ ),
    .ZN(u_multiplier_pp2_22 [4]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_22_0__21_  (.A1(u_multiplier_pp1_22 [13]),
    .A2(u_multiplier_pp1_22 [12]),
    .A3(u_multiplier_pp1_22 [14]),
    .ZN(u_multiplier_STAGE2_acci_pp2_22_0__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_22_0__22_  (.A(u_multiplier_pp1_22 [13]),
    .B(u_multiplier_pp1_22 [12]),
    .Z(u_multiplier_STAGE2_acci_pp2_22_0__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_22_0__23_  (.A(u_multiplier_pp1_22 [14]),
    .B(u_multiplier_pp1_22 [15]),
    .Z(u_multiplier_STAGE2_acci_pp2_22_0__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_22_0__24_  (.A1(u_multiplier_STAGE2_acci_pp2_22_0__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_22_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_22_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_22_0__25_  (.A(u_multiplier_STAGE2_acci_pp2_22_0__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_22_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_22_0__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_22_0__26_  (.A1(u_multiplier_STAGE2_acci_pp2_22_0__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_22_0__16_ ),
    .ZN(u_multiplier_pp2_22 [0]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_22_0__27_  (.A1(u_multiplier_pp1_22 [13]),
    .A2(u_multiplier_pp1_22 [12]),
    .B1(u_multiplier_pp1_22 [14]),
    .B2(u_multiplier_pp1_22 [15]),
    .ZN(u_multiplier_STAGE2_acci_pp2_22_0__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_22_0__28_  (.A1(u_multiplier_STAGE2_acci_pp2_22_0__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_22_0__17_ ),
    .ZN(u_multiplier_pp2_23 [7]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_22_1__21_  (.A1(u_multiplier_pp1_22 [9]),
    .A2(u_multiplier_pp1_22 [8]),
    .A3(u_multiplier_pp1_22 [10]),
    .ZN(u_multiplier_STAGE2_acci_pp2_22_1__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_22_1__22_  (.A(u_multiplier_pp1_22 [9]),
    .B(u_multiplier_pp1_22 [8]),
    .Z(u_multiplier_STAGE2_acci_pp2_22_1__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_22_1__23_  (.A(u_multiplier_pp1_22 [10]),
    .B(u_multiplier_pp1_22 [11]),
    .Z(u_multiplier_STAGE2_acci_pp2_22_1__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_22_1__24_  (.A1(u_multiplier_STAGE2_acci_pp2_22_1__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_22_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_22_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_22_1__25_  (.A(u_multiplier_STAGE2_acci_pp2_22_1__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_22_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_22_1__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_22_1__26_  (.A1(u_multiplier_STAGE2_acci_pp2_22_1__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_22_1__16_ ),
    .ZN(u_multiplier_pp2_22 [1]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_22_1__27_  (.A1(u_multiplier_pp1_22 [9]),
    .A2(u_multiplier_pp1_22 [8]),
    .B1(u_multiplier_pp1_22 [10]),
    .B2(u_multiplier_pp1_22 [11]),
    .ZN(u_multiplier_STAGE2_acci_pp2_22_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_22_1__28_  (.A1(u_multiplier_STAGE2_acci_pp2_22_1__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_22_1__17_ ),
    .ZN(u_multiplier_pp2_23 [6]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_22_2__21_  (.A1(u_multiplier_pp1_22 [5]),
    .A2(u_multiplier_pp1_22 [4]),
    .A3(u_multiplier_pp1_22 [6]),
    .ZN(u_multiplier_STAGE2_acci_pp2_22_2__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_22_2__22_  (.A(u_multiplier_pp1_22 [5]),
    .B(u_multiplier_pp1_22 [4]),
    .Z(u_multiplier_STAGE2_acci_pp2_22_2__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_22_2__23_  (.A(u_multiplier_pp1_22 [6]),
    .B(u_multiplier_pp1_22 [7]),
    .Z(u_multiplier_STAGE2_acci_pp2_22_2__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_22_2__24_  (.A1(u_multiplier_STAGE2_acci_pp2_22_2__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_22_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_22_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_22_2__25_  (.A(u_multiplier_STAGE2_acci_pp2_22_2__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_22_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_22_2__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_22_2__26_  (.A1(u_multiplier_STAGE2_acci_pp2_22_2__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_22_2__16_ ),
    .ZN(u_multiplier_pp2_22 [2]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_22_2__27_  (.A1(u_multiplier_pp1_22 [5]),
    .A2(u_multiplier_pp1_22 [4]),
    .B1(u_multiplier_pp1_22 [6]),
    .B2(u_multiplier_pp1_22 [7]),
    .ZN(u_multiplier_STAGE2_acci_pp2_22_2__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_22_2__28_  (.A1(u_multiplier_STAGE2_acci_pp2_22_2__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_22_2__17_ ),
    .ZN(u_multiplier_pp2_23 [5]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_22_3__21_  (.A1(u_multiplier_pp1_22 [1]),
    .A2(u_multiplier_pp1_22 [0]),
    .A3(u_multiplier_pp1_22 [2]),
    .ZN(u_multiplier_STAGE2_acci_pp2_22_3__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_22_3__22_  (.A(u_multiplier_pp1_22 [1]),
    .B(u_multiplier_pp1_22 [0]),
    .Z(u_multiplier_STAGE2_acci_pp2_22_3__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_22_3__23_  (.A(u_multiplier_pp1_22 [2]),
    .B(u_multiplier_pp1_22 [3]),
    .Z(u_multiplier_STAGE2_acci_pp2_22_3__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_22_3__24_  (.A1(u_multiplier_STAGE2_acci_pp2_22_3__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_22_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_22_3__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_22_3__25_  (.A(u_multiplier_STAGE2_acci_pp2_22_3__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_22_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_22_3__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_22_3__26_  (.A1(u_multiplier_STAGE2_acci_pp2_22_3__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_22_3__16_ ),
    .ZN(u_multiplier_pp2_22 [3]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_22_3__27_  (.A1(u_multiplier_pp1_22 [1]),
    .A2(u_multiplier_pp1_22 [0]),
    .B1(u_multiplier_pp1_22 [2]),
    .B2(u_multiplier_pp1_22 [3]),
    .ZN(u_multiplier_STAGE2_acci_pp2_22_3__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_22_3__28_  (.A1(u_multiplier_STAGE2_acci_pp2_22_3__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_22_3__17_ ),
    .ZN(u_multiplier_pp2_23 [4]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_23_0__21_  (.A1(u_multiplier_pp1_23 [13]),
    .A2(u_multiplier_pp1_23 [12]),
    .A3(u_multiplier_pp1_23 [14]),
    .ZN(u_multiplier_STAGE2_acci_pp2_23_0__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_23_0__22_  (.A(u_multiplier_pp1_23 [13]),
    .B(u_multiplier_pp1_23 [12]),
    .Z(u_multiplier_STAGE2_acci_pp2_23_0__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_23_0__23_  (.A(u_multiplier_pp1_23 [14]),
    .B(u_multiplier_pp1_23 [15]),
    .Z(u_multiplier_STAGE2_acci_pp2_23_0__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_23_0__24_  (.A1(u_multiplier_STAGE2_acci_pp2_23_0__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_23_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_23_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_23_0__25_  (.A(u_multiplier_STAGE2_acci_pp2_23_0__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_23_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_23_0__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_23_0__26_  (.A1(u_multiplier_STAGE2_acci_pp2_23_0__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_23_0__16_ ),
    .ZN(u_multiplier_pp2_23 [0]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_23_0__27_  (.A1(u_multiplier_pp1_23 [13]),
    .A2(u_multiplier_pp1_23 [12]),
    .B1(u_multiplier_pp1_23 [14]),
    .B2(u_multiplier_pp1_23 [15]),
    .ZN(u_multiplier_STAGE2_acci_pp2_23_0__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_23_0__28_  (.A1(u_multiplier_STAGE2_acci_pp2_23_0__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_23_0__17_ ),
    .ZN(u_multiplier_pp2_24 [7]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_23_1__21_  (.A1(u_multiplier_pp1_23 [9]),
    .A2(u_multiplier_pp1_23 [8]),
    .A3(u_multiplier_pp1_23 [10]),
    .ZN(u_multiplier_STAGE2_acci_pp2_23_1__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_23_1__22_  (.A(u_multiplier_pp1_23 [9]),
    .B(u_multiplier_pp1_23 [8]),
    .Z(u_multiplier_STAGE2_acci_pp2_23_1__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_23_1__23_  (.A(u_multiplier_pp1_23 [10]),
    .B(u_multiplier_pp1_23 [11]),
    .Z(u_multiplier_STAGE2_acci_pp2_23_1__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_23_1__24_  (.A1(u_multiplier_STAGE2_acci_pp2_23_1__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_23_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_23_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_23_1__25_  (.A(u_multiplier_STAGE2_acci_pp2_23_1__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_23_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_23_1__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_23_1__26_  (.A1(u_multiplier_STAGE2_acci_pp2_23_1__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_23_1__16_ ),
    .ZN(u_multiplier_pp2_23 [1]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_23_1__27_  (.A1(u_multiplier_pp1_23 [9]),
    .A2(u_multiplier_pp1_23 [8]),
    .B1(u_multiplier_pp1_23 [10]),
    .B2(u_multiplier_pp1_23 [11]),
    .ZN(u_multiplier_STAGE2_acci_pp2_23_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_23_1__28_  (.A1(u_multiplier_STAGE2_acci_pp2_23_1__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_23_1__17_ ),
    .ZN(u_multiplier_pp2_24 [6]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_23_2__21_  (.A1(u_multiplier_pp1_23 [5]),
    .A2(u_multiplier_pp1_23 [4]),
    .A3(u_multiplier_pp1_23 [6]),
    .ZN(u_multiplier_STAGE2_acci_pp2_23_2__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_23_2__22_  (.A(u_multiplier_pp1_23 [5]),
    .B(u_multiplier_pp1_23 [4]),
    .Z(u_multiplier_STAGE2_acci_pp2_23_2__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_23_2__23_  (.A(u_multiplier_pp1_23 [6]),
    .B(u_multiplier_pp1_23 [7]),
    .Z(u_multiplier_STAGE2_acci_pp2_23_2__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_23_2__24_  (.A1(u_multiplier_STAGE2_acci_pp2_23_2__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_23_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_23_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_23_2__25_  (.A(u_multiplier_STAGE2_acci_pp2_23_2__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_23_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_23_2__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_23_2__26_  (.A1(u_multiplier_STAGE2_acci_pp2_23_2__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_23_2__16_ ),
    .ZN(u_multiplier_pp2_23 [2]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_23_2__27_  (.A1(u_multiplier_pp1_23 [5]),
    .A2(u_multiplier_pp1_23 [4]),
    .B1(u_multiplier_pp1_23 [6]),
    .B2(u_multiplier_pp1_23 [7]),
    .ZN(u_multiplier_STAGE2_acci_pp2_23_2__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_23_2__28_  (.A1(u_multiplier_STAGE2_acci_pp2_23_2__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_23_2__17_ ),
    .ZN(u_multiplier_pp2_24 [5]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_23_3__21_  (.A1(u_multiplier_pp1_23 [1]),
    .A2(u_multiplier_pp1_23 [0]),
    .A3(u_multiplier_pp1_23 [2]),
    .ZN(u_multiplier_STAGE2_acci_pp2_23_3__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_23_3__22_  (.A(u_multiplier_pp1_23 [1]),
    .B(u_multiplier_pp1_23 [0]),
    .Z(u_multiplier_STAGE2_acci_pp2_23_3__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_23_3__23_  (.A(u_multiplier_pp1_23 [2]),
    .B(u_multiplier_pp1_23 [3]),
    .Z(u_multiplier_STAGE2_acci_pp2_23_3__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_23_3__24_  (.A1(u_multiplier_STAGE2_acci_pp2_23_3__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_23_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_23_3__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_23_3__25_  (.A(u_multiplier_STAGE2_acci_pp2_23_3__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_23_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_23_3__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_23_3__26_  (.A1(u_multiplier_STAGE2_acci_pp2_23_3__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_23_3__16_ ),
    .ZN(u_multiplier_pp2_23 [3]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_23_3__27_  (.A1(u_multiplier_pp1_23 [1]),
    .A2(u_multiplier_pp1_23 [0]),
    .B1(u_multiplier_pp1_23 [2]),
    .B2(u_multiplier_pp1_23 [3]),
    .ZN(u_multiplier_STAGE2_acci_pp2_23_3__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_23_3__28_  (.A1(u_multiplier_STAGE2_acci_pp2_23_3__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_23_3__17_ ),
    .ZN(u_multiplier_pp2_24 [4]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_24_0__21_  (.A1(u_multiplier_pp1_24 [13]),
    .A2(u_multiplier_pp1_24 [12]),
    .A3(u_multiplier_pp1_24 [14]),
    .ZN(u_multiplier_STAGE2_acci_pp2_24_0__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_24_0__22_  (.A(u_multiplier_pp1_24 [13]),
    .B(u_multiplier_pp1_24 [12]),
    .Z(u_multiplier_STAGE2_acci_pp2_24_0__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_24_0__23_  (.A(u_multiplier_pp1_24 [14]),
    .B(u_multiplier_pp1_24 [15]),
    .Z(u_multiplier_STAGE2_acci_pp2_24_0__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_24_0__24_  (.A1(u_multiplier_STAGE2_acci_pp2_24_0__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_24_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_24_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_24_0__25_  (.A(u_multiplier_STAGE2_acci_pp2_24_0__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_24_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_24_0__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_24_0__26_  (.A1(u_multiplier_STAGE2_acci_pp2_24_0__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_24_0__16_ ),
    .ZN(u_multiplier_pp2_24 [0]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_24_0__27_  (.A1(u_multiplier_pp1_24 [13]),
    .A2(u_multiplier_pp1_24 [12]),
    .B1(u_multiplier_pp1_24 [14]),
    .B2(u_multiplier_pp1_24 [15]),
    .ZN(u_multiplier_STAGE2_acci_pp2_24_0__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_24_0__28_  (.A1(u_multiplier_STAGE2_acci_pp2_24_0__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_24_0__17_ ),
    .ZN(u_multiplier_pp2_25 [7]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_24_1__21_  (.A1(u_multiplier_pp1_24 [9]),
    .A2(u_multiplier_pp1_24 [8]),
    .A3(u_multiplier_pp1_24 [10]),
    .ZN(u_multiplier_STAGE2_acci_pp2_24_1__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_24_1__22_  (.A(u_multiplier_pp1_24 [9]),
    .B(u_multiplier_pp1_24 [8]),
    .Z(u_multiplier_STAGE2_acci_pp2_24_1__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_24_1__23_  (.A(u_multiplier_pp1_24 [10]),
    .B(u_multiplier_pp1_24 [11]),
    .Z(u_multiplier_STAGE2_acci_pp2_24_1__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_24_1__24_  (.A1(u_multiplier_STAGE2_acci_pp2_24_1__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_24_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_24_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_24_1__25_  (.A(u_multiplier_STAGE2_acci_pp2_24_1__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_24_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_24_1__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_24_1__26_  (.A1(u_multiplier_STAGE2_acci_pp2_24_1__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_24_1__16_ ),
    .ZN(u_multiplier_pp2_24 [1]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_24_1__27_  (.A1(u_multiplier_pp1_24 [9]),
    .A2(u_multiplier_pp1_24 [8]),
    .B1(u_multiplier_pp1_24 [10]),
    .B2(u_multiplier_pp1_24 [11]),
    .ZN(u_multiplier_STAGE2_acci_pp2_24_1__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_24_1__28_  (.A1(u_multiplier_STAGE2_acci_pp2_24_1__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_24_1__17_ ),
    .ZN(u_multiplier_pp2_25 [6]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_24_2__21_  (.A1(u_multiplier_pp1_24 [5]),
    .A2(u_multiplier_pp1_24 [4]),
    .A3(u_multiplier_pp1_24 [6]),
    .ZN(u_multiplier_STAGE2_acci_pp2_24_2__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_24_2__22_  (.A(u_multiplier_pp1_24 [5]),
    .B(u_multiplier_pp1_24 [4]),
    .Z(u_multiplier_STAGE2_acci_pp2_24_2__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_24_2__23_  (.A(u_multiplier_pp1_24 [6]),
    .B(u_multiplier_pp1_24 [7]),
    .Z(u_multiplier_STAGE2_acci_pp2_24_2__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_24_2__24_  (.A1(u_multiplier_STAGE2_acci_pp2_24_2__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_24_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_24_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_24_2__25_  (.A(u_multiplier_STAGE2_acci_pp2_24_2__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_24_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_24_2__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_24_2__26_  (.A1(u_multiplier_STAGE2_acci_pp2_24_2__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_24_2__16_ ),
    .ZN(u_multiplier_pp2_24 [2]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_24_2__27_  (.A1(u_multiplier_pp1_24 [5]),
    .A2(u_multiplier_pp1_24 [4]),
    .B1(u_multiplier_pp1_24 [6]),
    .B2(u_multiplier_pp1_24 [7]),
    .ZN(u_multiplier_STAGE2_acci_pp2_24_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_24_2__28_  (.A1(u_multiplier_STAGE2_acci_pp2_24_2__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_24_2__17_ ),
    .ZN(u_multiplier_pp2_25 [5]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_24_3__21_  (.A1(u_multiplier_pp1_24 [1]),
    .A2(u_multiplier_pp1_24 [0]),
    .A3(u_multiplier_pp1_24 [2]),
    .ZN(u_multiplier_STAGE2_acci_pp2_24_3__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_24_3__22_  (.A(u_multiplier_pp1_24 [1]),
    .B(u_multiplier_pp1_24 [0]),
    .Z(u_multiplier_STAGE2_acci_pp2_24_3__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_24_3__23_  (.A(u_multiplier_pp1_24 [2]),
    .B(u_multiplier_pp1_24 [3]),
    .Z(u_multiplier_STAGE2_acci_pp2_24_3__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_24_3__24_  (.A1(u_multiplier_STAGE2_acci_pp2_24_3__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_24_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_24_3__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_24_3__25_  (.A(u_multiplier_STAGE2_acci_pp2_24_3__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_24_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_24_3__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_24_3__26_  (.A1(u_multiplier_STAGE2_acci_pp2_24_3__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_24_3__16_ ),
    .ZN(u_multiplier_pp2_24 [3]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_24_3__27_  (.A1(u_multiplier_pp1_24 [1]),
    .A2(u_multiplier_pp1_24 [0]),
    .B1(u_multiplier_pp1_24 [2]),
    .B2(u_multiplier_pp1_24 [3]),
    .ZN(u_multiplier_STAGE2_acci_pp2_24_3__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_24_3__28_  (.A1(u_multiplier_STAGE2_acci_pp2_24_3__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_24_3__17_ ),
    .ZN(u_multiplier_pp2_25 [4]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_25_0__21_  (.A1(u_multiplier_pp1_25 [13]),
    .A2(u_multiplier_pp1_25 [12]),
    .A3(u_multiplier_pp1_25 [14]),
    .ZN(u_multiplier_STAGE2_acci_pp2_25_0__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_25_0__22_  (.A(u_multiplier_pp1_25 [13]),
    .B(u_multiplier_pp1_25 [12]),
    .Z(u_multiplier_STAGE2_acci_pp2_25_0__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_25_0__23_  (.A(u_multiplier_pp1_25 [14]),
    .B(u_multiplier_pp1_25 [15]),
    .Z(u_multiplier_STAGE2_acci_pp2_25_0__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_25_0__24_  (.A1(u_multiplier_STAGE2_acci_pp2_25_0__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_25_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_25_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_25_0__25_  (.A(u_multiplier_STAGE2_acci_pp2_25_0__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_25_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_25_0__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_25_0__26_  (.A1(u_multiplier_STAGE2_acci_pp2_25_0__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_25_0__16_ ),
    .ZN(u_multiplier_pp2_25 [0]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_25_0__27_  (.A1(u_multiplier_pp1_25 [13]),
    .A2(u_multiplier_pp1_25 [12]),
    .B1(u_multiplier_pp1_25 [14]),
    .B2(u_multiplier_pp1_25 [15]),
    .ZN(u_multiplier_STAGE2_acci_pp2_25_0__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_25_0__28_  (.A1(u_multiplier_STAGE2_acci_pp2_25_0__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_25_0__17_ ),
    .ZN(u_multiplier_pp2_26 [7]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_25_1__21_  (.A1(u_multiplier_pp1_25 [9]),
    .A2(u_multiplier_pp1_25 [8]),
    .A3(u_multiplier_pp1_25 [10]),
    .ZN(u_multiplier_STAGE2_acci_pp2_25_1__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_25_1__22_  (.A(u_multiplier_pp1_25 [9]),
    .B(u_multiplier_pp1_25 [8]),
    .Z(u_multiplier_STAGE2_acci_pp2_25_1__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_25_1__23_  (.A(u_multiplier_pp1_25 [10]),
    .B(u_multiplier_pp1_25 [11]),
    .Z(u_multiplier_STAGE2_acci_pp2_25_1__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_25_1__24_  (.A1(u_multiplier_STAGE2_acci_pp2_25_1__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_25_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_25_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_25_1__25_  (.A(u_multiplier_STAGE2_acci_pp2_25_1__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_25_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_25_1__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_25_1__26_  (.A1(u_multiplier_STAGE2_acci_pp2_25_1__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_25_1__16_ ),
    .ZN(u_multiplier_pp2_25 [1]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_25_1__27_  (.A1(u_multiplier_pp1_25 [9]),
    .A2(u_multiplier_pp1_25 [8]),
    .B1(u_multiplier_pp1_25 [10]),
    .B2(u_multiplier_pp1_25 [11]),
    .ZN(u_multiplier_STAGE2_acci_pp2_25_1__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_25_1__28_  (.A1(u_multiplier_STAGE2_acci_pp2_25_1__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_25_1__17_ ),
    .ZN(u_multiplier_pp2_26 [6]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_25_2__21_  (.A1(u_multiplier_pp1_25 [5]),
    .A2(u_multiplier_pp1_25 [4]),
    .A3(u_multiplier_pp1_25 [6]),
    .ZN(u_multiplier_STAGE2_acci_pp2_25_2__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_25_2__22_  (.A(u_multiplier_pp1_25 [5]),
    .B(u_multiplier_pp1_25 [4]),
    .Z(u_multiplier_STAGE2_acci_pp2_25_2__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_25_2__23_  (.A(u_multiplier_pp1_25 [6]),
    .B(u_multiplier_pp1_25 [7]),
    .Z(u_multiplier_STAGE2_acci_pp2_25_2__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_25_2__24_  (.A1(u_multiplier_STAGE2_acci_pp2_25_2__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_25_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_25_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_25_2__25_  (.A(u_multiplier_STAGE2_acci_pp2_25_2__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_25_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_25_2__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_25_2__26_  (.A1(u_multiplier_STAGE2_acci_pp2_25_2__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_25_2__16_ ),
    .ZN(u_multiplier_pp2_25 [2]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_25_2__27_  (.A1(u_multiplier_pp1_25 [5]),
    .A2(u_multiplier_pp1_25 [4]),
    .B1(u_multiplier_pp1_25 [6]),
    .B2(u_multiplier_pp1_25 [7]),
    .ZN(u_multiplier_STAGE2_acci_pp2_25_2__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_25_2__28_  (.A1(u_multiplier_STAGE2_acci_pp2_25_2__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_25_2__17_ ),
    .ZN(u_multiplier_pp2_26 [5]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_25_3__21_  (.A1(u_multiplier_pp1_25 [1]),
    .A2(u_multiplier_pp1_25 [0]),
    .A3(u_multiplier_pp1_25 [2]),
    .ZN(u_multiplier_STAGE2_acci_pp2_25_3__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_25_3__22_  (.A(u_multiplier_pp1_25 [1]),
    .B(u_multiplier_pp1_25 [0]),
    .Z(u_multiplier_STAGE2_acci_pp2_25_3__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_25_3__23_  (.A(u_multiplier_pp1_25 [2]),
    .B(u_multiplier_pp1_25 [3]),
    .Z(u_multiplier_STAGE2_acci_pp2_25_3__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_25_3__24_  (.A1(u_multiplier_STAGE2_acci_pp2_25_3__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_25_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_25_3__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_25_3__25_  (.A(u_multiplier_STAGE2_acci_pp2_25_3__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_25_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_25_3__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_25_3__26_  (.A1(u_multiplier_STAGE2_acci_pp2_25_3__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_25_3__16_ ),
    .ZN(u_multiplier_pp2_25 [3]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_25_3__27_  (.A1(u_multiplier_pp1_25 [1]),
    .A2(u_multiplier_pp1_25 [0]),
    .B1(u_multiplier_pp1_25 [2]),
    .B2(u_multiplier_pp1_25 [3]),
    .ZN(u_multiplier_STAGE2_acci_pp2_25_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_25_3__28_  (.A1(u_multiplier_STAGE2_acci_pp2_25_3__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_25_3__17_ ),
    .ZN(u_multiplier_pp2_26 [4]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_26_0__21_  (.A1(u_multiplier_pp1_26 [13]),
    .A2(u_multiplier_pp1_26 [12]),
    .A3(u_multiplier_pp1_26 [14]),
    .ZN(u_multiplier_STAGE2_acci_pp2_26_0__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_26_0__22_  (.A(u_multiplier_pp1_26 [13]),
    .B(u_multiplier_pp1_26 [12]),
    .Z(u_multiplier_STAGE2_acci_pp2_26_0__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_26_0__23_  (.A(u_multiplier_pp1_26 [14]),
    .B(u_multiplier_pp1_26 [15]),
    .Z(u_multiplier_STAGE2_acci_pp2_26_0__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_26_0__24_  (.A1(u_multiplier_STAGE2_acci_pp2_26_0__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_26_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_26_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_26_0__25_  (.A(u_multiplier_STAGE2_acci_pp2_26_0__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_26_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_26_0__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_26_0__26_  (.A1(u_multiplier_STAGE2_acci_pp2_26_0__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_26_0__16_ ),
    .ZN(u_multiplier_pp2_26 [0]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_26_0__27_  (.A1(u_multiplier_pp1_26 [13]),
    .A2(u_multiplier_pp1_26 [12]),
    .B1(u_multiplier_pp1_26 [14]),
    .B2(u_multiplier_pp1_26 [15]),
    .ZN(u_multiplier_STAGE2_acci_pp2_26_0__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_26_0__28_  (.A1(u_multiplier_STAGE2_acci_pp2_26_0__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_26_0__17_ ),
    .ZN(u_multiplier_pp2_27 [7]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_26_1__21_  (.A1(u_multiplier_pp1_26 [9]),
    .A2(u_multiplier_pp1_26 [8]),
    .A3(u_multiplier_pp1_26 [10]),
    .ZN(u_multiplier_STAGE2_acci_pp2_26_1__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_26_1__22_  (.A(u_multiplier_pp1_26 [9]),
    .B(u_multiplier_pp1_26 [8]),
    .Z(u_multiplier_STAGE2_acci_pp2_26_1__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_26_1__23_  (.A(u_multiplier_pp1_26 [10]),
    .B(u_multiplier_pp1_26 [11]),
    .Z(u_multiplier_STAGE2_acci_pp2_26_1__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_26_1__24_  (.A1(u_multiplier_STAGE2_acci_pp2_26_1__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_26_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_26_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_26_1__25_  (.A(u_multiplier_STAGE2_acci_pp2_26_1__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_26_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_26_1__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_26_1__26_  (.A1(u_multiplier_STAGE2_acci_pp2_26_1__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_26_1__16_ ),
    .ZN(u_multiplier_pp2_26 [1]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_26_1__27_  (.A1(u_multiplier_pp1_26 [9]),
    .A2(u_multiplier_pp1_26 [8]),
    .B1(u_multiplier_pp1_26 [10]),
    .B2(u_multiplier_pp1_26 [11]),
    .ZN(u_multiplier_STAGE2_acci_pp2_26_1__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_26_1__28_  (.A1(u_multiplier_STAGE2_acci_pp2_26_1__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_26_1__17_ ),
    .ZN(u_multiplier_pp2_27 [6]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_26_2__21_  (.A1(u_multiplier_pp1_26 [5]),
    .A2(u_multiplier_pp1_26 [4]),
    .A3(u_multiplier_pp1_26 [6]),
    .ZN(u_multiplier_STAGE2_acci_pp2_26_2__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_26_2__22_  (.A(u_multiplier_pp1_26 [5]),
    .B(u_multiplier_pp1_26 [4]),
    .Z(u_multiplier_STAGE2_acci_pp2_26_2__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_26_2__23_  (.A(u_multiplier_pp1_26 [6]),
    .B(u_multiplier_pp1_26 [7]),
    .Z(u_multiplier_STAGE2_acci_pp2_26_2__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_26_2__24_  (.A1(u_multiplier_STAGE2_acci_pp2_26_2__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_26_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_26_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_26_2__25_  (.A(u_multiplier_STAGE2_acci_pp2_26_2__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_26_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_26_2__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_26_2__26_  (.A1(u_multiplier_STAGE2_acci_pp2_26_2__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_26_2__16_ ),
    .ZN(u_multiplier_pp2_26 [2]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_26_2__27_  (.A1(u_multiplier_pp1_26 [5]),
    .A2(u_multiplier_pp1_26 [4]),
    .B1(u_multiplier_pp1_26 [6]),
    .B2(u_multiplier_pp1_26 [7]),
    .ZN(u_multiplier_STAGE2_acci_pp2_26_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_26_2__28_  (.A1(u_multiplier_STAGE2_acci_pp2_26_2__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_26_2__17_ ),
    .ZN(u_multiplier_pp2_27 [5]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_26_3__21_  (.A1(u_multiplier_pp1_26 [1]),
    .A2(u_multiplier_pp1_26 [0]),
    .A3(u_multiplier_pp1_26 [2]),
    .ZN(u_multiplier_STAGE2_acci_pp2_26_3__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_26_3__22_  (.A(u_multiplier_pp1_26 [1]),
    .B(u_multiplier_pp1_26 [0]),
    .Z(u_multiplier_STAGE2_acci_pp2_26_3__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_26_3__23_  (.A(u_multiplier_pp1_26 [2]),
    .B(u_multiplier_pp1_26 [3]),
    .Z(u_multiplier_STAGE2_acci_pp2_26_3__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_26_3__24_  (.A1(u_multiplier_STAGE2_acci_pp2_26_3__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_26_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_26_3__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_26_3__25_  (.A(u_multiplier_STAGE2_acci_pp2_26_3__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_26_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_26_3__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_26_3__26_  (.A1(u_multiplier_STAGE2_acci_pp2_26_3__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_26_3__16_ ),
    .ZN(u_multiplier_pp2_26 [3]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_26_3__27_  (.A1(u_multiplier_pp1_26 [1]),
    .A2(u_multiplier_pp1_26 [0]),
    .B1(u_multiplier_pp1_26 [2]),
    .B2(u_multiplier_pp1_26 [3]),
    .ZN(u_multiplier_STAGE2_acci_pp2_26_3__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_26_3__28_  (.A1(u_multiplier_STAGE2_acci_pp2_26_3__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_26_3__17_ ),
    .ZN(u_multiplier_pp2_27 [4]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_27_0__21_  (.A1(u_multiplier_pp1_27 [13]),
    .A2(u_multiplier_pp1_27 [12]),
    .A3(u_multiplier_pp1_27 [14]),
    .ZN(u_multiplier_STAGE2_acci_pp2_27_0__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_27_0__22_  (.A(u_multiplier_pp1_27 [13]),
    .B(u_multiplier_pp1_27 [12]),
    .Z(u_multiplier_STAGE2_acci_pp2_27_0__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_27_0__23_  (.A(u_multiplier_pp1_27 [14]),
    .B(u_multiplier_pp1_27 [15]),
    .Z(u_multiplier_STAGE2_acci_pp2_27_0__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_27_0__24_  (.A1(u_multiplier_STAGE2_acci_pp2_27_0__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_27_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_27_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_27_0__25_  (.A(u_multiplier_STAGE2_acci_pp2_27_0__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_27_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_27_0__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_27_0__26_  (.A1(u_multiplier_STAGE2_acci_pp2_27_0__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_27_0__16_ ),
    .ZN(u_multiplier_pp2_27 [0]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_27_0__27_  (.A1(u_multiplier_pp1_27 [13]),
    .A2(u_multiplier_pp1_27 [12]),
    .B1(u_multiplier_pp1_27 [14]),
    .B2(u_multiplier_pp1_27 [15]),
    .ZN(u_multiplier_STAGE2_acci_pp2_27_0__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_27_0__28_  (.A1(u_multiplier_STAGE2_acci_pp2_27_0__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_27_0__17_ ),
    .ZN(u_multiplier_pp2_28 [7]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_27_1__21_  (.A1(u_multiplier_pp1_27 [9]),
    .A2(u_multiplier_pp1_27 [8]),
    .A3(u_multiplier_pp1_27 [10]),
    .ZN(u_multiplier_STAGE2_acci_pp2_27_1__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_27_1__22_  (.A(u_multiplier_pp1_27 [9]),
    .B(u_multiplier_pp1_27 [8]),
    .Z(u_multiplier_STAGE2_acci_pp2_27_1__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_27_1__23_  (.A(u_multiplier_pp1_27 [10]),
    .B(u_multiplier_pp1_27 [11]),
    .Z(u_multiplier_STAGE2_acci_pp2_27_1__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_27_1__24_  (.A1(u_multiplier_STAGE2_acci_pp2_27_1__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_27_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_27_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_27_1__25_  (.A(u_multiplier_STAGE2_acci_pp2_27_1__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_27_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_27_1__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_27_1__26_  (.A1(u_multiplier_STAGE2_acci_pp2_27_1__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_27_1__16_ ),
    .ZN(u_multiplier_pp2_27 [1]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_27_1__27_  (.A1(u_multiplier_pp1_27 [9]),
    .A2(u_multiplier_pp1_27 [8]),
    .B1(u_multiplier_pp1_27 [10]),
    .B2(u_multiplier_pp1_27 [11]),
    .ZN(u_multiplier_STAGE2_acci_pp2_27_1__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_27_1__28_  (.A1(u_multiplier_STAGE2_acci_pp2_27_1__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_27_1__17_ ),
    .ZN(u_multiplier_pp2_28 [6]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_27_2__21_  (.A1(u_multiplier_pp1_27 [5]),
    .A2(u_multiplier_pp1_27 [4]),
    .A3(u_multiplier_pp1_27 [6]),
    .ZN(u_multiplier_STAGE2_acci_pp2_27_2__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_27_2__22_  (.A(u_multiplier_pp1_27 [5]),
    .B(u_multiplier_pp1_27 [4]),
    .Z(u_multiplier_STAGE2_acci_pp2_27_2__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_27_2__23_  (.A(u_multiplier_pp1_27 [6]),
    .B(u_multiplier_pp1_27 [7]),
    .Z(u_multiplier_STAGE2_acci_pp2_27_2__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_27_2__24_  (.A1(u_multiplier_STAGE2_acci_pp2_27_2__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_27_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_27_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_27_2__25_  (.A(u_multiplier_STAGE2_acci_pp2_27_2__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_27_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_27_2__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_27_2__26_  (.A1(u_multiplier_STAGE2_acci_pp2_27_2__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_27_2__16_ ),
    .ZN(u_multiplier_pp2_27 [2]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_27_2__27_  (.A1(u_multiplier_pp1_27 [5]),
    .A2(u_multiplier_pp1_27 [4]),
    .B1(u_multiplier_pp1_27 [6]),
    .B2(u_multiplier_pp1_27 [7]),
    .ZN(u_multiplier_STAGE2_acci_pp2_27_2__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_27_2__28_  (.A1(u_multiplier_STAGE2_acci_pp2_27_2__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_27_2__17_ ),
    .ZN(u_multiplier_pp2_28 [5]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_27_3__21_  (.A1(u_multiplier_pp1_27 [1]),
    .A2(u_multiplier_pp1_27 [0]),
    .A3(u_multiplier_pp1_27 [2]),
    .ZN(u_multiplier_STAGE2_acci_pp2_27_3__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_27_3__22_  (.A(u_multiplier_pp1_27 [1]),
    .B(u_multiplier_pp1_27 [0]),
    .Z(u_multiplier_STAGE2_acci_pp2_27_3__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_27_3__23_  (.A(u_multiplier_pp1_27 [2]),
    .B(u_multiplier_pp1_27 [3]),
    .Z(u_multiplier_STAGE2_acci_pp2_27_3__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_27_3__24_  (.A1(u_multiplier_STAGE2_acci_pp2_27_3__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_27_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_27_3__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_27_3__25_  (.A(u_multiplier_STAGE2_acci_pp2_27_3__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_27_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_27_3__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_27_3__26_  (.A1(u_multiplier_STAGE2_acci_pp2_27_3__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_27_3__16_ ),
    .ZN(u_multiplier_pp2_27 [3]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_27_3__27_  (.A1(u_multiplier_pp1_27 [1]),
    .A2(u_multiplier_pp1_27 [0]),
    .B1(u_multiplier_pp1_27 [2]),
    .B2(u_multiplier_pp1_27 [3]),
    .ZN(u_multiplier_STAGE2_acci_pp2_27_3__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_27_3__28_  (.A1(u_multiplier_STAGE2_acci_pp2_27_3__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_27_3__17_ ),
    .ZN(u_multiplier_pp2_28 [4]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_28_0__21_  (.A1(u_multiplier_pp1_28 [13]),
    .A2(u_multiplier_pp1_28 [12]),
    .A3(u_multiplier_pp1_28 [14]),
    .ZN(u_multiplier_STAGE2_acci_pp2_28_0__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_28_0__22_  (.A(u_multiplier_pp1_28 [13]),
    .B(u_multiplier_pp1_28 [12]),
    .Z(u_multiplier_STAGE2_acci_pp2_28_0__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_28_0__23_  (.A(u_multiplier_pp1_28 [14]),
    .B(u_multiplier_pp1_28 [15]),
    .Z(u_multiplier_STAGE2_acci_pp2_28_0__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_28_0__24_  (.A1(u_multiplier_STAGE2_acci_pp2_28_0__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_28_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_28_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_28_0__25_  (.A(u_multiplier_STAGE2_acci_pp2_28_0__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_28_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_28_0__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_28_0__26_  (.A1(u_multiplier_STAGE2_acci_pp2_28_0__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_28_0__16_ ),
    .ZN(u_multiplier_pp2_28 [0]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_28_0__27_  (.A1(u_multiplier_pp1_28 [13]),
    .A2(u_multiplier_pp1_28 [12]),
    .B1(u_multiplier_pp1_28 [14]),
    .B2(u_multiplier_pp1_28 [15]),
    .ZN(u_multiplier_STAGE2_acci_pp2_28_0__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_28_0__28_  (.A1(u_multiplier_STAGE2_acci_pp2_28_0__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_28_0__17_ ),
    .ZN(u_multiplier_pp2_29 [7]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_28_1__21_  (.A1(u_multiplier_pp1_28 [9]),
    .A2(u_multiplier_pp1_28 [8]),
    .A3(u_multiplier_pp1_28 [10]),
    .ZN(u_multiplier_STAGE2_acci_pp2_28_1__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_28_1__22_  (.A(u_multiplier_pp1_28 [9]),
    .B(u_multiplier_pp1_28 [8]),
    .Z(u_multiplier_STAGE2_acci_pp2_28_1__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_28_1__23_  (.A(u_multiplier_pp1_28 [10]),
    .B(u_multiplier_pp1_28 [11]),
    .Z(u_multiplier_STAGE2_acci_pp2_28_1__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_28_1__24_  (.A1(u_multiplier_STAGE2_acci_pp2_28_1__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_28_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_28_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_28_1__25_  (.A(u_multiplier_STAGE2_acci_pp2_28_1__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_28_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_28_1__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_28_1__26_  (.A1(u_multiplier_STAGE2_acci_pp2_28_1__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_28_1__16_ ),
    .ZN(u_multiplier_pp2_28 [1]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_28_1__27_  (.A1(u_multiplier_pp1_28 [9]),
    .A2(u_multiplier_pp1_28 [8]),
    .B1(u_multiplier_pp1_28 [10]),
    .B2(u_multiplier_pp1_28 [11]),
    .ZN(u_multiplier_STAGE2_acci_pp2_28_1__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_28_1__28_  (.A1(u_multiplier_STAGE2_acci_pp2_28_1__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_28_1__17_ ),
    .ZN(u_multiplier_pp2_29 [6]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_28_2__21_  (.A1(u_multiplier_pp1_28 [5]),
    .A2(u_multiplier_pp1_28 [4]),
    .A3(u_multiplier_pp1_28 [6]),
    .ZN(u_multiplier_STAGE2_acci_pp2_28_2__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_28_2__22_  (.A(u_multiplier_pp1_28 [5]),
    .B(u_multiplier_pp1_28 [4]),
    .Z(u_multiplier_STAGE2_acci_pp2_28_2__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_28_2__23_  (.A(u_multiplier_pp1_28 [6]),
    .B(u_multiplier_pp1_28 [7]),
    .Z(u_multiplier_STAGE2_acci_pp2_28_2__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_28_2__24_  (.A1(u_multiplier_STAGE2_acci_pp2_28_2__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_28_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_28_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_28_2__25_  (.A(u_multiplier_STAGE2_acci_pp2_28_2__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_28_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_28_2__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_28_2__26_  (.A1(u_multiplier_STAGE2_acci_pp2_28_2__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_28_2__16_ ),
    .ZN(u_multiplier_pp2_28 [2]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_28_2__27_  (.A1(u_multiplier_pp1_28 [5]),
    .A2(u_multiplier_pp1_28 [4]),
    .B1(u_multiplier_pp1_28 [6]),
    .B2(u_multiplier_pp1_28 [7]),
    .ZN(u_multiplier_STAGE2_acci_pp2_28_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_28_2__28_  (.A1(u_multiplier_STAGE2_acci_pp2_28_2__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_28_2__17_ ),
    .ZN(u_multiplier_pp2_29 [5]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_28_3__21_  (.A1(u_multiplier_pp1_28 [1]),
    .A2(u_multiplier_pp1_28 [0]),
    .A3(u_multiplier_pp1_28 [2]),
    .ZN(u_multiplier_STAGE2_acci_pp2_28_3__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_28_3__22_  (.A(u_multiplier_pp1_28 [1]),
    .B(u_multiplier_pp1_28 [0]),
    .Z(u_multiplier_STAGE2_acci_pp2_28_3__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_28_3__23_  (.A(u_multiplier_pp1_28 [2]),
    .B(u_multiplier_pp1_28 [3]),
    .Z(u_multiplier_STAGE2_acci_pp2_28_3__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_28_3__24_  (.A1(u_multiplier_STAGE2_acci_pp2_28_3__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_28_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_28_3__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_28_3__25_  (.A(u_multiplier_STAGE2_acci_pp2_28_3__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_28_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_28_3__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_28_3__26_  (.A1(u_multiplier_STAGE2_acci_pp2_28_3__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_28_3__16_ ),
    .ZN(u_multiplier_pp2_28 [3]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_28_3__27_  (.A1(u_multiplier_pp1_28 [1]),
    .A2(u_multiplier_pp1_28 [0]),
    .B1(u_multiplier_pp1_28 [2]),
    .B2(u_multiplier_pp1_28 [3]),
    .ZN(u_multiplier_STAGE2_acci_pp2_28_3__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_28_3__28_  (.A1(u_multiplier_STAGE2_acci_pp2_28_3__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_28_3__17_ ),
    .ZN(u_multiplier_pp2_29 [4]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_29_0__21_  (.A1(u_multiplier_pp1_29 [13]),
    .A2(u_multiplier_pp1_29 [12]),
    .A3(u_multiplier_pp1_29 [14]),
    .ZN(u_multiplier_STAGE2_acci_pp2_29_0__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_29_0__22_  (.A(u_multiplier_pp1_29 [13]),
    .B(u_multiplier_pp1_29 [12]),
    .Z(u_multiplier_STAGE2_acci_pp2_29_0__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_29_0__23_  (.A(u_multiplier_pp1_29 [14]),
    .B(u_multiplier_pp1_29 [15]),
    .Z(u_multiplier_STAGE2_acci_pp2_29_0__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_29_0__24_  (.A1(u_multiplier_STAGE2_acci_pp2_29_0__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_29_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_29_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_29_0__25_  (.A(u_multiplier_STAGE2_acci_pp2_29_0__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_29_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_29_0__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_29_0__26_  (.A1(u_multiplier_STAGE2_acci_pp2_29_0__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_29_0__16_ ),
    .ZN(u_multiplier_pp2_29 [0]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_29_0__27_  (.A1(u_multiplier_pp1_29 [13]),
    .A2(u_multiplier_pp1_29 [12]),
    .B1(u_multiplier_pp1_29 [14]),
    .B2(u_multiplier_pp1_29 [15]),
    .ZN(u_multiplier_STAGE2_acci_pp2_29_0__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_29_0__28_  (.A1(u_multiplier_STAGE2_acci_pp2_29_0__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_29_0__17_ ),
    .ZN(u_multiplier_pp2_30 [7]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_29_1__21_  (.A1(u_multiplier_pp1_29 [9]),
    .A2(u_multiplier_pp1_29 [8]),
    .A3(u_multiplier_pp1_29 [10]),
    .ZN(u_multiplier_STAGE2_acci_pp2_29_1__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_29_1__22_  (.A(u_multiplier_pp1_29 [9]),
    .B(u_multiplier_pp1_29 [8]),
    .Z(u_multiplier_STAGE2_acci_pp2_29_1__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_29_1__23_  (.A(u_multiplier_pp1_29 [10]),
    .B(u_multiplier_pp1_29 [11]),
    .Z(u_multiplier_STAGE2_acci_pp2_29_1__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_29_1__24_  (.A1(u_multiplier_STAGE2_acci_pp2_29_1__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_29_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_29_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_29_1__25_  (.A(u_multiplier_STAGE2_acci_pp2_29_1__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_29_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_29_1__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_29_1__26_  (.A1(u_multiplier_STAGE2_acci_pp2_29_1__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_29_1__16_ ),
    .ZN(u_multiplier_pp2_29 [1]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_29_1__27_  (.A1(u_multiplier_pp1_29 [9]),
    .A2(u_multiplier_pp1_29 [8]),
    .B1(u_multiplier_pp1_29 [10]),
    .B2(u_multiplier_pp1_29 [11]),
    .ZN(u_multiplier_STAGE2_acci_pp2_29_1__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_29_1__28_  (.A1(u_multiplier_STAGE2_acci_pp2_29_1__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_29_1__17_ ),
    .ZN(u_multiplier_pp2_30 [6]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_29_2__21_  (.A1(u_multiplier_pp1_29 [5]),
    .A2(u_multiplier_pp1_29 [4]),
    .A3(u_multiplier_pp1_29 [6]),
    .ZN(u_multiplier_STAGE2_acci_pp2_29_2__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_29_2__22_  (.A(u_multiplier_pp1_29 [5]),
    .B(u_multiplier_pp1_29 [4]),
    .Z(u_multiplier_STAGE2_acci_pp2_29_2__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_29_2__23_  (.A(u_multiplier_pp1_29 [6]),
    .B(u_multiplier_pp1_29 [7]),
    .Z(u_multiplier_STAGE2_acci_pp2_29_2__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_29_2__24_  (.A1(u_multiplier_STAGE2_acci_pp2_29_2__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_29_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_29_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_29_2__25_  (.A(u_multiplier_STAGE2_acci_pp2_29_2__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_29_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_29_2__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_29_2__26_  (.A1(u_multiplier_STAGE2_acci_pp2_29_2__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_29_2__16_ ),
    .ZN(u_multiplier_pp2_29 [2]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_29_2__27_  (.A1(u_multiplier_pp1_29 [5]),
    .A2(u_multiplier_pp1_29 [4]),
    .B1(u_multiplier_pp1_29 [6]),
    .B2(u_multiplier_pp1_29 [7]),
    .ZN(u_multiplier_STAGE2_acci_pp2_29_2__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_29_2__28_  (.A1(u_multiplier_STAGE2_acci_pp2_29_2__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_29_2__17_ ),
    .ZN(u_multiplier_pp2_30 [5]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_29_3__21_  (.A1(u_multiplier_pp1_29 [1]),
    .A2(u_multiplier_pp1_29 [0]),
    .A3(u_multiplier_pp1_29 [2]),
    .ZN(u_multiplier_STAGE2_acci_pp2_29_3__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_29_3__22_  (.A(u_multiplier_pp1_29 [1]),
    .B(u_multiplier_pp1_29 [0]),
    .Z(u_multiplier_STAGE2_acci_pp2_29_3__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_29_3__23_  (.A(u_multiplier_pp1_29 [2]),
    .B(u_multiplier_pp1_29 [3]),
    .Z(u_multiplier_STAGE2_acci_pp2_29_3__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_29_3__24_  (.A1(u_multiplier_STAGE2_acci_pp2_29_3__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_29_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_29_3__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_29_3__25_  (.A(u_multiplier_STAGE2_acci_pp2_29_3__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_29_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_29_3__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_29_3__26_  (.A1(u_multiplier_STAGE2_acci_pp2_29_3__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_29_3__16_ ),
    .ZN(u_multiplier_pp2_29 [3]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_29_3__27_  (.A1(u_multiplier_pp1_29 [1]),
    .A2(u_multiplier_pp1_29 [0]),
    .B1(u_multiplier_pp1_29 [2]),
    .B2(u_multiplier_pp1_29 [3]),
    .ZN(u_multiplier_STAGE2_acci_pp2_29_3__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_29_3__28_  (.A1(u_multiplier_STAGE2_acci_pp2_29_3__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_29_3__17_ ),
    .ZN(u_multiplier_pp2_30 [4]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_30_0__21_  (.A1(u_multiplier_pp1_30 [13]),
    .A2(u_multiplier_pp1_30 [12]),
    .A3(u_multiplier_pp1_30 [14]),
    .ZN(u_multiplier_STAGE2_acci_pp2_30_0__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_30_0__22_  (.A(u_multiplier_pp1_30 [13]),
    .B(u_multiplier_pp1_30 [12]),
    .Z(u_multiplier_STAGE2_acci_pp2_30_0__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_30_0__23_  (.A(u_multiplier_pp1_30 [14]),
    .B(u_multiplier_pp1_30 [15]),
    .Z(u_multiplier_STAGE2_acci_pp2_30_0__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_30_0__24_  (.A1(u_multiplier_STAGE2_acci_pp2_30_0__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_30_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_30_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_30_0__25_  (.A(u_multiplier_STAGE2_acci_pp2_30_0__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_30_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_30_0__16_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_30_0__26_  (.A1(u_multiplier_STAGE2_acci_pp2_30_0__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_30_0__16_ ),
    .ZN(u_multiplier_pp2_30 [0]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_30_0__27_  (.A1(u_multiplier_pp1_30 [13]),
    .A2(u_multiplier_pp1_30 [12]),
    .B1(u_multiplier_pp1_30 [14]),
    .B2(u_multiplier_pp1_30 [15]),
    .ZN(u_multiplier_STAGE2_acci_pp2_30_0__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_30_0__28_  (.A1(u_multiplier_STAGE2_acci_pp2_30_0__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_30_0__17_ ),
    .ZN(u_multiplier_pp2_31 [7]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_30_1__21_  (.A1(u_multiplier_pp1_30 [9]),
    .A2(u_multiplier_pp1_30 [8]),
    .A3(u_multiplier_pp1_30 [10]),
    .ZN(u_multiplier_STAGE2_acci_pp2_30_1__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_30_1__22_  (.A(u_multiplier_pp1_30 [9]),
    .B(u_multiplier_pp1_30 [8]),
    .Z(u_multiplier_STAGE2_acci_pp2_30_1__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_30_1__23_  (.A(u_multiplier_pp1_30 [10]),
    .B(u_multiplier_pp1_30 [11]),
    .Z(u_multiplier_STAGE2_acci_pp2_30_1__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_30_1__24_  (.A1(u_multiplier_STAGE2_acci_pp2_30_1__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_30_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_30_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_30_1__25_  (.A(u_multiplier_STAGE2_acci_pp2_30_1__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_30_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_30_1__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_30_1__26_  (.A1(u_multiplier_STAGE2_acci_pp2_30_1__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_30_1__16_ ),
    .ZN(u_multiplier_pp2_30 [1]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_30_1__27_  (.A1(u_multiplier_pp1_30 [9]),
    .A2(u_multiplier_pp1_30 [8]),
    .B1(u_multiplier_pp1_30 [10]),
    .B2(u_multiplier_pp1_30 [11]),
    .ZN(u_multiplier_STAGE2_acci_pp2_30_1__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_30_1__28_  (.A1(u_multiplier_STAGE2_acci_pp2_30_1__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_30_1__17_ ),
    .ZN(u_multiplier_pp2_31 [6]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_30_2__21_  (.A1(u_multiplier_pp1_30 [5]),
    .A2(u_multiplier_pp1_30 [4]),
    .A3(u_multiplier_pp1_30 [6]),
    .ZN(u_multiplier_STAGE2_acci_pp2_30_2__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_30_2__22_  (.A(u_multiplier_pp1_30 [5]),
    .B(u_multiplier_pp1_30 [4]),
    .Z(u_multiplier_STAGE2_acci_pp2_30_2__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_30_2__23_  (.A(u_multiplier_pp1_30 [6]),
    .B(u_multiplier_pp1_30 [7]),
    .Z(u_multiplier_STAGE2_acci_pp2_30_2__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_30_2__24_  (.A1(u_multiplier_STAGE2_acci_pp2_30_2__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_30_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_30_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_30_2__25_  (.A(u_multiplier_STAGE2_acci_pp2_30_2__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_30_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_30_2__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_30_2__26_  (.A1(u_multiplier_STAGE2_acci_pp2_30_2__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_30_2__16_ ),
    .ZN(u_multiplier_pp2_30 [2]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_30_2__27_  (.A1(u_multiplier_pp1_30 [5]),
    .A2(u_multiplier_pp1_30 [4]),
    .B1(u_multiplier_pp1_30 [6]),
    .B2(u_multiplier_pp1_30 [7]),
    .ZN(u_multiplier_STAGE2_acci_pp2_30_2__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_30_2__28_  (.A1(u_multiplier_STAGE2_acci_pp2_30_2__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_30_2__17_ ),
    .ZN(u_multiplier_pp2_31 [5]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_30_3__21_  (.A1(u_multiplier_pp1_30 [1]),
    .A2(u_multiplier_pp1_30 [0]),
    .A3(u_multiplier_pp1_30 [2]),
    .ZN(u_multiplier_STAGE2_acci_pp2_30_3__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_30_3__22_  (.A(u_multiplier_pp1_30 [1]),
    .B(u_multiplier_pp1_30 [0]),
    .Z(u_multiplier_STAGE2_acci_pp2_30_3__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_30_3__23_  (.A(u_multiplier_pp1_30 [2]),
    .B(u_multiplier_pp1_30 [3]),
    .Z(u_multiplier_STAGE2_acci_pp2_30_3__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_30_3__24_  (.A1(u_multiplier_STAGE2_acci_pp2_30_3__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_30_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_30_3__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_30_3__25_  (.A(u_multiplier_STAGE2_acci_pp2_30_3__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_30_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_30_3__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_30_3__26_  (.A1(u_multiplier_STAGE2_acci_pp2_30_3__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_30_3__16_ ),
    .ZN(u_multiplier_pp2_30 [3]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_30_3__27_  (.A1(u_multiplier_pp1_30 [1]),
    .A2(u_multiplier_pp1_30 [0]),
    .B1(u_multiplier_pp1_30 [2]),
    .B2(u_multiplier_pp1_30 [3]),
    .ZN(u_multiplier_STAGE2_acci_pp2_30_3__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_30_3__28_  (.A1(u_multiplier_STAGE2_acci_pp2_30_3__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_30_3__17_ ),
    .ZN(u_multiplier_pp2_31 [4]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_31_0__21_  (.A1(u_multiplier_pp1_31 [13]),
    .A2(u_multiplier_pp1_31 [12]),
    .A3(u_multiplier_pp1_31 [14]),
    .ZN(u_multiplier_STAGE2_acci_pp2_31_0__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_31_0__22_  (.A(u_multiplier_pp1_31 [13]),
    .B(u_multiplier_pp1_31 [12]),
    .Z(u_multiplier_STAGE2_acci_pp2_31_0__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_31_0__23_  (.A(u_multiplier_pp1_31 [14]),
    .B(u_multiplier_pp1_31 [15]),
    .Z(u_multiplier_STAGE2_acci_pp2_31_0__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_31_0__24_  (.A1(u_multiplier_STAGE2_acci_pp2_31_0__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_31_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_31_0__15_ ));
 XNOR2_X2 u_multiplier_STAGE2_acci_pp2_31_0__25_  (.A(u_multiplier_STAGE2_acci_pp2_31_0__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_31_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_31_0__16_ ));
 NAND2_X4 u_multiplier_STAGE2_acci_pp2_31_0__26_  (.A1(u_multiplier_STAGE2_acci_pp2_31_0__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_31_0__16_ ),
    .ZN(u_multiplier_pp2_31 [0]));
 AOI22_X4 u_multiplier_STAGE2_acci_pp2_31_0__27_  (.A1(u_multiplier_pp1_31 [13]),
    .A2(u_multiplier_pp1_31 [12]),
    .B1(u_multiplier_pp1_31 [14]),
    .B2(u_multiplier_pp1_31 [15]),
    .ZN(u_multiplier_STAGE2_acci_pp2_31_0__17_ ));
 NAND2_X4 u_multiplier_STAGE2_acci_pp2_31_0__28_  (.A1(u_multiplier_STAGE2_acci_pp2_31_0__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_31_0__17_ ),
    .ZN(u_multiplier_pp2_32 [7]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_31_1__21_  (.A1(u_multiplier_pp1_31 [9]),
    .A2(u_multiplier_pp1_31 [8]),
    .A3(u_multiplier_pp1_31 [10]),
    .ZN(u_multiplier_STAGE2_acci_pp2_31_1__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_31_1__22_  (.A(u_multiplier_pp1_31 [9]),
    .B(u_multiplier_pp1_31 [8]),
    .Z(u_multiplier_STAGE2_acci_pp2_31_1__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_31_1__23_  (.A(u_multiplier_pp1_31 [10]),
    .B(u_multiplier_pp1_31 [11]),
    .Z(u_multiplier_STAGE2_acci_pp2_31_1__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_31_1__24_  (.A1(u_multiplier_STAGE2_acci_pp2_31_1__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_31_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_31_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_31_1__25_  (.A(u_multiplier_STAGE2_acci_pp2_31_1__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_31_1__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_31_1__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_31_1__26_  (.A1(u_multiplier_STAGE2_acci_pp2_31_1__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_31_1__16_ ),
    .ZN(u_multiplier_pp2_31 [1]));
 AOI22_X2 u_multiplier_STAGE2_acci_pp2_31_1__27_  (.A1(u_multiplier_pp1_31 [9]),
    .A2(u_multiplier_pp1_31 [8]),
    .B1(u_multiplier_pp1_31 [10]),
    .B2(u_multiplier_pp1_31 [11]),
    .ZN(u_multiplier_STAGE2_acci_pp2_31_1__17_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_31_1__28_  (.A1(u_multiplier_STAGE2_acci_pp2_31_1__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_31_1__17_ ),
    .ZN(u_multiplier_pp2_32 [6]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_31_2__21_  (.A1(u_multiplier_pp1_31 [5]),
    .A2(u_multiplier_pp1_31 [4]),
    .A3(u_multiplier_pp1_31 [6]),
    .ZN(u_multiplier_STAGE2_acci_pp2_31_2__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_31_2__22_  (.A(u_multiplier_pp1_31 [5]),
    .B(u_multiplier_pp1_31 [4]),
    .Z(u_multiplier_STAGE2_acci_pp2_31_2__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_31_2__23_  (.A(u_multiplier_pp1_31 [6]),
    .B(u_multiplier_pp1_31 [7]),
    .Z(u_multiplier_STAGE2_acci_pp2_31_2__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_31_2__24_  (.A1(u_multiplier_STAGE2_acci_pp2_31_2__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_31_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_31_2__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_31_2__25_  (.A(u_multiplier_STAGE2_acci_pp2_31_2__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_31_2__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_31_2__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_31_2__26_  (.A1(u_multiplier_STAGE2_acci_pp2_31_2__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_31_2__16_ ),
    .ZN(u_multiplier_pp2_31 [2]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_31_2__27_  (.A1(u_multiplier_pp1_31 [5]),
    .A2(u_multiplier_pp1_31 [4]),
    .B1(u_multiplier_pp1_31 [6]),
    .B2(u_multiplier_pp1_31 [7]),
    .ZN(u_multiplier_STAGE2_acci_pp2_31_2__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_31_2__28_  (.A1(u_multiplier_STAGE2_acci_pp2_31_2__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_31_2__17_ ),
    .ZN(u_multiplier_pp2_32 [5]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_31_3__21_  (.A1(u_multiplier_pp1_31 [1]),
    .A2(u_multiplier_pp1_31 [0]),
    .A3(u_multiplier_pp1_31 [2]),
    .ZN(u_multiplier_STAGE2_acci_pp2_31_3__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_31_3__22_  (.A(u_multiplier_pp1_31 [1]),
    .B(u_multiplier_pp1_31 [0]),
    .Z(u_multiplier_STAGE2_acci_pp2_31_3__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_31_3__23_  (.A(u_multiplier_pp1_31 [2]),
    .B(u_multiplier_pp1_31 [3]),
    .Z(u_multiplier_STAGE2_acci_pp2_31_3__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_31_3__24_  (.A1(u_multiplier_STAGE2_acci_pp2_31_3__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_31_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_31_3__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_31_3__25_  (.A(u_multiplier_STAGE2_acci_pp2_31_3__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_31_3__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_31_3__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_31_3__26_  (.A1(u_multiplier_STAGE2_acci_pp2_31_3__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_31_3__16_ ),
    .ZN(u_multiplier_pp2_31 [3]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_31_3__27_  (.A1(u_multiplier_pp1_31 [1]),
    .A2(u_multiplier_pp1_31 [0]),
    .B1(u_multiplier_pp1_31 [2]),
    .B2(u_multiplier_pp1_31 [3]),
    .ZN(u_multiplier_STAGE2_acci_pp2_31_3__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_31_3__28_  (.A1(u_multiplier_STAGE2_acci_pp2_31_3__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_31_3__17_ ),
    .ZN(u_multiplier_pp2_32 [4]));
 NAND3_X1 u_multiplier_STAGE2_acci_pp2_9_0__21_  (.A1(u_multiplier_pp1_9 [7]),
    .A2(u_multiplier_pp1_9 [6]),
    .A3(u_multiplier_pp1_9 [8]),
    .ZN(u_multiplier_STAGE2_acci_pp2_9_0__18_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_9_0__22_  (.A(u_multiplier_pp1_9 [7]),
    .B(u_multiplier_pp1_9 [6]),
    .Z(u_multiplier_STAGE2_acci_pp2_9_0__19_ ));
 XOR2_X2 u_multiplier_STAGE2_acci_pp2_9_0__23_  (.A(u_multiplier_pp1_9 [8]),
    .B(u_multiplier_pp1_9 [9]),
    .Z(u_multiplier_STAGE2_acci_pp2_9_0__20_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_9_0__24_  (.A1(u_multiplier_STAGE2_acci_pp2_9_0__19_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_9_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_9_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE2_acci_pp2_9_0__25_  (.A(u_multiplier_STAGE2_acci_pp2_9_0__19_ ),
    .B(u_multiplier_STAGE2_acci_pp2_9_0__20_ ),
    .ZN(u_multiplier_STAGE2_acci_pp2_9_0__16_ ));
 NAND2_X2 u_multiplier_STAGE2_acci_pp2_9_0__26_  (.A1(u_multiplier_STAGE2_acci_pp2_9_0__18_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_9_0__16_ ),
    .ZN(u_multiplier_pp2_9 [0]));
 AOI22_X1 u_multiplier_STAGE2_acci_pp2_9_0__27_  (.A1(u_multiplier_pp1_9 [7]),
    .A2(u_multiplier_pp1_9 [6]),
    .B1(u_multiplier_pp1_9 [8]),
    .B2(u_multiplier_pp1_9 [9]),
    .ZN(u_multiplier_STAGE2_acci_pp2_9_0__17_ ));
 NAND2_X1 u_multiplier_STAGE2_acci_pp2_9_0__28_  (.A1(u_multiplier_STAGE2_acci_pp2_9_0__15_ ),
    .A2(u_multiplier_STAGE2_acci_pp2_9_0__17_ ),
    .ZN(u_multiplier_pp2_10 [2]));
 LOGIC0_X1 u_multiplier_STAGE3_E_4_2_pp3_32_1__18__133  (.Z(net133));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_32_1__18_  (.A(net133),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_32_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_32_1__19_  (.A1(u_multiplier_pp2_32 [1]),
    .A2(u_multiplier_pp2_32 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_32_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_32_1__20_  (.A(u_multiplier_pp2_32 [1]),
    .B(u_multiplier_pp2_32 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_32_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_32_1__21_  (.A1(u_multiplier_pp2_32 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_32_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_32_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_32_1__22_  (.A(u_multiplier_pp2_32 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_32_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_32_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_32_1__23_  (.A1(u_multiplier_pp2_32 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_32_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_32_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_32_1__24_  (.A(u_multiplier_pp2_32 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_32_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_32_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_32_1__25_  (.A(net134),
    .B(u_multiplier_STAGE3_E_4_2_pp3_32_1__16_ ),
    .ZN(u_multiplier_pp3_32 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_32_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_32_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_32_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_32_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_32_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_32_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_32_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_32_1__17_ ),
    .ZN(u_multiplier_pp3_33 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_32_2__18_  (.A(net135),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_32_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_32_2__19_  (.A1(u_multiplier_pp2_32 [5]),
    .A2(u_multiplier_pp2_32 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_32_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_32_2__20_  (.A(u_multiplier_pp2_32 [5]),
    .B(u_multiplier_pp2_32 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_32_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_32_2__21_  (.A1(u_multiplier_pp2_32 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_32_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_32_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_32_2__22_  (.A(u_multiplier_pp2_32 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_32_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_32_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_32_2__23_  (.A1(u_multiplier_pp2_32 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_32_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_32_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_32_2__24_  (.A(u_multiplier_pp2_32 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_32_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_32_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_32_2__25_  (.A(net136),
    .B(u_multiplier_STAGE3_E_4_2_pp3_32_2__16_ ),
    .ZN(u_multiplier_pp3_32 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_32_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_32_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_32_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_32_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_32_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_32_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_32_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_32_2__17_ ),
    .ZN(u_multiplier_pp3_33 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_33_1__18_  (.A(u_multiplier_STAGE3_pp3_32_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_33_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_33_1__19_  (.A1(u_multiplier_pp2_33 [1]),
    .A2(u_multiplier_pp2_33 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_33_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_33_1__20_  (.A(u_multiplier_pp2_33 [1]),
    .B(u_multiplier_pp2_33 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_33_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_33_1__21_  (.A1(u_multiplier_pp2_33 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_33_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_33_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_33_1__22_  (.A(u_multiplier_pp2_33 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_33_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_33_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_33_1__23_  (.A1(u_multiplier_pp2_33 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_33_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_33_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_33_1__24_  (.A(u_multiplier_pp2_33 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_33_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_33_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_33_1__25_  (.A(u_multiplier_STAGE3_pp3_32_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_33_1__16_ ),
    .ZN(u_multiplier_pp3_33 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_33_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_33_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_33_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_33_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_33_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_33_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_33_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_33_1__17_ ),
    .ZN(u_multiplier_pp3_34 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_33_2__18_  (.A(u_multiplier_STAGE3_pp3_32_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_33_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_33_2__19_  (.A1(u_multiplier_pp2_33 [5]),
    .A2(u_multiplier_pp2_33 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_33_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_33_2__20_  (.A(u_multiplier_pp2_33 [5]),
    .B(u_multiplier_pp2_33 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_33_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_33_2__21_  (.A1(u_multiplier_pp2_33 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_33_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_33_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_33_2__22_  (.A(u_multiplier_pp2_33 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_33_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_33_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_33_2__23_  (.A1(u_multiplier_pp2_33 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_33_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_33_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_33_2__24_  (.A(u_multiplier_pp2_33 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_33_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_33_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_33_2__25_  (.A(u_multiplier_STAGE3_pp3_32_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_33_2__16_ ),
    .ZN(u_multiplier_pp3_33 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_33_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_33_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_33_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_33_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_33_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_33_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_33_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_33_2__17_ ),
    .ZN(u_multiplier_pp3_34 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_34_1__18_  (.A(u_multiplier_STAGE3_pp3_33_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_34_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_34_1__19_  (.A1(u_multiplier_pp2_34 [1]),
    .A2(u_multiplier_pp2_34 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_34_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_34_1__20_  (.A(u_multiplier_pp2_34 [1]),
    .B(u_multiplier_pp2_34 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_34_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_34_1__21_  (.A1(u_multiplier_pp2_34 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_34_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_34_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_34_1__22_  (.A(u_multiplier_pp2_34 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_34_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_34_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_34_1__23_  (.A1(u_multiplier_pp2_34 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_34_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_34_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_34_1__24_  (.A(u_multiplier_pp2_34 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_34_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_34_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_34_1__25_  (.A(u_multiplier_STAGE3_pp3_33_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_34_1__16_ ),
    .ZN(u_multiplier_pp3_34 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_34_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_34_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_34_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_34_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_34_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_34_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_34_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_34_1__17_ ),
    .ZN(u_multiplier_pp3_35 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_34_2__18_  (.A(u_multiplier_STAGE3_pp3_33_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_34_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_34_2__19_  (.A1(u_multiplier_pp2_34 [5]),
    .A2(u_multiplier_pp2_34 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_34_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_34_2__20_  (.A(u_multiplier_pp2_34 [5]),
    .B(u_multiplier_pp2_34 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_34_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_34_2__21_  (.A1(u_multiplier_pp2_34 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_34_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_34_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_34_2__22_  (.A(u_multiplier_pp2_34 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_34_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_34_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_34_2__23_  (.A1(u_multiplier_pp2_34 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_34_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_34_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_34_2__24_  (.A(u_multiplier_pp2_34 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_34_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_34_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_34_2__25_  (.A(u_multiplier_STAGE3_pp3_33_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_34_2__16_ ),
    .ZN(u_multiplier_pp3_34 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_34_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_34_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_34_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_34_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_34_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_34_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_34_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_34_2__17_ ),
    .ZN(u_multiplier_pp3_35 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_35_1__18_  (.A(u_multiplier_STAGE3_pp3_34_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_35_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_35_1__19_  (.A1(u_multiplier_pp2_35 [1]),
    .A2(u_multiplier_pp2_35 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_35_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_35_1__20_  (.A(u_multiplier_pp2_35 [1]),
    .B(u_multiplier_pp2_35 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_35_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_35_1__21_  (.A1(u_multiplier_pp2_35 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_35_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_35_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_35_1__22_  (.A(u_multiplier_pp2_35 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_35_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_35_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_35_1__23_  (.A1(u_multiplier_pp2_35 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_35_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_35_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_35_1__24_  (.A(u_multiplier_pp2_35 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_35_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_35_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_35_1__25_  (.A(u_multiplier_STAGE3_pp3_34_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_35_1__16_ ),
    .ZN(u_multiplier_pp3_35 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_35_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_35_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_35_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_35_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_35_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_35_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_35_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_35_1__17_ ),
    .ZN(u_multiplier_pp3_36 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_35_2__18_  (.A(u_multiplier_STAGE3_pp3_34_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_35_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_35_2__19_  (.A1(u_multiplier_pp2_35 [5]),
    .A2(u_multiplier_pp2_35 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_35_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_35_2__20_  (.A(u_multiplier_pp2_35 [5]),
    .B(u_multiplier_pp2_35 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_35_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_35_2__21_  (.A1(u_multiplier_pp2_35 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_35_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_35_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_35_2__22_  (.A(u_multiplier_pp2_35 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_35_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_35_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_35_2__23_  (.A1(u_multiplier_pp2_35 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_35_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_35_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_35_2__24_  (.A(u_multiplier_pp2_35 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_35_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_35_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_35_2__25_  (.A(u_multiplier_STAGE3_pp3_34_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_35_2__16_ ),
    .ZN(u_multiplier_pp3_35 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_35_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_35_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_35_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_35_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_35_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_35_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_35_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_35_2__17_ ),
    .ZN(u_multiplier_pp3_36 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_36_1__18_  (.A(u_multiplier_STAGE3_pp3_35_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_36_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_36_1__19_  (.A1(u_multiplier_pp2_36 [1]),
    .A2(u_multiplier_pp2_36 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_36_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_36_1__20_  (.A(u_multiplier_pp2_36 [1]),
    .B(u_multiplier_pp2_36 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_36_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_36_1__21_  (.A1(u_multiplier_pp2_36 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_36_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_36_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_36_1__22_  (.A(u_multiplier_pp2_36 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_36_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_36_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_36_1__23_  (.A1(u_multiplier_pp2_36 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_36_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_36_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_36_1__24_  (.A(u_multiplier_pp2_36 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_36_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_36_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_36_1__25_  (.A(u_multiplier_STAGE3_pp3_35_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_36_1__16_ ),
    .ZN(u_multiplier_pp3_36 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_36_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_36_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_36_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_36_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_36_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_36_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_36_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_36_1__17_ ),
    .ZN(u_multiplier_pp3_37 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_36_2__18_  (.A(u_multiplier_STAGE3_pp3_35_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_36_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_36_2__19_  (.A1(u_multiplier_pp2_36 [5]),
    .A2(u_multiplier_pp2_36 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_36_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_36_2__20_  (.A(u_multiplier_pp2_36 [5]),
    .B(u_multiplier_pp2_36 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_36_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_36_2__21_  (.A1(u_multiplier_pp2_36 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_36_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_36_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_36_2__22_  (.A(u_multiplier_pp2_36 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_36_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_36_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_36_2__23_  (.A1(u_multiplier_pp2_36 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_36_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_36_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_36_2__24_  (.A(u_multiplier_pp2_36 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_36_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_36_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_36_2__25_  (.A(u_multiplier_STAGE3_pp3_35_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_36_2__16_ ),
    .ZN(u_multiplier_pp3_36 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_36_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_36_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_36_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_36_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_36_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_36_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_36_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_36_2__17_ ),
    .ZN(u_multiplier_pp3_37 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_37_1__18_  (.A(u_multiplier_STAGE3_pp3_36_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_37_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_37_1__19_  (.A1(u_multiplier_pp2_37 [1]),
    .A2(u_multiplier_pp2_37 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_37_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_37_1__20_  (.A(u_multiplier_pp2_37 [1]),
    .B(u_multiplier_pp2_37 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_37_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_37_1__21_  (.A1(u_multiplier_pp2_37 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_37_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_37_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_37_1__22_  (.A(u_multiplier_pp2_37 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_37_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_37_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_37_1__23_  (.A1(u_multiplier_pp2_37 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_37_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_37_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_37_1__24_  (.A(u_multiplier_pp2_37 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_37_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_37_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_37_1__25_  (.A(u_multiplier_STAGE3_pp3_36_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_37_1__16_ ),
    .ZN(u_multiplier_pp3_37 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_37_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_37_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_37_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_37_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_37_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_37_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_37_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_37_1__17_ ),
    .ZN(u_multiplier_pp3_38 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_37_2__18_  (.A(u_multiplier_STAGE3_pp3_36_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_37_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_37_2__19_  (.A1(u_multiplier_pp2_37 [5]),
    .A2(u_multiplier_pp2_37 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_37_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_37_2__20_  (.A(u_multiplier_pp2_37 [5]),
    .B(u_multiplier_pp2_37 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_37_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_37_2__21_  (.A1(u_multiplier_pp2_37 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_37_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_37_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_37_2__22_  (.A(u_multiplier_pp2_37 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_37_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_37_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_37_2__23_  (.A1(u_multiplier_pp2_37 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_37_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_37_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_37_2__24_  (.A(u_multiplier_pp2_37 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_37_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_37_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_37_2__25_  (.A(u_multiplier_STAGE3_pp3_36_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_37_2__16_ ),
    .ZN(u_multiplier_pp3_37 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_37_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_37_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_37_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_37_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_37_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_37_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_37_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_37_2__17_ ),
    .ZN(u_multiplier_pp3_38 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_38_1__18_  (.A(u_multiplier_STAGE3_pp3_37_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_38_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_38_1__19_  (.A1(u_multiplier_pp2_38 [1]),
    .A2(u_multiplier_pp2_38 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_38_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_38_1__20_  (.A(u_multiplier_pp2_38 [1]),
    .B(u_multiplier_pp2_38 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_38_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_38_1__21_  (.A1(u_multiplier_pp2_38 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_38_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_38_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_38_1__22_  (.A(u_multiplier_pp2_38 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_38_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_38_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_38_1__23_  (.A1(u_multiplier_pp2_38 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_38_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_38_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_38_1__24_  (.A(u_multiplier_pp2_38 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_38_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_38_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_38_1__25_  (.A(u_multiplier_STAGE3_pp3_37_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_38_1__16_ ),
    .ZN(u_multiplier_pp3_38 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_38_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_38_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_38_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_38_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_38_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_38_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_38_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_38_1__17_ ),
    .ZN(u_multiplier_pp3_39 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_38_2__18_  (.A(u_multiplier_STAGE3_pp3_37_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_38_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_38_2__19_  (.A1(u_multiplier_pp2_38 [5]),
    .A2(u_multiplier_pp2_38 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_38_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_38_2__20_  (.A(u_multiplier_pp2_38 [5]),
    .B(u_multiplier_pp2_38 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_38_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_38_2__21_  (.A1(u_multiplier_pp2_38 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_38_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_38_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_38_2__22_  (.A(u_multiplier_pp2_38 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_38_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_38_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_38_2__23_  (.A1(u_multiplier_pp2_38 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_38_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_38_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_38_2__24_  (.A(u_multiplier_pp2_38 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_38_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_38_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_38_2__25_  (.A(u_multiplier_STAGE3_pp3_37_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_38_2__16_ ),
    .ZN(u_multiplier_pp3_38 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_38_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_38_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_38_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_38_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_38_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_38_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_38_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_38_2__17_ ),
    .ZN(u_multiplier_pp3_39 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_39_1__18_  (.A(u_multiplier_STAGE3_pp3_38_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_39_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_39_1__19_  (.A1(u_multiplier_pp2_39 [1]),
    .A2(u_multiplier_pp2_39 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_39_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_39_1__20_  (.A(u_multiplier_pp2_39 [1]),
    .B(u_multiplier_pp2_39 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_39_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_39_1__21_  (.A1(u_multiplier_pp2_39 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_39_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_39_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_39_1__22_  (.A(u_multiplier_pp2_39 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_39_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_39_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_39_1__23_  (.A1(u_multiplier_pp2_39 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_39_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_39_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_39_1__24_  (.A(u_multiplier_pp2_39 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_39_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_39_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_39_1__25_  (.A(u_multiplier_STAGE3_pp3_38_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_39_1__16_ ),
    .ZN(u_multiplier_pp3_39 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_39_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_39_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_39_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_39_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_39_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_39_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_39_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_39_1__17_ ),
    .ZN(u_multiplier_pp3_40 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_39_2__18_  (.A(u_multiplier_STAGE3_pp3_38_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_39_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_39_2__19_  (.A1(u_multiplier_pp2_39 [5]),
    .A2(u_multiplier_pp2_39 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_39_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_39_2__20_  (.A(u_multiplier_pp2_39 [5]),
    .B(u_multiplier_pp2_39 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_39_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_39_2__21_  (.A1(u_multiplier_pp2_39 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_39_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_39_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_39_2__22_  (.A(u_multiplier_pp2_39 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_39_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_39_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_39_2__23_  (.A1(u_multiplier_pp2_39 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_39_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_39_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_39_2__24_  (.A(u_multiplier_pp2_39 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_39_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_39_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_39_2__25_  (.A(u_multiplier_STAGE3_pp3_38_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_39_2__16_ ),
    .ZN(u_multiplier_pp3_39 [0]));
 NAND2_X2 u_multiplier_STAGE3_E_4_2_pp3_39_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_39_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_39_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_39_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_39_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_39_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_39_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_39_2__17_ ),
    .ZN(u_multiplier_pp3_40 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_40_1__18_  (.A(u_multiplier_STAGE3_pp3_39_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_40_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_40_1__19_  (.A1(u_multiplier_pp2_40 [1]),
    .A2(u_multiplier_pp2_40 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_40_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_40_1__20_  (.A(u_multiplier_pp2_40 [1]),
    .B(u_multiplier_pp2_40 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_40_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_40_1__21_  (.A1(u_multiplier_pp2_40 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_40_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_40_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_40_1__22_  (.A(u_multiplier_pp2_40 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_40_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_40_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_40_1__23_  (.A1(u_multiplier_pp2_40 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_40_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_40_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_40_1__24_  (.A(u_multiplier_pp2_40 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_40_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_40_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_40_1__25_  (.A(u_multiplier_STAGE3_pp3_39_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_40_1__16_ ),
    .ZN(u_multiplier_pp3_40 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_40_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_40_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_40_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_40_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_40_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_40_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_40_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_40_1__17_ ),
    .ZN(u_multiplier_pp3_41 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_40_2__18_  (.A(u_multiplier_STAGE3_pp3_39_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_40_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_40_2__19_  (.A1(u_multiplier_pp2_40 [5]),
    .A2(u_multiplier_pp2_40 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_40_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_40_2__20_  (.A(u_multiplier_pp2_40 [5]),
    .B(u_multiplier_pp2_40 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_40_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_40_2__21_  (.A1(u_multiplier_pp2_40 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_40_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_40_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_40_2__22_  (.A(u_multiplier_pp2_40 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_40_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_40_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_40_2__23_  (.A1(u_multiplier_pp2_40 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_40_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_40_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_40_2__24_  (.A(u_multiplier_pp2_40 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_40_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_40_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_40_2__25_  (.A(u_multiplier_STAGE3_pp3_39_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_40_2__16_ ),
    .ZN(u_multiplier_pp3_40 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_40_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_40_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_40_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_40_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_40_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_40_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_40_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_40_2__17_ ),
    .ZN(u_multiplier_pp3_41 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_41_1__18_  (.A(u_multiplier_STAGE3_pp3_40_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_41_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_41_1__19_  (.A1(u_multiplier_pp2_41 [1]),
    .A2(u_multiplier_pp2_41 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_41_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_41_1__20_  (.A(u_multiplier_pp2_41 [1]),
    .B(u_multiplier_pp2_41 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_41_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_41_1__21_  (.A1(u_multiplier_pp2_41 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_41_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_41_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_41_1__22_  (.A(u_multiplier_pp2_41 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_41_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_41_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_41_1__23_  (.A1(u_multiplier_pp2_41 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_41_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_41_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_41_1__24_  (.A(u_multiplier_pp2_41 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_41_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_41_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_41_1__25_  (.A(u_multiplier_STAGE3_pp3_40_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_41_1__16_ ),
    .ZN(u_multiplier_pp3_41 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_41_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_41_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_41_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_41_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_41_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_41_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_41_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_41_1__17_ ),
    .ZN(u_multiplier_pp3_42 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_41_2__18_  (.A(u_multiplier_STAGE3_pp3_40_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_41_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_41_2__19_  (.A1(u_multiplier_pp2_41 [5]),
    .A2(u_multiplier_pp2_41 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_41_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_41_2__20_  (.A(u_multiplier_pp2_41 [5]),
    .B(u_multiplier_pp2_41 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_41_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_41_2__21_  (.A1(u_multiplier_pp2_41 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_41_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_41_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_41_2__22_  (.A(u_multiplier_pp2_41 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_41_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_41_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_41_2__23_  (.A1(u_multiplier_pp2_41 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_41_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_41_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_41_2__24_  (.A(u_multiplier_pp2_41 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_41_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_41_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_41_2__25_  (.A(u_multiplier_STAGE3_pp3_40_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_41_2__16_ ),
    .ZN(u_multiplier_pp3_41 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_41_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_41_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_41_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_41_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_41_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_41_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_41_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_41_2__17_ ),
    .ZN(u_multiplier_pp3_42 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_42_1__18_  (.A(u_multiplier_STAGE3_pp3_41_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_42_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_42_1__19_  (.A1(u_multiplier_pp2_42 [1]),
    .A2(u_multiplier_pp2_42 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_42_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_42_1__20_  (.A(u_multiplier_pp2_42 [1]),
    .B(u_multiplier_pp2_42 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_42_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_42_1__21_  (.A1(u_multiplier_pp2_42 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_42_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_42_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_42_1__22_  (.A(u_multiplier_pp2_42 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_42_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_42_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_42_1__23_  (.A1(u_multiplier_pp2_42 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_42_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_42_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_42_1__24_  (.A(u_multiplier_pp2_42 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_42_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_42_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_42_1__25_  (.A(u_multiplier_STAGE3_pp3_41_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_42_1__16_ ),
    .ZN(u_multiplier_pp3_42 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_42_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_42_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_42_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_42_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_42_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_42_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_42_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_42_1__17_ ),
    .ZN(u_multiplier_pp3_43 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_42_2__18_  (.A(u_multiplier_STAGE3_pp3_41_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_42_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_42_2__19_  (.A1(u_multiplier_pp2_42 [5]),
    .A2(u_multiplier_pp2_42 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_42_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_42_2__20_  (.A(u_multiplier_pp2_42 [5]),
    .B(u_multiplier_pp2_42 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_42_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_42_2__21_  (.A1(u_multiplier_pp2_42 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_42_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_42_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_42_2__22_  (.A(u_multiplier_pp2_42 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_42_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_42_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_42_2__23_  (.A1(u_multiplier_pp2_42 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_42_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_42_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_42_2__24_  (.A(u_multiplier_pp2_42 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_42_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_42_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_42_2__25_  (.A(u_multiplier_STAGE3_pp3_41_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_42_2__16_ ),
    .ZN(u_multiplier_pp3_42 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_42_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_42_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_42_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_42_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_42_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_42_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_42_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_42_2__17_ ),
    .ZN(u_multiplier_pp3_43 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_43_1__18_  (.A(u_multiplier_STAGE3_pp3_42_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_43_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_43_1__19_  (.A1(u_multiplier_pp2_43 [1]),
    .A2(u_multiplier_pp2_43 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_43_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_43_1__20_  (.A(u_multiplier_pp2_43 [1]),
    .B(u_multiplier_pp2_43 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_43_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_43_1__21_  (.A1(u_multiplier_pp2_43 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_43_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_43_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_43_1__22_  (.A(u_multiplier_pp2_43 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_43_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_43_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_43_1__23_  (.A1(u_multiplier_pp2_43 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_43_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_43_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_43_1__24_  (.A(u_multiplier_pp2_43 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_43_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_43_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_43_1__25_  (.A(u_multiplier_STAGE3_pp3_42_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_43_1__16_ ),
    .ZN(u_multiplier_pp3_43 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_43_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_43_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_43_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_43_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_43_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_43_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_43_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_43_1__17_ ),
    .ZN(u_multiplier_pp3_44 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_43_2__18_  (.A(u_multiplier_STAGE3_pp3_42_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_43_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_43_2__19_  (.A1(u_multiplier_pp2_43 [5]),
    .A2(u_multiplier_pp2_43 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_43_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_43_2__20_  (.A(u_multiplier_pp2_43 [5]),
    .B(u_multiplier_pp2_43 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_43_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_43_2__21_  (.A1(u_multiplier_pp2_43 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_43_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_43_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_43_2__22_  (.A(u_multiplier_pp2_43 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_43_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_43_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_43_2__23_  (.A1(u_multiplier_pp2_43 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_43_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_43_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_43_2__24_  (.A(u_multiplier_pp2_43 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_43_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_43_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_43_2__25_  (.A(u_multiplier_STAGE3_pp3_42_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_43_2__16_ ),
    .ZN(u_multiplier_pp3_43 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_43_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_43_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_43_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_43_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_43_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_43_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_43_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_43_2__17_ ),
    .ZN(u_multiplier_pp3_44 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_44_1__18_  (.A(u_multiplier_STAGE3_pp3_43_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_44_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_44_1__19_  (.A1(u_multiplier_pp2_44 [1]),
    .A2(u_multiplier_pp2_44 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_44_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_44_1__20_  (.A(u_multiplier_pp2_44 [1]),
    .B(u_multiplier_pp2_44 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_44_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_44_1__21_  (.A1(u_multiplier_pp2_44 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_44_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_44_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_44_1__22_  (.A(u_multiplier_pp2_44 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_44_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_44_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_44_1__23_  (.A1(u_multiplier_pp2_44 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_44_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_44_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_44_1__24_  (.A(u_multiplier_pp2_44 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_44_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_44_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_44_1__25_  (.A(u_multiplier_STAGE3_pp3_43_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_44_1__16_ ),
    .ZN(u_multiplier_pp3_44 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_44_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_44_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_44_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_44_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_44_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_44_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_44_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_44_1__17_ ),
    .ZN(u_multiplier_pp3_45 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_44_2__18_  (.A(u_multiplier_STAGE3_pp3_43_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_44_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_44_2__19_  (.A1(u_multiplier_pp2_44 [5]),
    .A2(u_multiplier_pp2_44 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_44_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_44_2__20_  (.A(u_multiplier_pp2_44 [5]),
    .B(u_multiplier_pp2_44 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_44_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_44_2__21_  (.A1(u_multiplier_pp2_44 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_44_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_44_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_44_2__22_  (.A(u_multiplier_pp2_44 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_44_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_44_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_44_2__23_  (.A1(u_multiplier_pp2_44 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_44_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_44_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_44_2__24_  (.A(u_multiplier_pp2_44 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_44_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_44_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_44_2__25_  (.A(u_multiplier_STAGE3_pp3_43_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_44_2__16_ ),
    .ZN(u_multiplier_pp3_44 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_44_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_44_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_44_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_44_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_44_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_44_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_44_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_44_2__17_ ),
    .ZN(u_multiplier_pp3_45 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_45_1__18_  (.A(u_multiplier_STAGE3_pp3_44_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_45_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_45_1__19_  (.A1(u_multiplier_pp2_45 [1]),
    .A2(u_multiplier_pp2_45 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_45_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_45_1__20_  (.A(u_multiplier_pp2_45 [1]),
    .B(u_multiplier_pp2_45 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_45_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_45_1__21_  (.A1(u_multiplier_pp2_45 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_45_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_45_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_45_1__22_  (.A(u_multiplier_pp2_45 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_45_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_45_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_45_1__23_  (.A1(u_multiplier_pp2_45 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_45_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_45_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_45_1__24_  (.A(u_multiplier_pp2_45 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_45_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_45_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_45_1__25_  (.A(u_multiplier_STAGE3_pp3_44_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_45_1__16_ ),
    .ZN(u_multiplier_pp3_45 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_45_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_45_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_45_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_45_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_45_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_45_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_45_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_45_1__17_ ),
    .ZN(u_multiplier_pp3_46 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_45_2__18_  (.A(u_multiplier_STAGE3_pp3_44_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_45_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_45_2__19_  (.A1(u_multiplier_pp2_45 [5]),
    .A2(u_multiplier_pp2_45 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_45_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_45_2__20_  (.A(u_multiplier_pp2_45 [5]),
    .B(u_multiplier_pp2_45 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_45_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_45_2__21_  (.A1(u_multiplier_pp2_45 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_45_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_45_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_45_2__22_  (.A(u_multiplier_pp2_45 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_45_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_45_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_45_2__23_  (.A1(u_multiplier_pp2_45 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_45_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_45_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_45_2__24_  (.A(u_multiplier_pp2_45 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_45_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_45_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_45_2__25_  (.A(u_multiplier_STAGE3_pp3_44_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_45_2__16_ ),
    .ZN(u_multiplier_pp3_45 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_45_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_45_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_45_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_45_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_45_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_45_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_45_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_45_2__17_ ),
    .ZN(u_multiplier_pp3_46 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_46_1__18_  (.A(u_multiplier_STAGE3_pp3_45_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_46_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_46_1__19_  (.A1(u_multiplier_pp2_46 [1]),
    .A2(u_multiplier_pp2_46 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_46_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_46_1__20_  (.A(u_multiplier_pp2_46 [1]),
    .B(u_multiplier_pp2_46 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_46_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_46_1__21_  (.A1(u_multiplier_pp2_46 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_46_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_46_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_46_1__22_  (.A(u_multiplier_pp2_46 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_46_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_46_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_46_1__23_  (.A1(u_multiplier_pp2_46 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_46_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_46_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_46_1__24_  (.A(u_multiplier_pp2_46 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_46_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_46_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_46_1__25_  (.A(u_multiplier_STAGE3_pp3_45_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_46_1__16_ ),
    .ZN(u_multiplier_pp3_46 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_46_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_46_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_46_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_46_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_46_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_46_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_46_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_46_1__17_ ),
    .ZN(u_multiplier_pp3_47 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_46_2__18_  (.A(u_multiplier_STAGE3_pp3_45_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_46_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_46_2__19_  (.A1(u_multiplier_pp2_46 [5]),
    .A2(u_multiplier_pp2_46 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_46_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_46_2__20_  (.A(u_multiplier_pp2_46 [5]),
    .B(u_multiplier_pp2_46 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_46_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_46_2__21_  (.A1(u_multiplier_pp2_46 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_46_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_46_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_46_2__22_  (.A(u_multiplier_pp2_46 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_46_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_46_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_46_2__23_  (.A1(u_multiplier_pp2_46 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_46_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_46_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_46_2__24_  (.A(u_multiplier_pp2_46 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_46_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_46_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_46_2__25_  (.A(u_multiplier_STAGE3_pp3_45_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_46_2__16_ ),
    .ZN(u_multiplier_pp3_46 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_46_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_46_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_46_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_46_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_46_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_46_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_46_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_46_2__17_ ),
    .ZN(u_multiplier_pp3_47 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_47_1__18_  (.A(u_multiplier_STAGE3_pp3_46_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_47_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_47_1__19_  (.A1(u_multiplier_pp2_47 [1]),
    .A2(u_multiplier_pp2_47 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_47_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_47_1__20_  (.A(u_multiplier_pp2_47 [1]),
    .B(u_multiplier_pp2_47 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_47_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_47_1__21_  (.A1(u_multiplier_pp2_47 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_47_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_47_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_47_1__22_  (.A(u_multiplier_pp2_47 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_47_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_47_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_47_1__23_  (.A1(u_multiplier_pp2_47 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_47_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_47_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_47_1__24_  (.A(u_multiplier_pp2_47 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_47_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_47_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_47_1__25_  (.A(u_multiplier_STAGE3_pp3_46_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_47_1__16_ ),
    .ZN(u_multiplier_pp3_47 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_47_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_47_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_47_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_47_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_47_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_47_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_47_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_47_1__17_ ),
    .ZN(u_multiplier_pp3_48 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_47_2__18_  (.A(u_multiplier_STAGE3_pp3_46_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_47_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_47_2__19_  (.A1(u_multiplier_pp2_47 [5]),
    .A2(u_multiplier_pp2_47 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_47_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_47_2__20_  (.A(u_multiplier_pp2_47 [5]),
    .B(u_multiplier_pp2_47 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_47_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_47_2__21_  (.A1(u_multiplier_pp2_47 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_47_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_47_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_47_2__22_  (.A(u_multiplier_pp2_47 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_47_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_47_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_47_2__23_  (.A1(u_multiplier_pp2_47 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_47_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_47_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_47_2__24_  (.A(u_multiplier_pp2_47 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_47_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_47_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_47_2__25_  (.A(u_multiplier_STAGE3_pp3_46_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_47_2__16_ ),
    .ZN(u_multiplier_pp3_47 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_47_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_47_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_47_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_47_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_47_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_47_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_47_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_47_2__17_ ),
    .ZN(u_multiplier_pp3_48 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_48_1__18_  (.A(u_multiplier_STAGE3_pp3_47_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_48_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_48_1__19_  (.A1(u_multiplier_pp2_48 [1]),
    .A2(u_multiplier_pp2_48 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_48_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_48_1__20_  (.A(u_multiplier_pp2_48 [1]),
    .B(u_multiplier_pp2_48 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_48_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_48_1__21_  (.A1(u_multiplier_pp2_48 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_48_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_48_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_48_1__22_  (.A(u_multiplier_pp2_48 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_48_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_48_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_48_1__23_  (.A1(u_multiplier_pp2_48 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_48_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_48_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_48_1__24_  (.A(u_multiplier_pp2_48 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_48_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_48_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_48_1__25_  (.A(u_multiplier_STAGE3_pp3_47_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_48_1__16_ ),
    .ZN(u_multiplier_pp3_48 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_48_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_48_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_48_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_48_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_48_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_48_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_48_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_48_1__17_ ),
    .ZN(u_multiplier_pp3_49 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_48_2__18_  (.A(u_multiplier_STAGE3_pp3_47_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_48_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_48_2__19_  (.A1(u_multiplier_pp2_48 [5]),
    .A2(u_multiplier_pp2_48 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_48_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_48_2__20_  (.A(u_multiplier_pp2_48 [5]),
    .B(u_multiplier_pp2_48 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_48_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_48_2__21_  (.A1(u_multiplier_pp2_48 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_48_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_48_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_48_2__22_  (.A(u_multiplier_pp2_48 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_48_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_48_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_48_2__23_  (.A1(u_multiplier_pp2_48 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_48_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_48_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_48_2__24_  (.A(u_multiplier_pp2_48 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_48_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_48_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_48_2__25_  (.A(u_multiplier_STAGE3_pp3_47_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_48_2__16_ ),
    .ZN(u_multiplier_pp3_48 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_48_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_48_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_48_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_48_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_48_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_48_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_48_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_48_2__17_ ),
    .ZN(u_multiplier_pp3_49 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_49_1__18_  (.A(u_multiplier_STAGE3_pp3_48_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_49_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_49_1__19_  (.A1(u_multiplier_pp2_49 [1]),
    .A2(u_multiplier_pp2_49 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_49_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_49_1__20_  (.A(u_multiplier_pp2_49 [1]),
    .B(u_multiplier_pp2_49 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_49_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_49_1__21_  (.A1(u_multiplier_pp2_49 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_49_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_49_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_49_1__22_  (.A(u_multiplier_pp2_49 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_49_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_49_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_49_1__23_  (.A1(u_multiplier_pp2_49 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_49_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_49_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_49_1__24_  (.A(u_multiplier_pp2_49 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_49_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_49_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_49_1__25_  (.A(u_multiplier_STAGE3_pp3_48_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_49_1__16_ ),
    .ZN(u_multiplier_pp3_49 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_49_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_49_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_49_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_49_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_49_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_49_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_49_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_49_1__17_ ),
    .ZN(u_multiplier_pp3_50 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_49_2__18_  (.A(u_multiplier_STAGE3_pp3_48_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_49_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_49_2__19_  (.A1(u_multiplier_pp2_49 [5]),
    .A2(u_multiplier_pp2_49 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_49_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_49_2__20_  (.A(u_multiplier_pp2_49 [5]),
    .B(u_multiplier_pp2_49 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_49_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_49_2__21_  (.A1(u_multiplier_pp2_49 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_49_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_49_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_49_2__22_  (.A(u_multiplier_pp2_49 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_49_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_49_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_49_2__23_  (.A1(u_multiplier_pp2_49 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_49_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_49_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_49_2__24_  (.A(u_multiplier_pp2_49 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_49_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_49_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_49_2__25_  (.A(u_multiplier_STAGE3_pp3_48_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_49_2__16_ ),
    .ZN(u_multiplier_pp3_49 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_49_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_49_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_49_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_49_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_49_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_49_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_49_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_49_2__17_ ),
    .ZN(u_multiplier_pp3_50 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_50_1__18_  (.A(u_multiplier_STAGE3_pp3_49_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_50_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_50_1__19_  (.A1(u_multiplier_pp2_50 [1]),
    .A2(u_multiplier_pp2_50 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_50_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_50_1__20_  (.A(u_multiplier_pp2_50 [1]),
    .B(u_multiplier_pp2_50 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_50_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_50_1__21_  (.A1(u_multiplier_pp2_50 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_50_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_50_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_50_1__22_  (.A(u_multiplier_pp2_50 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_50_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_50_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_50_1__23_  (.A1(u_multiplier_pp2_50 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_50_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_50_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_50_1__24_  (.A(u_multiplier_pp2_50 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_50_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_50_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_50_1__25_  (.A(u_multiplier_STAGE3_pp3_49_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_50_1__16_ ),
    .ZN(u_multiplier_pp3_50 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_50_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_50_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_50_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_50_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_50_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_50_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_50_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_50_1__17_ ),
    .ZN(u_multiplier_pp3_51 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_50_2__18_  (.A(u_multiplier_STAGE3_pp3_49_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_50_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_50_2__19_  (.A1(u_multiplier_pp2_50 [5]),
    .A2(u_multiplier_pp2_50 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_50_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_50_2__20_  (.A(u_multiplier_pp2_50 [5]),
    .B(u_multiplier_pp2_50 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_50_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_50_2__21_  (.A1(u_multiplier_pp2_50 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_50_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_50_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_50_2__22_  (.A(u_multiplier_pp2_50 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_50_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_50_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_50_2__23_  (.A1(u_multiplier_pp2_50 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_50_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_50_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_50_2__24_  (.A(u_multiplier_pp2_50 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_50_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_50_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_50_2__25_  (.A(u_multiplier_STAGE3_pp3_49_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_50_2__16_ ),
    .ZN(u_multiplier_pp3_50 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_50_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_50_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_50_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_50_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_50_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_50_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_50_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_50_2__17_ ),
    .ZN(u_multiplier_pp3_51 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_51_1__18_  (.A(u_multiplier_STAGE3_pp3_50_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_51_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_51_1__19_  (.A1(u_multiplier_pp2_51 [1]),
    .A2(u_multiplier_pp2_51 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_51_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_51_1__20_  (.A(u_multiplier_pp2_51 [1]),
    .B(u_multiplier_pp2_51 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_51_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_51_1__21_  (.A1(u_multiplier_pp2_51 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_51_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_51_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_51_1__22_  (.A(u_multiplier_pp2_51 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_51_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_51_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_51_1__23_  (.A1(u_multiplier_pp2_51 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_51_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_51_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_51_1__24_  (.A(u_multiplier_pp2_51 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_51_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_51_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_51_1__25_  (.A(u_multiplier_STAGE3_pp3_50_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_51_1__16_ ),
    .ZN(u_multiplier_pp3_51 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_51_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_51_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_51_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_51_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_51_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_51_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_51_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_51_1__17_ ),
    .ZN(u_multiplier_pp3_52 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_51_2__18_  (.A(u_multiplier_STAGE3_pp3_50_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_51_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_51_2__19_  (.A1(u_multiplier_pp2_51 [5]),
    .A2(u_multiplier_pp2_51 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_51_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_51_2__20_  (.A(u_multiplier_pp2_51 [5]),
    .B(u_multiplier_pp2_51 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_51_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_51_2__21_  (.A1(u_multiplier_pp2_51 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_51_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_51_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_51_2__22_  (.A(u_multiplier_pp2_51 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_51_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_51_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_51_2__23_  (.A1(u_multiplier_pp2_51 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_51_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_51_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_51_2__24_  (.A(u_multiplier_pp2_51 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_51_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_51_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_51_2__25_  (.A(u_multiplier_STAGE3_pp3_50_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_51_2__16_ ),
    .ZN(u_multiplier_pp3_51 [0]));
 NAND2_X2 u_multiplier_STAGE3_E_4_2_pp3_51_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_51_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_51_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_51_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_51_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_51_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_51_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_51_2__17_ ),
    .ZN(u_multiplier_pp3_52 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_52_1__18_  (.A(u_multiplier_STAGE3_pp3_51_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_52_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_52_1__19_  (.A1(u_multiplier_pp2_52 [1]),
    .A2(u_multiplier_pp2_52 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_52_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_52_1__20_  (.A(u_multiplier_pp2_52 [1]),
    .B(u_multiplier_pp2_52 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_52_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_52_1__21_  (.A1(u_multiplier_pp2_52 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_52_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_52_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_52_1__22_  (.A(u_multiplier_pp2_52 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_52_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_52_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_52_1__23_  (.A1(u_multiplier_pp2_52 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_52_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_52_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_52_1__24_  (.A(u_multiplier_pp2_52 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_52_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_52_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_52_1__25_  (.A(u_multiplier_STAGE3_pp3_51_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_52_1__16_ ),
    .ZN(u_multiplier_pp3_52 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_52_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_52_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_52_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_52_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_52_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_52_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_52_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_52_1__17_ ),
    .ZN(u_multiplier_pp3_53 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_52_2__18_  (.A(u_multiplier_STAGE3_pp3_51_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_52_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_52_2__19_  (.A1(u_multiplier_pp2_52 [5]),
    .A2(u_multiplier_pp2_52 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_52_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_52_2__20_  (.A(u_multiplier_pp2_52 [5]),
    .B(u_multiplier_pp2_52 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_52_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_52_2__21_  (.A1(u_multiplier_pp2_52 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_52_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_52_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_52_2__22_  (.A(u_multiplier_pp2_52 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_52_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_52_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_52_2__23_  (.A1(u_multiplier_pp2_52 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_52_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_52_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_52_2__24_  (.A(u_multiplier_pp2_52 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_52_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_52_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_52_2__25_  (.A(u_multiplier_STAGE3_pp3_51_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_52_2__16_ ),
    .ZN(u_multiplier_pp3_52 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_52_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_52_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_52_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_52_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_52_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_52_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_52_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_52_2__17_ ),
    .ZN(u_multiplier_pp3_53 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_53_1__18_  (.A(u_multiplier_STAGE3_pp3_52_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_53_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_53_1__19_  (.A1(u_multiplier_pp2_53 [1]),
    .A2(u_multiplier_pp2_53 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_53_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_53_1__20_  (.A(u_multiplier_pp2_53 [1]),
    .B(u_multiplier_pp2_53 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_53_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_53_1__21_  (.A1(u_multiplier_pp2_53 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_53_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_53_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_53_1__22_  (.A(u_multiplier_pp2_53 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_53_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_53_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_53_1__23_  (.A1(u_multiplier_pp2_53 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_53_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_53_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_53_1__24_  (.A(u_multiplier_pp2_53 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_53_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_53_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_53_1__25_  (.A(u_multiplier_STAGE3_pp3_52_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_53_1__16_ ),
    .ZN(u_multiplier_pp3_53 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_53_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_53_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_53_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_53_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_53_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_53_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_53_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_53_1__17_ ),
    .ZN(u_multiplier_pp3_54 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_53_2__18_  (.A(u_multiplier_STAGE3_pp3_52_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_53_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_53_2__19_  (.A1(u_multiplier_pp2_53 [5]),
    .A2(u_multiplier_pp2_53 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_53_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_53_2__20_  (.A(u_multiplier_pp2_53 [5]),
    .B(u_multiplier_pp2_53 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_53_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_53_2__21_  (.A1(u_multiplier_pp2_53 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_53_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_53_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_53_2__22_  (.A(u_multiplier_pp2_53 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_53_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_53_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_53_2__23_  (.A1(u_multiplier_pp2_53 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_53_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_53_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_53_2__24_  (.A(u_multiplier_pp2_53 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_53_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_53_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_53_2__25_  (.A(u_multiplier_STAGE3_pp3_52_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_53_2__16_ ),
    .ZN(u_multiplier_pp3_53 [0]));
 NAND2_X2 u_multiplier_STAGE3_E_4_2_pp3_53_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_53_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_53_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_53_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_53_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_53_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_53_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_53_2__17_ ),
    .ZN(u_multiplier_pp3_54 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_54_1__18_  (.A(u_multiplier_STAGE3_pp3_53_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_54_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_54_1__19_  (.A1(u_multiplier_pp2_54 [1]),
    .A2(u_multiplier_pp2_54 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_54_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_54_1__20_  (.A(u_multiplier_pp2_54 [1]),
    .B(u_multiplier_pp2_54 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_54_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_54_1__21_  (.A1(u_multiplier_pp2_54 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_54_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_54_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_54_1__22_  (.A(u_multiplier_pp2_54 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_54_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_54_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_54_1__23_  (.A1(u_multiplier_pp2_54 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_54_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_54_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_54_1__24_  (.A(u_multiplier_pp2_54 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_54_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_54_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_54_1__25_  (.A(u_multiplier_STAGE3_pp3_53_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_54_1__16_ ),
    .ZN(u_multiplier_pp3_54 [1]));
 NAND2_X2 u_multiplier_STAGE3_E_4_2_pp3_54_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_54_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_54_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_54_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_54_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_54_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_54_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_54_1__17_ ),
    .ZN(u_multiplier_pp3_55 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_54_2__18_  (.A(u_multiplier_STAGE3_pp3_53_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_54_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_54_2__19_  (.A1(u_multiplier_pp2_54 [5]),
    .A2(u_multiplier_pp2_54 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_54_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_54_2__20_  (.A(u_multiplier_pp2_54 [5]),
    .B(u_multiplier_pp2_54 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_54_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_54_2__21_  (.A1(u_multiplier_pp2_54 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_54_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_54_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_54_2__22_  (.A(u_multiplier_pp2_54 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_54_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_54_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_54_2__23_  (.A1(u_multiplier_pp2_54 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_54_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_54_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_54_2__24_  (.A(u_multiplier_pp2_54 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_54_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_54_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_54_2__25_  (.A(u_multiplier_STAGE3_pp3_53_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_54_2__16_ ),
    .ZN(u_multiplier_pp3_54 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_54_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_54_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_54_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_54_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_54_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_54_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_54_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_54_2__17_ ),
    .ZN(u_multiplier_pp3_55 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_55_1__18_  (.A(u_multiplier_STAGE3_pp3_54_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_55_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_55_1__19_  (.A1(u_multiplier_pp2_55 [1]),
    .A2(u_multiplier_pp2_55 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_55_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_55_1__20_  (.A(u_multiplier_pp2_55 [1]),
    .B(u_multiplier_pp2_55 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_55_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_55_1__21_  (.A1(u_multiplier_pp2_55 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_55_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_55_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_55_1__22_  (.A(u_multiplier_pp2_55 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_55_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_55_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_55_1__23_  (.A1(u_multiplier_pp2_55 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_55_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_55_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_55_1__24_  (.A(u_multiplier_pp2_55 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_55_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_55_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_55_1__25_  (.A(u_multiplier_STAGE3_pp3_54_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_55_1__16_ ),
    .ZN(u_multiplier_pp3_55 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_55_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_55_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_55_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_55_e42_1_cout ));
 OAI21_X1 u_multiplier_STAGE3_E_4_2_pp3_55_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_55_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_55_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_55_1__17_ ),
    .ZN(u_multiplier_pp3_56 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_55_2__18_  (.A(u_multiplier_STAGE3_pp3_54_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_55_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_55_2__19_  (.A1(u_multiplier_pp2_55 [5]),
    .A2(u_multiplier_pp2_55 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_55_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_55_2__20_  (.A(u_multiplier_pp2_55 [5]),
    .B(u_multiplier_pp2_55 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_55_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_55_2__21_  (.A1(u_multiplier_pp2_55 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_55_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_55_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_55_2__22_  (.A(u_multiplier_pp2_55 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_55_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_55_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_55_2__23_  (.A1(u_multiplier_pp2_55 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_55_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_55_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_55_2__24_  (.A(u_multiplier_pp2_55 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_55_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_55_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_55_2__25_  (.A(u_multiplier_STAGE3_pp3_54_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_55_2__16_ ),
    .ZN(u_multiplier_pp3_55 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_55_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_55_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_55_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_55_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_55_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_55_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_55_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_55_2__17_ ),
    .ZN(u_multiplier_pp3_56 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_56_1__18_  (.A(u_multiplier_STAGE3_pp3_55_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_56_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_56_1__19_  (.A1(u_multiplier_pp2_56 [1]),
    .A2(u_multiplier_pp2_56 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_56_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_56_1__20_  (.A(u_multiplier_pp2_56 [1]),
    .B(u_multiplier_pp2_56 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_56_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_56_1__21_  (.A1(u_multiplier_pp2_56 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_56_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_56_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_56_1__22_  (.A(u_multiplier_pp2_56 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_56_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_56_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_56_1__23_  (.A1(u_multiplier_pp2_56 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_56_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_56_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_56_1__24_  (.A(u_multiplier_pp2_56 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_56_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_56_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_56_1__25_  (.A(u_multiplier_STAGE3_pp3_55_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_56_1__16_ ),
    .ZN(u_multiplier_pp3_56 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_56_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_56_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_56_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_56_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_56_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_56_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_56_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_56_1__17_ ),
    .ZN(u_multiplier_pp3_57 [3]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_56_2__18_  (.A(u_multiplier_STAGE3_pp3_55_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_56_2__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_56_2__19_  (.A1(u_multiplier_pp2_56 [5]),
    .A2(u_multiplier_pp2_56 [4]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_56_2__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_56_2__20_  (.A(u_multiplier_pp2_56 [5]),
    .B(u_multiplier_pp2_56 [4]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_56_2__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_56_2__21_  (.A1(u_multiplier_pp2_56 [6]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_56_2__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_56_2__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_56_2__22_  (.A(u_multiplier_pp2_56 [6]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_56_2__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_56_2__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_56_2__23_  (.A1(u_multiplier_pp2_56 [7]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_56_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_56_2__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_56_2__24_  (.A(u_multiplier_pp2_56 [7]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_56_2__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_56_2__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_56_2__25_  (.A(u_multiplier_STAGE3_pp3_55_e42_2_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_56_2__16_ ),
    .ZN(u_multiplier_pp3_56 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_56_2__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_56_2__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_56_2__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_56_e42_2_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_56_2__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_56_2__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_56_2__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_56_2__17_ ),
    .ZN(u_multiplier_pp3_57 [2]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_57_1__18_  (.A(u_multiplier_STAGE3_pp3_56_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_57_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_57_1__19_  (.A1(u_multiplier_pp2_57 [1]),
    .A2(u_multiplier_pp2_57 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_57_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_57_1__20_  (.A(u_multiplier_pp2_57 [1]),
    .B(u_multiplier_pp2_57 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_57_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_57_1__21_  (.A1(u_multiplier_pp2_57 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_57_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_57_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_57_1__22_  (.A(u_multiplier_pp2_57 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_57_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_57_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_57_1__23_  (.A1(u_multiplier_pp2_57 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_57_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_57_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_57_1__24_  (.A(u_multiplier_pp2_57 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_57_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_57_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_57_1__25_  (.A(u_multiplier_STAGE3_pp3_56_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_57_1__16_ ),
    .ZN(u_multiplier_pp3_57 [1]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_57_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_57_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_57_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_57_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_57_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_57_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_57_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_57_1__17_ ),
    .ZN(u_multiplier_pp3_58 [1]));
 INV_X1 u_multiplier_STAGE3_E_4_2_pp3_58_1__18_  (.A(u_multiplier_STAGE3_pp3_57_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_58_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_58_1__19_  (.A1(u_multiplier_pp2_58 [1]),
    .A2(u_multiplier_pp2_58 [0]),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_58_1__11_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_58_1__20_  (.A(u_multiplier_pp2_58 [1]),
    .B(u_multiplier_pp2_58 [0]),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_58_1__12_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_58_1__21_  (.A1(u_multiplier_pp2_58 [2]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_58_1__12_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_58_1__13_ ));
 XOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_58_1__22_  (.A(u_multiplier_pp2_58 [2]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_58_1__12_ ),
    .Z(u_multiplier_STAGE3_E_4_2_pp3_58_1__14_ ));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_58_1__23_  (.A1(u_multiplier_pp2_58 [3]),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_58_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_58_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_58_1__24_  (.A(u_multiplier_pp2_58 [3]),
    .B(u_multiplier_STAGE3_E_4_2_pp3_58_1__14_ ),
    .ZN(u_multiplier_STAGE3_E_4_2_pp3_58_1__16_ ));
 XNOR2_X2 u_multiplier_STAGE3_E_4_2_pp3_58_1__25_  (.A(u_multiplier_STAGE3_pp3_57_e42_1_cout ),
    .B(u_multiplier_STAGE3_E_4_2_pp3_58_1__16_ ),
    .ZN(u_multiplier_pp3_58 [0]));
 NAND2_X1 u_multiplier_STAGE3_E_4_2_pp3_58_1__26_  (.A1(u_multiplier_STAGE3_E_4_2_pp3_58_1__11_ ),
    .A2(u_multiplier_STAGE3_E_4_2_pp3_58_1__13_ ),
    .ZN(u_multiplier_STAGE3_pp3_58_e42_1_cout ));
 OAI21_X2 u_multiplier_STAGE3_E_4_2_pp3_58_1__27_  (.A(u_multiplier_STAGE3_E_4_2_pp3_58_1__15_ ),
    .B1(u_multiplier_STAGE3_E_4_2_pp3_58_1__16_ ),
    .B2(u_multiplier_STAGE3_E_4_2_pp3_58_1__17_ ),
    .ZN(u_multiplier_pp3_59 [1]));
 INV_X1 u_multiplier_STAGE3_Full_adder_pp3_57_1__12_  (.A(u_multiplier_STAGE3_pp3_56_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_Full_adder_pp3_57_1__08_ ));
 NAND3_X2 u_multiplier_STAGE3_Full_adder_pp3_57_1__13_  (.A1(u_multiplier_pp2_57 [5]),
    .A2(u_multiplier_pp2_57 [4]),
    .A3(u_multiplier_STAGE3_pp3_56_e42_2_cout ),
    .ZN(u_multiplier_STAGE3_Full_adder_pp3_57_1__09_ ));
 NOR2_X2 u_multiplier_STAGE3_Full_adder_pp3_57_1__14_  (.A1(u_multiplier_pp2_57 [5]),
    .A2(u_multiplier_pp2_57 [4]),
    .ZN(u_multiplier_STAGE3_Full_adder_pp3_57_1__10_ ));
 AOI21_X1 u_multiplier_STAGE3_Full_adder_pp3_57_1__15_  (.A(u_multiplier_STAGE3_pp3_56_e42_2_cout ),
    .B1(u_multiplier_pp2_57 [4]),
    .B2(u_multiplier_pp2_57 [5]),
    .ZN(u_multiplier_STAGE3_Full_adder_pp3_57_1__11_ ));
 NOR2_X2 u_multiplier_STAGE3_Full_adder_pp3_57_1__16_  (.A1(u_multiplier_STAGE3_Full_adder_pp3_57_1__10_ ),
    .A2(u_multiplier_STAGE3_Full_adder_pp3_57_1__11_ ),
    .ZN(u_multiplier_pp3_58 [2]));
 AOI22_X4 u_multiplier_STAGE3_Full_adder_pp3_57_1__17_  (.A1(u_multiplier_STAGE3_Full_adder_pp3_57_1__08_ ),
    .A2(u_multiplier_STAGE3_Full_adder_pp3_57_1__10_ ),
    .B1(u_multiplier_pp3_58 [2]),
    .B2(u_multiplier_STAGE3_Full_adder_pp3_57_1__09_ ),
    .ZN(u_multiplier_pp3_57 [0]));
 INV_X1 u_multiplier_STAGE3_Full_adder_pp3_59_1__12_  (.A(u_multiplier_STAGE3_pp3_58_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_Full_adder_pp3_59_1__08_ ));
 NAND3_X1 u_multiplier_STAGE3_Full_adder_pp3_59_1__13_  (.A1(u_multiplier_pp2_59 [1]),
    .A2(u_multiplier_pp2_59 [0]),
    .A3(u_multiplier_STAGE3_pp3_58_e42_1_cout ),
    .ZN(u_multiplier_STAGE3_Full_adder_pp3_59_1__09_ ));
 NOR2_X2 u_multiplier_STAGE3_Full_adder_pp3_59_1__14_  (.A1(u_multiplier_pp2_59 [1]),
    .A2(u_multiplier_pp2_59 [0]),
    .ZN(u_multiplier_STAGE3_Full_adder_pp3_59_1__10_ ));
 AOI21_X1 u_multiplier_STAGE3_Full_adder_pp3_59_1__15_  (.A(u_multiplier_STAGE3_pp3_58_e42_1_cout ),
    .B1(u_multiplier_pp2_59 [0]),
    .B2(u_multiplier_pp2_59 [1]),
    .ZN(u_multiplier_STAGE3_Full_adder_pp3_59_1__11_ ));
 NOR2_X2 u_multiplier_STAGE3_Full_adder_pp3_59_1__16_  (.A1(u_multiplier_STAGE3_Full_adder_pp3_59_1__10_ ),
    .A2(u_multiplier_STAGE3_Full_adder_pp3_59_1__11_ ),
    .ZN(u_multiplier_pp3_60 [0]));
 AOI22_X2 u_multiplier_STAGE3_Full_adder_pp3_59_1__17_  (.A1(u_multiplier_STAGE3_Full_adder_pp3_59_1__08_ ),
    .A2(u_multiplier_STAGE3_Full_adder_pp3_59_1__10_ ),
    .B1(u_multiplier_pp3_60 [0]),
    .B2(u_multiplier_STAGE3_Full_adder_pp3_59_1__09_ ),
    .ZN(u_multiplier_pp3_59 [0]));
 AND2_X1 u_multiplier_STAGE3_Half_adder_pp3_4__4_  (.A1(u_multiplier_pp2_4 [4]),
    .A2(u_multiplier_pp2_4 [3]),
    .ZN(u_multiplier_pp3_5 [1]));
 XOR2_X2 u_multiplier_STAGE3_Half_adder_pp3_4__5_  (.A(u_multiplier_pp2_4 [4]),
    .B(u_multiplier_pp2_4 [3]),
    .Z(u_multiplier_pp3_4 [0]));
 AND2_X1 u_multiplier_STAGE3_Half_adder_pp3_6__4_  (.A1(u_multiplier_pp2_6 [2]),
    .A2(u_multiplier_pp2_6 [1]),
    .ZN(u_multiplier_pp3_7 [2]));
 XOR2_X2 u_multiplier_STAGE3_Half_adder_pp3_6__5_  (.A(u_multiplier_pp2_6 [2]),
    .B(u_multiplier_pp2_6 [1]),
    .Z(u_multiplier_pp3_6 [1]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_10_0__21_  (.A1(u_multiplier_pp2_10 [5]),
    .A2(u_multiplier_pp2_10 [4]),
    .A3(u_multiplier_pp2_10 [6]),
    .ZN(u_multiplier_STAGE3_acci_pp3_10_0__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_10_0__22_  (.A(u_multiplier_pp2_10 [5]),
    .B(u_multiplier_pp2_10 [4]),
    .Z(u_multiplier_STAGE3_acci_pp3_10_0__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_10_0__23_  (.A(u_multiplier_pp2_10 [6]),
    .B(u_multiplier_pp2_10 [7]),
    .Z(u_multiplier_STAGE3_acci_pp3_10_0__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_10_0__24_  (.A1(u_multiplier_STAGE3_acci_pp3_10_0__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_10_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_10_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_10_0__25_  (.A(u_multiplier_STAGE3_acci_pp3_10_0__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_10_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_10_0__16_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_10_0__26_  (.A1(u_multiplier_STAGE3_acci_pp3_10_0__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_10_0__16_ ),
    .ZN(u_multiplier_pp3_10 [0]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_10_0__27_  (.A1(u_multiplier_pp2_10 [5]),
    .A2(u_multiplier_pp2_10 [4]),
    .B1(u_multiplier_pp2_10 [6]),
    .B2(u_multiplier_pp2_10 [7]),
    .ZN(u_multiplier_STAGE3_acci_pp3_10_0__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_10_0__28_  (.A1(u_multiplier_STAGE3_acci_pp3_10_0__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_10_0__17_ ),
    .ZN(u_multiplier_pp3_11 [3]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_10_1__21_  (.A1(u_multiplier_pp2_10 [1]),
    .A2(u_multiplier_pp2_10 [0]),
    .A3(u_multiplier_pp2_10 [2]),
    .ZN(u_multiplier_STAGE3_acci_pp3_10_1__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_10_1__22_  (.A(u_multiplier_pp2_10 [1]),
    .B(u_multiplier_pp2_10 [0]),
    .Z(u_multiplier_STAGE3_acci_pp3_10_1__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_10_1__23_  (.A(u_multiplier_pp2_10 [2]),
    .B(u_multiplier_pp2_10 [3]),
    .Z(u_multiplier_STAGE3_acci_pp3_10_1__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_10_1__24_  (.A1(u_multiplier_STAGE3_acci_pp3_10_1__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_10_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_10_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_10_1__25_  (.A(u_multiplier_STAGE3_acci_pp3_10_1__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_10_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_10_1__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_10_1__26_  (.A1(u_multiplier_STAGE3_acci_pp3_10_1__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_10_1__16_ ),
    .ZN(u_multiplier_pp3_10 [1]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_10_1__27_  (.A1(u_multiplier_pp2_10 [1]),
    .A2(u_multiplier_pp2_10 [0]),
    .B1(u_multiplier_pp2_10 [2]),
    .B2(u_multiplier_pp2_10 [3]),
    .ZN(u_multiplier_STAGE3_acci_pp3_10_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_10_1__28_  (.A1(u_multiplier_STAGE3_acci_pp3_10_1__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_10_1__17_ ),
    .ZN(u_multiplier_pp3_11 [2]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_11_0__21_  (.A1(u_multiplier_pp2_11 [5]),
    .A2(u_multiplier_pp2_11 [4]),
    .A3(u_multiplier_pp2_11 [6]),
    .ZN(u_multiplier_STAGE3_acci_pp3_11_0__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_11_0__22_  (.A(u_multiplier_pp2_11 [5]),
    .B(u_multiplier_pp2_11 [4]),
    .Z(u_multiplier_STAGE3_acci_pp3_11_0__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_11_0__23_  (.A(u_multiplier_pp2_11 [6]),
    .B(u_multiplier_pp2_11 [7]),
    .Z(u_multiplier_STAGE3_acci_pp3_11_0__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_11_0__24_  (.A1(u_multiplier_STAGE3_acci_pp3_11_0__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_11_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_11_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_11_0__25_  (.A(u_multiplier_STAGE3_acci_pp3_11_0__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_11_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_11_0__16_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_11_0__26_  (.A1(u_multiplier_STAGE3_acci_pp3_11_0__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_11_0__16_ ),
    .ZN(u_multiplier_pp3_11 [0]));
 AOI22_X2 u_multiplier_STAGE3_acci_pp3_11_0__27_  (.A1(u_multiplier_pp2_11 [5]),
    .A2(u_multiplier_pp2_11 [4]),
    .B1(u_multiplier_pp2_11 [6]),
    .B2(u_multiplier_pp2_11 [7]),
    .ZN(u_multiplier_STAGE3_acci_pp3_11_0__17_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_11_0__28_  (.A1(u_multiplier_STAGE3_acci_pp3_11_0__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_11_0__17_ ),
    .ZN(u_multiplier_pp3_12 [3]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_11_1__21_  (.A1(u_multiplier_pp2_11 [1]),
    .A2(u_multiplier_pp2_11 [0]),
    .A3(u_multiplier_pp2_11 [2]),
    .ZN(u_multiplier_STAGE3_acci_pp3_11_1__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_11_1__22_  (.A(u_multiplier_pp2_11 [1]),
    .B(u_multiplier_pp2_11 [0]),
    .Z(u_multiplier_STAGE3_acci_pp3_11_1__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_11_1__23_  (.A(u_multiplier_pp2_11 [2]),
    .B(u_multiplier_pp2_11 [3]),
    .Z(u_multiplier_STAGE3_acci_pp3_11_1__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_11_1__24_  (.A1(u_multiplier_STAGE3_acci_pp3_11_1__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_11_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_11_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_11_1__25_  (.A(u_multiplier_STAGE3_acci_pp3_11_1__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_11_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_11_1__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_11_1__26_  (.A1(u_multiplier_STAGE3_acci_pp3_11_1__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_11_1__16_ ),
    .ZN(u_multiplier_pp3_11 [1]));
 AOI22_X2 u_multiplier_STAGE3_acci_pp3_11_1__27_  (.A1(u_multiplier_pp2_11 [1]),
    .A2(u_multiplier_pp2_11 [0]),
    .B1(u_multiplier_pp2_11 [2]),
    .B2(u_multiplier_pp2_11 [3]),
    .ZN(u_multiplier_STAGE3_acci_pp3_11_1__17_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_11_1__28_  (.A1(u_multiplier_STAGE3_acci_pp3_11_1__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_11_1__17_ ),
    .ZN(u_multiplier_pp3_12 [2]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_12_0__21_  (.A1(u_multiplier_pp2_12 [5]),
    .A2(u_multiplier_pp2_12 [4]),
    .A3(u_multiplier_pp2_12 [6]),
    .ZN(u_multiplier_STAGE3_acci_pp3_12_0__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_12_0__22_  (.A(u_multiplier_pp2_12 [5]),
    .B(u_multiplier_pp2_12 [4]),
    .Z(u_multiplier_STAGE3_acci_pp3_12_0__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_12_0__23_  (.A(u_multiplier_pp2_12 [6]),
    .B(u_multiplier_pp2_12 [7]),
    .Z(u_multiplier_STAGE3_acci_pp3_12_0__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_12_0__24_  (.A1(u_multiplier_STAGE3_acci_pp3_12_0__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_12_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_12_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_12_0__25_  (.A(u_multiplier_STAGE3_acci_pp3_12_0__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_12_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_12_0__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_12_0__26_  (.A1(u_multiplier_STAGE3_acci_pp3_12_0__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_12_0__16_ ),
    .ZN(u_multiplier_pp3_12 [0]));
 AOI22_X2 u_multiplier_STAGE3_acci_pp3_12_0__27_  (.A1(u_multiplier_pp2_12 [5]),
    .A2(u_multiplier_pp2_12 [4]),
    .B1(u_multiplier_pp2_12 [6]),
    .B2(u_multiplier_pp2_12 [7]),
    .ZN(u_multiplier_STAGE3_acci_pp3_12_0__17_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_12_0__28_  (.A1(u_multiplier_STAGE3_acci_pp3_12_0__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_12_0__17_ ),
    .ZN(u_multiplier_pp3_13 [3]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_12_1__21_  (.A1(u_multiplier_pp2_12 [1]),
    .A2(u_multiplier_pp2_12 [0]),
    .A3(u_multiplier_pp2_12 [2]),
    .ZN(u_multiplier_STAGE3_acci_pp3_12_1__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_12_1__22_  (.A(u_multiplier_pp2_12 [1]),
    .B(u_multiplier_pp2_12 [0]),
    .Z(u_multiplier_STAGE3_acci_pp3_12_1__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_12_1__23_  (.A(u_multiplier_pp2_12 [2]),
    .B(u_multiplier_pp2_12 [3]),
    .Z(u_multiplier_STAGE3_acci_pp3_12_1__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_12_1__24_  (.A1(u_multiplier_STAGE3_acci_pp3_12_1__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_12_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_12_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_12_1__25_  (.A(u_multiplier_STAGE3_acci_pp3_12_1__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_12_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_12_1__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_12_1__26_  (.A1(u_multiplier_STAGE3_acci_pp3_12_1__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_12_1__16_ ),
    .ZN(u_multiplier_pp3_12 [1]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_12_1__27_  (.A1(u_multiplier_pp2_12 [1]),
    .A2(u_multiplier_pp2_12 [0]),
    .B1(u_multiplier_pp2_12 [2]),
    .B2(u_multiplier_pp2_12 [3]),
    .ZN(u_multiplier_STAGE3_acci_pp3_12_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_12_1__28_  (.A1(u_multiplier_STAGE3_acci_pp3_12_1__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_12_1__17_ ),
    .ZN(u_multiplier_pp3_13 [2]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_13_0__21_  (.A1(u_multiplier_pp2_13 [5]),
    .A2(u_multiplier_pp2_13 [4]),
    .A3(u_multiplier_pp2_13 [6]),
    .ZN(u_multiplier_STAGE3_acci_pp3_13_0__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_13_0__22_  (.A(u_multiplier_pp2_13 [5]),
    .B(u_multiplier_pp2_13 [4]),
    .Z(u_multiplier_STAGE3_acci_pp3_13_0__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_13_0__23_  (.A(u_multiplier_pp2_13 [6]),
    .B(u_multiplier_pp2_13 [7]),
    .Z(u_multiplier_STAGE3_acci_pp3_13_0__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_13_0__24_  (.A1(u_multiplier_STAGE3_acci_pp3_13_0__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_13_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_13_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_13_0__25_  (.A(u_multiplier_STAGE3_acci_pp3_13_0__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_13_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_13_0__16_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_13_0__26_  (.A1(u_multiplier_STAGE3_acci_pp3_13_0__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_13_0__16_ ),
    .ZN(u_multiplier_pp3_13 [0]));
 AOI22_X2 u_multiplier_STAGE3_acci_pp3_13_0__27_  (.A1(u_multiplier_pp2_13 [5]),
    .A2(u_multiplier_pp2_13 [4]),
    .B1(u_multiplier_pp2_13 [6]),
    .B2(u_multiplier_pp2_13 [7]),
    .ZN(u_multiplier_STAGE3_acci_pp3_13_0__17_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_13_0__28_  (.A1(u_multiplier_STAGE3_acci_pp3_13_0__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_13_0__17_ ),
    .ZN(u_multiplier_pp3_14 [3]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_13_1__21_  (.A1(u_multiplier_pp2_13 [1]),
    .A2(u_multiplier_pp2_13 [0]),
    .A3(u_multiplier_pp2_13 [2]),
    .ZN(u_multiplier_STAGE3_acci_pp3_13_1__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_13_1__22_  (.A(u_multiplier_pp2_13 [1]),
    .B(u_multiplier_pp2_13 [0]),
    .Z(u_multiplier_STAGE3_acci_pp3_13_1__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_13_1__23_  (.A(u_multiplier_pp2_13 [2]),
    .B(u_multiplier_pp2_13 [3]),
    .Z(u_multiplier_STAGE3_acci_pp3_13_1__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_13_1__24_  (.A1(u_multiplier_STAGE3_acci_pp3_13_1__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_13_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_13_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_13_1__25_  (.A(u_multiplier_STAGE3_acci_pp3_13_1__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_13_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_13_1__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_13_1__26_  (.A1(u_multiplier_STAGE3_acci_pp3_13_1__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_13_1__16_ ),
    .ZN(u_multiplier_pp3_13 [1]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_13_1__27_  (.A1(u_multiplier_pp2_13 [1]),
    .A2(u_multiplier_pp2_13 [0]),
    .B1(u_multiplier_pp2_13 [2]),
    .B2(u_multiplier_pp2_13 [3]),
    .ZN(u_multiplier_STAGE3_acci_pp3_13_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_13_1__28_  (.A1(u_multiplier_STAGE3_acci_pp3_13_1__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_13_1__17_ ),
    .ZN(u_multiplier_pp3_14 [2]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_14_0__21_  (.A1(u_multiplier_pp2_14 [5]),
    .A2(u_multiplier_pp2_14 [4]),
    .A3(u_multiplier_pp2_14 [6]),
    .ZN(u_multiplier_STAGE3_acci_pp3_14_0__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_14_0__22_  (.A(u_multiplier_pp2_14 [5]),
    .B(u_multiplier_pp2_14 [4]),
    .Z(u_multiplier_STAGE3_acci_pp3_14_0__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_14_0__23_  (.A(u_multiplier_pp2_14 [6]),
    .B(u_multiplier_pp2_14 [7]),
    .Z(u_multiplier_STAGE3_acci_pp3_14_0__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_14_0__24_  (.A1(u_multiplier_STAGE3_acci_pp3_14_0__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_14_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_14_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_14_0__25_  (.A(u_multiplier_STAGE3_acci_pp3_14_0__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_14_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_14_0__16_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_14_0__26_  (.A1(u_multiplier_STAGE3_acci_pp3_14_0__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_14_0__16_ ),
    .ZN(u_multiplier_pp3_14 [0]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_14_0__27_  (.A1(u_multiplier_pp2_14 [5]),
    .A2(u_multiplier_pp2_14 [4]),
    .B1(u_multiplier_pp2_14 [6]),
    .B2(u_multiplier_pp2_14 [7]),
    .ZN(u_multiplier_STAGE3_acci_pp3_14_0__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_14_0__28_  (.A1(u_multiplier_STAGE3_acci_pp3_14_0__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_14_0__17_ ),
    .ZN(u_multiplier_pp3_15 [3]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_14_1__21_  (.A1(u_multiplier_pp2_14 [1]),
    .A2(u_multiplier_pp2_14 [0]),
    .A3(u_multiplier_pp2_14 [2]),
    .ZN(u_multiplier_STAGE3_acci_pp3_14_1__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_14_1__22_  (.A(u_multiplier_pp2_14 [1]),
    .B(u_multiplier_pp2_14 [0]),
    .Z(u_multiplier_STAGE3_acci_pp3_14_1__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_14_1__23_  (.A(u_multiplier_pp2_14 [2]),
    .B(u_multiplier_pp2_14 [3]),
    .Z(u_multiplier_STAGE3_acci_pp3_14_1__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_14_1__24_  (.A1(u_multiplier_STAGE3_acci_pp3_14_1__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_14_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_14_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_14_1__25_  (.A(u_multiplier_STAGE3_acci_pp3_14_1__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_14_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_14_1__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_14_1__26_  (.A1(u_multiplier_STAGE3_acci_pp3_14_1__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_14_1__16_ ),
    .ZN(u_multiplier_pp3_14 [1]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_14_1__27_  (.A1(u_multiplier_pp2_14 [1]),
    .A2(u_multiplier_pp2_14 [0]),
    .B1(u_multiplier_pp2_14 [2]),
    .B2(u_multiplier_pp2_14 [3]),
    .ZN(u_multiplier_STAGE3_acci_pp3_14_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_14_1__28_  (.A1(u_multiplier_STAGE3_acci_pp3_14_1__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_14_1__17_ ),
    .ZN(u_multiplier_pp3_15 [2]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_15_0__21_  (.A1(u_multiplier_pp2_15 [5]),
    .A2(u_multiplier_pp2_15 [4]),
    .A3(u_multiplier_pp2_15 [6]),
    .ZN(u_multiplier_STAGE3_acci_pp3_15_0__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_15_0__22_  (.A(u_multiplier_pp2_15 [5]),
    .B(u_multiplier_pp2_15 [4]),
    .Z(u_multiplier_STAGE3_acci_pp3_15_0__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_15_0__23_  (.A(u_multiplier_pp2_15 [6]),
    .B(u_multiplier_pp2_15 [7]),
    .Z(u_multiplier_STAGE3_acci_pp3_15_0__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_15_0__24_  (.A1(u_multiplier_STAGE3_acci_pp3_15_0__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_15_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_15_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_15_0__25_  (.A(u_multiplier_STAGE3_acci_pp3_15_0__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_15_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_15_0__16_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_15_0__26_  (.A1(u_multiplier_STAGE3_acci_pp3_15_0__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_15_0__16_ ),
    .ZN(u_multiplier_pp3_15 [0]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_15_0__27_  (.A1(u_multiplier_pp2_15 [5]),
    .A2(u_multiplier_pp2_15 [4]),
    .B1(u_multiplier_pp2_15 [6]),
    .B2(u_multiplier_pp2_15 [7]),
    .ZN(u_multiplier_STAGE3_acci_pp3_15_0__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_15_0__28_  (.A1(u_multiplier_STAGE3_acci_pp3_15_0__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_15_0__17_ ),
    .ZN(u_multiplier_pp3_16 [3]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_15_1__21_  (.A1(u_multiplier_pp2_15 [1]),
    .A2(u_multiplier_pp2_15 [0]),
    .A3(u_multiplier_pp2_15 [2]),
    .ZN(u_multiplier_STAGE3_acci_pp3_15_1__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_15_1__22_  (.A(u_multiplier_pp2_15 [1]),
    .B(u_multiplier_pp2_15 [0]),
    .Z(u_multiplier_STAGE3_acci_pp3_15_1__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_15_1__23_  (.A(u_multiplier_pp2_15 [2]),
    .B(u_multiplier_pp2_15 [3]),
    .Z(u_multiplier_STAGE3_acci_pp3_15_1__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_15_1__24_  (.A1(u_multiplier_STAGE3_acci_pp3_15_1__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_15_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_15_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_15_1__25_  (.A(u_multiplier_STAGE3_acci_pp3_15_1__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_15_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_15_1__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_15_1__26_  (.A1(u_multiplier_STAGE3_acci_pp3_15_1__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_15_1__16_ ),
    .ZN(u_multiplier_pp3_15 [1]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_15_1__27_  (.A1(u_multiplier_pp2_15 [1]),
    .A2(u_multiplier_pp2_15 [0]),
    .B1(u_multiplier_pp2_15 [2]),
    .B2(u_multiplier_pp2_15 [3]),
    .ZN(u_multiplier_STAGE3_acci_pp3_15_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_15_1__28_  (.A1(u_multiplier_STAGE3_acci_pp3_15_1__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_15_1__17_ ),
    .ZN(u_multiplier_pp3_16 [2]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_16_0__21_  (.A1(u_multiplier_pp2_16 [5]),
    .A2(u_multiplier_pp2_16 [4]),
    .A3(u_multiplier_pp2_16 [6]),
    .ZN(u_multiplier_STAGE3_acci_pp3_16_0__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_16_0__22_  (.A(u_multiplier_pp2_16 [5]),
    .B(u_multiplier_pp2_16 [4]),
    .Z(u_multiplier_STAGE3_acci_pp3_16_0__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_16_0__23_  (.A(u_multiplier_pp2_16 [6]),
    .B(u_multiplier_pp2_16 [7]),
    .Z(u_multiplier_STAGE3_acci_pp3_16_0__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_16_0__24_  (.A1(u_multiplier_STAGE3_acci_pp3_16_0__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_16_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_16_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_16_0__25_  (.A(u_multiplier_STAGE3_acci_pp3_16_0__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_16_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_16_0__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_16_0__26_  (.A1(u_multiplier_STAGE3_acci_pp3_16_0__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_16_0__16_ ),
    .ZN(u_multiplier_pp3_16 [0]));
 AOI22_X2 u_multiplier_STAGE3_acci_pp3_16_0__27_  (.A1(u_multiplier_pp2_16 [5]),
    .A2(u_multiplier_pp2_16 [4]),
    .B1(u_multiplier_pp2_16 [6]),
    .B2(u_multiplier_pp2_16 [7]),
    .ZN(u_multiplier_STAGE3_acci_pp3_16_0__17_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_16_0__28_  (.A1(u_multiplier_STAGE3_acci_pp3_16_0__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_16_0__17_ ),
    .ZN(u_multiplier_pp3_17 [3]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_16_1__21_  (.A1(u_multiplier_pp2_16 [1]),
    .A2(u_multiplier_pp2_16 [0]),
    .A3(u_multiplier_pp2_16 [2]),
    .ZN(u_multiplier_STAGE3_acci_pp3_16_1__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_16_1__22_  (.A(u_multiplier_pp2_16 [1]),
    .B(u_multiplier_pp2_16 [0]),
    .Z(u_multiplier_STAGE3_acci_pp3_16_1__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_16_1__23_  (.A(u_multiplier_pp2_16 [2]),
    .B(u_multiplier_pp2_16 [3]),
    .Z(u_multiplier_STAGE3_acci_pp3_16_1__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_16_1__24_  (.A1(u_multiplier_STAGE3_acci_pp3_16_1__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_16_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_16_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_16_1__25_  (.A(u_multiplier_STAGE3_acci_pp3_16_1__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_16_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_16_1__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_16_1__26_  (.A1(u_multiplier_STAGE3_acci_pp3_16_1__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_16_1__16_ ),
    .ZN(u_multiplier_pp3_16 [1]));
 AOI22_X2 u_multiplier_STAGE3_acci_pp3_16_1__27_  (.A1(u_multiplier_pp2_16 [1]),
    .A2(u_multiplier_pp2_16 [0]),
    .B1(u_multiplier_pp2_16 [2]),
    .B2(u_multiplier_pp2_16 [3]),
    .ZN(u_multiplier_STAGE3_acci_pp3_16_1__17_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_16_1__28_  (.A1(u_multiplier_STAGE3_acci_pp3_16_1__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_16_1__17_ ),
    .ZN(u_multiplier_pp3_17 [2]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_17_0__21_  (.A1(u_multiplier_pp2_17 [5]),
    .A2(u_multiplier_pp2_17 [4]),
    .A3(u_multiplier_pp2_17 [6]),
    .ZN(u_multiplier_STAGE3_acci_pp3_17_0__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_17_0__22_  (.A(u_multiplier_pp2_17 [5]),
    .B(u_multiplier_pp2_17 [4]),
    .Z(u_multiplier_STAGE3_acci_pp3_17_0__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_17_0__23_  (.A(u_multiplier_pp2_17 [6]),
    .B(u_multiplier_pp2_17 [7]),
    .Z(u_multiplier_STAGE3_acci_pp3_17_0__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_17_0__24_  (.A1(u_multiplier_STAGE3_acci_pp3_17_0__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_17_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_17_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_17_0__25_  (.A(u_multiplier_STAGE3_acci_pp3_17_0__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_17_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_17_0__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_17_0__26_  (.A1(u_multiplier_STAGE3_acci_pp3_17_0__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_17_0__16_ ),
    .ZN(u_multiplier_pp3_17 [0]));
 AOI22_X2 u_multiplier_STAGE3_acci_pp3_17_0__27_  (.A1(u_multiplier_pp2_17 [5]),
    .A2(u_multiplier_pp2_17 [4]),
    .B1(u_multiplier_pp2_17 [6]),
    .B2(u_multiplier_pp2_17 [7]),
    .ZN(u_multiplier_STAGE3_acci_pp3_17_0__17_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_17_0__28_  (.A1(u_multiplier_STAGE3_acci_pp3_17_0__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_17_0__17_ ),
    .ZN(u_multiplier_pp3_18 [3]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_17_1__21_  (.A1(u_multiplier_pp2_17 [1]),
    .A2(u_multiplier_pp2_17 [0]),
    .A3(u_multiplier_pp2_17 [2]),
    .ZN(u_multiplier_STAGE3_acci_pp3_17_1__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_17_1__22_  (.A(u_multiplier_pp2_17 [1]),
    .B(u_multiplier_pp2_17 [0]),
    .Z(u_multiplier_STAGE3_acci_pp3_17_1__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_17_1__23_  (.A(u_multiplier_pp2_17 [2]),
    .B(u_multiplier_pp2_17 [3]),
    .Z(u_multiplier_STAGE3_acci_pp3_17_1__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_17_1__24_  (.A1(u_multiplier_STAGE3_acci_pp3_17_1__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_17_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_17_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_17_1__25_  (.A(u_multiplier_STAGE3_acci_pp3_17_1__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_17_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_17_1__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_17_1__26_  (.A1(u_multiplier_STAGE3_acci_pp3_17_1__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_17_1__16_ ),
    .ZN(u_multiplier_pp3_17 [1]));
 AOI22_X2 u_multiplier_STAGE3_acci_pp3_17_1__27_  (.A1(u_multiplier_pp2_17 [1]),
    .A2(u_multiplier_pp2_17 [0]),
    .B1(u_multiplier_pp2_17 [2]),
    .B2(u_multiplier_pp2_17 [3]),
    .ZN(u_multiplier_STAGE3_acci_pp3_17_1__17_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_17_1__28_  (.A1(u_multiplier_STAGE3_acci_pp3_17_1__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_17_1__17_ ),
    .ZN(u_multiplier_pp3_18 [2]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_18_0__21_  (.A1(u_multiplier_pp2_18 [5]),
    .A2(u_multiplier_pp2_18 [4]),
    .A3(u_multiplier_pp2_18 [6]),
    .ZN(u_multiplier_STAGE3_acci_pp3_18_0__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_18_0__22_  (.A(u_multiplier_pp2_18 [5]),
    .B(u_multiplier_pp2_18 [4]),
    .Z(u_multiplier_STAGE3_acci_pp3_18_0__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_18_0__23_  (.A(u_multiplier_pp2_18 [6]),
    .B(u_multiplier_pp2_18 [7]),
    .Z(u_multiplier_STAGE3_acci_pp3_18_0__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_18_0__24_  (.A1(u_multiplier_STAGE3_acci_pp3_18_0__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_18_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_18_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_18_0__25_  (.A(u_multiplier_STAGE3_acci_pp3_18_0__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_18_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_18_0__16_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_18_0__26_  (.A1(u_multiplier_STAGE3_acci_pp3_18_0__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_18_0__16_ ),
    .ZN(u_multiplier_pp3_18 [0]));
 AOI22_X2 u_multiplier_STAGE3_acci_pp3_18_0__27_  (.A1(u_multiplier_pp2_18 [5]),
    .A2(u_multiplier_pp2_18 [4]),
    .B1(u_multiplier_pp2_18 [6]),
    .B2(u_multiplier_pp2_18 [7]),
    .ZN(u_multiplier_STAGE3_acci_pp3_18_0__17_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_18_0__28_  (.A1(u_multiplier_STAGE3_acci_pp3_18_0__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_18_0__17_ ),
    .ZN(u_multiplier_pp3_19 [3]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_18_1__21_  (.A1(u_multiplier_pp2_18 [1]),
    .A2(u_multiplier_pp2_18 [0]),
    .A3(u_multiplier_pp2_18 [2]),
    .ZN(u_multiplier_STAGE3_acci_pp3_18_1__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_18_1__22_  (.A(u_multiplier_pp2_18 [1]),
    .B(u_multiplier_pp2_18 [0]),
    .Z(u_multiplier_STAGE3_acci_pp3_18_1__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_18_1__23_  (.A(u_multiplier_pp2_18 [2]),
    .B(u_multiplier_pp2_18 [3]),
    .Z(u_multiplier_STAGE3_acci_pp3_18_1__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_18_1__24_  (.A1(u_multiplier_STAGE3_acci_pp3_18_1__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_18_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_18_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_18_1__25_  (.A(u_multiplier_STAGE3_acci_pp3_18_1__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_18_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_18_1__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_18_1__26_  (.A1(u_multiplier_STAGE3_acci_pp3_18_1__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_18_1__16_ ),
    .ZN(u_multiplier_pp3_18 [1]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_18_1__27_  (.A1(u_multiplier_pp2_18 [1]),
    .A2(u_multiplier_pp2_18 [0]),
    .B1(u_multiplier_pp2_18 [2]),
    .B2(u_multiplier_pp2_18 [3]),
    .ZN(u_multiplier_STAGE3_acci_pp3_18_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_18_1__28_  (.A1(u_multiplier_STAGE3_acci_pp3_18_1__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_18_1__17_ ),
    .ZN(u_multiplier_pp3_19 [2]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_19_0__21_  (.A1(u_multiplier_pp2_19 [5]),
    .A2(u_multiplier_pp2_19 [4]),
    .A3(u_multiplier_pp2_19 [6]),
    .ZN(u_multiplier_STAGE3_acci_pp3_19_0__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_19_0__22_  (.A(u_multiplier_pp2_19 [5]),
    .B(u_multiplier_pp2_19 [4]),
    .Z(u_multiplier_STAGE3_acci_pp3_19_0__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_19_0__23_  (.A(u_multiplier_pp2_19 [6]),
    .B(u_multiplier_pp2_19 [7]),
    .Z(u_multiplier_STAGE3_acci_pp3_19_0__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_19_0__24_  (.A1(u_multiplier_STAGE3_acci_pp3_19_0__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_19_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_19_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_19_0__25_  (.A(u_multiplier_STAGE3_acci_pp3_19_0__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_19_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_19_0__16_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_19_0__26_  (.A1(u_multiplier_STAGE3_acci_pp3_19_0__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_19_0__16_ ),
    .ZN(u_multiplier_pp3_19 [0]));
 AOI22_X2 u_multiplier_STAGE3_acci_pp3_19_0__27_  (.A1(u_multiplier_pp2_19 [5]),
    .A2(u_multiplier_pp2_19 [4]),
    .B1(u_multiplier_pp2_19 [6]),
    .B2(u_multiplier_pp2_19 [7]),
    .ZN(u_multiplier_STAGE3_acci_pp3_19_0__17_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_19_0__28_  (.A1(u_multiplier_STAGE3_acci_pp3_19_0__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_19_0__17_ ),
    .ZN(u_multiplier_pp3_20 [3]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_19_1__21_  (.A1(u_multiplier_pp2_19 [1]),
    .A2(u_multiplier_pp2_19 [0]),
    .A3(u_multiplier_pp2_19 [2]),
    .ZN(u_multiplier_STAGE3_acci_pp3_19_1__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_19_1__22_  (.A(u_multiplier_pp2_19 [1]),
    .B(u_multiplier_pp2_19 [0]),
    .Z(u_multiplier_STAGE3_acci_pp3_19_1__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_19_1__23_  (.A(u_multiplier_pp2_19 [2]),
    .B(u_multiplier_pp2_19 [3]),
    .Z(u_multiplier_STAGE3_acci_pp3_19_1__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_19_1__24_  (.A1(u_multiplier_STAGE3_acci_pp3_19_1__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_19_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_19_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_19_1__25_  (.A(u_multiplier_STAGE3_acci_pp3_19_1__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_19_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_19_1__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_19_1__26_  (.A1(u_multiplier_STAGE3_acci_pp3_19_1__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_19_1__16_ ),
    .ZN(u_multiplier_pp3_19 [1]));
 AOI22_X2 u_multiplier_STAGE3_acci_pp3_19_1__27_  (.A1(u_multiplier_pp2_19 [1]),
    .A2(u_multiplier_pp2_19 [0]),
    .B1(u_multiplier_pp2_19 [2]),
    .B2(u_multiplier_pp2_19 [3]),
    .ZN(u_multiplier_STAGE3_acci_pp3_19_1__17_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_19_1__28_  (.A1(u_multiplier_STAGE3_acci_pp3_19_1__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_19_1__17_ ),
    .ZN(u_multiplier_pp3_20 [2]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_20_0__21_  (.A1(u_multiplier_pp2_20 [5]),
    .A2(u_multiplier_pp2_20 [4]),
    .A3(u_multiplier_pp2_20 [6]),
    .ZN(u_multiplier_STAGE3_acci_pp3_20_0__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_20_0__22_  (.A(u_multiplier_pp2_20 [5]),
    .B(u_multiplier_pp2_20 [4]),
    .Z(u_multiplier_STAGE3_acci_pp3_20_0__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_20_0__23_  (.A(u_multiplier_pp2_20 [6]),
    .B(u_multiplier_pp2_20 [7]),
    .Z(u_multiplier_STAGE3_acci_pp3_20_0__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_20_0__24_  (.A1(u_multiplier_STAGE3_acci_pp3_20_0__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_20_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_20_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_20_0__25_  (.A(u_multiplier_STAGE3_acci_pp3_20_0__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_20_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_20_0__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_20_0__26_  (.A1(u_multiplier_STAGE3_acci_pp3_20_0__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_20_0__16_ ),
    .ZN(u_multiplier_pp3_20 [0]));
 AOI22_X2 u_multiplier_STAGE3_acci_pp3_20_0__27_  (.A1(u_multiplier_pp2_20 [5]),
    .A2(u_multiplier_pp2_20 [4]),
    .B1(u_multiplier_pp2_20 [6]),
    .B2(u_multiplier_pp2_20 [7]),
    .ZN(u_multiplier_STAGE3_acci_pp3_20_0__17_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_20_0__28_  (.A1(u_multiplier_STAGE3_acci_pp3_20_0__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_20_0__17_ ),
    .ZN(u_multiplier_pp3_21 [3]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_20_1__21_  (.A1(u_multiplier_pp2_20 [1]),
    .A2(u_multiplier_pp2_20 [0]),
    .A3(u_multiplier_pp2_20 [2]),
    .ZN(u_multiplier_STAGE3_acci_pp3_20_1__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_20_1__22_  (.A(u_multiplier_pp2_20 [1]),
    .B(u_multiplier_pp2_20 [0]),
    .Z(u_multiplier_STAGE3_acci_pp3_20_1__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_20_1__23_  (.A(u_multiplier_pp2_20 [2]),
    .B(u_multiplier_pp2_20 [3]),
    .Z(u_multiplier_STAGE3_acci_pp3_20_1__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_20_1__24_  (.A1(u_multiplier_STAGE3_acci_pp3_20_1__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_20_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_20_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_20_1__25_  (.A(u_multiplier_STAGE3_acci_pp3_20_1__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_20_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_20_1__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_20_1__26_  (.A1(u_multiplier_STAGE3_acci_pp3_20_1__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_20_1__16_ ),
    .ZN(u_multiplier_pp3_20 [1]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_20_1__27_  (.A1(u_multiplier_pp2_20 [1]),
    .A2(u_multiplier_pp2_20 [0]),
    .B1(u_multiplier_pp2_20 [2]),
    .B2(u_multiplier_pp2_20 [3]),
    .ZN(u_multiplier_STAGE3_acci_pp3_20_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_20_1__28_  (.A1(u_multiplier_STAGE3_acci_pp3_20_1__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_20_1__17_ ),
    .ZN(u_multiplier_pp3_21 [2]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_21_0__21_  (.A1(u_multiplier_pp2_21 [5]),
    .A2(u_multiplier_pp2_21 [4]),
    .A3(u_multiplier_pp2_21 [6]),
    .ZN(u_multiplier_STAGE3_acci_pp3_21_0__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_21_0__22_  (.A(u_multiplier_pp2_21 [5]),
    .B(u_multiplier_pp2_21 [4]),
    .Z(u_multiplier_STAGE3_acci_pp3_21_0__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_21_0__23_  (.A(u_multiplier_pp2_21 [6]),
    .B(u_multiplier_pp2_21 [7]),
    .Z(u_multiplier_STAGE3_acci_pp3_21_0__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_21_0__24_  (.A1(u_multiplier_STAGE3_acci_pp3_21_0__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_21_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_21_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_21_0__25_  (.A(u_multiplier_STAGE3_acci_pp3_21_0__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_21_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_21_0__16_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_21_0__26_  (.A1(u_multiplier_STAGE3_acci_pp3_21_0__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_21_0__16_ ),
    .ZN(u_multiplier_pp3_21 [0]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_21_0__27_  (.A1(u_multiplier_pp2_21 [5]),
    .A2(u_multiplier_pp2_21 [4]),
    .B1(u_multiplier_pp2_21 [6]),
    .B2(u_multiplier_pp2_21 [7]),
    .ZN(u_multiplier_STAGE3_acci_pp3_21_0__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_21_0__28_  (.A1(u_multiplier_STAGE3_acci_pp3_21_0__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_21_0__17_ ),
    .ZN(u_multiplier_pp3_22 [3]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_21_1__21_  (.A1(u_multiplier_pp2_21 [1]),
    .A2(u_multiplier_pp2_21 [0]),
    .A3(u_multiplier_pp2_21 [2]),
    .ZN(u_multiplier_STAGE3_acci_pp3_21_1__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_21_1__22_  (.A(u_multiplier_pp2_21 [1]),
    .B(u_multiplier_pp2_21 [0]),
    .Z(u_multiplier_STAGE3_acci_pp3_21_1__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_21_1__23_  (.A(u_multiplier_pp2_21 [2]),
    .B(u_multiplier_pp2_21 [3]),
    .Z(u_multiplier_STAGE3_acci_pp3_21_1__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_21_1__24_  (.A1(u_multiplier_STAGE3_acci_pp3_21_1__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_21_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_21_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_21_1__25_  (.A(u_multiplier_STAGE3_acci_pp3_21_1__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_21_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_21_1__16_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_21_1__26_  (.A1(u_multiplier_STAGE3_acci_pp3_21_1__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_21_1__16_ ),
    .ZN(u_multiplier_pp3_21 [1]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_21_1__27_  (.A1(u_multiplier_pp2_21 [1]),
    .A2(u_multiplier_pp2_21 [0]),
    .B1(u_multiplier_pp2_21 [2]),
    .B2(u_multiplier_pp2_21 [3]),
    .ZN(u_multiplier_STAGE3_acci_pp3_21_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_21_1__28_  (.A1(u_multiplier_STAGE3_acci_pp3_21_1__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_21_1__17_ ),
    .ZN(u_multiplier_pp3_22 [2]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_22_0__21_  (.A1(u_multiplier_pp2_22 [5]),
    .A2(u_multiplier_pp2_22 [4]),
    .A3(u_multiplier_pp2_22 [6]),
    .ZN(u_multiplier_STAGE3_acci_pp3_22_0__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_22_0__22_  (.A(u_multiplier_pp2_22 [5]),
    .B(u_multiplier_pp2_22 [4]),
    .Z(u_multiplier_STAGE3_acci_pp3_22_0__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_22_0__23_  (.A(u_multiplier_pp2_22 [6]),
    .B(u_multiplier_pp2_22 [7]),
    .Z(u_multiplier_STAGE3_acci_pp3_22_0__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_22_0__24_  (.A1(u_multiplier_STAGE3_acci_pp3_22_0__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_22_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_22_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_22_0__25_  (.A(u_multiplier_STAGE3_acci_pp3_22_0__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_22_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_22_0__16_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_22_0__26_  (.A1(u_multiplier_STAGE3_acci_pp3_22_0__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_22_0__16_ ),
    .ZN(u_multiplier_pp3_22 [0]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_22_0__27_  (.A1(u_multiplier_pp2_22 [5]),
    .A2(u_multiplier_pp2_22 [4]),
    .B1(u_multiplier_pp2_22 [6]),
    .B2(u_multiplier_pp2_22 [7]),
    .ZN(u_multiplier_STAGE3_acci_pp3_22_0__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_22_0__28_  (.A1(u_multiplier_STAGE3_acci_pp3_22_0__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_22_0__17_ ),
    .ZN(u_multiplier_pp3_23 [3]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_22_1__21_  (.A1(u_multiplier_pp2_22 [1]),
    .A2(u_multiplier_pp2_22 [0]),
    .A3(u_multiplier_pp2_22 [2]),
    .ZN(u_multiplier_STAGE3_acci_pp3_22_1__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_22_1__22_  (.A(u_multiplier_pp2_22 [1]),
    .B(u_multiplier_pp2_22 [0]),
    .Z(u_multiplier_STAGE3_acci_pp3_22_1__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_22_1__23_  (.A(u_multiplier_pp2_22 [2]),
    .B(u_multiplier_pp2_22 [3]),
    .Z(u_multiplier_STAGE3_acci_pp3_22_1__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_22_1__24_  (.A1(u_multiplier_STAGE3_acci_pp3_22_1__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_22_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_22_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_22_1__25_  (.A(u_multiplier_STAGE3_acci_pp3_22_1__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_22_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_22_1__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_22_1__26_  (.A1(u_multiplier_STAGE3_acci_pp3_22_1__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_22_1__16_ ),
    .ZN(u_multiplier_pp3_22 [1]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_22_1__27_  (.A1(u_multiplier_pp2_22 [1]),
    .A2(u_multiplier_pp2_22 [0]),
    .B1(u_multiplier_pp2_22 [2]),
    .B2(u_multiplier_pp2_22 [3]),
    .ZN(u_multiplier_STAGE3_acci_pp3_22_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_22_1__28_  (.A1(u_multiplier_STAGE3_acci_pp3_22_1__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_22_1__17_ ),
    .ZN(u_multiplier_pp3_23 [2]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_23_0__21_  (.A1(u_multiplier_pp2_23 [5]),
    .A2(u_multiplier_pp2_23 [4]),
    .A3(u_multiplier_pp2_23 [6]),
    .ZN(u_multiplier_STAGE3_acci_pp3_23_0__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_23_0__22_  (.A(u_multiplier_pp2_23 [5]),
    .B(u_multiplier_pp2_23 [4]),
    .Z(u_multiplier_STAGE3_acci_pp3_23_0__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_23_0__23_  (.A(u_multiplier_pp2_23 [6]),
    .B(u_multiplier_pp2_23 [7]),
    .Z(u_multiplier_STAGE3_acci_pp3_23_0__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_23_0__24_  (.A1(u_multiplier_STAGE3_acci_pp3_23_0__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_23_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_23_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_23_0__25_  (.A(u_multiplier_STAGE3_acci_pp3_23_0__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_23_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_23_0__16_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_23_0__26_  (.A1(u_multiplier_STAGE3_acci_pp3_23_0__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_23_0__16_ ),
    .ZN(u_multiplier_pp3_23 [0]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_23_0__27_  (.A1(u_multiplier_pp2_23 [5]),
    .A2(u_multiplier_pp2_23 [4]),
    .B1(u_multiplier_pp2_23 [6]),
    .B2(u_multiplier_pp2_23 [7]),
    .ZN(u_multiplier_STAGE3_acci_pp3_23_0__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_23_0__28_  (.A1(u_multiplier_STAGE3_acci_pp3_23_0__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_23_0__17_ ),
    .ZN(u_multiplier_pp3_24 [3]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_23_1__21_  (.A1(u_multiplier_pp2_23 [1]),
    .A2(u_multiplier_pp2_23 [0]),
    .A3(u_multiplier_pp2_23 [2]),
    .ZN(u_multiplier_STAGE3_acci_pp3_23_1__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_23_1__22_  (.A(u_multiplier_pp2_23 [1]),
    .B(u_multiplier_pp2_23 [0]),
    .Z(u_multiplier_STAGE3_acci_pp3_23_1__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_23_1__23_  (.A(u_multiplier_pp2_23 [2]),
    .B(u_multiplier_pp2_23 [3]),
    .Z(u_multiplier_STAGE3_acci_pp3_23_1__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_23_1__24_  (.A1(u_multiplier_STAGE3_acci_pp3_23_1__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_23_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_23_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_23_1__25_  (.A(u_multiplier_STAGE3_acci_pp3_23_1__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_23_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_23_1__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_23_1__26_  (.A1(u_multiplier_STAGE3_acci_pp3_23_1__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_23_1__16_ ),
    .ZN(u_multiplier_pp3_23 [1]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_23_1__27_  (.A1(u_multiplier_pp2_23 [1]),
    .A2(u_multiplier_pp2_23 [0]),
    .B1(u_multiplier_pp2_23 [2]),
    .B2(u_multiplier_pp2_23 [3]),
    .ZN(u_multiplier_STAGE3_acci_pp3_23_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_23_1__28_  (.A1(u_multiplier_STAGE3_acci_pp3_23_1__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_23_1__17_ ),
    .ZN(u_multiplier_pp3_24 [2]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_24_0__21_  (.A1(u_multiplier_pp2_24 [5]),
    .A2(u_multiplier_pp2_24 [4]),
    .A3(u_multiplier_pp2_24 [6]),
    .ZN(u_multiplier_STAGE3_acci_pp3_24_0__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_24_0__22_  (.A(u_multiplier_pp2_24 [5]),
    .B(u_multiplier_pp2_24 [4]),
    .Z(u_multiplier_STAGE3_acci_pp3_24_0__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_24_0__23_  (.A(u_multiplier_pp2_24 [6]),
    .B(u_multiplier_pp2_24 [7]),
    .Z(u_multiplier_STAGE3_acci_pp3_24_0__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_24_0__24_  (.A1(u_multiplier_STAGE3_acci_pp3_24_0__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_24_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_24_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_24_0__25_  (.A(u_multiplier_STAGE3_acci_pp3_24_0__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_24_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_24_0__16_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_24_0__26_  (.A1(u_multiplier_STAGE3_acci_pp3_24_0__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_24_0__16_ ),
    .ZN(u_multiplier_pp3_24 [0]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_24_0__27_  (.A1(u_multiplier_pp2_24 [5]),
    .A2(u_multiplier_pp2_24 [4]),
    .B1(u_multiplier_pp2_24 [6]),
    .B2(u_multiplier_pp2_24 [7]),
    .ZN(u_multiplier_STAGE3_acci_pp3_24_0__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_24_0__28_  (.A1(u_multiplier_STAGE3_acci_pp3_24_0__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_24_0__17_ ),
    .ZN(u_multiplier_pp3_25 [3]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_24_1__21_  (.A1(u_multiplier_pp2_24 [1]),
    .A2(u_multiplier_pp2_24 [0]),
    .A3(u_multiplier_pp2_24 [2]),
    .ZN(u_multiplier_STAGE3_acci_pp3_24_1__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_24_1__22_  (.A(u_multiplier_pp2_24 [1]),
    .B(u_multiplier_pp2_24 [0]),
    .Z(u_multiplier_STAGE3_acci_pp3_24_1__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_24_1__23_  (.A(u_multiplier_pp2_24 [2]),
    .B(u_multiplier_pp2_24 [3]),
    .Z(u_multiplier_STAGE3_acci_pp3_24_1__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_24_1__24_  (.A1(u_multiplier_STAGE3_acci_pp3_24_1__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_24_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_24_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_24_1__25_  (.A(u_multiplier_STAGE3_acci_pp3_24_1__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_24_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_24_1__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_24_1__26_  (.A1(u_multiplier_STAGE3_acci_pp3_24_1__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_24_1__16_ ),
    .ZN(u_multiplier_pp3_24 [1]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_24_1__27_  (.A1(u_multiplier_pp2_24 [1]),
    .A2(u_multiplier_pp2_24 [0]),
    .B1(u_multiplier_pp2_24 [2]),
    .B2(u_multiplier_pp2_24 [3]),
    .ZN(u_multiplier_STAGE3_acci_pp3_24_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_24_1__28_  (.A1(u_multiplier_STAGE3_acci_pp3_24_1__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_24_1__17_ ),
    .ZN(u_multiplier_pp3_25 [2]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_25_0__21_  (.A1(u_multiplier_pp2_25 [5]),
    .A2(u_multiplier_pp2_25 [4]),
    .A3(u_multiplier_pp2_25 [6]),
    .ZN(u_multiplier_STAGE3_acci_pp3_25_0__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_25_0__22_  (.A(u_multiplier_pp2_25 [5]),
    .B(u_multiplier_pp2_25 [4]),
    .Z(u_multiplier_STAGE3_acci_pp3_25_0__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_25_0__23_  (.A(u_multiplier_pp2_25 [6]),
    .B(u_multiplier_pp2_25 [7]),
    .Z(u_multiplier_STAGE3_acci_pp3_25_0__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_25_0__24_  (.A1(u_multiplier_STAGE3_acci_pp3_25_0__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_25_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_25_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_25_0__25_  (.A(u_multiplier_STAGE3_acci_pp3_25_0__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_25_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_25_0__16_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_25_0__26_  (.A1(u_multiplier_STAGE3_acci_pp3_25_0__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_25_0__16_ ),
    .ZN(u_multiplier_pp3_25 [0]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_25_0__27_  (.A1(u_multiplier_pp2_25 [5]),
    .A2(u_multiplier_pp2_25 [4]),
    .B1(u_multiplier_pp2_25 [6]),
    .B2(u_multiplier_pp2_25 [7]),
    .ZN(u_multiplier_STAGE3_acci_pp3_25_0__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_25_0__28_  (.A1(u_multiplier_STAGE3_acci_pp3_25_0__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_25_0__17_ ),
    .ZN(u_multiplier_pp3_26 [3]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_25_1__21_  (.A1(u_multiplier_pp2_25 [1]),
    .A2(u_multiplier_pp2_25 [0]),
    .A3(u_multiplier_pp2_25 [2]),
    .ZN(u_multiplier_STAGE3_acci_pp3_25_1__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_25_1__22_  (.A(u_multiplier_pp2_25 [1]),
    .B(u_multiplier_pp2_25 [0]),
    .Z(u_multiplier_STAGE3_acci_pp3_25_1__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_25_1__23_  (.A(u_multiplier_pp2_25 [2]),
    .B(u_multiplier_pp2_25 [3]),
    .Z(u_multiplier_STAGE3_acci_pp3_25_1__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_25_1__24_  (.A1(u_multiplier_STAGE3_acci_pp3_25_1__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_25_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_25_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_25_1__25_  (.A(u_multiplier_STAGE3_acci_pp3_25_1__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_25_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_25_1__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_25_1__26_  (.A1(u_multiplier_STAGE3_acci_pp3_25_1__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_25_1__16_ ),
    .ZN(u_multiplier_pp3_25 [1]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_25_1__27_  (.A1(u_multiplier_pp2_25 [1]),
    .A2(u_multiplier_pp2_25 [0]),
    .B1(u_multiplier_pp2_25 [2]),
    .B2(u_multiplier_pp2_25 [3]),
    .ZN(u_multiplier_STAGE3_acci_pp3_25_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_25_1__28_  (.A1(u_multiplier_STAGE3_acci_pp3_25_1__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_25_1__17_ ),
    .ZN(u_multiplier_pp3_26 [2]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_26_0__21_  (.A1(u_multiplier_pp2_26 [5]),
    .A2(u_multiplier_pp2_26 [4]),
    .A3(u_multiplier_pp2_26 [6]),
    .ZN(u_multiplier_STAGE3_acci_pp3_26_0__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_26_0__22_  (.A(u_multiplier_pp2_26 [5]),
    .B(u_multiplier_pp2_26 [4]),
    .Z(u_multiplier_STAGE3_acci_pp3_26_0__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_26_0__23_  (.A(u_multiplier_pp2_26 [6]),
    .B(u_multiplier_pp2_26 [7]),
    .Z(u_multiplier_STAGE3_acci_pp3_26_0__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_26_0__24_  (.A1(u_multiplier_STAGE3_acci_pp3_26_0__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_26_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_26_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_26_0__25_  (.A(u_multiplier_STAGE3_acci_pp3_26_0__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_26_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_26_0__16_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_26_0__26_  (.A1(u_multiplier_STAGE3_acci_pp3_26_0__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_26_0__16_ ),
    .ZN(u_multiplier_pp3_26 [0]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_26_0__27_  (.A1(u_multiplier_pp2_26 [5]),
    .A2(u_multiplier_pp2_26 [4]),
    .B1(u_multiplier_pp2_26 [6]),
    .B2(u_multiplier_pp2_26 [7]),
    .ZN(u_multiplier_STAGE3_acci_pp3_26_0__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_26_0__28_  (.A1(u_multiplier_STAGE3_acci_pp3_26_0__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_26_0__17_ ),
    .ZN(u_multiplier_pp3_27 [3]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_26_1__21_  (.A1(u_multiplier_pp2_26 [1]),
    .A2(u_multiplier_pp2_26 [0]),
    .A3(u_multiplier_pp2_26 [2]),
    .ZN(u_multiplier_STAGE3_acci_pp3_26_1__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_26_1__22_  (.A(u_multiplier_pp2_26 [1]),
    .B(u_multiplier_pp2_26 [0]),
    .Z(u_multiplier_STAGE3_acci_pp3_26_1__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_26_1__23_  (.A(u_multiplier_pp2_26 [2]),
    .B(u_multiplier_pp2_26 [3]),
    .Z(u_multiplier_STAGE3_acci_pp3_26_1__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_26_1__24_  (.A1(u_multiplier_STAGE3_acci_pp3_26_1__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_26_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_26_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_26_1__25_  (.A(u_multiplier_STAGE3_acci_pp3_26_1__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_26_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_26_1__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_26_1__26_  (.A1(u_multiplier_STAGE3_acci_pp3_26_1__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_26_1__16_ ),
    .ZN(u_multiplier_pp3_26 [1]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_26_1__27_  (.A1(u_multiplier_pp2_26 [1]),
    .A2(u_multiplier_pp2_26 [0]),
    .B1(u_multiplier_pp2_26 [2]),
    .B2(u_multiplier_pp2_26 [3]),
    .ZN(u_multiplier_STAGE3_acci_pp3_26_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_26_1__28_  (.A1(u_multiplier_STAGE3_acci_pp3_26_1__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_26_1__17_ ),
    .ZN(u_multiplier_pp3_27 [2]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_27_0__21_  (.A1(u_multiplier_pp2_27 [5]),
    .A2(u_multiplier_pp2_27 [4]),
    .A3(u_multiplier_pp2_27 [6]),
    .ZN(u_multiplier_STAGE3_acci_pp3_27_0__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_27_0__22_  (.A(u_multiplier_pp2_27 [5]),
    .B(u_multiplier_pp2_27 [4]),
    .Z(u_multiplier_STAGE3_acci_pp3_27_0__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_27_0__23_  (.A(u_multiplier_pp2_27 [6]),
    .B(u_multiplier_pp2_27 [7]),
    .Z(u_multiplier_STAGE3_acci_pp3_27_0__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_27_0__24_  (.A1(u_multiplier_STAGE3_acci_pp3_27_0__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_27_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_27_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_27_0__25_  (.A(u_multiplier_STAGE3_acci_pp3_27_0__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_27_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_27_0__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_27_0__26_  (.A1(u_multiplier_STAGE3_acci_pp3_27_0__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_27_0__16_ ),
    .ZN(u_multiplier_pp3_27 [0]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_27_0__27_  (.A1(u_multiplier_pp2_27 [5]),
    .A2(u_multiplier_pp2_27 [4]),
    .B1(u_multiplier_pp2_27 [6]),
    .B2(u_multiplier_pp2_27 [7]),
    .ZN(u_multiplier_STAGE3_acci_pp3_27_0__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_27_0__28_  (.A1(u_multiplier_STAGE3_acci_pp3_27_0__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_27_0__17_ ),
    .ZN(u_multiplier_pp3_28 [3]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_27_1__21_  (.A1(u_multiplier_pp2_27 [1]),
    .A2(u_multiplier_pp2_27 [0]),
    .A3(u_multiplier_pp2_27 [2]),
    .ZN(u_multiplier_STAGE3_acci_pp3_27_1__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_27_1__22_  (.A(u_multiplier_pp2_27 [1]),
    .B(u_multiplier_pp2_27 [0]),
    .Z(u_multiplier_STAGE3_acci_pp3_27_1__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_27_1__23_  (.A(u_multiplier_pp2_27 [2]),
    .B(u_multiplier_pp2_27 [3]),
    .Z(u_multiplier_STAGE3_acci_pp3_27_1__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_27_1__24_  (.A1(u_multiplier_STAGE3_acci_pp3_27_1__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_27_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_27_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_27_1__25_  (.A(u_multiplier_STAGE3_acci_pp3_27_1__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_27_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_27_1__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_27_1__26_  (.A1(u_multiplier_STAGE3_acci_pp3_27_1__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_27_1__16_ ),
    .ZN(u_multiplier_pp3_27 [1]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_27_1__27_  (.A1(u_multiplier_pp2_27 [1]),
    .A2(u_multiplier_pp2_27 [0]),
    .B1(u_multiplier_pp2_27 [2]),
    .B2(u_multiplier_pp2_27 [3]),
    .ZN(u_multiplier_STAGE3_acci_pp3_27_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_27_1__28_  (.A1(u_multiplier_STAGE3_acci_pp3_27_1__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_27_1__17_ ),
    .ZN(u_multiplier_pp3_28 [2]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_28_0__21_  (.A1(u_multiplier_pp2_28 [5]),
    .A2(u_multiplier_pp2_28 [4]),
    .A3(u_multiplier_pp2_28 [6]),
    .ZN(u_multiplier_STAGE3_acci_pp3_28_0__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_28_0__22_  (.A(u_multiplier_pp2_28 [5]),
    .B(u_multiplier_pp2_28 [4]),
    .Z(u_multiplier_STAGE3_acci_pp3_28_0__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_28_0__23_  (.A(u_multiplier_pp2_28 [6]),
    .B(u_multiplier_pp2_28 [7]),
    .Z(u_multiplier_STAGE3_acci_pp3_28_0__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_28_0__24_  (.A1(u_multiplier_STAGE3_acci_pp3_28_0__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_28_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_28_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_28_0__25_  (.A(u_multiplier_STAGE3_acci_pp3_28_0__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_28_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_28_0__16_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_28_0__26_  (.A1(u_multiplier_STAGE3_acci_pp3_28_0__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_28_0__16_ ),
    .ZN(u_multiplier_pp3_28 [0]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_28_0__27_  (.A1(u_multiplier_pp2_28 [5]),
    .A2(u_multiplier_pp2_28 [4]),
    .B1(u_multiplier_pp2_28 [6]),
    .B2(u_multiplier_pp2_28 [7]),
    .ZN(u_multiplier_STAGE3_acci_pp3_28_0__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_28_0__28_  (.A1(u_multiplier_STAGE3_acci_pp3_28_0__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_28_0__17_ ),
    .ZN(u_multiplier_pp3_29 [3]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_28_1__21_  (.A1(u_multiplier_pp2_28 [1]),
    .A2(u_multiplier_pp2_28 [0]),
    .A3(u_multiplier_pp2_28 [2]),
    .ZN(u_multiplier_STAGE3_acci_pp3_28_1__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_28_1__22_  (.A(u_multiplier_pp2_28 [1]),
    .B(u_multiplier_pp2_28 [0]),
    .Z(u_multiplier_STAGE3_acci_pp3_28_1__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_28_1__23_  (.A(u_multiplier_pp2_28 [2]),
    .B(u_multiplier_pp2_28 [3]),
    .Z(u_multiplier_STAGE3_acci_pp3_28_1__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_28_1__24_  (.A1(u_multiplier_STAGE3_acci_pp3_28_1__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_28_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_28_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_28_1__25_  (.A(u_multiplier_STAGE3_acci_pp3_28_1__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_28_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_28_1__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_28_1__26_  (.A1(u_multiplier_STAGE3_acci_pp3_28_1__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_28_1__16_ ),
    .ZN(u_multiplier_pp3_28 [1]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_28_1__27_  (.A1(u_multiplier_pp2_28 [1]),
    .A2(u_multiplier_pp2_28 [0]),
    .B1(u_multiplier_pp2_28 [2]),
    .B2(u_multiplier_pp2_28 [3]),
    .ZN(u_multiplier_STAGE3_acci_pp3_28_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_28_1__28_  (.A1(u_multiplier_STAGE3_acci_pp3_28_1__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_28_1__17_ ),
    .ZN(u_multiplier_pp3_29 [2]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_29_0__21_  (.A1(u_multiplier_pp2_29 [5]),
    .A2(u_multiplier_pp2_29 [4]),
    .A3(u_multiplier_pp2_29 [6]),
    .ZN(u_multiplier_STAGE3_acci_pp3_29_0__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_29_0__22_  (.A(u_multiplier_pp2_29 [5]),
    .B(u_multiplier_pp2_29 [4]),
    .Z(u_multiplier_STAGE3_acci_pp3_29_0__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_29_0__23_  (.A(u_multiplier_pp2_29 [6]),
    .B(u_multiplier_pp2_29 [7]),
    .Z(u_multiplier_STAGE3_acci_pp3_29_0__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_29_0__24_  (.A1(u_multiplier_STAGE3_acci_pp3_29_0__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_29_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_29_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_29_0__25_  (.A(u_multiplier_STAGE3_acci_pp3_29_0__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_29_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_29_0__16_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_29_0__26_  (.A1(u_multiplier_STAGE3_acci_pp3_29_0__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_29_0__16_ ),
    .ZN(u_multiplier_pp3_29 [0]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_29_0__27_  (.A1(u_multiplier_pp2_29 [5]),
    .A2(u_multiplier_pp2_29 [4]),
    .B1(u_multiplier_pp2_29 [6]),
    .B2(u_multiplier_pp2_29 [7]),
    .ZN(u_multiplier_STAGE3_acci_pp3_29_0__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_29_0__28_  (.A1(u_multiplier_STAGE3_acci_pp3_29_0__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_29_0__17_ ),
    .ZN(u_multiplier_pp3_30 [3]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_29_1__21_  (.A1(u_multiplier_pp2_29 [1]),
    .A2(u_multiplier_pp2_29 [0]),
    .A3(u_multiplier_pp2_29 [2]),
    .ZN(u_multiplier_STAGE3_acci_pp3_29_1__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_29_1__22_  (.A(u_multiplier_pp2_29 [1]),
    .B(u_multiplier_pp2_29 [0]),
    .Z(u_multiplier_STAGE3_acci_pp3_29_1__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_29_1__23_  (.A(u_multiplier_pp2_29 [2]),
    .B(u_multiplier_pp2_29 [3]),
    .Z(u_multiplier_STAGE3_acci_pp3_29_1__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_29_1__24_  (.A1(u_multiplier_STAGE3_acci_pp3_29_1__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_29_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_29_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_29_1__25_  (.A(u_multiplier_STAGE3_acci_pp3_29_1__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_29_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_29_1__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_29_1__26_  (.A1(u_multiplier_STAGE3_acci_pp3_29_1__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_29_1__16_ ),
    .ZN(u_multiplier_pp3_29 [1]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_29_1__27_  (.A1(u_multiplier_pp2_29 [1]),
    .A2(u_multiplier_pp2_29 [0]),
    .B1(u_multiplier_pp2_29 [2]),
    .B2(u_multiplier_pp2_29 [3]),
    .ZN(u_multiplier_STAGE3_acci_pp3_29_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_29_1__28_  (.A1(u_multiplier_STAGE3_acci_pp3_29_1__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_29_1__17_ ),
    .ZN(u_multiplier_pp3_30 [2]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_30_0__21_  (.A1(u_multiplier_pp2_30 [5]),
    .A2(u_multiplier_pp2_30 [4]),
    .A3(u_multiplier_pp2_30 [6]),
    .ZN(u_multiplier_STAGE3_acci_pp3_30_0__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_30_0__22_  (.A(u_multiplier_pp2_30 [5]),
    .B(u_multiplier_pp2_30 [4]),
    .Z(u_multiplier_STAGE3_acci_pp3_30_0__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_30_0__23_  (.A(u_multiplier_pp2_30 [6]),
    .B(u_multiplier_pp2_30 [7]),
    .Z(u_multiplier_STAGE3_acci_pp3_30_0__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_30_0__24_  (.A1(u_multiplier_STAGE3_acci_pp3_30_0__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_30_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_30_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_30_0__25_  (.A(u_multiplier_STAGE3_acci_pp3_30_0__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_30_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_30_0__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_30_0__26_  (.A1(u_multiplier_STAGE3_acci_pp3_30_0__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_30_0__16_ ),
    .ZN(u_multiplier_pp3_30 [0]));
 AOI22_X2 u_multiplier_STAGE3_acci_pp3_30_0__27_  (.A1(u_multiplier_pp2_30 [5]),
    .A2(u_multiplier_pp2_30 [4]),
    .B1(u_multiplier_pp2_30 [6]),
    .B2(u_multiplier_pp2_30 [7]),
    .ZN(u_multiplier_STAGE3_acci_pp3_30_0__17_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_30_0__28_  (.A1(u_multiplier_STAGE3_acci_pp3_30_0__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_30_0__17_ ),
    .ZN(u_multiplier_pp3_31 [3]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_30_1__21_  (.A1(u_multiplier_pp2_30 [1]),
    .A2(u_multiplier_pp2_30 [0]),
    .A3(u_multiplier_pp2_30 [2]),
    .ZN(u_multiplier_STAGE3_acci_pp3_30_1__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_30_1__22_  (.A(u_multiplier_pp2_30 [1]),
    .B(u_multiplier_pp2_30 [0]),
    .Z(u_multiplier_STAGE3_acci_pp3_30_1__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_30_1__23_  (.A(u_multiplier_pp2_30 [2]),
    .B(u_multiplier_pp2_30 [3]),
    .Z(u_multiplier_STAGE3_acci_pp3_30_1__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_30_1__24_  (.A1(u_multiplier_STAGE3_acci_pp3_30_1__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_30_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_30_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_30_1__25_  (.A(u_multiplier_STAGE3_acci_pp3_30_1__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_30_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_30_1__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_30_1__26_  (.A1(u_multiplier_STAGE3_acci_pp3_30_1__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_30_1__16_ ),
    .ZN(u_multiplier_pp3_30 [1]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_30_1__27_  (.A1(u_multiplier_pp2_30 [1]),
    .A2(u_multiplier_pp2_30 [0]),
    .B1(u_multiplier_pp2_30 [2]),
    .B2(u_multiplier_pp2_30 [3]),
    .ZN(u_multiplier_STAGE3_acci_pp3_30_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_30_1__28_  (.A1(u_multiplier_STAGE3_acci_pp3_30_1__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_30_1__17_ ),
    .ZN(u_multiplier_pp3_31 [2]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_31_0__21_  (.A1(u_multiplier_pp2_31 [5]),
    .A2(u_multiplier_pp2_31 [4]),
    .A3(u_multiplier_pp2_31 [6]),
    .ZN(u_multiplier_STAGE3_acci_pp3_31_0__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_31_0__22_  (.A(u_multiplier_pp2_31 [5]),
    .B(u_multiplier_pp2_31 [4]),
    .Z(u_multiplier_STAGE3_acci_pp3_31_0__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_31_0__23_  (.A(u_multiplier_pp2_31 [6]),
    .B(u_multiplier_pp2_31 [7]),
    .Z(u_multiplier_STAGE3_acci_pp3_31_0__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_31_0__24_  (.A1(u_multiplier_STAGE3_acci_pp3_31_0__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_31_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_31_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_31_0__25_  (.A(u_multiplier_STAGE3_acci_pp3_31_0__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_31_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_31_0__16_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_31_0__26_  (.A1(u_multiplier_STAGE3_acci_pp3_31_0__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_31_0__16_ ),
    .ZN(u_multiplier_pp3_31 [0]));
 AOI22_X4 u_multiplier_STAGE3_acci_pp3_31_0__27_  (.A1(u_multiplier_pp2_31 [5]),
    .A2(u_multiplier_pp2_31 [4]),
    .B1(u_multiplier_pp2_31 [6]),
    .B2(u_multiplier_pp2_31 [7]),
    .ZN(u_multiplier_STAGE3_acci_pp3_31_0__17_ ));
 NAND2_X4 u_multiplier_STAGE3_acci_pp3_31_0__28_  (.A1(u_multiplier_STAGE3_acci_pp3_31_0__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_31_0__17_ ),
    .ZN(u_multiplier_pp3_32 [3]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_31_1__21_  (.A1(u_multiplier_pp2_31 [1]),
    .A2(u_multiplier_pp2_31 [0]),
    .A3(u_multiplier_pp2_31 [2]),
    .ZN(u_multiplier_STAGE3_acci_pp3_31_1__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_31_1__22_  (.A(u_multiplier_pp2_31 [1]),
    .B(u_multiplier_pp2_31 [0]),
    .Z(u_multiplier_STAGE3_acci_pp3_31_1__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_31_1__23_  (.A(u_multiplier_pp2_31 [2]),
    .B(u_multiplier_pp2_31 [3]),
    .Z(u_multiplier_STAGE3_acci_pp3_31_1__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_31_1__24_  (.A1(u_multiplier_STAGE3_acci_pp3_31_1__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_31_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_31_1__15_ ));
 XNOR2_X2 u_multiplier_STAGE3_acci_pp3_31_1__25_  (.A(u_multiplier_STAGE3_acci_pp3_31_1__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_31_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_31_1__16_ ));
 NAND2_X4 u_multiplier_STAGE3_acci_pp3_31_1__26_  (.A1(u_multiplier_STAGE3_acci_pp3_31_1__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_31_1__16_ ),
    .ZN(u_multiplier_pp3_31 [1]));
 AOI22_X2 u_multiplier_STAGE3_acci_pp3_31_1__27_  (.A1(u_multiplier_pp2_31 [1]),
    .A2(u_multiplier_pp2_31 [0]),
    .B1(u_multiplier_pp2_31 [2]),
    .B2(u_multiplier_pp2_31 [3]),
    .ZN(u_multiplier_STAGE3_acci_pp3_31_1__17_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_31_1__28_  (.A1(u_multiplier_STAGE3_acci_pp3_31_1__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_31_1__17_ ),
    .ZN(u_multiplier_pp3_32 [2]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_5_0__21_  (.A1(u_multiplier_pp2_5 [3]),
    .A2(u_multiplier_pp2_5 [2]),
    .A3(u_multiplier_pp2_5 [4]),
    .ZN(u_multiplier_STAGE3_acci_pp3_5_0__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_5_0__22_  (.A(u_multiplier_pp2_5 [3]),
    .B(u_multiplier_pp2_5 [2]),
    .Z(u_multiplier_STAGE3_acci_pp3_5_0__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_5_0__23_  (.A(u_multiplier_pp2_5 [4]),
    .B(u_multiplier_pp2_5 [5]),
    .Z(u_multiplier_STAGE3_acci_pp3_5_0__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_5_0__24_  (.A1(u_multiplier_STAGE3_acci_pp3_5_0__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_5_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_5_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_5_0__25_  (.A(u_multiplier_STAGE3_acci_pp3_5_0__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_5_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_5_0__16_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_5_0__26_  (.A1(u_multiplier_STAGE3_acci_pp3_5_0__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_5_0__16_ ),
    .ZN(u_multiplier_pp3_5 [0]));
 AOI22_X2 u_multiplier_STAGE3_acci_pp3_5_0__27_  (.A1(u_multiplier_pp2_5 [3]),
    .A2(u_multiplier_pp2_5 [2]),
    .B1(u_multiplier_pp2_5 [4]),
    .B2(u_multiplier_pp2_5 [5]),
    .ZN(u_multiplier_STAGE3_acci_pp3_5_0__17_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_5_0__28_  (.A1(u_multiplier_STAGE3_acci_pp3_5_0__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_5_0__17_ ),
    .ZN(u_multiplier_pp3_6 [2]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_6_0__21_  (.A1(u_multiplier_pp2_6 [4]),
    .A2(u_multiplier_pp2_6 [3]),
    .A3(u_multiplier_pp2_6 [5]),
    .ZN(u_multiplier_STAGE3_acci_pp3_6_0__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_6_0__22_  (.A(u_multiplier_pp2_6 [4]),
    .B(u_multiplier_pp2_6 [3]),
    .Z(u_multiplier_STAGE3_acci_pp3_6_0__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_6_0__23_  (.A(u_multiplier_pp2_6 [5]),
    .B(u_multiplier_pp2_6 [6]),
    .Z(u_multiplier_STAGE3_acci_pp3_6_0__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_6_0__24_  (.A1(u_multiplier_STAGE3_acci_pp3_6_0__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_6_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_6_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_6_0__25_  (.A(u_multiplier_STAGE3_acci_pp3_6_0__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_6_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_6_0__16_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_6_0__26_  (.A1(u_multiplier_STAGE3_acci_pp3_6_0__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_6_0__16_ ),
    .ZN(u_multiplier_pp3_6 [0]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_6_0__27_  (.A1(u_multiplier_pp2_6 [4]),
    .A2(u_multiplier_pp2_6 [3]),
    .B1(u_multiplier_pp2_6 [5]),
    .B2(u_multiplier_pp2_6 [6]),
    .ZN(u_multiplier_STAGE3_acci_pp3_6_0__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_6_0__28_  (.A1(u_multiplier_STAGE3_acci_pp3_6_0__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_6_0__17_ ),
    .ZN(u_multiplier_pp3_7 [3]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_7_0__21_  (.A1(u_multiplier_pp2_7 [5]),
    .A2(u_multiplier_pp2_7 [4]),
    .A3(u_multiplier_pp2_7 [6]),
    .ZN(u_multiplier_STAGE3_acci_pp3_7_0__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_7_0__22_  (.A(u_multiplier_pp2_7 [5]),
    .B(u_multiplier_pp2_7 [4]),
    .Z(u_multiplier_STAGE3_acci_pp3_7_0__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_7_0__23_  (.A(u_multiplier_pp2_7 [6]),
    .B(u_multiplier_pp2_7 [7]),
    .Z(u_multiplier_STAGE3_acci_pp3_7_0__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_7_0__24_  (.A1(u_multiplier_STAGE3_acci_pp3_7_0__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_7_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_7_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_7_0__25_  (.A(u_multiplier_STAGE3_acci_pp3_7_0__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_7_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_7_0__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_7_0__26_  (.A1(u_multiplier_STAGE3_acci_pp3_7_0__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_7_0__16_ ),
    .ZN(u_multiplier_pp3_7 [0]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_7_0__27_  (.A1(u_multiplier_pp2_7 [5]),
    .A2(u_multiplier_pp2_7 [4]),
    .B1(u_multiplier_pp2_7 [6]),
    .B2(u_multiplier_pp2_7 [7]),
    .ZN(u_multiplier_STAGE3_acci_pp3_7_0__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_7_0__28_  (.A1(u_multiplier_STAGE3_acci_pp3_7_0__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_7_0__17_ ),
    .ZN(u_multiplier_pp3_8 [3]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_7_1__21_  (.A1(u_multiplier_pp2_7 [1]),
    .A2(u_multiplier_pp2_7 [0]),
    .A3(u_multiplier_pp2_7 [2]),
    .ZN(u_multiplier_STAGE3_acci_pp3_7_1__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_7_1__22_  (.A(u_multiplier_pp2_7 [1]),
    .B(u_multiplier_pp2_7 [0]),
    .Z(u_multiplier_STAGE3_acci_pp3_7_1__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_7_1__23_  (.A(u_multiplier_pp2_7 [2]),
    .B(u_multiplier_pp2_7 [3]),
    .Z(u_multiplier_STAGE3_acci_pp3_7_1__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_7_1__24_  (.A1(u_multiplier_STAGE3_acci_pp3_7_1__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_7_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_7_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_7_1__25_  (.A(u_multiplier_STAGE3_acci_pp3_7_1__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_7_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_7_1__16_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_7_1__26_  (.A1(u_multiplier_STAGE3_acci_pp3_7_1__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_7_1__16_ ),
    .ZN(u_multiplier_pp3_7 [1]));
 AOI22_X2 u_multiplier_STAGE3_acci_pp3_7_1__27_  (.A1(u_multiplier_pp2_7 [1]),
    .A2(u_multiplier_pp2_7 [0]),
    .B1(u_multiplier_pp2_7 [2]),
    .B2(u_multiplier_pp2_7 [3]),
    .ZN(u_multiplier_STAGE3_acci_pp3_7_1__17_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_7_1__28_  (.A1(u_multiplier_STAGE3_acci_pp3_7_1__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_7_1__17_ ),
    .ZN(u_multiplier_pp3_8 [2]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_8_0__21_  (.A1(u_multiplier_pp2_8 [5]),
    .A2(u_multiplier_pp2_8 [4]),
    .A3(u_multiplier_pp2_8 [6]),
    .ZN(u_multiplier_STAGE3_acci_pp3_8_0__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_8_0__22_  (.A(u_multiplier_pp2_8 [5]),
    .B(u_multiplier_pp2_8 [4]),
    .Z(u_multiplier_STAGE3_acci_pp3_8_0__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_8_0__23_  (.A(u_multiplier_pp2_8 [6]),
    .B(u_multiplier_pp2_8 [7]),
    .Z(u_multiplier_STAGE3_acci_pp3_8_0__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_8_0__24_  (.A1(u_multiplier_STAGE3_acci_pp3_8_0__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_8_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_8_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_8_0__25_  (.A(u_multiplier_STAGE3_acci_pp3_8_0__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_8_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_8_0__16_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_8_0__26_  (.A1(u_multiplier_STAGE3_acci_pp3_8_0__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_8_0__16_ ),
    .ZN(u_multiplier_pp3_8 [0]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_8_0__27_  (.A1(u_multiplier_pp2_8 [5]),
    .A2(u_multiplier_pp2_8 [4]),
    .B1(u_multiplier_pp2_8 [6]),
    .B2(u_multiplier_pp2_8 [7]),
    .ZN(u_multiplier_STAGE3_acci_pp3_8_0__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_8_0__28_  (.A1(u_multiplier_STAGE3_acci_pp3_8_0__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_8_0__17_ ),
    .ZN(u_multiplier_pp3_9 [3]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_8_1__21_  (.A1(u_multiplier_pp2_8 [1]),
    .A2(u_multiplier_pp2_8 [0]),
    .A3(u_multiplier_pp2_8 [2]),
    .ZN(u_multiplier_STAGE3_acci_pp3_8_1__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_8_1__22_  (.A(u_multiplier_pp2_8 [1]),
    .B(u_multiplier_pp2_8 [0]),
    .Z(u_multiplier_STAGE3_acci_pp3_8_1__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_8_1__23_  (.A(u_multiplier_pp2_8 [2]),
    .B(u_multiplier_pp2_8 [3]),
    .Z(u_multiplier_STAGE3_acci_pp3_8_1__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_8_1__24_  (.A1(u_multiplier_STAGE3_acci_pp3_8_1__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_8_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_8_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_8_1__25_  (.A(u_multiplier_STAGE3_acci_pp3_8_1__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_8_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_8_1__16_ ));
 NAND2_X2 u_multiplier_STAGE3_acci_pp3_8_1__26_  (.A1(u_multiplier_STAGE3_acci_pp3_8_1__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_8_1__16_ ),
    .ZN(u_multiplier_pp3_8 [1]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_8_1__27_  (.A1(u_multiplier_pp2_8 [1]),
    .A2(u_multiplier_pp2_8 [0]),
    .B1(u_multiplier_pp2_8 [2]),
    .B2(u_multiplier_pp2_8 [3]),
    .ZN(u_multiplier_STAGE3_acci_pp3_8_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_8_1__28_  (.A1(u_multiplier_STAGE3_acci_pp3_8_1__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_8_1__17_ ),
    .ZN(u_multiplier_pp3_9 [2]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_9_0__21_  (.A1(u_multiplier_pp2_9 [5]),
    .A2(u_multiplier_pp2_9 [4]),
    .A3(u_multiplier_pp2_9 [6]),
    .ZN(u_multiplier_STAGE3_acci_pp3_9_0__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_9_0__22_  (.A(u_multiplier_pp2_9 [5]),
    .B(u_multiplier_pp2_9 [4]),
    .Z(u_multiplier_STAGE3_acci_pp3_9_0__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_9_0__23_  (.A(u_multiplier_pp2_9 [6]),
    .B(u_multiplier_pp2_9 [7]),
    .Z(u_multiplier_STAGE3_acci_pp3_9_0__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_9_0__24_  (.A1(u_multiplier_STAGE3_acci_pp3_9_0__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_9_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_9_0__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_9_0__25_  (.A(u_multiplier_STAGE3_acci_pp3_9_0__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_9_0__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_9_0__16_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_9_0__26_  (.A1(u_multiplier_STAGE3_acci_pp3_9_0__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_9_0__16_ ),
    .ZN(u_multiplier_pp3_9 [0]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_9_0__27_  (.A1(u_multiplier_pp2_9 [5]),
    .A2(u_multiplier_pp2_9 [4]),
    .B1(u_multiplier_pp2_9 [6]),
    .B2(u_multiplier_pp2_9 [7]),
    .ZN(u_multiplier_STAGE3_acci_pp3_9_0__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_9_0__28_  (.A1(u_multiplier_STAGE3_acci_pp3_9_0__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_9_0__17_ ),
    .ZN(u_multiplier_pp3_10 [3]));
 NAND3_X1 u_multiplier_STAGE3_acci_pp3_9_1__21_  (.A1(u_multiplier_pp2_9 [1]),
    .A2(u_multiplier_pp2_9 [0]),
    .A3(u_multiplier_pp2_9 [2]),
    .ZN(u_multiplier_STAGE3_acci_pp3_9_1__18_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_9_1__22_  (.A(u_multiplier_pp2_9 [1]),
    .B(u_multiplier_pp2_9 [0]),
    .Z(u_multiplier_STAGE3_acci_pp3_9_1__19_ ));
 XOR2_X2 u_multiplier_STAGE3_acci_pp3_9_1__23_  (.A(u_multiplier_pp2_9 [2]),
    .B(u_multiplier_pp2_9 [3]),
    .Z(u_multiplier_STAGE3_acci_pp3_9_1__20_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_9_1__24_  (.A1(u_multiplier_STAGE3_acci_pp3_9_1__19_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_9_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_9_1__15_ ));
 XNOR2_X1 u_multiplier_STAGE3_acci_pp3_9_1__25_  (.A(u_multiplier_STAGE3_acci_pp3_9_1__19_ ),
    .B(u_multiplier_STAGE3_acci_pp3_9_1__20_ ),
    .ZN(u_multiplier_STAGE3_acci_pp3_9_1__16_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_9_1__26_  (.A1(u_multiplier_STAGE3_acci_pp3_9_1__18_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_9_1__16_ ),
    .ZN(u_multiplier_pp3_9 [1]));
 AOI22_X1 u_multiplier_STAGE3_acci_pp3_9_1__27_  (.A1(u_multiplier_pp2_9 [1]),
    .A2(u_multiplier_pp2_9 [0]),
    .B1(u_multiplier_pp2_9 [2]),
    .B2(u_multiplier_pp2_9 [3]),
    .ZN(u_multiplier_STAGE3_acci_pp3_9_1__17_ ));
 NAND2_X1 u_multiplier_STAGE3_acci_pp3_9_1__28_  (.A1(u_multiplier_STAGE3_acci_pp3_9_1__15_ ),
    .A2(u_multiplier_STAGE3_acci_pp3_9_1__17_ ),
    .ZN(u_multiplier_pp3_10 [2]));
 LOGIC0_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__40__137  (.Z(net137));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_10__21_  (.A1(u_multiplier_pp3_10 [1]),
    .A2(u_multiplier_pp3_10 [0]),
    .A3(u_multiplier_pp3_10 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_10__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_10__22_  (.A(u_multiplier_pp3_10 [1]),
    .B(u_multiplier_pp3_10 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_10__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_10__23_  (.A(u_multiplier_pp3_10 [2]),
    .B(u_multiplier_pp3_10 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_10__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_10__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_10__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_10__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_10__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_10__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_10__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_10__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_10__16_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_10__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_10__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_10__16_ ),
    .ZN(u_multiplier_A [10]));
 AOI22_X1 u_multiplier_STAGE4_ACCI_pp4_10__27_  (.A1(u_multiplier_pp3_10 [1]),
    .A2(u_multiplier_pp3_10 [0]),
    .B1(u_multiplier_pp3_10 [2]),
    .B2(u_multiplier_pp3_10 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_10__17_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_10__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_10__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_10__17_ ),
    .ZN(u_multiplier_B [11]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_11__21_  (.A1(u_multiplier_pp3_11 [1]),
    .A2(u_multiplier_pp3_11 [0]),
    .A3(u_multiplier_pp3_11 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_11__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_11__22_  (.A(u_multiplier_pp3_11 [1]),
    .B(u_multiplier_pp3_11 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_11__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_11__23_  (.A(u_multiplier_pp3_11 [2]),
    .B(u_multiplier_pp3_11 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_11__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_11__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_11__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_11__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_11__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_11__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_11__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_11__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_11__16_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_11__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_11__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_11__16_ ),
    .ZN(u_multiplier_A [11]));
 AOI22_X1 u_multiplier_STAGE4_ACCI_pp4_11__27_  (.A1(u_multiplier_pp3_11 [1]),
    .A2(u_multiplier_pp3_11 [0]),
    .B1(u_multiplier_pp3_11 [2]),
    .B2(u_multiplier_pp3_11 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_11__17_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_11__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_11__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_11__17_ ),
    .ZN(u_multiplier_B [12]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_12__21_  (.A1(u_multiplier_pp3_12 [1]),
    .A2(u_multiplier_pp3_12 [0]),
    .A3(u_multiplier_pp3_12 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_12__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_12__22_  (.A(u_multiplier_pp3_12 [1]),
    .B(u_multiplier_pp3_12 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_12__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_12__23_  (.A(u_multiplier_pp3_12 [2]),
    .B(u_multiplier_pp3_12 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_12__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_12__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_12__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_12__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_12__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_12__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_12__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_12__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_12__16_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_12__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_12__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_12__16_ ),
    .ZN(u_multiplier_A [12]));
 AOI22_X2 u_multiplier_STAGE4_ACCI_pp4_12__27_  (.A1(u_multiplier_pp3_12 [1]),
    .A2(u_multiplier_pp3_12 [0]),
    .B1(u_multiplier_pp3_12 [2]),
    .B2(u_multiplier_pp3_12 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_12__17_ ));
 NAND2_X2 u_multiplier_STAGE4_ACCI_pp4_12__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_12__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_12__17_ ),
    .ZN(u_multiplier_B [13]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_13__21_  (.A1(u_multiplier_pp3_13 [1]),
    .A2(u_multiplier_pp3_13 [0]),
    .A3(u_multiplier_pp3_13 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_13__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_13__22_  (.A(u_multiplier_pp3_13 [1]),
    .B(u_multiplier_pp3_13 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_13__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_13__23_  (.A(u_multiplier_pp3_13 [2]),
    .B(u_multiplier_pp3_13 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_13__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_13__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_13__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_13__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_13__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_13__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_13__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_13__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_13__16_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_13__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_13__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_13__16_ ),
    .ZN(u_multiplier_A [13]));
 AOI22_X1 u_multiplier_STAGE4_ACCI_pp4_13__27_  (.A1(u_multiplier_pp3_13 [1]),
    .A2(u_multiplier_pp3_13 [0]),
    .B1(u_multiplier_pp3_13 [2]),
    .B2(u_multiplier_pp3_13 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_13__17_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_13__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_13__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_13__17_ ),
    .ZN(u_multiplier_B [14]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_14__21_  (.A1(u_multiplier_pp3_14 [1]),
    .A2(u_multiplier_pp3_14 [0]),
    .A3(u_multiplier_pp3_14 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_14__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_14__22_  (.A(u_multiplier_pp3_14 [1]),
    .B(u_multiplier_pp3_14 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_14__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_14__23_  (.A(u_multiplier_pp3_14 [2]),
    .B(u_multiplier_pp3_14 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_14__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_14__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_14__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_14__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_14__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_14__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_14__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_14__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_14__16_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_14__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_14__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_14__16_ ),
    .ZN(u_multiplier_A [14]));
 AOI22_X1 u_multiplier_STAGE4_ACCI_pp4_14__27_  (.A1(u_multiplier_pp3_14 [1]),
    .A2(u_multiplier_pp3_14 [0]),
    .B1(u_multiplier_pp3_14 [2]),
    .B2(u_multiplier_pp3_14 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_14__17_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_14__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_14__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_14__17_ ),
    .ZN(u_multiplier_B [15]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_15__21_  (.A1(u_multiplier_pp3_15 [1]),
    .A2(u_multiplier_pp3_15 [0]),
    .A3(u_multiplier_pp3_15 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_15__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_15__22_  (.A(u_multiplier_pp3_15 [1]),
    .B(u_multiplier_pp3_15 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_15__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_15__23_  (.A(u_multiplier_pp3_15 [2]),
    .B(u_multiplier_pp3_15 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_15__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_15__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_15__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_15__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_15__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_15__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_15__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_15__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_15__16_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_15__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_15__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_15__16_ ),
    .ZN(u_multiplier_A [15]));
 AOI22_X1 u_multiplier_STAGE4_ACCI_pp4_15__27_  (.A1(u_multiplier_pp3_15 [1]),
    .A2(u_multiplier_pp3_15 [0]),
    .B1(u_multiplier_pp3_15 [2]),
    .B2(u_multiplier_pp3_15 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_15__17_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_15__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_15__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_15__17_ ),
    .ZN(u_multiplier_B [16]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_16__21_  (.A1(u_multiplier_pp3_16 [1]),
    .A2(u_multiplier_pp3_16 [0]),
    .A3(u_multiplier_pp3_16 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_16__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_16__22_  (.A(u_multiplier_pp3_16 [1]),
    .B(u_multiplier_pp3_16 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_16__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_16__23_  (.A(u_multiplier_pp3_16 [2]),
    .B(u_multiplier_pp3_16 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_16__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_16__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_16__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_16__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_16__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_16__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_16__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_16__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_16__16_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_16__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_16__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_16__16_ ),
    .ZN(u_multiplier_A [16]));
 AOI22_X1 u_multiplier_STAGE4_ACCI_pp4_16__27_  (.A1(u_multiplier_pp3_16 [1]),
    .A2(u_multiplier_pp3_16 [0]),
    .B1(u_multiplier_pp3_16 [2]),
    .B2(u_multiplier_pp3_16 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_16__17_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_16__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_16__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_16__17_ ),
    .ZN(u_multiplier_B [17]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_17__21_  (.A1(u_multiplier_pp3_17 [1]),
    .A2(u_multiplier_pp3_17 [0]),
    .A3(u_multiplier_pp3_17 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_17__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_17__22_  (.A(u_multiplier_pp3_17 [1]),
    .B(u_multiplier_pp3_17 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_17__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_17__23_  (.A(u_multiplier_pp3_17 [2]),
    .B(u_multiplier_pp3_17 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_17__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_17__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_17__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_17__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_17__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_17__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_17__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_17__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_17__16_ ));
 NAND2_X2 u_multiplier_STAGE4_ACCI_pp4_17__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_17__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_17__16_ ),
    .ZN(u_multiplier_A [17]));
 AOI22_X1 u_multiplier_STAGE4_ACCI_pp4_17__27_  (.A1(u_multiplier_pp3_17 [1]),
    .A2(u_multiplier_pp3_17 [0]),
    .B1(u_multiplier_pp3_17 [2]),
    .B2(u_multiplier_pp3_17 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_17__17_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_17__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_17__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_17__17_ ),
    .ZN(u_multiplier_B [18]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_18__21_  (.A1(u_multiplier_pp3_18 [1]),
    .A2(u_multiplier_pp3_18 [0]),
    .A3(u_multiplier_pp3_18 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_18__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_18__22_  (.A(u_multiplier_pp3_18 [1]),
    .B(u_multiplier_pp3_18 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_18__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_18__23_  (.A(u_multiplier_pp3_18 [2]),
    .B(u_multiplier_pp3_18 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_18__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_18__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_18__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_18__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_18__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_18__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_18__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_18__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_18__16_ ));
 NAND2_X2 u_multiplier_STAGE4_ACCI_pp4_18__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_18__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_18__16_ ),
    .ZN(u_multiplier_A [18]));
 AOI22_X1 u_multiplier_STAGE4_ACCI_pp4_18__27_  (.A1(u_multiplier_pp3_18 [1]),
    .A2(u_multiplier_pp3_18 [0]),
    .B1(u_multiplier_pp3_18 [2]),
    .B2(u_multiplier_pp3_18 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_18__17_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_18__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_18__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_18__17_ ),
    .ZN(u_multiplier_B [19]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_19__21_  (.A1(u_multiplier_pp3_19 [1]),
    .A2(u_multiplier_pp3_19 [0]),
    .A3(u_multiplier_pp3_19 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_19__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_19__22_  (.A(u_multiplier_pp3_19 [1]),
    .B(u_multiplier_pp3_19 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_19__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_19__23_  (.A(u_multiplier_pp3_19 [2]),
    .B(u_multiplier_pp3_19 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_19__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_19__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_19__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_19__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_19__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_19__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_19__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_19__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_19__16_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_19__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_19__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_19__16_ ),
    .ZN(u_multiplier_A [19]));
 AOI22_X1 u_multiplier_STAGE4_ACCI_pp4_19__27_  (.A1(u_multiplier_pp3_19 [1]),
    .A2(u_multiplier_pp3_19 [0]),
    .B1(u_multiplier_pp3_19 [2]),
    .B2(u_multiplier_pp3_19 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_19__17_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_19__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_19__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_19__17_ ),
    .ZN(u_multiplier_B [20]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_20__21_  (.A1(u_multiplier_pp3_20 [1]),
    .A2(u_multiplier_pp3_20 [0]),
    .A3(u_multiplier_pp3_20 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_20__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_20__22_  (.A(u_multiplier_pp3_20 [1]),
    .B(u_multiplier_pp3_20 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_20__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_20__23_  (.A(u_multiplier_pp3_20 [2]),
    .B(u_multiplier_pp3_20 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_20__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_20__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_20__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_20__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_20__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_20__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_20__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_20__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_20__16_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_20__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_20__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_20__16_ ),
    .ZN(u_multiplier_A [20]));
 AOI22_X2 u_multiplier_STAGE4_ACCI_pp4_20__27_  (.A1(u_multiplier_pp3_20 [1]),
    .A2(u_multiplier_pp3_20 [0]),
    .B1(u_multiplier_pp3_20 [2]),
    .B2(u_multiplier_pp3_20 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_20__17_ ));
 NAND2_X2 u_multiplier_STAGE4_ACCI_pp4_20__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_20__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_20__17_ ),
    .ZN(u_multiplier_B [21]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_21__21_  (.A1(u_multiplier_pp3_21 [1]),
    .A2(u_multiplier_pp3_21 [0]),
    .A3(u_multiplier_pp3_21 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_21__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_21__22_  (.A(u_multiplier_pp3_21 [1]),
    .B(u_multiplier_pp3_21 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_21__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_21__23_  (.A(u_multiplier_pp3_21 [2]),
    .B(u_multiplier_pp3_21 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_21__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_21__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_21__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_21__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_21__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_21__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_21__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_21__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_21__16_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_21__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_21__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_21__16_ ),
    .ZN(u_multiplier_A [21]));
 AOI22_X1 u_multiplier_STAGE4_ACCI_pp4_21__27_  (.A1(u_multiplier_pp3_21 [1]),
    .A2(u_multiplier_pp3_21 [0]),
    .B1(u_multiplier_pp3_21 [2]),
    .B2(u_multiplier_pp3_21 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_21__17_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_21__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_21__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_21__17_ ),
    .ZN(u_multiplier_B [22]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_22__21_  (.A1(u_multiplier_pp3_22 [1]),
    .A2(u_multiplier_pp3_22 [0]),
    .A3(u_multiplier_pp3_22 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_22__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_22__22_  (.A(u_multiplier_pp3_22 [1]),
    .B(u_multiplier_pp3_22 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_22__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_22__23_  (.A(u_multiplier_pp3_22 [2]),
    .B(u_multiplier_pp3_22 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_22__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_22__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_22__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_22__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_22__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_22__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_22__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_22__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_22__16_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_22__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_22__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_22__16_ ),
    .ZN(u_multiplier_A [22]));
 AOI22_X1 u_multiplier_STAGE4_ACCI_pp4_22__27_  (.A1(u_multiplier_pp3_22 [1]),
    .A2(u_multiplier_pp3_22 [0]),
    .B1(u_multiplier_pp3_22 [2]),
    .B2(u_multiplier_pp3_22 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_22__17_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_22__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_22__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_22__17_ ),
    .ZN(u_multiplier_B [23]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_23__21_  (.A1(u_multiplier_pp3_23 [1]),
    .A2(u_multiplier_pp3_23 [0]),
    .A3(u_multiplier_pp3_23 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_23__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_23__22_  (.A(u_multiplier_pp3_23 [1]),
    .B(u_multiplier_pp3_23 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_23__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_23__23_  (.A(u_multiplier_pp3_23 [2]),
    .B(u_multiplier_pp3_23 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_23__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_23__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_23__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_23__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_23__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_23__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_23__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_23__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_23__16_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_23__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_23__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_23__16_ ),
    .ZN(u_multiplier_A [23]));
 AOI22_X1 u_multiplier_STAGE4_ACCI_pp4_23__27_  (.A1(u_multiplier_pp3_23 [1]),
    .A2(u_multiplier_pp3_23 [0]),
    .B1(u_multiplier_pp3_23 [2]),
    .B2(u_multiplier_pp3_23 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_23__17_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_23__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_23__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_23__17_ ),
    .ZN(u_multiplier_B [24]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_24__21_  (.A1(u_multiplier_pp3_24 [1]),
    .A2(u_multiplier_pp3_24 [0]),
    .A3(u_multiplier_pp3_24 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_24__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_24__22_  (.A(u_multiplier_pp3_24 [1]),
    .B(u_multiplier_pp3_24 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_24__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_24__23_  (.A(u_multiplier_pp3_24 [2]),
    .B(u_multiplier_pp3_24 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_24__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_24__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_24__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_24__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_24__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_24__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_24__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_24__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_24__16_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_24__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_24__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_24__16_ ),
    .ZN(u_multiplier_A [24]));
 AOI22_X1 u_multiplier_STAGE4_ACCI_pp4_24__27_  (.A1(u_multiplier_pp3_24 [1]),
    .A2(u_multiplier_pp3_24 [0]),
    .B1(u_multiplier_pp3_24 [2]),
    .B2(u_multiplier_pp3_24 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_24__17_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_24__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_24__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_24__17_ ),
    .ZN(u_multiplier_B [25]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_25__21_  (.A1(u_multiplier_pp3_25 [1]),
    .A2(u_multiplier_pp3_25 [0]),
    .A3(u_multiplier_pp3_25 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_25__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_25__22_  (.A(u_multiplier_pp3_25 [1]),
    .B(u_multiplier_pp3_25 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_25__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_25__23_  (.A(u_multiplier_pp3_25 [2]),
    .B(u_multiplier_pp3_25 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_25__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_25__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_25__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_25__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_25__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_25__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_25__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_25__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_25__16_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_25__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_25__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_25__16_ ),
    .ZN(u_multiplier_A [25]));
 AOI22_X1 u_multiplier_STAGE4_ACCI_pp4_25__27_  (.A1(u_multiplier_pp3_25 [1]),
    .A2(u_multiplier_pp3_25 [0]),
    .B1(u_multiplier_pp3_25 [2]),
    .B2(u_multiplier_pp3_25 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_25__17_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_25__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_25__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_25__17_ ),
    .ZN(u_multiplier_B [26]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_26__21_  (.A1(u_multiplier_pp3_26 [1]),
    .A2(u_multiplier_pp3_26 [0]),
    .A3(u_multiplier_pp3_26 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_26__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_26__22_  (.A(u_multiplier_pp3_26 [1]),
    .B(u_multiplier_pp3_26 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_26__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_26__23_  (.A(u_multiplier_pp3_26 [2]),
    .B(u_multiplier_pp3_26 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_26__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_26__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_26__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_26__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_26__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_26__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_26__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_26__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_26__16_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_26__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_26__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_26__16_ ),
    .ZN(u_multiplier_A [26]));
 AOI22_X1 u_multiplier_STAGE4_ACCI_pp4_26__27_  (.A1(u_multiplier_pp3_26 [1]),
    .A2(u_multiplier_pp3_26 [0]),
    .B1(u_multiplier_pp3_26 [2]),
    .B2(u_multiplier_pp3_26 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_26__17_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_26__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_26__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_26__17_ ),
    .ZN(u_multiplier_B [27]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_27__21_  (.A1(u_multiplier_pp3_27 [1]),
    .A2(u_multiplier_pp3_27 [0]),
    .A3(u_multiplier_pp3_27 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_27__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_27__22_  (.A(u_multiplier_pp3_27 [1]),
    .B(u_multiplier_pp3_27 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_27__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_27__23_  (.A(u_multiplier_pp3_27 [2]),
    .B(u_multiplier_pp3_27 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_27__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_27__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_27__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_27__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_27__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_27__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_27__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_27__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_27__16_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_27__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_27__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_27__16_ ),
    .ZN(u_multiplier_A [27]));
 AOI22_X1 u_multiplier_STAGE4_ACCI_pp4_27__27_  (.A1(u_multiplier_pp3_27 [1]),
    .A2(u_multiplier_pp3_27 [0]),
    .B1(u_multiplier_pp3_27 [2]),
    .B2(u_multiplier_pp3_27 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_27__17_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_27__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_27__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_27__17_ ),
    .ZN(u_multiplier_B [28]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_28__21_  (.A1(u_multiplier_pp3_28 [1]),
    .A2(u_multiplier_pp3_28 [0]),
    .A3(u_multiplier_pp3_28 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_28__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_28__22_  (.A(u_multiplier_pp3_28 [1]),
    .B(u_multiplier_pp3_28 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_28__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_28__23_  (.A(u_multiplier_pp3_28 [2]),
    .B(u_multiplier_pp3_28 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_28__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_28__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_28__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_28__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_28__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_28__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_28__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_28__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_28__16_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_28__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_28__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_28__16_ ),
    .ZN(u_multiplier_A [28]));
 AOI22_X1 u_multiplier_STAGE4_ACCI_pp4_28__27_  (.A1(u_multiplier_pp3_28 [1]),
    .A2(u_multiplier_pp3_28 [0]),
    .B1(u_multiplier_pp3_28 [2]),
    .B2(u_multiplier_pp3_28 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_28__17_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_28__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_28__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_28__17_ ),
    .ZN(u_multiplier_B [29]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_29__21_  (.A1(u_multiplier_pp3_29 [1]),
    .A2(u_multiplier_pp3_29 [0]),
    .A3(u_multiplier_pp3_29 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_29__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_29__22_  (.A(u_multiplier_pp3_29 [1]),
    .B(u_multiplier_pp3_29 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_29__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_29__23_  (.A(u_multiplier_pp3_29 [2]),
    .B(u_multiplier_pp3_29 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_29__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_29__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_29__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_29__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_29__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_29__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_29__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_29__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_29__16_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_29__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_29__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_29__16_ ),
    .ZN(u_multiplier_A [29]));
 AOI22_X1 u_multiplier_STAGE4_ACCI_pp4_29__27_  (.A1(u_multiplier_pp3_29 [1]),
    .A2(u_multiplier_pp3_29 [0]),
    .B1(u_multiplier_pp3_29 [2]),
    .B2(u_multiplier_pp3_29 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_29__17_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_29__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_29__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_29__17_ ),
    .ZN(u_multiplier_B [30]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_3__21_  (.A1(u_multiplier_pp3_3 [1]),
    .A2(u_multiplier_pp3_3 [0]),
    .A3(u_multiplier_pp3_3 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_3__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_3__22_  (.A(u_multiplier_pp3_3 [1]),
    .B(u_multiplier_pp3_3 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_3__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_3__23_  (.A(u_multiplier_pp3_3 [2]),
    .B(u_multiplier_pp3_3 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_3__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_3__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_3__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_3__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_3__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_3__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_3__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_3__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_3__16_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_3__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_3__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_3__16_ ),
    .ZN(u_multiplier_A [3]));
 AOI22_X4 u_multiplier_STAGE4_ACCI_pp4_3__27_  (.A1(u_multiplier_pp3_3 [1]),
    .A2(u_multiplier_pp3_3 [0]),
    .B1(u_multiplier_pp3_3 [2]),
    .B2(u_multiplier_pp3_3 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_3__17_ ));
 NAND2_X4 u_multiplier_STAGE4_ACCI_pp4_3__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_3__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_3__17_ ),
    .ZN(u_multiplier_B [4]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_30__21_  (.A1(u_multiplier_pp3_30 [1]),
    .A2(u_multiplier_pp3_30 [0]),
    .A3(u_multiplier_pp3_30 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_30__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_30__22_  (.A(u_multiplier_pp3_30 [1]),
    .B(u_multiplier_pp3_30 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_30__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_30__23_  (.A(u_multiplier_pp3_30 [2]),
    .B(u_multiplier_pp3_30 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_30__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_30__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_30__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_30__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_30__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_30__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_30__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_30__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_30__16_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_30__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_30__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_30__16_ ),
    .ZN(u_multiplier_A [30]));
 AOI22_X1 u_multiplier_STAGE4_ACCI_pp4_30__27_  (.A1(u_multiplier_pp3_30 [1]),
    .A2(u_multiplier_pp3_30 [0]),
    .B1(u_multiplier_pp3_30 [2]),
    .B2(u_multiplier_pp3_30 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_30__17_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_30__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_30__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_30__17_ ),
    .ZN(u_multiplier_B [31]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_31__21_  (.A1(u_multiplier_pp3_31 [1]),
    .A2(u_multiplier_pp3_31 [0]),
    .A3(u_multiplier_pp3_31 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_31__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_31__22_  (.A(u_multiplier_pp3_31 [1]),
    .B(u_multiplier_pp3_31 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_31__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_31__23_  (.A(u_multiplier_pp3_31 [2]),
    .B(u_multiplier_pp3_31 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_31__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_31__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_31__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_31__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_31__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_31__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_31__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_31__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_31__16_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_31__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_31__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_31__16_ ),
    .ZN(u_multiplier_A [31]));
 AOI22_X1 u_multiplier_STAGE4_ACCI_pp4_31__27_  (.A1(u_multiplier_pp3_31 [1]),
    .A2(u_multiplier_pp3_31 [0]),
    .B1(u_multiplier_pp3_31 [2]),
    .B2(u_multiplier_pp3_31 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_31__17_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_31__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_31__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_31__17_ ),
    .ZN(u_multiplier_B [32]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_4__21_  (.A1(u_multiplier_pp3_4 [1]),
    .A2(u_multiplier_pp3_4 [0]),
    .A3(u_multiplier_pp3_4 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_4__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_4__22_  (.A(u_multiplier_pp3_4 [1]),
    .B(u_multiplier_pp3_4 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_4__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_4__23_  (.A(u_multiplier_pp3_4 [2]),
    .B(u_multiplier_pp3_4 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_4__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_4__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_4__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_4__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_4__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_4__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_4__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_4__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_4__16_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_4__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_4__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_4__16_ ),
    .ZN(u_multiplier_A [4]));
 AOI22_X1 u_multiplier_STAGE4_ACCI_pp4_4__27_  (.A1(u_multiplier_pp3_4 [1]),
    .A2(u_multiplier_pp3_4 [0]),
    .B1(u_multiplier_pp3_4 [2]),
    .B2(u_multiplier_pp3_4 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_4__17_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_4__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_4__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_4__17_ ),
    .ZN(u_multiplier_B [5]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_5__21_  (.A1(u_multiplier_pp3_5 [1]),
    .A2(u_multiplier_pp3_5 [0]),
    .A3(u_multiplier_pp3_5 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_5__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_5__22_  (.A(u_multiplier_pp3_5 [1]),
    .B(u_multiplier_pp3_5 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_5__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_5__23_  (.A(u_multiplier_pp3_5 [2]),
    .B(u_multiplier_pp3_5 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_5__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_5__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_5__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_5__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_5__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_5__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_5__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_5__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_5__16_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_5__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_5__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_5__16_ ),
    .ZN(u_multiplier_A [5]));
 AOI22_X1 u_multiplier_STAGE4_ACCI_pp4_5__27_  (.A1(u_multiplier_pp3_5 [1]),
    .A2(u_multiplier_pp3_5 [0]),
    .B1(u_multiplier_pp3_5 [2]),
    .B2(u_multiplier_pp3_5 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_5__17_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_5__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_5__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_5__17_ ),
    .ZN(u_multiplier_B [6]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_6__21_  (.A1(u_multiplier_pp3_6 [1]),
    .A2(u_multiplier_pp3_6 [0]),
    .A3(u_multiplier_pp3_6 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_6__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_6__22_  (.A(u_multiplier_pp3_6 [1]),
    .B(u_multiplier_pp3_6 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_6__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_6__23_  (.A(u_multiplier_pp3_6 [2]),
    .B(u_multiplier_pp3_6 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_6__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_6__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_6__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_6__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_6__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_6__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_6__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_6__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_6__16_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_6__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_6__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_6__16_ ),
    .ZN(u_multiplier_A [6]));
 AOI22_X1 u_multiplier_STAGE4_ACCI_pp4_6__27_  (.A1(u_multiplier_pp3_6 [1]),
    .A2(u_multiplier_pp3_6 [0]),
    .B1(u_multiplier_pp3_6 [2]),
    .B2(u_multiplier_pp3_6 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_6__17_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_6__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_6__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_6__17_ ),
    .ZN(u_multiplier_B [7]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_7__21_  (.A1(u_multiplier_pp3_7 [1]),
    .A2(u_multiplier_pp3_7 [0]),
    .A3(u_multiplier_pp3_7 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_7__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_7__22_  (.A(u_multiplier_pp3_7 [1]),
    .B(u_multiplier_pp3_7 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_7__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_7__23_  (.A(u_multiplier_pp3_7 [2]),
    .B(u_multiplier_pp3_7 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_7__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_7__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_7__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_7__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_7__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_7__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_7__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_7__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_7__16_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_7__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_7__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_7__16_ ),
    .ZN(u_multiplier_A [7]));
 AOI22_X1 u_multiplier_STAGE4_ACCI_pp4_7__27_  (.A1(u_multiplier_pp3_7 [1]),
    .A2(u_multiplier_pp3_7 [0]),
    .B1(u_multiplier_pp3_7 [2]),
    .B2(u_multiplier_pp3_7 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_7__17_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_7__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_7__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_7__17_ ),
    .ZN(u_multiplier_B [8]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_8__21_  (.A1(u_multiplier_pp3_8 [1]),
    .A2(u_multiplier_pp3_8 [0]),
    .A3(u_multiplier_pp3_8 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_8__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_8__22_  (.A(u_multiplier_pp3_8 [1]),
    .B(u_multiplier_pp3_8 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_8__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_8__23_  (.A(u_multiplier_pp3_8 [2]),
    .B(u_multiplier_pp3_8 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_8__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_8__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_8__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_8__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_8__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_8__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_8__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_8__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_8__16_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_8__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_8__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_8__16_ ),
    .ZN(u_multiplier_A [8]));
 AOI22_X1 u_multiplier_STAGE4_ACCI_pp4_8__27_  (.A1(u_multiplier_pp3_8 [1]),
    .A2(u_multiplier_pp3_8 [0]),
    .B1(u_multiplier_pp3_8 [2]),
    .B2(u_multiplier_pp3_8 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_8__17_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_8__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_8__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_8__17_ ),
    .ZN(u_multiplier_B [9]));
 NAND3_X1 u_multiplier_STAGE4_ACCI_pp4_9__21_  (.A1(u_multiplier_pp3_9 [1]),
    .A2(u_multiplier_pp3_9 [0]),
    .A3(u_multiplier_pp3_9 [2]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_9__18_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_9__22_  (.A(u_multiplier_pp3_9 [1]),
    .B(u_multiplier_pp3_9 [0]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_9__19_ ));
 XOR2_X2 u_multiplier_STAGE4_ACCI_pp4_9__23_  (.A(u_multiplier_pp3_9 [2]),
    .B(u_multiplier_pp3_9 [3]),
    .Z(u_multiplier_STAGE4_ACCI_pp4_9__20_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_9__24_  (.A1(u_multiplier_STAGE4_ACCI_pp4_9__19_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_9__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_9__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_ACCI_pp4_9__25_  (.A(u_multiplier_STAGE4_ACCI_pp4_9__19_ ),
    .B(u_multiplier_STAGE4_ACCI_pp4_9__20_ ),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_9__16_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_9__26_  (.A1(u_multiplier_STAGE4_ACCI_pp4_9__18_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_9__16_ ),
    .ZN(u_multiplier_A [9]));
 AOI22_X1 u_multiplier_STAGE4_ACCI_pp4_9__27_  (.A1(u_multiplier_pp3_9 [1]),
    .A2(u_multiplier_pp3_9 [0]),
    .B1(u_multiplier_pp3_9 [2]),
    .B2(u_multiplier_pp3_9 [3]),
    .ZN(u_multiplier_STAGE4_ACCI_pp4_9__17_ ));
 NAND2_X1 u_multiplier_STAGE4_ACCI_pp4_9__28_  (.A1(u_multiplier_STAGE4_ACCI_pp4_9__15_ ),
    .A2(u_multiplier_STAGE4_ACCI_pp4_9__17_ ),
    .ZN(u_multiplier_B [10]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_32__18_  (.A(net140),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_32__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_32__19_  (.A1(u_multiplier_pp3_32 [1]),
    .A2(u_multiplier_pp3_32 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_32__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_32__20_  (.A(u_multiplier_pp3_32 [1]),
    .B(u_multiplier_pp3_32 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_32__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_32__21_  (.A1(u_multiplier_pp3_32 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_32__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_32__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_32__22_  (.A(u_multiplier_pp3_32 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_32__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_32__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_32__23_  (.A1(u_multiplier_pp3_32 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_32__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_32__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_32__24_  (.A(u_multiplier_pp3_32 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_32__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_32__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_32__25_  (.A(net141),
    .B(u_multiplier_STAGE4_E_4_2_pp4_32__16_ ),
    .ZN(u_multiplier_A [32]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_32__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_32__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_32__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_32_c2 ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_32__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_32__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_32__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_32__17_ ),
    .ZN(u_multiplier_B [33]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_33__18_  (.A(u_multiplier_STAGE4_pp4_32_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_33__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_33__19_  (.A1(u_multiplier_pp3_33 [1]),
    .A2(u_multiplier_pp3_33 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_33__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_33__20_  (.A(u_multiplier_pp3_33 [1]),
    .B(u_multiplier_pp3_33 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_33__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_33__21_  (.A1(u_multiplier_pp3_33 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_33__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_33__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_33__22_  (.A(u_multiplier_pp3_33 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_33__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_33__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_33__23_  (.A1(u_multiplier_pp3_33 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_33__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_33__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_33__24_  (.A(u_multiplier_pp3_33 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_33__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_33__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_33__25_  (.A(u_multiplier_STAGE4_pp4_32_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_33__16_ ),
    .ZN(u_multiplier_A [33]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_33__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_33__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_33__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_33_c2 ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_33__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_33__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_33__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_33__17_ ),
    .ZN(u_multiplier_B [34]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_34__18_  (.A(u_multiplier_STAGE4_pp4_33_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_34__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_34__19_  (.A1(u_multiplier_pp3_34 [1]),
    .A2(u_multiplier_pp3_34 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_34__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_34__20_  (.A(u_multiplier_pp3_34 [1]),
    .B(u_multiplier_pp3_34 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_34__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_34__21_  (.A1(u_multiplier_pp3_34 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_34__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_34__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_34__22_  (.A(u_multiplier_pp3_34 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_34__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_34__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_34__23_  (.A1(u_multiplier_pp3_34 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_34__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_34__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_34__24_  (.A(u_multiplier_pp3_34 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_34__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_34__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_34__25_  (.A(u_multiplier_STAGE4_pp4_33_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_34__16_ ),
    .ZN(u_multiplier_A [34]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_34__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_34__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_34__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_34_c2 ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_34__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_34__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_34__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_34__17_ ),
    .ZN(u_multiplier_B [35]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_35__18_  (.A(u_multiplier_STAGE4_pp4_34_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_35__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_35__19_  (.A1(u_multiplier_pp3_35 [1]),
    .A2(u_multiplier_pp3_35 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_35__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_35__20_  (.A(u_multiplier_pp3_35 [1]),
    .B(u_multiplier_pp3_35 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_35__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_35__21_  (.A1(u_multiplier_pp3_35 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_35__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_35__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_35__22_  (.A(u_multiplier_pp3_35 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_35__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_35__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_35__23_  (.A1(u_multiplier_pp3_35 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_35__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_35__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_35__24_  (.A(u_multiplier_pp3_35 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_35__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_35__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_35__25_  (.A(u_multiplier_STAGE4_pp4_34_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_35__16_ ),
    .ZN(u_multiplier_A [35]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_35__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_35__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_35__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_35_c2 ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_35__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_35__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_35__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_35__17_ ),
    .ZN(u_multiplier_B [36]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_36__18_  (.A(u_multiplier_STAGE4_pp4_35_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_36__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_36__19_  (.A1(u_multiplier_pp3_36 [1]),
    .A2(u_multiplier_pp3_36 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_36__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_36__20_  (.A(u_multiplier_pp3_36 [1]),
    .B(u_multiplier_pp3_36 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_36__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_36__21_  (.A1(u_multiplier_pp3_36 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_36__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_36__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_36__22_  (.A(u_multiplier_pp3_36 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_36__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_36__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_36__23_  (.A1(u_multiplier_pp3_36 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_36__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_36__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_36__24_  (.A(u_multiplier_pp3_36 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_36__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_36__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_36__25_  (.A(u_multiplier_STAGE4_pp4_35_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_36__16_ ),
    .ZN(u_multiplier_A [36]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_36__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_36__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_36__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_36_c2 ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_36__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_36__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_36__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_36__17_ ),
    .ZN(u_multiplier_B [37]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_37__18_  (.A(u_multiplier_STAGE4_pp4_36_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_37__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_37__19_  (.A1(u_multiplier_pp3_37 [1]),
    .A2(u_multiplier_pp3_37 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_37__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_37__20_  (.A(u_multiplier_pp3_37 [1]),
    .B(u_multiplier_pp3_37 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_37__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_37__21_  (.A1(u_multiplier_pp3_37 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_37__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_37__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_37__22_  (.A(u_multiplier_pp3_37 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_37__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_37__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_37__23_  (.A1(u_multiplier_pp3_37 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_37__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_37__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_37__24_  (.A(u_multiplier_pp3_37 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_37__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_37__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_37__25_  (.A(u_multiplier_STAGE4_pp4_36_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_37__16_ ),
    .ZN(u_multiplier_A [37]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_37__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_37__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_37__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_37_c2 ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_37__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_37__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_37__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_37__17_ ),
    .ZN(u_multiplier_B [38]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_38__18_  (.A(u_multiplier_STAGE4_pp4_37_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_38__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_38__19_  (.A1(u_multiplier_pp3_38 [1]),
    .A2(u_multiplier_pp3_38 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_38__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_38__20_  (.A(u_multiplier_pp3_38 [1]),
    .B(u_multiplier_pp3_38 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_38__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_38__21_  (.A1(u_multiplier_pp3_38 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_38__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_38__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_38__22_  (.A(u_multiplier_pp3_38 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_38__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_38__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_38__23_  (.A1(u_multiplier_pp3_38 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_38__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_38__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_38__24_  (.A(u_multiplier_pp3_38 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_38__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_38__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_38__25_  (.A(u_multiplier_STAGE4_pp4_37_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_38__16_ ),
    .ZN(u_multiplier_A [38]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_38__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_38__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_38__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_38_c2 ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_38__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_38__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_38__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_38__17_ ),
    .ZN(u_multiplier_B [39]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_39__18_  (.A(u_multiplier_STAGE4_pp4_38_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_39__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_39__19_  (.A1(u_multiplier_pp3_39 [1]),
    .A2(u_multiplier_pp3_39 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_39__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_39__20_  (.A(u_multiplier_pp3_39 [1]),
    .B(u_multiplier_pp3_39 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_39__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_39__21_  (.A1(u_multiplier_pp3_39 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_39__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_39__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_39__22_  (.A(u_multiplier_pp3_39 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_39__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_39__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_39__23_  (.A1(u_multiplier_pp3_39 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_39__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_39__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_39__24_  (.A(u_multiplier_pp3_39 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_39__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_39__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_39__25_  (.A(u_multiplier_STAGE4_pp4_38_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_39__16_ ),
    .ZN(u_multiplier_A [39]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_39__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_39__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_39__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_39_c2 ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_39__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_39__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_39__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_39__17_ ),
    .ZN(u_multiplier_B [40]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_40__18_  (.A(u_multiplier_STAGE4_pp4_39_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_40__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_40__19_  (.A1(u_multiplier_pp3_40 [1]),
    .A2(u_multiplier_pp3_40 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_40__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_40__20_  (.A(u_multiplier_pp3_40 [1]),
    .B(u_multiplier_pp3_40 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_40__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_40__21_  (.A1(u_multiplier_pp3_40 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_40__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_40__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_40__22_  (.A(u_multiplier_pp3_40 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_40__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_40__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_40__23_  (.A1(u_multiplier_pp3_40 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_40__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_40__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_40__24_  (.A(u_multiplier_pp3_40 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_40__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_40__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_40__25_  (.A(u_multiplier_STAGE4_pp4_39_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_40__16_ ),
    .ZN(u_multiplier_A [40]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_40__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_40__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_40__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_40_c2 ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_40__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_40__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_40__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_40__17_ ),
    .ZN(u_multiplier_B [41]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_41__18_  (.A(u_multiplier_STAGE4_pp4_40_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_41__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_41__19_  (.A1(u_multiplier_pp3_41 [1]),
    .A2(u_multiplier_pp3_41 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_41__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_41__20_  (.A(u_multiplier_pp3_41 [1]),
    .B(u_multiplier_pp3_41 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_41__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_41__21_  (.A1(u_multiplier_pp3_41 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_41__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_41__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_41__22_  (.A(u_multiplier_pp3_41 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_41__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_41__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_41__23_  (.A1(u_multiplier_pp3_41 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_41__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_41__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_41__24_  (.A(u_multiplier_pp3_41 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_41__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_41__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_41__25_  (.A(u_multiplier_STAGE4_pp4_40_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_41__16_ ),
    .ZN(u_multiplier_A [41]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_41__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_41__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_41__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_41_c2 ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_41__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_41__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_41__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_41__17_ ),
    .ZN(u_multiplier_B [42]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_42__18_  (.A(u_multiplier_STAGE4_pp4_41_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_42__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_42__19_  (.A1(u_multiplier_pp3_42 [1]),
    .A2(u_multiplier_pp3_42 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_42__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_42__20_  (.A(u_multiplier_pp3_42 [1]),
    .B(u_multiplier_pp3_42 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_42__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_42__21_  (.A1(u_multiplier_pp3_42 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_42__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_42__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_42__22_  (.A(u_multiplier_pp3_42 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_42__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_42__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_42__23_  (.A1(u_multiplier_pp3_42 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_42__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_42__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_42__24_  (.A(u_multiplier_pp3_42 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_42__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_42__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_42__25_  (.A(u_multiplier_STAGE4_pp4_41_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_42__16_ ),
    .ZN(u_multiplier_A [42]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_42__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_42__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_42__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_42_c2 ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_42__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_42__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_42__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_42__17_ ),
    .ZN(u_multiplier_B [43]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_43__18_  (.A(u_multiplier_STAGE4_pp4_42_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_43__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_43__19_  (.A1(u_multiplier_pp3_43 [1]),
    .A2(u_multiplier_pp3_43 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_43__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_43__20_  (.A(u_multiplier_pp3_43 [1]),
    .B(u_multiplier_pp3_43 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_43__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_43__21_  (.A1(u_multiplier_pp3_43 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_43__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_43__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_43__22_  (.A(u_multiplier_pp3_43 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_43__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_43__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_43__23_  (.A1(u_multiplier_pp3_43 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_43__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_43__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_43__24_  (.A(u_multiplier_pp3_43 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_43__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_43__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_43__25_  (.A(u_multiplier_STAGE4_pp4_42_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_43__16_ ),
    .ZN(u_multiplier_A [43]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_43__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_43__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_43__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_43_c2 ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_43__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_43__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_43__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_43__17_ ),
    .ZN(u_multiplier_B [44]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_44__18_  (.A(u_multiplier_STAGE4_pp4_43_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_44__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_44__19_  (.A1(u_multiplier_pp3_44 [1]),
    .A2(u_multiplier_pp3_44 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_44__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_44__20_  (.A(u_multiplier_pp3_44 [1]),
    .B(u_multiplier_pp3_44 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_44__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_44__21_  (.A1(u_multiplier_pp3_44 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_44__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_44__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_44__22_  (.A(u_multiplier_pp3_44 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_44__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_44__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_44__23_  (.A1(u_multiplier_pp3_44 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_44__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_44__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_44__24_  (.A(u_multiplier_pp3_44 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_44__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_44__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_44__25_  (.A(u_multiplier_STAGE4_pp4_43_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_44__16_ ),
    .ZN(u_multiplier_A [44]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_44__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_44__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_44__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_44_c2 ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_44__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_44__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_44__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_44__17_ ),
    .ZN(u_multiplier_B [45]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_45__18_  (.A(u_multiplier_STAGE4_pp4_44_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_45__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_45__19_  (.A1(u_multiplier_pp3_45 [1]),
    .A2(u_multiplier_pp3_45 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_45__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_45__20_  (.A(u_multiplier_pp3_45 [1]),
    .B(u_multiplier_pp3_45 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_45__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_45__21_  (.A1(u_multiplier_pp3_45 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_45__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_45__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_45__22_  (.A(u_multiplier_pp3_45 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_45__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_45__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_45__23_  (.A1(u_multiplier_pp3_45 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_45__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_45__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_45__24_  (.A(u_multiplier_pp3_45 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_45__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_45__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_45__25_  (.A(u_multiplier_STAGE4_pp4_44_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_45__16_ ),
    .ZN(u_multiplier_A [45]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_45__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_45__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_45__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_45_c2 ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_45__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_45__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_45__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_45__17_ ),
    .ZN(u_multiplier_B [46]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_46__18_  (.A(u_multiplier_STAGE4_pp4_45_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_46__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_46__19_  (.A1(u_multiplier_pp3_46 [1]),
    .A2(u_multiplier_pp3_46 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_46__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_46__20_  (.A(u_multiplier_pp3_46 [1]),
    .B(u_multiplier_pp3_46 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_46__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_46__21_  (.A1(u_multiplier_pp3_46 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_46__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_46__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_46__22_  (.A(u_multiplier_pp3_46 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_46__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_46__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_46__23_  (.A1(u_multiplier_pp3_46 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_46__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_46__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_46__24_  (.A(u_multiplier_pp3_46 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_46__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_46__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_46__25_  (.A(u_multiplier_STAGE4_pp4_45_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_46__16_ ),
    .ZN(u_multiplier_A [46]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_46__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_46__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_46__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_46_c2 ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_46__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_46__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_46__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_46__17_ ),
    .ZN(u_multiplier_B [47]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_47__18_  (.A(u_multiplier_STAGE4_pp4_46_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_47__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_47__19_  (.A1(u_multiplier_pp3_47 [1]),
    .A2(u_multiplier_pp3_47 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_47__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_47__20_  (.A(u_multiplier_pp3_47 [1]),
    .B(u_multiplier_pp3_47 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_47__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_47__21_  (.A1(u_multiplier_pp3_47 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_47__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_47__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_47__22_  (.A(u_multiplier_pp3_47 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_47__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_47__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_47__23_  (.A1(u_multiplier_pp3_47 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_47__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_47__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_47__24_  (.A(u_multiplier_pp3_47 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_47__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_47__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_47__25_  (.A(u_multiplier_STAGE4_pp4_46_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_47__16_ ),
    .ZN(u_multiplier_A [47]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_47__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_47__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_47__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_47_c2 ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_47__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_47__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_47__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_47__17_ ),
    .ZN(u_multiplier_B [48]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_48__18_  (.A(u_multiplier_STAGE4_pp4_47_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_48__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_48__19_  (.A1(u_multiplier_pp3_48 [1]),
    .A2(u_multiplier_pp3_48 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_48__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_48__20_  (.A(u_multiplier_pp3_48 [1]),
    .B(u_multiplier_pp3_48 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_48__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_48__21_  (.A1(u_multiplier_pp3_48 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_48__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_48__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_48__22_  (.A(u_multiplier_pp3_48 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_48__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_48__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_48__23_  (.A1(u_multiplier_pp3_48 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_48__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_48__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_48__24_  (.A(u_multiplier_pp3_48 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_48__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_48__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_48__25_  (.A(u_multiplier_STAGE4_pp4_47_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_48__16_ ),
    .ZN(u_multiplier_A [48]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_48__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_48__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_48__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_48_c2 ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_48__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_48__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_48__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_48__17_ ),
    .ZN(u_multiplier_B [49]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_49__18_  (.A(u_multiplier_STAGE4_pp4_48_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_49__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_49__19_  (.A1(u_multiplier_pp3_49 [1]),
    .A2(u_multiplier_pp3_49 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_49__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_49__20_  (.A(u_multiplier_pp3_49 [1]),
    .B(u_multiplier_pp3_49 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_49__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_49__21_  (.A1(u_multiplier_pp3_49 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_49__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_49__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_49__22_  (.A(u_multiplier_pp3_49 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_49__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_49__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_49__23_  (.A1(u_multiplier_pp3_49 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_49__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_49__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_49__24_  (.A(u_multiplier_pp3_49 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_49__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_49__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_49__25_  (.A(u_multiplier_STAGE4_pp4_48_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_49__16_ ),
    .ZN(u_multiplier_A [49]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_49__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_49__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_49__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_49_c2 ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_49__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_49__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_49__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_49__17_ ),
    .ZN(u_multiplier_B [50]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_50__18_  (.A(u_multiplier_STAGE4_pp4_49_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_50__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_50__19_  (.A1(u_multiplier_pp3_50 [1]),
    .A2(u_multiplier_pp3_50 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_50__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_50__20_  (.A(u_multiplier_pp3_50 [1]),
    .B(u_multiplier_pp3_50 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_50__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_50__21_  (.A1(u_multiplier_pp3_50 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_50__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_50__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_50__22_  (.A(u_multiplier_pp3_50 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_50__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_50__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_50__23_  (.A1(u_multiplier_pp3_50 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_50__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_50__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_50__24_  (.A(u_multiplier_pp3_50 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_50__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_50__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_50__25_  (.A(u_multiplier_STAGE4_pp4_49_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_50__16_ ),
    .ZN(u_multiplier_A [50]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_50__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_50__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_50__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_50_c2 ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_50__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_50__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_50__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_50__17_ ),
    .ZN(u_multiplier_B [51]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_51__18_  (.A(u_multiplier_STAGE4_pp4_50_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_51__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_51__19_  (.A1(u_multiplier_pp3_51 [1]),
    .A2(u_multiplier_pp3_51 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_51__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_51__20_  (.A(u_multiplier_pp3_51 [1]),
    .B(u_multiplier_pp3_51 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_51__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_51__21_  (.A1(u_multiplier_pp3_51 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_51__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_51__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_51__22_  (.A(u_multiplier_pp3_51 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_51__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_51__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_51__23_  (.A1(u_multiplier_pp3_51 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_51__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_51__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_51__24_  (.A(u_multiplier_pp3_51 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_51__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_51__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_51__25_  (.A(u_multiplier_STAGE4_pp4_50_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_51__16_ ),
    .ZN(u_multiplier_A [51]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_51__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_51__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_51__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_51_c2 ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_51__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_51__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_51__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_51__17_ ),
    .ZN(u_multiplier_B [52]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_52__18_  (.A(u_multiplier_STAGE4_pp4_51_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_52__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_52__19_  (.A1(u_multiplier_pp3_52 [1]),
    .A2(u_multiplier_pp3_52 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_52__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_52__20_  (.A(u_multiplier_pp3_52 [1]),
    .B(u_multiplier_pp3_52 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_52__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_52__21_  (.A1(u_multiplier_pp3_52 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_52__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_52__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_52__22_  (.A(u_multiplier_pp3_52 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_52__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_52__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_52__23_  (.A1(u_multiplier_pp3_52 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_52__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_52__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_52__24_  (.A(u_multiplier_pp3_52 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_52__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_52__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_52__25_  (.A(u_multiplier_STAGE4_pp4_51_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_52__16_ ),
    .ZN(u_multiplier_A [52]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_52__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_52__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_52__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_52_c2 ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_52__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_52__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_52__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_52__17_ ),
    .ZN(u_multiplier_B [53]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_53__18_  (.A(u_multiplier_STAGE4_pp4_52_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_53__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_53__19_  (.A1(u_multiplier_pp3_53 [1]),
    .A2(u_multiplier_pp3_53 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_53__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_53__20_  (.A(u_multiplier_pp3_53 [1]),
    .B(u_multiplier_pp3_53 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_53__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_53__21_  (.A1(u_multiplier_pp3_53 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_53__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_53__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_53__22_  (.A(u_multiplier_pp3_53 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_53__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_53__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_53__23_  (.A1(u_multiplier_pp3_53 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_53__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_53__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_53__24_  (.A(u_multiplier_pp3_53 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_53__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_53__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_53__25_  (.A(u_multiplier_STAGE4_pp4_52_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_53__16_ ),
    .ZN(u_multiplier_A [53]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_53__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_53__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_53__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_53_c2 ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_53__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_53__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_53__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_53__17_ ),
    .ZN(u_multiplier_B [54]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_54__18_  (.A(u_multiplier_STAGE4_pp4_53_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_54__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_54__19_  (.A1(u_multiplier_pp3_54 [1]),
    .A2(u_multiplier_pp3_54 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_54__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_54__20_  (.A(u_multiplier_pp3_54 [1]),
    .B(u_multiplier_pp3_54 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_54__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_54__21_  (.A1(u_multiplier_pp3_54 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_54__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_54__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_54__22_  (.A(u_multiplier_pp3_54 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_54__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_54__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_54__23_  (.A1(u_multiplier_pp3_54 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_54__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_54__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_54__24_  (.A(u_multiplier_pp3_54 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_54__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_54__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_54__25_  (.A(u_multiplier_STAGE4_pp4_53_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_54__16_ ),
    .ZN(u_multiplier_A [54]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_54__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_54__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_54__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_54_c2 ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_54__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_54__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_54__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_54__17_ ),
    .ZN(u_multiplier_B [55]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_55__18_  (.A(u_multiplier_STAGE4_pp4_54_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_55__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_55__19_  (.A1(u_multiplier_pp3_55 [1]),
    .A2(u_multiplier_pp3_55 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_55__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_55__20_  (.A(u_multiplier_pp3_55 [1]),
    .B(u_multiplier_pp3_55 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_55__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_55__21_  (.A1(u_multiplier_pp3_55 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_55__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_55__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_55__22_  (.A(u_multiplier_pp3_55 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_55__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_55__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_55__23_  (.A1(u_multiplier_pp3_55 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_55__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_55__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_55__24_  (.A(u_multiplier_pp3_55 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_55__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_55__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_55__25_  (.A(u_multiplier_STAGE4_pp4_54_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_55__16_ ),
    .ZN(u_multiplier_A [55]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_55__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_55__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_55__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_55_c2 ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_55__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_55__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_55__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_55__17_ ),
    .ZN(u_multiplier_B [56]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_56__18_  (.A(u_multiplier_STAGE4_pp4_55_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_56__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_56__19_  (.A1(u_multiplier_pp3_56 [1]),
    .A2(u_multiplier_pp3_56 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_56__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_56__20_  (.A(u_multiplier_pp3_56 [1]),
    .B(u_multiplier_pp3_56 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_56__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_56__21_  (.A1(u_multiplier_pp3_56 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_56__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_56__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_56__22_  (.A(u_multiplier_pp3_56 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_56__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_56__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_56__23_  (.A1(u_multiplier_pp3_56 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_56__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_56__15_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_56__24_  (.A(u_multiplier_pp3_56 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_56__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_56__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_56__25_  (.A(u_multiplier_STAGE4_pp4_55_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_56__16_ ),
    .ZN(u_multiplier_A [56]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_56__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_56__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_56__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_56_c2 ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_56__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_56__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_56__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_56__17_ ),
    .ZN(u_multiplier_B [57]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_57__18_  (.A(u_multiplier_STAGE4_pp4_56_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_57__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_57__19_  (.A1(u_multiplier_pp3_57 [1]),
    .A2(u_multiplier_pp3_57 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_57__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_57__20_  (.A(u_multiplier_pp3_57 [1]),
    .B(u_multiplier_pp3_57 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_57__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_57__21_  (.A1(u_multiplier_pp3_57 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_57__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_57__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_57__22_  (.A(u_multiplier_pp3_57 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_57__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_57__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_57__23_  (.A1(u_multiplier_pp3_57 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_57__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_57__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_57__24_  (.A(u_multiplier_pp3_57 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_57__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_57__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_57__25_  (.A(u_multiplier_STAGE4_pp4_56_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_57__16_ ),
    .ZN(u_multiplier_A [57]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_57__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_57__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_57__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_57_c2 ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_57__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_57__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_57__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_57__17_ ),
    .ZN(u_multiplier_B [58]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_58__18_  (.A(u_multiplier_STAGE4_pp4_57_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_58__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_58__19_  (.A1(u_multiplier_pp3_58 [1]),
    .A2(u_multiplier_pp3_58 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_58__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_58__20_  (.A(u_multiplier_pp3_58 [1]),
    .B(u_multiplier_pp3_58 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_58__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_58__21_  (.A1(u_multiplier_pp3_58 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_58__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_58__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_58__22_  (.A(u_multiplier_pp3_58 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_58__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_58__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_58__23_  (.A1(u_multiplier_pp3_58 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_58__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_58__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_58__24_  (.A(u_multiplier_pp3_58 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_58__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_58__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_58__25_  (.A(u_multiplier_STAGE4_pp4_57_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_58__16_ ),
    .ZN(u_multiplier_A [58]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_58__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_58__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_58__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_58_c2 ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_58__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_58__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_58__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_58__17_ ),
    .ZN(u_multiplier_B [59]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_59__18_  (.A(u_multiplier_STAGE4_pp4_58_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_59__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_59__19_  (.A1(u_multiplier_pp3_59 [1]),
    .A2(u_multiplier_pp3_59 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_59__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_59__20_  (.A(u_multiplier_pp3_59 [1]),
    .B(u_multiplier_pp3_59 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_59__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_59__21_  (.A1(u_multiplier_pp3_59 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_59__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_59__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_59__22_  (.A(u_multiplier_pp3_59 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_59__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_59__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_59__23_  (.A1(u_multiplier_pp3_59 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_59__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_59__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_59__24_  (.A(u_multiplier_pp3_59 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_59__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_59__16_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_59__25_  (.A(u_multiplier_STAGE4_pp4_58_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_59__16_ ),
    .ZN(u_multiplier_A [59]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_59__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_59__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_59__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_59_c2 ));
 OAI21_X1 u_multiplier_STAGE4_E_4_2_pp4_59__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_59__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_59__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_59__17_ ),
    .ZN(u_multiplier_B [60]));
 INV_X1 u_multiplier_STAGE4_E_4_2_pp4_60__18_  (.A(u_multiplier_STAGE4_pp4_59_c2 ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_60__17_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_60__19_  (.A1(u_multiplier_pp3_60 [1]),
    .A2(u_multiplier_pp3_60 [0]),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_60__11_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_60__20_  (.A(u_multiplier_pp3_60 [1]),
    .B(u_multiplier_pp3_60 [0]),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_60__12_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_60__21_  (.A1(u_multiplier_pp3_60 [2]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_60__12_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_60__13_ ));
 XOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_60__22_  (.A(u_multiplier_pp3_60 [2]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_60__12_ ),
    .Z(u_multiplier_STAGE4_E_4_2_pp4_60__14_ ));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_60__23_  (.A1(u_multiplier_pp3_60 [3]),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_60__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_60__15_ ));
 XNOR2_X2 u_multiplier_STAGE4_E_4_2_pp4_60__24_  (.A(u_multiplier_pp3_60 [3]),
    .B(u_multiplier_STAGE4_E_4_2_pp4_60__14_ ),
    .ZN(u_multiplier_STAGE4_E_4_2_pp4_60__16_ ));
 XNOR2_X1 u_multiplier_STAGE4_E_4_2_pp4_60__25_  (.A(u_multiplier_STAGE4_pp4_59_c2 ),
    .B(u_multiplier_STAGE4_E_4_2_pp4_60__16_ ),
    .ZN(u_multiplier_A [60]));
 NAND2_X1 u_multiplier_STAGE4_E_4_2_pp4_60__26_  (.A1(u_multiplier_STAGE4_E_4_2_pp4_60__11_ ),
    .A2(u_multiplier_STAGE4_E_4_2_pp4_60__13_ ),
    .ZN(u_multiplier_STAGE4_pp4_60_c2 ));
 OAI21_X2 u_multiplier_STAGE4_E_4_2_pp4_60__27_  (.A(u_multiplier_STAGE4_E_4_2_pp4_60__15_ ),
    .B1(u_multiplier_STAGE4_E_4_2_pp4_60__16_ ),
    .B2(u_multiplier_STAGE4_E_4_2_pp4_60__17_ ),
    .ZN(u_multiplier_B [61]));
 INV_X1 u_multiplier_STAGE4_Full_adder_pp4_61__12_  (.A(u_multiplier_STAGE4_pp4_60_c2 ),
    .ZN(u_multiplier_STAGE4_Full_adder_pp4_61__08_ ));
 NAND3_X2 u_multiplier_STAGE4_Full_adder_pp4_61__13_  (.A1(u_multiplier_pp3_61 [1]),
    .A2(u_multiplier_pp3_61 [0]),
    .A3(u_multiplier_STAGE4_pp4_60_c2 ),
    .ZN(u_multiplier_STAGE4_Full_adder_pp4_61__09_ ));
 NOR2_X2 u_multiplier_STAGE4_Full_adder_pp4_61__14_  (.A1(u_multiplier_pp3_61 [1]),
    .A2(u_multiplier_pp3_61 [0]),
    .ZN(u_multiplier_STAGE4_Full_adder_pp4_61__10_ ));
 AOI21_X1 u_multiplier_STAGE4_Full_adder_pp4_61__15_  (.A(u_multiplier_STAGE4_pp4_60_c2 ),
    .B1(u_multiplier_pp3_61 [0]),
    .B2(u_multiplier_pp3_61 [1]),
    .ZN(u_multiplier_STAGE4_Full_adder_pp4_61__11_ ));
 NOR2_X2 u_multiplier_STAGE4_Full_adder_pp4_61__16_  (.A1(u_multiplier_STAGE4_Full_adder_pp4_61__10_ ),
    .A2(u_multiplier_STAGE4_Full_adder_pp4_61__11_ ),
    .ZN(u_multiplier_B [62]));
 AOI22_X4 u_multiplier_STAGE4_Full_adder_pp4_61__17_  (.A1(u_multiplier_STAGE4_Full_adder_pp4_61__08_ ),
    .A2(u_multiplier_STAGE4_Full_adder_pp4_61__10_ ),
    .B1(u_multiplier_B [62]),
    .B2(u_multiplier_STAGE4_Full_adder_pp4_61__09_ ),
    .ZN(u_multiplier_A [61]));
 AND2_X1 u_multiplier_STAGE4_Half_adder_pp4_2__4_  (.A1(u_multiplier_pp3_2 [1]),
    .A2(u_multiplier_pp3_2 [0]),
    .ZN(u_multiplier_B [3]));
 XOR2_X2 u_multiplier_STAGE4_Half_adder_pp4_2__5_  (.A(u_multiplier_pp3_2 [1]),
    .B(u_multiplier_pp3_2 [0]),
    .Z(u_multiplier_A [2]));
 LOGIC0_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__43__142  (.Z(net142));
 CLKBUF_X1 hold150 (.A(net211),
    .Z(net150));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_219_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_220_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_221_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_222_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_223_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_224_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_225_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_226_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_227_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_228_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_229_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_230_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_231_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_232_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_233_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_234_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_235_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_236_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_237_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_2_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_2_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_2_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_2_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_2_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_2_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_2_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_2_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_2_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_2_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_2_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_2_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_2_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_2_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_2_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_2_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_2_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_2_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_2_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_2_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_2_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_2_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_2_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_2_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_2_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_2_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_2_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_2_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_2_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_2_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_2_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_2_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_2_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_2_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_2_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_2_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_2_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_2_Right_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_2_Right_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_2_Right_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_2_Right_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_2_Right_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_2_Right_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_2_Right_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_2_Right_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_2_Right_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_2_Right_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_2_Right_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_2_Right_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_2_Right_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_2_Right_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_2_Right_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_2_Right_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_2_Right_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_2_Right_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_2_Right_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_2_Right_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_2_Right_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_2_Right_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_2_Right_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_2_Right_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_2_Right_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_2_Right_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_2_Right_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_2_Right_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_2_Right_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_2_Right_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_2_Right_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_2_Right_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_2_Right_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_2_Right_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_2_Right_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_2_Right_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_2_Right_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_2_Right_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_2_Right_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_2_Right_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_2_Right_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_2_Right_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_2_Right_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_2_Right_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_2_Right_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_2_Right_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_2_Right_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_2_Right_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_2_Right_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_2_Right_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_2_Right_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_2_Right_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_2_Right_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_2_Right_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_2_Right_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_2_Right_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_2_Right_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_2_Right_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_2_Right_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_2_Right_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_2_Right_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_2_Right_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_2_Right_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_2_Right_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_2_Right_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_2_Right_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_2_Right_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_2_Right_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_2_Right_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_2_Right_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_2_Right_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_2_Right_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_2_Right_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_2_Right_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_2_Right_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_2_Right_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_2_Right_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_2_Right_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_2_Right_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_2_Right_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_2_Right_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_2_Right_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_2_Right_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_2_Right_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_2_Right_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_2_Right_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_2_Right_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_2_Right_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_2_Right_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_2_Right_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_2_Right_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_2_Right_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_2_Right_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_2_Right_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_2_Right_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_2_Right_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_2_Right_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_2_Right_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_2_Right_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_2_Right_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_2_Right_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_2_Right_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_2_Right_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_2_Right_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_2_Right_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_2_Right_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_2_Right_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_2_Right_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_2_Right_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_2_Right_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_2_Right_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_2_Right_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_2_Right_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_2_Right_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_2_Right_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_2_Right_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_2_Right_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_2_Right_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_2_Right_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_2_Right_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_2_Right_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_2_Right_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_2_Right_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_2_Right_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_2_Right_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_2_Right_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_2_Right_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_2_Right_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_2_Right_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_2_Right_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_2_Right_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_265 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_266 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_267 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_268 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_269 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_270 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_271 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_272 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_273 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_274 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_275 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_276 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_277 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_1_Left_278 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_1_Left_279 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_1_Left_280 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_1_Left_281 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_1_Left_282 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_1_Left_283 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_1_Left_284 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_1_Left_285 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_1_Left_286 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_1_Left_287 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_1_Left_288 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_1_Left_289 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_1_Left_290 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_1_Left_291 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_1_Left_292 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_1_Left_293 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_1_Left_294 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_1_Left_295 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_1_Left_296 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_1_Left_297 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_1_Left_298 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_1_Left_299 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_1_Left_300 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_1_Left_301 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_1_Left_302 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_1_Left_303 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_1_Left_304 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_1_Left_305 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_1_Left_306 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_1_Left_307 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_1_Left_308 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_1_Left_309 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_1_Left_310 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_1_Left_311 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_1_Left_312 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_1_Left_313 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_1_Left_314 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_1_Left_315 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_1_Left_316 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_1_Left_317 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_1_Left_318 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_1_Left_319 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_1_Left_320 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_1_Left_321 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_1_Left_322 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_1_Left_323 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_1_Left_324 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_1_Left_325 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_1_Left_326 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_1_Left_327 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_1_Left_328 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_1_Left_329 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_1_Left_330 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_1_Left_331 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_1_Left_332 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_1_Left_333 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_1_Left_334 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_1_Left_335 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_1_Left_336 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_1_Left_337 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_1_Left_338 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_1_Left_339 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_1_Left_340 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_1_Left_341 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_1_Left_342 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_1_Left_343 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_1_Left_344 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_1_Left_345 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_1_Left_346 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_1_Left_347 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_1_Left_348 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_1_Left_349 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_1_Left_350 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_1_Left_351 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_1_Left_352 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_1_Left_353 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_1_Left_354 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_1_Left_355 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_1_Left_356 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_1_Left_357 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_1_Left_358 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_1_Left_359 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_1_Left_360 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_1_Left_361 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_1_Left_362 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_1_Left_363 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_1_Left_364 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_1_Left_365 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_1_Left_366 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_1_Left_367 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_1_Left_368 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_1_Left_369 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_1_Left_370 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_1_Left_371 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_1_Left_372 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_1_Left_373 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_1_Left_374 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_1_Left_375 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_1_Left_376 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_1_Left_377 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_1_Left_378 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_1_Left_379 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_1_Left_380 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_1_Left_381 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_1_Left_382 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_1_Left_383 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_1_Left_384 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_1_Left_385 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_1_Left_386 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_1_Left_387 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_1_Left_388 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_1_Left_389 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_1_Left_390 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_1_Left_391 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_1_Left_392 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_1_Left_393 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_1_Left_394 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_1_Left_395 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_1_Left_396 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_1_Left_397 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_1_Left_398 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_1_Left_399 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_1_Left_400 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_1_Left_401 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_1_Left_402 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_1_Left_403 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_1_Left_404 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_1_Left_405 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_1_Left_406 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_1_Left_407 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_1_Left_408 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_1_Left_409 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_1_Left_410 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_1_Left_411 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_1_Left_412 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_1_Left_413 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_1_Left_414 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_1_Left_415 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_1_Left_416 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_1_Left_417 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_1_Left_418 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_1_Left_419 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_1_Left_420 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_1_Left_421 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_1_Left_422 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_1_Left_423 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_1_Left_424 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_1_Left_425 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_1_Left_426 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_1_Left_427 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_1_Left_428 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_1_Left_429 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_1_Left_430 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_1_Left_431 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_1_Left_432 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_1_Left_433 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_1_Left_434 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_1_Left_435 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_1_Left_436 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_1_Left_437 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_1_Left_438 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_1_Left_439 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_1_Left_440 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_1_Left_441 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_1_Left_442 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_1_Left_443 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_1_Left_444 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Left_445 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Left_446 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Left_447 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Left_448 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Left_449 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Left_450 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Left_451 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Left_452 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Left_453 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Left_454 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Left_455 ();
 TAPCELL_X1 PHY_EDGE_ROW_219_Left_456 ();
 TAPCELL_X1 PHY_EDGE_ROW_220_Left_457 ();
 TAPCELL_X1 PHY_EDGE_ROW_221_Left_458 ();
 TAPCELL_X1 PHY_EDGE_ROW_222_Left_459 ();
 TAPCELL_X1 PHY_EDGE_ROW_223_Left_460 ();
 TAPCELL_X1 PHY_EDGE_ROW_224_Left_461 ();
 TAPCELL_X1 PHY_EDGE_ROW_225_Left_462 ();
 TAPCELL_X1 PHY_EDGE_ROW_226_Left_463 ();
 TAPCELL_X1 PHY_EDGE_ROW_227_Left_464 ();
 TAPCELL_X1 PHY_EDGE_ROW_228_Left_465 ();
 TAPCELL_X1 PHY_EDGE_ROW_229_Left_466 ();
 TAPCELL_X1 PHY_EDGE_ROW_230_Left_467 ();
 TAPCELL_X1 PHY_EDGE_ROW_231_Left_468 ();
 TAPCELL_X1 PHY_EDGE_ROW_232_Left_469 ();
 TAPCELL_X1 PHY_EDGE_ROW_233_Left_470 ();
 TAPCELL_X1 PHY_EDGE_ROW_234_Left_471 ();
 TAPCELL_X1 PHY_EDGE_ROW_235_Left_472 ();
 TAPCELL_X1 PHY_EDGE_ROW_236_Left_473 ();
 TAPCELL_X1 PHY_EDGE_ROW_237_Left_474 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_1_Left_475 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_2_Left_476 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_2_Left_477 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_2_Left_478 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_2_Left_479 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_2_Left_480 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_2_Left_481 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_2_Left_482 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_2_Left_483 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_2_Left_484 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_2_Left_485 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_2_Left_486 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_2_Left_487 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_2_Left_488 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_2_Left_489 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_2_Left_490 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_2_Left_491 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_2_Left_492 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_2_Left_493 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_2_Left_494 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_2_Left_495 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_2_Left_496 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_2_Left_497 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_2_Left_498 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_2_Left_499 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_2_Left_500 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_2_Left_501 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_2_Left_502 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_2_Left_503 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_2_Left_504 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_2_Left_505 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_2_Left_506 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_2_Left_507 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_2_Left_508 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_2_Left_509 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_2_Left_510 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_2_Left_511 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_2_Left_512 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_2_Left_513 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_2_Left_514 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_2_Left_515 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_2_Left_516 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_2_Left_517 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_2_Left_518 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_2_Left_519 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_2_Left_520 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_2_Left_521 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_2_Left_522 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_2_Left_523 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_2_Left_524 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_2_Left_525 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_2_Left_526 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_2_Left_527 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_2_Left_528 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_2_Left_529 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_2_Left_530 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_2_Left_531 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_2_Left_532 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_2_Left_533 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_2_Left_534 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_2_Left_535 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_2_Left_536 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_2_Left_537 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_2_Left_538 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_2_Left_539 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_2_Left_540 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_2_Left_541 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_2_Left_542 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_2_Left_543 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_2_Left_544 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_2_Left_545 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_2_Left_546 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_2_Left_547 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_2_Left_548 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_2_Left_549 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_2_Left_550 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_2_Left_551 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_2_Left_552 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_2_Left_553 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_2_Left_554 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_2_Left_555 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_2_Left_556 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_2_Left_557 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_2_Left_558 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_2_Left_559 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_2_Left_560 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_2_Left_561 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_2_Left_562 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_2_Left_563 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_2_Left_564 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_2_Left_565 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_2_Left_566 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_2_Left_567 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_2_Left_568 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_2_Left_569 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_2_Left_570 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_2_Left_571 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_2_Left_572 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_2_Left_573 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_2_Left_574 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_2_Left_575 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_2_Left_576 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_2_Left_577 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_2_Left_578 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_2_Left_579 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_2_Left_580 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_2_Left_581 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_2_Left_582 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_2_Left_583 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_2_Left_584 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_2_Left_585 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_2_Left_586 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_2_Left_587 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_2_Left_588 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_2_Left_589 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_2_Left_590 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_2_Left_591 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_2_Left_592 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_2_Left_593 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_2_Left_594 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_2_Left_595 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_2_Left_596 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_2_Left_597 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_2_Left_598 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_2_Left_599 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_2_Left_600 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_2_Left_601 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_2_Left_602 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_2_Left_603 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_2_Left_604 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_2_Left_605 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_2_Left_606 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_2_Left_607 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_2_Left_608 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_2_Left_609 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_2_Left_610 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_2_Left_611 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_2_Left_612 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_2_Left_613 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_2_Left_614 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_2_Left_615 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_2_Left_616 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_2_Left_617 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_2_Left_618 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_2_Left_619 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_2_Left_620 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_2_Left_621 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_2_Left_622 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_2_Left_623 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_2_Left_624 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_2_Left_625 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_2_Left_626 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_2_Left_627 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_2_Left_628 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_2_Left_629 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_2_Left_630 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_2_Left_631 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_2_Left_632 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_2_Left_633 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_2_Left_634 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_2_Left_635 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_2_Left_636 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_2_Left_637 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_2_Left_638 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_2_Left_639 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_2_Left_640 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_2_Left_641 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_2_Left_642 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_2_Left_643 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_1_Right_644 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_1_Right_645 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_1_Right_646 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_1_Right_647 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_1_Right_648 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_1_Right_649 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_1_Right_650 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_1_Right_651 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_1_Right_652 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_1_Right_653 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_1_Right_654 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_1_Right_655 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_1_Right_656 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_1_Right_657 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_1_Right_658 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_1_Right_659 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_1_Right_660 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_1_Right_661 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_1_Right_662 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_1_Right_663 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_1_Right_664 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_1_Right_665 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_1_Right_666 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_1_Right_667 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_1_Right_668 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_1_Right_669 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_1_Right_670 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_1_Right_671 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_1_Right_672 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_1_Right_673 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_1_Right_674 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_1_Right_675 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_1_Right_676 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_1_Right_677 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_1_Right_678 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_1_Right_679 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_1_Right_680 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_1_Right_681 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_1_Right_682 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_1_Right_683 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_1_Right_684 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_1_Right_685 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_1_Right_686 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_1_Right_687 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_1_Right_688 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_1_Right_689 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_1_Right_690 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_1_Right_691 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_1_Right_692 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_1_Right_693 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_1_Right_694 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_1_Right_695 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_1_Right_696 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_1_Right_697 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_1_Right_698 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_1_Right_699 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_1_Right_700 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_1_Right_701 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_1_Right_702 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_1_Right_703 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_1_Right_704 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_1_Right_705 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_1_Right_706 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_1_Right_707 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_1_Right_708 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_1_Right_709 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_1_Right_710 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_1_Right_711 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_1_Right_712 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_1_Right_713 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_1_Right_714 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_1_Right_715 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_1_Right_716 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_1_Right_717 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_1_Right_718 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_1_Right_719 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_1_Right_720 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_1_Right_721 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_1_Right_722 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_1_Right_723 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_1_Right_724 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_1_Right_725 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_1_Right_726 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_1_Right_727 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_1_Right_728 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_1_Right_729 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_1_Right_730 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_1_Right_731 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_1_Right_732 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_1_Right_733 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_1_Right_734 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_1_Right_735 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_1_Right_736 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_1_Right_737 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_1_Right_738 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_1_Right_739 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_1_Right_740 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_1_Right_741 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_1_Right_742 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_1_Right_743 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_1_Right_744 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_1_Right_745 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_1_Right_746 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_1_Right_747 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_1_Right_748 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_1_Right_749 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_1_Right_750 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_1_Right_751 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_1_Right_752 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_1_Right_753 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_1_Right_754 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_1_Right_755 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_1_Right_756 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_1_Right_757 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_1_Right_758 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_1_Right_759 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_1_Right_760 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_1_Right_761 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_1_Right_762 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_1_Right_763 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_1_Right_764 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_1_Right_765 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_1_Right_766 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_1_Right_767 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_1_Right_768 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_1_Right_769 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_1_Right_770 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_1_Right_771 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_1_Right_772 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_1_Right_773 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_1_Right_774 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_1_Right_775 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_1_Right_776 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_1_Right_777 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_1_Right_778 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_1_Right_779 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_1_Right_780 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_1_Right_781 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_1_Right_782 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_1_Right_783 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_1_Right_784 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_1_Right_785 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_1_Right_786 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_1_Right_787 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_1_Right_788 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_1_Right_789 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_1_Right_790 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_1_Right_791 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_1_Right_792 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_1_Right_793 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_1_Right_794 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_1_Right_795 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_1_Right_796 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_1_Right_797 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_1_Right_798 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_1_Right_799 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_1_Right_800 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_1_Right_801 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_1_Right_802 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_1_Right_803 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_1_Right_804 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_1_Right_805 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_1_Right_806 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_1_Right_807 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_1_Right_808 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_1_Right_809 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_1_Right_810 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_1_Right_811 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_812 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_813 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_814 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_815 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_816 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_817 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_818 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_819 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_820 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_821 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_822 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_823 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_824 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_825 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_826 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_827 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_828 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_829 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_830 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_831 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_832 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_833 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_834 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_835 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_836 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_837 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_838 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_839 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_840 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_841 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_842 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_843 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_844 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_845 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_846 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_847 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_848 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_849 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_850 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_851 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_852 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_853 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_208_854 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_208_855 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_209_856 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_210_857 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_211_858 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_212_859 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_213_860 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_214_861 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_215_862 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_216_863 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_217_864 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_218_865 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_219_866 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_220_867 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_221_868 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_222_869 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_223_870 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_224_871 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_225_872 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_226_873 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_227_874 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_228_875 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_229_876 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_230_877 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_231_878 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_232_879 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_233_880 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_234_881 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_235_882 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_236_883 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_237_884 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_237_885 ();
 BUF_X16 max_length7 (.A(_0303_),
    .Z(net7));
 BUF_X16 max_length8 (.A(net9),
    .Z(net8));
 BUF_X16 max_length9 (.A(net44),
    .Z(net9));
 BUF_X4 input10 (.A(data_in[0]),
    .Z(net10));
 BUF_X4 input11 (.A(data_in[10]),
    .Z(net11));
 BUF_X1 input12 (.A(data_in[11]),
    .Z(net12));
 BUF_X1 input13 (.A(data_in[12]),
    .Z(net13));
 CLKBUF_X3 input14 (.A(data_in[13]),
    .Z(net14));
 BUF_X4 input15 (.A(data_in[14]),
    .Z(net15));
 BUF_X1 input16 (.A(data_in[15]),
    .Z(net16));
 BUF_X1 input17 (.A(data_in[16]),
    .Z(net17));
 BUF_X2 input18 (.A(data_in[17]),
    .Z(net18));
 BUF_X1 input19 (.A(data_in[18]),
    .Z(net19));
 BUF_X4 input20 (.A(data_in[19]),
    .Z(net20));
 BUF_X1 input21 (.A(data_in[1]),
    .Z(net21));
 BUF_X1 input22 (.A(data_in[20]),
    .Z(net22));
 BUF_X1 input23 (.A(data_in[21]),
    .Z(net23));
 BUF_X4 input24 (.A(data_in[22]),
    .Z(net24));
 BUF_X4 input25 (.A(data_in[23]),
    .Z(net25));
 BUF_X1 input26 (.A(data_in[24]),
    .Z(net26));
 CLKBUF_X2 input27 (.A(data_in[25]),
    .Z(net27));
 CLKBUF_X3 input28 (.A(data_in[26]),
    .Z(net28));
 BUF_X2 input29 (.A(data_in[27]),
    .Z(net29));
 BUF_X1 input30 (.A(data_in[28]),
    .Z(net30));
 BUF_X1 input31 (.A(data_in[29]),
    .Z(net31));
 CLKBUF_X2 input32 (.A(data_in[2]),
    .Z(net32));
 BUF_X1 input33 (.A(data_in[30]),
    .Z(net33));
 BUF_X2 input34 (.A(data_in[31]),
    .Z(net34));
 BUF_X4 input35 (.A(data_in[3]),
    .Z(net35));
 BUF_X4 input36 (.A(data_in[4]),
    .Z(net36));
 CLKBUF_X3 input37 (.A(data_in[5]),
    .Z(net37));
 BUF_X1 input38 (.A(data_in[6]),
    .Z(net38));
 BUF_X1 input39 (.A(data_in[7]),
    .Z(net39));
 BUF_X4 input40 (.A(data_in[8]),
    .Z(net40));
 BUF_X4 input41 (.A(data_in[9]),
    .Z(net41));
 BUF_X4 input42 (.A(init_enable),
    .Z(net42));
 BUF_X4 input43 (.A(pe_ce),
    .Z(net43));
 BUF_X8 input44 (.A(rst_n),
    .Z(net44));
 BUF_X1 output45 (.A(net45),
    .Z(curr_state[1]));
 BUF_X1 output46 (.A(net46),
    .Z(data_out[0]));
 BUF_X1 output47 (.A(net47),
    .Z(data_out[10]));
 BUF_X1 output48 (.A(net48),
    .Z(data_out[11]));
 BUF_X1 output49 (.A(net49),
    .Z(data_out[12]));
 BUF_X1 output50 (.A(net50),
    .Z(data_out[13]));
 BUF_X1 output51 (.A(net51),
    .Z(data_out[14]));
 BUF_X1 output52 (.A(net52),
    .Z(data_out[15]));
 BUF_X1 output53 (.A(net53),
    .Z(data_out[16]));
 BUF_X1 output54 (.A(net54),
    .Z(data_out[17]));
 BUF_X1 output55 (.A(net55),
    .Z(data_out[18]));
 BUF_X1 output56 (.A(net56),
    .Z(data_out[19]));
 BUF_X1 output57 (.A(net57),
    .Z(data_out[1]));
 BUF_X1 output58 (.A(net58),
    .Z(data_out[20]));
 BUF_X1 output59 (.A(net59),
    .Z(data_out[21]));
 BUF_X1 output60 (.A(net60),
    .Z(data_out[22]));
 BUF_X1 output61 (.A(net61),
    .Z(data_out[23]));
 BUF_X1 output62 (.A(net62),
    .Z(data_out[24]));
 BUF_X1 output63 (.A(net63),
    .Z(data_out[25]));
 BUF_X1 output64 (.A(net64),
    .Z(data_out[26]));
 BUF_X1 output65 (.A(net65),
    .Z(data_out[27]));
 BUF_X1 output66 (.A(net66),
    .Z(data_out[28]));
 BUF_X1 output67 (.A(net67),
    .Z(data_out[29]));
 BUF_X1 output68 (.A(net68),
    .Z(data_out[2]));
 BUF_X1 output69 (.A(net69),
    .Z(data_out[30]));
 BUF_X1 output70 (.A(net70),
    .Z(data_out[31]));
 BUF_X1 output71 (.A(net71),
    .Z(data_out[32]));
 BUF_X1 output72 (.A(net72),
    .Z(data_out[33]));
 BUF_X1 output73 (.A(net73),
    .Z(data_out[34]));
 BUF_X1 output74 (.A(net74),
    .Z(data_out[35]));
 BUF_X1 output75 (.A(net75),
    .Z(data_out[36]));
 BUF_X1 output76 (.A(net76),
    .Z(data_out[37]));
 BUF_X1 output77 (.A(net77),
    .Z(data_out[38]));
 BUF_X1 output78 (.A(net78),
    .Z(data_out[39]));
 BUF_X1 output79 (.A(net79),
    .Z(data_out[3]));
 BUF_X1 output80 (.A(net80),
    .Z(data_out[40]));
 BUF_X1 output81 (.A(net81),
    .Z(data_out[41]));
 BUF_X1 output82 (.A(net82),
    .Z(data_out[42]));
 BUF_X1 output83 (.A(net83),
    .Z(data_out[43]));
 BUF_X1 output84 (.A(net84),
    .Z(data_out[44]));
 BUF_X1 output85 (.A(net85),
    .Z(data_out[45]));
 BUF_X1 output86 (.A(net86),
    .Z(data_out[46]));
 BUF_X1 output87 (.A(net87),
    .Z(data_out[47]));
 BUF_X1 output88 (.A(net88),
    .Z(data_out[48]));
 BUF_X1 output89 (.A(net89),
    .Z(data_out[49]));
 BUF_X1 output90 (.A(net90),
    .Z(data_out[4]));
 BUF_X1 output91 (.A(net91),
    .Z(data_out[50]));
 BUF_X1 output92 (.A(net92),
    .Z(data_out[51]));
 BUF_X1 output93 (.A(net93),
    .Z(data_out[52]));
 BUF_X1 output94 (.A(net94),
    .Z(data_out[53]));
 BUF_X1 output95 (.A(net95),
    .Z(data_out[54]));
 BUF_X1 output96 (.A(net96),
    .Z(data_out[55]));
 BUF_X1 output97 (.A(net97),
    .Z(data_out[56]));
 BUF_X1 output98 (.A(net98),
    .Z(data_out[57]));
 BUF_X1 output99 (.A(net99),
    .Z(data_out[58]));
 BUF_X1 output100 (.A(net100),
    .Z(data_out[59]));
 BUF_X1 output101 (.A(net101),
    .Z(data_out[5]));
 BUF_X1 output102 (.A(net102),
    .Z(data_out[60]));
 BUF_X1 output103 (.A(net103),
    .Z(data_out[61]));
 BUF_X1 output104 (.A(net104),
    .Z(data_out[62]));
 BUF_X1 output105 (.A(net105),
    .Z(data_out[63]));
 BUF_X1 output106 (.A(net106),
    .Z(data_out[6]));
 BUF_X1 output107 (.A(net107),
    .Z(data_out[7]));
 BUF_X1 output108 (.A(net108),
    .Z(data_out[8]));
 BUF_X1 output109 (.A(net109),
    .Z(data_out[9]));
 BUF_X1 output110 (.A(net110),
    .Z(valid_reg_out));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_32_1__18__111  (.Z(net111));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_32_1__25__112  (.Z(net112));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_32_2__18__113  (.Z(net113));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_32_2__25__114  (.Z(net114));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_32_3__18__115  (.Z(net115));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_32_3__25__116  (.Z(net116));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_32_4__18__117  (.Z(net117));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_32_4__25__118  (.Z(net118));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_32_5__18__119  (.Z(net119));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_32_5__25__120  (.Z(net120));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_32_6__18__121  (.Z(net121));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_32_6__25__122  (.Z(net122));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_32_7__18__123  (.Z(net123));
 LOGIC0_X1 u_multiplier_STAGE1_E_4_2_pp_32_7__25__124  (.Z(net124));
 LOGIC0_X1 u_multiplier_STAGE2_E_4_2_pp2_32_1__25__126  (.Z(net126));
 LOGIC0_X1 u_multiplier_STAGE2_E_4_2_pp2_32_2__18__127  (.Z(net127));
 LOGIC0_X1 u_multiplier_STAGE2_E_4_2_pp2_32_2__25__128  (.Z(net128));
 LOGIC0_X1 u_multiplier_STAGE2_E_4_2_pp2_32_3__18__129  (.Z(net129));
 LOGIC0_X1 u_multiplier_STAGE2_E_4_2_pp2_32_3__25__130  (.Z(net130));
 LOGIC0_X1 u_multiplier_STAGE2_E_4_2_pp2_32_4__18__131  (.Z(net131));
 LOGIC0_X1 u_multiplier_STAGE2_E_4_2_pp2_32_4__25__132  (.Z(net132));
 LOGIC0_X1 u_multiplier_STAGE3_E_4_2_pp3_32_1__25__134  (.Z(net134));
 LOGIC0_X1 u_multiplier_STAGE3_E_4_2_pp3_32_2__18__135  (.Z(net135));
 LOGIC0_X1 u_multiplier_STAGE3_E_4_2_pp3_32_2__25__136  (.Z(net136));
 LOGIC0_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__41__138  (.Z(net138));
 LOGIC0_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__42__139  (.Z(net139));
 LOGIC0_X1 u_multiplier_STAGE4_E_4_2_pp4_32__18__140  (.Z(net140));
 LOGIC0_X1 u_multiplier_STAGE4_E_4_2_pp4_32__25__141  (.Z(net141));
 LOGIC0_X1 u_multiplier_Final_add_cla1_cla1_cla1_cla1__44__143  (.Z(net143));
 LOGIC0_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__55__144  (.Z(net144));
 LOGIC0_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__55__145  (.Z(net145));
 LOGIC0_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__56__146  (.Z(net146));
 LOGIC0_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__56__147  (.Z(net147));
 LOGIC0_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__57__148  (.Z(net148));
 LOGIC0_X1 u_multiplier_Final_add_cla2_cla2_cla2_cla2__57__149  (.Z(net149));
 CLKBUF_X1 hold151 (.A(_0268_),
    .Z(net151));
 CLKBUF_X1 hold152 (.A(net217),
    .Z(net152));
 CLKBUF_X1 hold153 (.A(_0304_),
    .Z(net153));
 CLKBUF_X1 hold154 (.A(net1),
    .Z(net154));
 CLKBUF_X1 hold155 (.A(net170),
    .Z(net155));
 CLKBUF_X1 hold156 (.A(net3),
    .Z(net156));
 CLKBUF_X1 hold157 (.A(net182),
    .Z(net157));
 CLKBUF_X1 hold158 (.A(net179),
    .Z(net158));
 CLKBUF_X1 hold159 (.A(net6),
    .Z(net159));
 CLKBUF_X1 hold160 (.A(net176),
    .Z(net160));
 CLKBUF_X1 hold161 (.A(net185),
    .Z(net161));
 CLKBUF_X1 hold162 (.A(net187),
    .Z(net162));
 CLKBUF_X1 hold163 (.A(net195),
    .Z(net163));
 CLKBUF_X1 hold164 (.A(net197),
    .Z(net164));
 CLKBUF_X1 hold165 (.A(net199),
    .Z(net165));
 CLKBUF_X1 hold166 (.A(net201),
    .Z(net166));
 CLKBUF_X1 hold167 (.A(net205),
    .Z(net167));
 CLKBUF_X1 hold168 (.A(net213),
    .Z(net168));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_1_0_0_clk));
 CLKBUF_X3 clkbuf_1_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_1_1_0_clk));
 CLKBUF_X3 clkbuf_2_0_0_clk (.A(clknet_1_0_0_clk),
    .Z(clknet_2_0_0_clk));
 CLKBUF_X3 clkbuf_2_1_0_clk (.A(clknet_1_0_0_clk),
    .Z(clknet_2_1_0_clk));
 CLKBUF_X3 clkbuf_2_2_0_clk (.A(clknet_1_1_0_clk),
    .Z(clknet_2_2_0_clk));
 CLKBUF_X3 clkbuf_2_3_0_clk (.A(clknet_1_1_0_clk),
    .Z(clknet_2_3_0_clk));
 CLKBUF_X3 clkbuf_3_0_0_clk (.A(clknet_2_0_0_clk),
    .Z(clknet_3_0_0_clk));
 CLKBUF_X3 clkbuf_3_1_0_clk (.A(clknet_2_0_0_clk),
    .Z(clknet_3_1_0_clk));
 CLKBUF_X3 clkbuf_3_2_0_clk (.A(clknet_2_1_0_clk),
    .Z(clknet_3_2_0_clk));
 CLKBUF_X3 clkbuf_3_3_0_clk (.A(clknet_2_1_0_clk),
    .Z(clknet_3_3_0_clk));
 CLKBUF_X3 clkbuf_3_4_0_clk (.A(clknet_2_2_0_clk),
    .Z(clknet_3_4_0_clk));
 CLKBUF_X3 clkbuf_3_5_0_clk (.A(clknet_2_2_0_clk),
    .Z(clknet_3_5_0_clk));
 CLKBUF_X3 clkbuf_3_6_0_clk (.A(clknet_2_3_0_clk),
    .Z(clknet_3_6_0_clk));
 CLKBUF_X3 clkbuf_3_7_0_clk (.A(clknet_2_3_0_clk),
    .Z(clknet_3_7_0_clk));
 CLKBUF_X3 clkbuf_4_0__f_clk (.A(clknet_3_0_0_clk),
    .Z(clknet_4_0__leaf_clk));
 CLKBUF_X3 clkbuf_4_1__f_clk (.A(clknet_3_0_0_clk),
    .Z(clknet_4_1__leaf_clk));
 CLKBUF_X3 clkbuf_4_2__f_clk (.A(clknet_3_1_0_clk),
    .Z(clknet_4_2__leaf_clk));
 CLKBUF_X3 clkbuf_4_3__f_clk (.A(clknet_3_1_0_clk),
    .Z(clknet_4_3__leaf_clk));
 CLKBUF_X3 clkbuf_4_4__f_clk (.A(clknet_3_2_0_clk),
    .Z(clknet_4_4__leaf_clk));
 CLKBUF_X3 clkbuf_4_5__f_clk (.A(clknet_3_2_0_clk),
    .Z(clknet_4_5__leaf_clk));
 CLKBUF_X3 clkbuf_4_6__f_clk (.A(clknet_3_3_0_clk),
    .Z(clknet_4_6__leaf_clk));
 CLKBUF_X3 clkbuf_4_7__f_clk (.A(clknet_3_3_0_clk),
    .Z(clknet_4_7__leaf_clk));
 CLKBUF_X3 clkbuf_4_8__f_clk (.A(clknet_3_4_0_clk),
    .Z(clknet_4_8__leaf_clk));
 CLKBUF_X3 clkbuf_4_9__f_clk (.A(clknet_3_4_0_clk),
    .Z(clknet_4_9__leaf_clk));
 CLKBUF_X3 clkbuf_4_10__f_clk (.A(clknet_3_5_0_clk),
    .Z(clknet_4_10__leaf_clk));
 CLKBUF_X3 clkbuf_4_11__f_clk (.A(clknet_3_5_0_clk),
    .Z(clknet_4_11__leaf_clk));
 CLKBUF_X3 clkbuf_4_12__f_clk (.A(clknet_3_6_0_clk),
    .Z(clknet_4_12__leaf_clk));
 CLKBUF_X3 clkbuf_4_13__f_clk (.A(clknet_3_6_0_clk),
    .Z(clknet_4_13__leaf_clk));
 CLKBUF_X3 clkbuf_4_14__f_clk (.A(clknet_3_7_0_clk),
    .Z(clknet_4_14__leaf_clk));
 CLKBUF_X3 clkbuf_4_15__f_clk (.A(clknet_3_7_0_clk),
    .Z(clknet_4_15__leaf_clk));
 CLKBUF_X1 clkload0 (.A(clknet_4_1__leaf_clk));
 INV_X1 clkload1 (.A(clknet_4_2__leaf_clk));
 CLKBUF_X1 clkload2 (.A(clknet_4_4__leaf_clk));
 INV_X1 clkload3 (.A(clknet_4_6__leaf_clk));
 INV_X1 clkload4 (.A(clknet_4_8__leaf_clk));
 INV_X1 clkload5 (.A(clknet_4_10__leaf_clk));
 INV_X2 clkload6 (.A(clknet_4_15__leaf_clk));
 CLKBUF_X1 hold1 (.A(_0651_),
    .Z(net1));
 CLKBUF_X1 hold2 (.A(net154),
    .Z(net2));
 CLKBUF_X1 hold3 (.A(_0650_),
    .Z(net3));
 CLKBUF_X1 hold4 (.A(_0405_),
    .Z(net4));
 CLKBUF_X1 hold5 (.A(_0163_),
    .Z(net5));
 CLKBUF_X1 hold6 (.A(addr_ptr[2]),
    .Z(net6));
 CLKBUF_X1 hold7 (.A(net159),
    .Z(net169));
 CLKBUF_X1 hold8 (.A(_0656_),
    .Z(net170));
 CLKBUF_X1 hold9 (.A(net155),
    .Z(net171));
 CLKBUF_X1 hold10 (.A(_0265_),
    .Z(net172));
 CLKBUF_X1 hold11 (.A(_0655_),
    .Z(net173));
 CLKBUF_X1 hold12 (.A(_0419_),
    .Z(net174));
 CLKBUF_X1 hold13 (.A(_0168_),
    .Z(net175));
 CLKBUF_X1 hold14 (.A(_0660_),
    .Z(net176));
 CLKBUF_X1 hold15 (.A(net160),
    .Z(net177));
 CLKBUF_X1 hold16 (.A(_0269_),
    .Z(net178));
 CLKBUF_X1 hold17 (.A(_0658_),
    .Z(net179));
 CLKBUF_X1 hold18 (.A(net158),
    .Z(net180));
 CLKBUF_X1 hold19 (.A(_0267_),
    .Z(net181));
 CLKBUF_X1 hold20 (.A(_0661_),
    .Z(net182));
 CLKBUF_X1 hold21 (.A(net157),
    .Z(net183));
 CLKBUF_X1 hold22 (.A(_0270_),
    .Z(net184));
 CLKBUF_X1 hold23 (.A(addr_ptr[3]),
    .Z(net185));
 CLKBUF_X1 hold24 (.A(net161),
    .Z(net186));
 CLKBUF_X1 hold25 (.A(_0657_),
    .Z(net187));
 CLKBUF_X1 hold26 (.A(net162),
    .Z(net188));
 CLKBUF_X1 hold27 (.A(_0654_),
    .Z(net189));
 CLKBUF_X1 hold28 (.A(_0418_),
    .Z(net190));
 CLKBUF_X1 hold29 (.A(_0167_),
    .Z(net191));
 CLKBUF_X1 hold30 (.A(curr_state[0]),
    .Z(net192));
 CLKBUF_X1 hold31 (.A(_0384_),
    .Z(net193));
 CLKBUF_X1 hold32 (.A(_0306_),
    .Z(net194));
 CLKBUF_X1 hold33 (.A(addr_ptr[4]),
    .Z(net195));
 CLKBUF_X1 hold34 (.A(net163),
    .Z(net196));
 CLKBUF_X1 hold35 (.A(addr_ptr[5]),
    .Z(net197));
 CLKBUF_X1 hold36 (.A(net164),
    .Z(net198));
 CLKBUF_X1 hold37 (.A(addr_ptr[1]),
    .Z(net199));
 CLKBUF_X1 hold38 (.A(net165),
    .Z(net200));
 CLKBUF_X1 hold39 (.A(addr_ptr[0]),
    .Z(net201));
 CLKBUF_X1 hold40 (.A(net166),
    .Z(net202));
 CLKBUF_X1 hold41 (.A(data_in_reg[24]),
    .Z(net203));
 CLKBUF_X1 hold42 (.A(data_in_reg[23]),
    .Z(net204));
 CLKBUF_X1 hold43 (.A(_0652_),
    .Z(net205));
 CLKBUF_X1 hold44 (.A(net167),
    .Z(net206));
 CLKBUF_X1 hold45 (.A(data_in_reg[15]),
    .Z(net207));
 CLKBUF_X1 hold46 (.A(data_in_reg[0]),
    .Z(net208));
 CLKBUF_X1 hold47 (.A(data_in_reg[12]),
    .Z(net209));
 CLKBUF_X1 hold48 (.A(data_in_reg[31]),
    .Z(net210));
 CLKBUF_X1 hold49 (.A(_0659_),
    .Z(net211));
 CLKBUF_X1 hold50 (.A(data_in_reg[22]),
    .Z(net212));
 CLKBUF_X1 hold51 (.A(_0653_),
    .Z(net213));
 CLKBUF_X1 hold52 (.A(data_in_reg[3]),
    .Z(net214));
 CLKBUF_X1 hold53 (.A(data_in_reg[28]),
    .Z(net215));
 CLKBUF_X1 hold54 (.A(data_in_reg[6]),
    .Z(net216));
 CLKBUF_X1 hold55 (.A(_0518_),
    .Z(net217));
 CLKBUF_X1 hold56 (.A(curr_state[2]),
    .Z(net218));
 CLKBUF_X1 hold57 (.A(data_in_reg[29]),
    .Z(net219));
 CLKBUF_X1 hold58 (.A(init_count[5]),
    .Z(net220));
 CLKBUF_X1 hold59 (.A(addr_ptr[1]),
    .Z(net221));
 CLKBUF_X1 hold60 (.A(init_count[4]),
    .Z(net222));
 FILLCELL_X4 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_8 ();
 FILLCELL_X4 FILLER_0_40 ();
 FILLCELL_X16 FILLER_0_47 ();
 FILLCELL_X8 FILLER_0_63 ();
 FILLCELL_X8 FILLER_0_80 ();
 FILLCELL_X2 FILLER_0_88 ();
 FILLCELL_X1 FILLER_0_90 ();
 FILLCELL_X4 FILLER_0_94 ();
 FILLCELL_X2 FILLER_0_98 ();
 FILLCELL_X1 FILLER_0_100 ();
 FILLCELL_X4 FILLER_0_104 ();
 FILLCELL_X4 FILLER_0_111 ();
 FILLCELL_X1 FILLER_0_115 ();
 FILLCELL_X4 FILLER_0_119 ();
 FILLCELL_X1 FILLER_0_123 ();
 FILLCELL_X8 FILLER_0_128 ();
 FILLCELL_X4 FILLER_0_136 ();
 FILLCELL_X1 FILLER_0_140 ();
 FILLCELL_X4 FILLER_0_145 ();
 FILLCELL_X8 FILLER_0_152 ();
 FILLCELL_X2 FILLER_0_160 ();
 FILLCELL_X1 FILLER_0_162 ();
 FILLCELL_X4 FILLER_0_167 ();
 FILLCELL_X2 FILLER_0_171 ();
 FILLCELL_X4 FILLER_0_180 ();
 FILLCELL_X2 FILLER_0_184 ();
 FILLCELL_X4 FILLER_0_189 ();
 FILLCELL_X8 FILLER_0_197 ();
 FILLCELL_X1 FILLER_0_205 ();
 FILLCELL_X8 FILLER_0_209 ();
 FILLCELL_X4 FILLER_0_221 ();
 FILLCELL_X4 FILLER_0_228 ();
 FILLCELL_X2 FILLER_0_232 ();
 FILLCELL_X1 FILLER_0_234 ();
 FILLCELL_X8 FILLER_0_239 ();
 FILLCELL_X2 FILLER_0_247 ();
 FILLCELL_X1 FILLER_0_249 ();
 FILLCELL_X4 FILLER_0_257 ();
 FILLCELL_X8 FILLER_0_264 ();
 FILLCELL_X4 FILLER_0_272 ();
 FILLCELL_X4 FILLER_0_280 ();
 FILLCELL_X4 FILLER_0_287 ();
 FILLCELL_X4 FILLER_0_294 ();
 FILLCELL_X2 FILLER_0_298 ();
 FILLCELL_X4 FILLER_0_304 ();
 FILLCELL_X1 FILLER_0_308 ();
 FILLCELL_X8 FILLER_0_312 ();
 FILLCELL_X4 FILLER_0_320 ();
 FILLCELL_X2 FILLER_0_324 ();
 FILLCELL_X1 FILLER_0_326 ();
 FILLCELL_X8 FILLER_0_330 ();
 FILLCELL_X4 FILLER_0_341 ();
 FILLCELL_X8 FILLER_0_352 ();
 FILLCELL_X4 FILLER_0_360 ();
 FILLCELL_X2 FILLER_0_364 ();
 FILLCELL_X1 FILLER_0_366 ();
 FILLCELL_X4 FILLER_0_371 ();
 FILLCELL_X4 FILLER_0_379 ();
 FILLCELL_X1 FILLER_0_383 ();
 FILLCELL_X4 FILLER_0_387 ();
 FILLCELL_X4 FILLER_0_394 ();
 FILLCELL_X4 FILLER_0_401 ();
 FILLCELL_X8 FILLER_0_409 ();
 FILLCELL_X2 FILLER_0_417 ();
 FILLCELL_X1 FILLER_0_419 ();
 FILLCELL_X4 FILLER_0_424 ();
 FILLCELL_X32 FILLER_0_432 ();
 FILLCELL_X8 FILLER_0_464 ();
 FILLCELL_X8 FILLER_0_476 ();
 FILLCELL_X2 FILLER_0_484 ();
 FILLCELL_X4 FILLER_0_489 ();
 FILLCELL_X4 FILLER_0_496 ();
 FILLCELL_X16 FILLER_0_504 ();
 FILLCELL_X1 FILLER_0_520 ();
 FILLCELL_X8 FILLER_0_525 ();
 FILLCELL_X2 FILLER_0_533 ();
 FILLCELL_X4 FILLER_0_540 ();
 FILLCELL_X4 FILLER_0_548 ();
 FILLCELL_X2 FILLER_0_552 ();
 FILLCELL_X4 FILLER_0_557 ();
 FILLCELL_X4 FILLER_0_564 ();
 FILLCELL_X8 FILLER_0_570 ();
 FILLCELL_X4 FILLER_0_578 ();
 FILLCELL_X2 FILLER_0_582 ();
 FILLCELL_X1 FILLER_0_584 ();
 FILLCELL_X8 FILLER_0_588 ();
 FILLCELL_X4 FILLER_0_600 ();
 FILLCELL_X1 FILLER_0_604 ();
 FILLCELL_X4 FILLER_0_608 ();
 FILLCELL_X4 FILLER_0_615 ();
 FILLCELL_X8 FILLER_0_623 ();
 FILLCELL_X4 FILLER_0_632 ();
 FILLCELL_X4 FILLER_0_639 ();
 FILLCELL_X4 FILLER_0_647 ();
 FILLCELL_X2 FILLER_0_651 ();
 FILLCELL_X8 FILLER_0_656 ();
 FILLCELL_X1 FILLER_0_664 ();
 FILLCELL_X8 FILLER_0_674 ();
 FILLCELL_X2 FILLER_0_682 ();
 FILLCELL_X4 FILLER_0_688 ();
 FILLCELL_X4 FILLER_0_695 ();
 FILLCELL_X4 FILLER_0_702 ();
 FILLCELL_X2 FILLER_0_706 ();
 FILLCELL_X4 FILLER_0_710 ();
 FILLCELL_X8 FILLER_0_721 ();
 FILLCELL_X2 FILLER_0_729 ();
 FILLCELL_X4 FILLER_0_734 ();
 FILLCELL_X4 FILLER_0_742 ();
 FILLCELL_X1 FILLER_0_746 ();
 FILLCELL_X8 FILLER_0_751 ();
 FILLCELL_X2 FILLER_0_759 ();
 FILLCELL_X4 FILLER_0_764 ();
 FILLCELL_X8 FILLER_0_771 ();
 FILLCELL_X8 FILLER_0_788 ();
 FILLCELL_X2 FILLER_0_796 ();
 FILLCELL_X8 FILLER_0_801 ();
 FILLCELL_X4 FILLER_0_809 ();
 FILLCELL_X2 FILLER_0_813 ();
 FILLCELL_X4 FILLER_0_818 ();
 FILLCELL_X4 FILLER_0_825 ();
 FILLCELL_X2 FILLER_0_829 ();
 FILLCELL_X1 FILLER_0_831 ();
 FILLCELL_X4 FILLER_0_842 ();
 FILLCELL_X2 FILLER_0_846 ();
 FILLCELL_X1 FILLER_0_848 ();
 FILLCELL_X4 FILLER_0_853 ();
 FILLCELL_X4 FILLER_0_861 ();
 FILLCELL_X2 FILLER_0_865 ();
 FILLCELL_X4 FILLER_0_870 ();
 FILLCELL_X2 FILLER_0_874 ();
 FILLCELL_X4 FILLER_0_883 ();
 FILLCELL_X4 FILLER_0_891 ();
 FILLCELL_X1 FILLER_0_895 ();
 FILLCELL_X4 FILLER_0_899 ();
 FILLCELL_X16 FILLER_0_906 ();
 FILLCELL_X4 FILLER_0_922 ();
 FILLCELL_X2 FILLER_0_926 ();
 FILLCELL_X8 FILLER_0_932 ();
 FILLCELL_X1 FILLER_0_940 ();
 FILLCELL_X4 FILLER_0_950 ();
 FILLCELL_X2 FILLER_0_954 ();
 FILLCELL_X8 FILLER_0_959 ();
 FILLCELL_X4 FILLER_0_971 ();
 FILLCELL_X4 FILLER_0_978 ();
 FILLCELL_X4 FILLER_0_985 ();
 FILLCELL_X4 FILLER_0_992 ();
 FILLCELL_X2 FILLER_0_996 ();
 FILLCELL_X4 FILLER_0_1002 ();
 FILLCELL_X4 FILLER_0_1009 ();
 FILLCELL_X2 FILLER_0_1013 ();
 FILLCELL_X4 FILLER_0_1019 ();
 FILLCELL_X4 FILLER_0_1026 ();
 FILLCELL_X4 FILLER_0_1033 ();
 FILLCELL_X8 FILLER_0_1041 ();
 FILLCELL_X1 FILLER_0_1049 ();
 FILLCELL_X4 FILLER_0_1054 ();
 FILLCELL_X16 FILLER_0_1061 ();
 FILLCELL_X4 FILLER_0_1086 ();
 FILLCELL_X2 FILLER_0_1090 ();
 FILLCELL_X4 FILLER_0_1101 ();
 FILLCELL_X4 FILLER_0_1108 ();
 FILLCELL_X2 FILLER_0_1112 ();
 FILLCELL_X4 FILLER_0_1118 ();
 FILLCELL_X8 FILLER_0_1125 ();
 FILLCELL_X4 FILLER_0_1133 ();
 FILLCELL_X2 FILLER_0_1137 ();
 FILLCELL_X4 FILLER_0_1143 ();
 FILLCELL_X8 FILLER_0_1150 ();
 FILLCELL_X4 FILLER_0_1158 ();
 FILLCELL_X1 FILLER_0_1162 ();
 FILLCELL_X4 FILLER_0_1167 ();
 FILLCELL_X4 FILLER_0_1174 ();
 FILLCELL_X4 FILLER_0_1181 ();
 FILLCELL_X4 FILLER_0_1187 ();
 FILLCELL_X4 FILLER_0_1195 ();
 FILLCELL_X8 FILLER_0_1206 ();
 FILLCELL_X2 FILLER_0_1214 ();
 FILLCELL_X8 FILLER_0_1220 ();
 FILLCELL_X2 FILLER_0_1228 ();
 FILLCELL_X4 FILLER_0_1234 ();
 FILLCELL_X4 FILLER_0_1245 ();
 FILLCELL_X4 FILLER_0_1258 ();
 FILLCELL_X4 FILLER_0_1263 ();
 FILLCELL_X4 FILLER_0_1270 ();
 FILLCELL_X4 FILLER_0_1277 ();
 FILLCELL_X4 FILLER_0_1284 ();
 FILLCELL_X4 FILLER_0_1297 ();
 FILLCELL_X4 FILLER_0_1304 ();
 FILLCELL_X4 FILLER_0_1310 ();
 FILLCELL_X2 FILLER_0_1314 ();
 FILLCELL_X4 FILLER_0_1323 ();
 FILLCELL_X4 FILLER_0_1330 ();
 FILLCELL_X1 FILLER_0_1334 ();
 FILLCELL_X4 FILLER_0_1339 ();
 FILLCELL_X4 FILLER_0_1346 ();
 FILLCELL_X16 FILLER_0_1353 ();
 FILLCELL_X4 FILLER_0_1373 ();
 FILLCELL_X2 FILLER_0_1377 ();
 FILLCELL_X1 FILLER_0_1379 ();
 FILLCELL_X4 FILLER_0_1384 ();
 FILLCELL_X32 FILLER_0_1391 ();
 FILLCELL_X32 FILLER_0_1423 ();
 FILLCELL_X4 FILLER_0_1455 ();
 FILLCELL_X32 FILLER_0_1462 ();
 FILLCELL_X32 FILLER_0_1494 ();
 FILLCELL_X4 FILLER_0_1526 ();
 FILLCELL_X32 FILLER_0_1533 ();
 FILLCELL_X32 FILLER_0_1565 ();
 FILLCELL_X2 FILLER_0_1597 ();
 FILLCELL_X1 FILLER_0_1599 ();
 FILLCELL_X32 FILLER_0_1603 ();
 FILLCELL_X32 FILLER_0_1635 ();
 FILLCELL_X4 FILLER_0_1667 ();
 FILLCELL_X32 FILLER_0_1674 ();
 FILLCELL_X32 FILLER_0_1706 ();
 FILLCELL_X4 FILLER_0_1738 ();
 FILLCELL_X8 FILLER_0_1745 ();
 FILLCELL_X2 FILLER_0_1753 ();
 FILLCELL_X1 FILLER_0_1755 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X16 FILLER_1_33 ();
 FILLCELL_X8 FILLER_1_49 ();
 FILLCELL_X4 FILLER_1_57 ();
 FILLCELL_X4 FILLER_1_64 ();
 FILLCELL_X4 FILLER_1_77 ();
 FILLCELL_X4 FILLER_1_85 ();
 FILLCELL_X4 FILLER_1_99 ();
 FILLCELL_X4 FILLER_1_107 ();
 FILLCELL_X2 FILLER_1_111 ();
 FILLCELL_X4 FILLER_1_122 ();
 FILLCELL_X1 FILLER_1_126 ();
 FILLCELL_X8 FILLER_1_136 ();
 FILLCELL_X2 FILLER_1_144 ();
 FILLCELL_X1 FILLER_1_146 ();
 FILLCELL_X8 FILLER_1_157 ();
 FILLCELL_X2 FILLER_1_165 ();
 FILLCELL_X4 FILLER_1_177 ();
 FILLCELL_X4 FILLER_1_191 ();
 FILLCELL_X2 FILLER_1_195 ();
 FILLCELL_X4 FILLER_1_201 ();
 FILLCELL_X8 FILLER_1_214 ();
 FILLCELL_X1 FILLER_1_222 ();
 FILLCELL_X4 FILLER_1_232 ();
 FILLCELL_X2 FILLER_1_236 ();
 FILLCELL_X8 FILLER_1_248 ();
 FILLCELL_X1 FILLER_1_256 ();
 FILLCELL_X4 FILLER_1_267 ();
 FILLCELL_X4 FILLER_1_275 ();
 FILLCELL_X4 FILLER_1_288 ();
 FILLCELL_X2 FILLER_1_292 ();
 FILLCELL_X4 FILLER_1_298 ();
 FILLCELL_X4 FILLER_1_311 ();
 FILLCELL_X2 FILLER_1_315 ();
 FILLCELL_X4 FILLER_1_326 ();
 FILLCELL_X4 FILLER_1_334 ();
 FILLCELL_X4 FILLER_1_348 ();
 FILLCELL_X2 FILLER_1_352 ();
 FILLCELL_X8 FILLER_1_364 ();
 FILLCELL_X1 FILLER_1_372 ();
 FILLCELL_X4 FILLER_1_382 ();
 FILLCELL_X1 FILLER_1_386 ();
 FILLCELL_X4 FILLER_1_391 ();
 FILLCELL_X4 FILLER_1_404 ();
 FILLCELL_X8 FILLER_1_417 ();
 FILLCELL_X1 FILLER_1_425 ();
 FILLCELL_X16 FILLER_1_445 ();
 FILLCELL_X1 FILLER_1_461 ();
 FILLCELL_X4 FILLER_1_465 ();
 FILLCELL_X4 FILLER_1_478 ();
 FILLCELL_X4 FILLER_1_486 ();
 FILLCELL_X4 FILLER_1_493 ();
 FILLCELL_X4 FILLER_1_506 ();
 FILLCELL_X4 FILLER_1_514 ();
 FILLCELL_X2 FILLER_1_518 ();
 FILLCELL_X1 FILLER_1_520 ();
 FILLCELL_X4 FILLER_1_526 ();
 FILLCELL_X4 FILLER_1_539 ();
 FILLCELL_X4 FILLER_1_552 ();
 FILLCELL_X8 FILLER_1_566 ();
 FILLCELL_X1 FILLER_1_574 ();
 FILLCELL_X4 FILLER_1_579 ();
 FILLCELL_X1 FILLER_1_583 ();
 FILLCELL_X8 FILLER_1_594 ();
 FILLCELL_X1 FILLER_1_602 ();
 FILLCELL_X4 FILLER_1_612 ();
 FILLCELL_X4 FILLER_1_625 ();
 FILLCELL_X4 FILLER_1_638 ();
 FILLCELL_X8 FILLER_1_661 ();
 FILLCELL_X4 FILLER_1_679 ();
 FILLCELL_X2 FILLER_1_683 ();
 FILLCELL_X4 FILLER_1_695 ();
 FILLCELL_X4 FILLER_1_709 ();
 FILLCELL_X4 FILLER_1_723 ();
 FILLCELL_X2 FILLER_1_727 ();
 FILLCELL_X4 FILLER_1_732 ();
 FILLCELL_X8 FILLER_1_745 ();
 FILLCELL_X1 FILLER_1_753 ();
 FILLCELL_X4 FILLER_1_763 ();
 FILLCELL_X4 FILLER_1_771 ();
 FILLCELL_X8 FILLER_1_794 ();
 FILLCELL_X4 FILLER_1_807 ();
 FILLCELL_X4 FILLER_1_820 ();
 FILLCELL_X2 FILLER_1_824 ();
 FILLCELL_X1 FILLER_1_826 ();
 FILLCELL_X4 FILLER_1_830 ();
 FILLCELL_X2 FILLER_1_834 ();
 FILLCELL_X8 FILLER_1_846 ();
 FILLCELL_X1 FILLER_1_854 ();
 FILLCELL_X4 FILLER_1_865 ();
 FILLCELL_X2 FILLER_1_869 ();
 FILLCELL_X4 FILLER_1_880 ();
 FILLCELL_X4 FILLER_1_894 ();
 FILLCELL_X1 FILLER_1_898 ();
 FILLCELL_X4 FILLER_1_903 ();
 FILLCELL_X4 FILLER_1_911 ();
 FILLCELL_X4 FILLER_1_918 ();
 FILLCELL_X4 FILLER_1_926 ();
 FILLCELL_X4 FILLER_1_939 ();
 FILLCELL_X8 FILLER_1_947 ();
 FILLCELL_X4 FILLER_1_965 ();
 FILLCELL_X2 FILLER_1_969 ();
 FILLCELL_X1 FILLER_1_971 ();
 FILLCELL_X4 FILLER_1_976 ();
 FILLCELL_X2 FILLER_1_980 ();
 FILLCELL_X4 FILLER_1_986 ();
 FILLCELL_X2 FILLER_1_990 ();
 FILLCELL_X8 FILLER_1_996 ();
 FILLCELL_X8 FILLER_1_1013 ();
 FILLCELL_X4 FILLER_1_1030 ();
 FILLCELL_X2 FILLER_1_1034 ();
 FILLCELL_X8 FILLER_1_1046 ();
 FILLCELL_X2 FILLER_1_1054 ();
 FILLCELL_X8 FILLER_1_1075 ();
 FILLCELL_X1 FILLER_1_1083 ();
 FILLCELL_X4 FILLER_1_1087 ();
 FILLCELL_X4 FILLER_1_1110 ();
 FILLCELL_X4 FILLER_1_1124 ();
 FILLCELL_X4 FILLER_1_1138 ();
 FILLCELL_X4 FILLER_1_1151 ();
 FILLCELL_X4 FILLER_1_1164 ();
 FILLCELL_X1 FILLER_1_1168 ();
 FILLCELL_X4 FILLER_1_1178 ();
 FILLCELL_X4 FILLER_1_1191 ();
 FILLCELL_X2 FILLER_1_1195 ();
 FILLCELL_X4 FILLER_1_1207 ();
 FILLCELL_X4 FILLER_1_1230 ();
 FILLCELL_X8 FILLER_1_1253 ();
 FILLCELL_X2 FILLER_1_1261 ();
 FILLCELL_X4 FILLER_1_1264 ();
 FILLCELL_X4 FILLER_1_1277 ();
 FILLCELL_X8 FILLER_1_1290 ();
 FILLCELL_X1 FILLER_1_1298 ();
 FILLCELL_X8 FILLER_1_1309 ();
 FILLCELL_X4 FILLER_1_1327 ();
 FILLCELL_X4 FILLER_1_1335 ();
 FILLCELL_X1 FILLER_1_1339 ();
 FILLCELL_X4 FILLER_1_1349 ();
 FILLCELL_X4 FILLER_1_1362 ();
 FILLCELL_X8 FILLER_1_1370 ();
 FILLCELL_X2 FILLER_1_1378 ();
 FILLCELL_X4 FILLER_1_1389 ();
 FILLCELL_X4 FILLER_1_1396 ();
 FILLCELL_X32 FILLER_1_1403 ();
 FILLCELL_X32 FILLER_1_1435 ();
 FILLCELL_X32 FILLER_1_1467 ();
 FILLCELL_X32 FILLER_1_1499 ();
 FILLCELL_X32 FILLER_1_1531 ();
 FILLCELL_X32 FILLER_1_1563 ();
 FILLCELL_X32 FILLER_1_1595 ();
 FILLCELL_X32 FILLER_1_1627 ();
 FILLCELL_X32 FILLER_1_1659 ();
 FILLCELL_X32 FILLER_1_1691 ();
 FILLCELL_X16 FILLER_1_1723 ();
 FILLCELL_X8 FILLER_1_1739 ();
 FILLCELL_X1 FILLER_1_1747 ();
 FILLCELL_X4 FILLER_1_1752 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X16 FILLER_2_33 ();
 FILLCELL_X8 FILLER_2_49 ();
 FILLCELL_X4 FILLER_2_57 ();
 FILLCELL_X1 FILLER_2_61 ();
 FILLCELL_X4 FILLER_2_65 ();
 FILLCELL_X4 FILLER_2_72 ();
 FILLCELL_X4 FILLER_2_80 ();
 FILLCELL_X4 FILLER_2_88 ();
 FILLCELL_X2 FILLER_2_92 ();
 FILLCELL_X4 FILLER_2_101 ();
 FILLCELL_X2 FILLER_2_105 ();
 FILLCELL_X4 FILLER_2_111 ();
 FILLCELL_X4 FILLER_2_119 ();
 FILLCELL_X4 FILLER_2_126 ();
 FILLCELL_X2 FILLER_2_130 ();
 FILLCELL_X4 FILLER_2_136 ();
 FILLCELL_X4 FILLER_2_149 ();
 FILLCELL_X2 FILLER_2_153 ();
 FILLCELL_X1 FILLER_2_155 ();
 FILLCELL_X4 FILLER_2_163 ();
 FILLCELL_X1 FILLER_2_167 ();
 FILLCELL_X4 FILLER_2_171 ();
 FILLCELL_X4 FILLER_2_185 ();
 FILLCELL_X8 FILLER_2_192 ();
 FILLCELL_X2 FILLER_2_200 ();
 FILLCELL_X1 FILLER_2_202 ();
 FILLCELL_X4 FILLER_2_206 ();
 FILLCELL_X4 FILLER_2_213 ();
 FILLCELL_X8 FILLER_2_221 ();
 FILLCELL_X4 FILLER_2_233 ();
 FILLCELL_X2 FILLER_2_237 ();
 FILLCELL_X1 FILLER_2_239 ();
 FILLCELL_X8 FILLER_2_243 ();
 FILLCELL_X2 FILLER_2_251 ();
 FILLCELL_X4 FILLER_2_255 ();
 FILLCELL_X1 FILLER_2_259 ();
 FILLCELL_X4 FILLER_2_263 ();
 FILLCELL_X4 FILLER_2_270 ();
 FILLCELL_X4 FILLER_2_277 ();
 FILLCELL_X4 FILLER_2_285 ();
 FILLCELL_X8 FILLER_2_298 ();
 FILLCELL_X4 FILLER_2_310 ();
 FILLCELL_X4 FILLER_2_318 ();
 FILLCELL_X16 FILLER_2_332 ();
 FILLCELL_X2 FILLER_2_348 ();
 FILLCELL_X4 FILLER_2_352 ();
 FILLCELL_X1 FILLER_2_356 ();
 FILLCELL_X4 FILLER_2_360 ();
 FILLCELL_X4 FILLER_2_367 ();
 FILLCELL_X4 FILLER_2_374 ();
 FILLCELL_X4 FILLER_2_382 ();
 FILLCELL_X4 FILLER_2_389 ();
 FILLCELL_X1 FILLER_2_393 ();
 FILLCELL_X4 FILLER_2_398 ();
 FILLCELL_X8 FILLER_2_405 ();
 FILLCELL_X2 FILLER_2_413 ();
 FILLCELL_X4 FILLER_2_418 ();
 FILLCELL_X16 FILLER_2_432 ();
 FILLCELL_X1 FILLER_2_448 ();
 FILLCELL_X4 FILLER_2_453 ();
 FILLCELL_X8 FILLER_2_466 ();
 FILLCELL_X1 FILLER_2_474 ();
 FILLCELL_X8 FILLER_2_478 ();
 FILLCELL_X4 FILLER_2_486 ();
 FILLCELL_X2 FILLER_2_490 ();
 FILLCELL_X1 FILLER_2_492 ();
 FILLCELL_X4 FILLER_2_496 ();
 FILLCELL_X1 FILLER_2_500 ();
 FILLCELL_X16 FILLER_2_504 ();
 FILLCELL_X2 FILLER_2_520 ();
 FILLCELL_X1 FILLER_2_522 ();
 FILLCELL_X4 FILLER_2_527 ();
 FILLCELL_X4 FILLER_2_535 ();
 FILLCELL_X16 FILLER_2_541 ();
 FILLCELL_X2 FILLER_2_557 ();
 FILLCELL_X8 FILLER_2_562 ();
 FILLCELL_X2 FILLER_2_570 ();
 FILLCELL_X4 FILLER_2_574 ();
 FILLCELL_X4 FILLER_2_588 ();
 FILLCELL_X8 FILLER_2_595 ();
 FILLCELL_X2 FILLER_2_603 ();
 FILLCELL_X8 FILLER_2_609 ();
 FILLCELL_X2 FILLER_2_617 ();
 FILLCELL_X8 FILLER_2_623 ();
 FILLCELL_X4 FILLER_2_632 ();
 FILLCELL_X8 FILLER_2_639 ();
 FILLCELL_X4 FILLER_2_647 ();
 FILLCELL_X4 FILLER_2_654 ();
 FILLCELL_X2 FILLER_2_658 ();
 FILLCELL_X4 FILLER_2_663 ();
 FILLCELL_X8 FILLER_2_670 ();
 FILLCELL_X1 FILLER_2_678 ();
 FILLCELL_X4 FILLER_2_681 ();
 FILLCELL_X4 FILLER_2_689 ();
 FILLCELL_X1 FILLER_2_693 ();
 FILLCELL_X8 FILLER_2_704 ();
 FILLCELL_X4 FILLER_2_716 ();
 FILLCELL_X4 FILLER_2_724 ();
 FILLCELL_X4 FILLER_2_737 ();
 FILLCELL_X4 FILLER_2_744 ();
 FILLCELL_X2 FILLER_2_748 ();
 FILLCELL_X4 FILLER_2_754 ();
 FILLCELL_X8 FILLER_2_767 ();
 FILLCELL_X4 FILLER_2_779 ();
 FILLCELL_X4 FILLER_2_787 ();
 FILLCELL_X4 FILLER_2_795 ();
 FILLCELL_X4 FILLER_2_804 ();
 FILLCELL_X4 FILLER_2_817 ();
 FILLCELL_X2 FILLER_2_821 ();
 FILLCELL_X1 FILLER_2_823 ();
 FILLCELL_X4 FILLER_2_826 ();
 FILLCELL_X4 FILLER_2_839 ();
 FILLCELL_X16 FILLER_2_846 ();
 FILLCELL_X2 FILLER_2_862 ();
 FILLCELL_X1 FILLER_2_864 ();
 FILLCELL_X8 FILLER_2_867 ();
 FILLCELL_X4 FILLER_2_875 ();
 FILLCELL_X1 FILLER_2_879 ();
 FILLCELL_X4 FILLER_2_883 ();
 FILLCELL_X4 FILLER_2_890 ();
 FILLCELL_X1 FILLER_2_894 ();
 FILLCELL_X4 FILLER_2_899 ();
 FILLCELL_X2 FILLER_2_903 ();
 FILLCELL_X4 FILLER_2_914 ();
 FILLCELL_X4 FILLER_2_923 ();
 FILLCELL_X1 FILLER_2_927 ();
 FILLCELL_X4 FILLER_2_931 ();
 FILLCELL_X8 FILLER_2_938 ();
 FILLCELL_X1 FILLER_2_946 ();
 FILLCELL_X4 FILLER_2_954 ();
 FILLCELL_X8 FILLER_2_968 ();
 FILLCELL_X2 FILLER_2_976 ();
 FILLCELL_X4 FILLER_2_987 ();
 FILLCELL_X4 FILLER_2_1000 ();
 FILLCELL_X8 FILLER_2_1007 ();
 FILLCELL_X2 FILLER_2_1015 ();
 FILLCELL_X16 FILLER_2_1020 ();
 FILLCELL_X4 FILLER_2_1036 ();
 FILLCELL_X4 FILLER_2_1047 ();
 FILLCELL_X8 FILLER_2_1053 ();
 FILLCELL_X2 FILLER_2_1061 ();
 FILLCELL_X1 FILLER_2_1063 ();
 FILLCELL_X4 FILLER_2_1067 ();
 FILLCELL_X4 FILLER_2_1075 ();
 FILLCELL_X4 FILLER_2_1083 ();
 FILLCELL_X2 FILLER_2_1087 ();
 FILLCELL_X1 FILLER_2_1089 ();
 FILLCELL_X4 FILLER_2_1094 ();
 FILLCELL_X8 FILLER_2_1102 ();
 FILLCELL_X4 FILLER_2_1117 ();
 FILLCELL_X16 FILLER_2_1131 ();
 FILLCELL_X1 FILLER_2_1147 ();
 FILLCELL_X4 FILLER_2_1152 ();
 FILLCELL_X8 FILLER_2_1159 ();
 FILLCELL_X1 FILLER_2_1167 ();
 FILLCELL_X4 FILLER_2_1172 ();
 FILLCELL_X1 FILLER_2_1176 ();
 FILLCELL_X4 FILLER_2_1180 ();
 FILLCELL_X1 FILLER_2_1184 ();
 FILLCELL_X4 FILLER_2_1188 ();
 FILLCELL_X4 FILLER_2_1195 ();
 FILLCELL_X4 FILLER_2_1203 ();
 FILLCELL_X16 FILLER_2_1210 ();
 FILLCELL_X4 FILLER_2_1226 ();
 FILLCELL_X1 FILLER_2_1230 ();
 FILLCELL_X8 FILLER_2_1235 ();
 FILLCELL_X4 FILLER_2_1243 ();
 FILLCELL_X1 FILLER_2_1247 ();
 FILLCELL_X4 FILLER_2_1252 ();
 FILLCELL_X4 FILLER_2_1260 ();
 FILLCELL_X4 FILLER_2_1268 ();
 FILLCELL_X8 FILLER_2_1275 ();
 FILLCELL_X1 FILLER_2_1283 ();
 FILLCELL_X4 FILLER_2_1294 ();
 FILLCELL_X8 FILLER_2_1301 ();
 FILLCELL_X2 FILLER_2_1309 ();
 FILLCELL_X4 FILLER_2_1315 ();
 FILLCELL_X1 FILLER_2_1319 ();
 FILLCELL_X16 FILLER_2_1323 ();
 FILLCELL_X8 FILLER_2_1339 ();
 FILLCELL_X4 FILLER_2_1347 ();
 FILLCELL_X4 FILLER_2_1354 ();
 FILLCELL_X1 FILLER_2_1358 ();
 FILLCELL_X4 FILLER_2_1361 ();
 FILLCELL_X8 FILLER_2_1372 ();
 FILLCELL_X4 FILLER_2_1389 ();
 FILLCELL_X4 FILLER_2_1397 ();
 FILLCELL_X32 FILLER_2_1404 ();
 FILLCELL_X32 FILLER_2_1436 ();
 FILLCELL_X32 FILLER_2_1468 ();
 FILLCELL_X32 FILLER_2_1500 ();
 FILLCELL_X32 FILLER_2_1532 ();
 FILLCELL_X32 FILLER_2_1564 ();
 FILLCELL_X32 FILLER_2_1596 ();
 FILLCELL_X32 FILLER_2_1628 ();
 FILLCELL_X32 FILLER_2_1660 ();
 FILLCELL_X32 FILLER_2_1692 ();
 FILLCELL_X32 FILLER_2_1724 ();
 FILLCELL_X16 FILLER_3_1 ();
 FILLCELL_X2 FILLER_3_17 ();
 FILLCELL_X1 FILLER_3_19 ();
 FILLCELL_X16 FILLER_3_24 ();
 FILLCELL_X8 FILLER_3_40 ();
 FILLCELL_X2 FILLER_3_48 ();
 FILLCELL_X1 FILLER_3_50 ();
 FILLCELL_X32 FILLER_3_54 ();
 FILLCELL_X8 FILLER_3_86 ();
 FILLCELL_X4 FILLER_3_96 ();
 FILLCELL_X16 FILLER_3_110 ();
 FILLCELL_X2 FILLER_3_126 ();
 FILLCELL_X1 FILLER_3_128 ();
 FILLCELL_X4 FILLER_3_138 ();
 FILLCELL_X4 FILLER_3_145 ();
 FILLCELL_X1 FILLER_3_149 ();
 FILLCELL_X4 FILLER_3_153 ();
 FILLCELL_X4 FILLER_3_166 ();
 FILLCELL_X8 FILLER_3_172 ();
 FILLCELL_X2 FILLER_3_180 ();
 FILLCELL_X4 FILLER_3_184 ();
 FILLCELL_X2 FILLER_3_188 ();
 FILLCELL_X4 FILLER_3_193 ();
 FILLCELL_X4 FILLER_3_201 ();
 FILLCELL_X4 FILLER_3_214 ();
 FILLCELL_X4 FILLER_3_227 ();
 FILLCELL_X4 FILLER_3_241 ();
 FILLCELL_X2 FILLER_3_245 ();
 FILLCELL_X4 FILLER_3_249 ();
 FILLCELL_X4 FILLER_3_263 ();
 FILLCELL_X16 FILLER_3_276 ();
 FILLCELL_X8 FILLER_3_292 ();
 FILLCELL_X1 FILLER_3_300 ();
 FILLCELL_X16 FILLER_3_304 ();
 FILLCELL_X4 FILLER_3_320 ();
 FILLCELL_X4 FILLER_3_327 ();
 FILLCELL_X2 FILLER_3_331 ();
 FILLCELL_X4 FILLER_3_340 ();
 FILLCELL_X1 FILLER_3_344 ();
 FILLCELL_X4 FILLER_3_347 ();
 FILLCELL_X4 FILLER_3_361 ();
 FILLCELL_X4 FILLER_3_374 ();
 FILLCELL_X2 FILLER_3_378 ();
 FILLCELL_X1 FILLER_3_380 ();
 FILLCELL_X16 FILLER_3_390 ();
 FILLCELL_X4 FILLER_3_406 ();
 FILLCELL_X16 FILLER_3_413 ();
 FILLCELL_X8 FILLER_3_429 ();
 FILLCELL_X16 FILLER_3_439 ();
 FILLCELL_X16 FILLER_3_459 ();
 FILLCELL_X4 FILLER_3_479 ();
 FILLCELL_X8 FILLER_3_492 ();
 FILLCELL_X32 FILLER_3_504 ();
 FILLCELL_X2 FILLER_3_536 ();
 FILLCELL_X16 FILLER_3_541 ();
 FILLCELL_X8 FILLER_3_560 ();
 FILLCELL_X2 FILLER_3_568 ();
 FILLCELL_X8 FILLER_3_580 ();
 FILLCELL_X4 FILLER_3_588 ();
 FILLCELL_X1 FILLER_3_592 ();
 FILLCELL_X8 FILLER_3_600 ();
 FILLCELL_X4 FILLER_3_612 ();
 FILLCELL_X4 FILLER_3_619 ();
 FILLCELL_X2 FILLER_3_623 ();
 FILLCELL_X4 FILLER_3_628 ();
 FILLCELL_X4 FILLER_3_636 ();
 FILLCELL_X8 FILLER_3_649 ();
 FILLCELL_X1 FILLER_3_657 ();
 FILLCELL_X16 FILLER_3_661 ();
 FILLCELL_X4 FILLER_3_677 ();
 FILLCELL_X2 FILLER_3_681 ();
 FILLCELL_X1 FILLER_3_683 ();
 FILLCELL_X8 FILLER_3_686 ();
 FILLCELL_X4 FILLER_3_701 ();
 FILLCELL_X1 FILLER_3_705 ();
 FILLCELL_X16 FILLER_3_709 ();
 FILLCELL_X4 FILLER_3_728 ();
 FILLCELL_X2 FILLER_3_732 ();
 FILLCELL_X32 FILLER_3_737 ();
 FILLCELL_X16 FILLER_3_772 ();
 FILLCELL_X4 FILLER_3_788 ();
 FILLCELL_X4 FILLER_3_796 ();
 FILLCELL_X1 FILLER_3_800 ();
 FILLCELL_X4 FILLER_3_805 ();
 FILLCELL_X16 FILLER_3_811 ();
 FILLCELL_X4 FILLER_3_827 ();
 FILLCELL_X16 FILLER_3_834 ();
 FILLCELL_X4 FILLER_3_850 ();
 FILLCELL_X2 FILLER_3_854 ();
 FILLCELL_X4 FILLER_3_866 ();
 FILLCELL_X4 FILLER_3_873 ();
 FILLCELL_X4 FILLER_3_886 ();
 FILLCELL_X4 FILLER_3_895 ();
 FILLCELL_X2 FILLER_3_899 ();
 FILLCELL_X4 FILLER_3_910 ();
 FILLCELL_X8 FILLER_3_917 ();
 FILLCELL_X2 FILLER_3_925 ();
 FILLCELL_X4 FILLER_3_931 ();
 FILLCELL_X2 FILLER_3_935 ();
 FILLCELL_X1 FILLER_3_937 ();
 FILLCELL_X16 FILLER_3_941 ();
 FILLCELL_X2 FILLER_3_957 ();
 FILLCELL_X8 FILLER_3_961 ();
 FILLCELL_X4 FILLER_3_969 ();
 FILLCELL_X2 FILLER_3_973 ();
 FILLCELL_X4 FILLER_3_979 ();
 FILLCELL_X4 FILLER_3_986 ();
 FILLCELL_X1 FILLER_3_990 ();
 FILLCELL_X4 FILLER_3_995 ();
 FILLCELL_X4 FILLER_3_1002 ();
 FILLCELL_X2 FILLER_3_1006 ();
 FILLCELL_X4 FILLER_3_1012 ();
 FILLCELL_X16 FILLER_3_1026 ();
 FILLCELL_X2 FILLER_3_1042 ();
 FILLCELL_X8 FILLER_3_1054 ();
 FILLCELL_X4 FILLER_3_1062 ();
 FILLCELL_X1 FILLER_3_1066 ();
 FILLCELL_X4 FILLER_3_1070 ();
 FILLCELL_X32 FILLER_3_1077 ();
 FILLCELL_X8 FILLER_3_1109 ();
 FILLCELL_X4 FILLER_3_1117 ();
 FILLCELL_X1 FILLER_3_1121 ();
 FILLCELL_X16 FILLER_3_1124 ();
 FILLCELL_X4 FILLER_3_1140 ();
 FILLCELL_X2 FILLER_3_1144 ();
 FILLCELL_X8 FILLER_3_1150 ();
 FILLCELL_X1 FILLER_3_1158 ();
 FILLCELL_X8 FILLER_3_1162 ();
 FILLCELL_X4 FILLER_3_1170 ();
 FILLCELL_X4 FILLER_3_1178 ();
 FILLCELL_X2 FILLER_3_1182 ();
 FILLCELL_X8 FILLER_3_1194 ();
 FILLCELL_X4 FILLER_3_1202 ();
 FILLCELL_X2 FILLER_3_1206 ();
 FILLCELL_X4 FILLER_3_1218 ();
 FILLCELL_X4 FILLER_3_1224 ();
 FILLCELL_X1 FILLER_3_1228 ();
 FILLCELL_X4 FILLER_3_1239 ();
 FILLCELL_X16 FILLER_3_1246 ();
 FILLCELL_X1 FILLER_3_1262 ();
 FILLCELL_X16 FILLER_3_1264 ();
 FILLCELL_X4 FILLER_3_1280 ();
 FILLCELL_X2 FILLER_3_1284 ();
 FILLCELL_X8 FILLER_3_1288 ();
 FILLCELL_X1 FILLER_3_1296 ();
 FILLCELL_X4 FILLER_3_1301 ();
 FILLCELL_X2 FILLER_3_1305 ();
 FILLCELL_X1 FILLER_3_1307 ();
 FILLCELL_X8 FILLER_3_1310 ();
 FILLCELL_X4 FILLER_3_1318 ();
 FILLCELL_X8 FILLER_3_1331 ();
 FILLCELL_X2 FILLER_3_1339 ();
 FILLCELL_X8 FILLER_3_1344 ();
 FILLCELL_X2 FILLER_3_1352 ();
 FILLCELL_X1 FILLER_3_1354 ();
 FILLCELL_X4 FILLER_3_1365 ();
 FILLCELL_X8 FILLER_3_1379 ();
 FILLCELL_X32 FILLER_3_1391 ();
 FILLCELL_X32 FILLER_3_1423 ();
 FILLCELL_X32 FILLER_3_1455 ();
 FILLCELL_X32 FILLER_3_1487 ();
 FILLCELL_X32 FILLER_3_1519 ();
 FILLCELL_X32 FILLER_3_1551 ();
 FILLCELL_X32 FILLER_3_1583 ();
 FILLCELL_X32 FILLER_3_1615 ();
 FILLCELL_X32 FILLER_3_1647 ();
 FILLCELL_X32 FILLER_3_1679 ();
 FILLCELL_X32 FILLER_3_1711 ();
 FILLCELL_X8 FILLER_3_1743 ();
 FILLCELL_X4 FILLER_3_1751 ();
 FILLCELL_X1 FILLER_3_1755 ();
 FILLCELL_X16 FILLER_4_1 ();
 FILLCELL_X1 FILLER_4_17 ();
 FILLCELL_X8 FILLER_4_37 ();
 FILLCELL_X4 FILLER_4_49 ();
 FILLCELL_X2 FILLER_4_53 ();
 FILLCELL_X1 FILLER_4_55 ();
 FILLCELL_X8 FILLER_4_60 ();
 FILLCELL_X4 FILLER_4_68 ();
 FILLCELL_X2 FILLER_4_72 ();
 FILLCELL_X1 FILLER_4_74 ();
 FILLCELL_X4 FILLER_4_79 ();
 FILLCELL_X4 FILLER_4_86 ();
 FILLCELL_X2 FILLER_4_90 ();
 FILLCELL_X4 FILLER_4_99 ();
 FILLCELL_X8 FILLER_4_105 ();
 FILLCELL_X4 FILLER_4_113 ();
 FILLCELL_X1 FILLER_4_117 ();
 FILLCELL_X4 FILLER_4_121 ();
 FILLCELL_X4 FILLER_4_129 ();
 FILLCELL_X8 FILLER_4_137 ();
 FILLCELL_X4 FILLER_4_145 ();
 FILLCELL_X1 FILLER_4_149 ();
 FILLCELL_X16 FILLER_4_153 ();
 FILLCELL_X4 FILLER_4_169 ();
 FILLCELL_X1 FILLER_4_173 ();
 FILLCELL_X4 FILLER_4_177 ();
 FILLCELL_X8 FILLER_4_190 ();
 FILLCELL_X4 FILLER_4_198 ();
 FILLCELL_X16 FILLER_4_206 ();
 FILLCELL_X8 FILLER_4_222 ();
 FILLCELL_X2 FILLER_4_230 ();
 FILLCELL_X1 FILLER_4_232 ();
 FILLCELL_X4 FILLER_4_236 ();
 FILLCELL_X2 FILLER_4_240 ();
 FILLCELL_X1 FILLER_4_242 ();
 FILLCELL_X8 FILLER_4_250 ();
 FILLCELL_X2 FILLER_4_258 ();
 FILLCELL_X4 FILLER_4_263 ();
 FILLCELL_X2 FILLER_4_267 ();
 FILLCELL_X4 FILLER_4_272 ();
 FILLCELL_X1 FILLER_4_276 ();
 FILLCELL_X16 FILLER_4_286 ();
 FILLCELL_X4 FILLER_4_302 ();
 FILLCELL_X1 FILLER_4_306 ();
 FILLCELL_X4 FILLER_4_311 ();
 FILLCELL_X8 FILLER_4_317 ();
 FILLCELL_X2 FILLER_4_325 ();
 FILLCELL_X1 FILLER_4_327 ();
 FILLCELL_X4 FILLER_4_331 ();
 FILLCELL_X8 FILLER_4_344 ();
 FILLCELL_X4 FILLER_4_352 ();
 FILLCELL_X1 FILLER_4_356 ();
 FILLCELL_X16 FILLER_4_360 ();
 FILLCELL_X4 FILLER_4_376 ();
 FILLCELL_X2 FILLER_4_380 ();
 FILLCELL_X1 FILLER_4_382 ();
 FILLCELL_X4 FILLER_4_387 ();
 FILLCELL_X4 FILLER_4_395 ();
 FILLCELL_X1 FILLER_4_399 ();
 FILLCELL_X4 FILLER_4_404 ();
 FILLCELL_X4 FILLER_4_418 ();
 FILLCELL_X2 FILLER_4_422 ();
 FILLCELL_X4 FILLER_4_431 ();
 FILLCELL_X4 FILLER_4_445 ();
 FILLCELL_X2 FILLER_4_449 ();
 FILLCELL_X1 FILLER_4_451 ();
 FILLCELL_X4 FILLER_4_456 ();
 FILLCELL_X4 FILLER_4_463 ();
 FILLCELL_X4 FILLER_4_471 ();
 FILLCELL_X8 FILLER_4_478 ();
 FILLCELL_X2 FILLER_4_486 ();
 FILLCELL_X1 FILLER_4_488 ();
 FILLCELL_X4 FILLER_4_492 ();
 FILLCELL_X4 FILLER_4_500 ();
 FILLCELL_X4 FILLER_4_513 ();
 FILLCELL_X4 FILLER_4_521 ();
 FILLCELL_X2 FILLER_4_525 ();
 FILLCELL_X1 FILLER_4_527 ();
 FILLCELL_X4 FILLER_4_532 ();
 FILLCELL_X4 FILLER_4_540 ();
 FILLCELL_X1 FILLER_4_544 ();
 FILLCELL_X4 FILLER_4_548 ();
 FILLCELL_X4 FILLER_4_561 ();
 FILLCELL_X2 FILLER_4_565 ();
 FILLCELL_X1 FILLER_4_567 ();
 FILLCELL_X8 FILLER_4_571 ();
 FILLCELL_X2 FILLER_4_579 ();
 FILLCELL_X1 FILLER_4_581 ();
 FILLCELL_X4 FILLER_4_589 ();
 FILLCELL_X1 FILLER_4_593 ();
 FILLCELL_X8 FILLER_4_604 ();
 FILLCELL_X2 FILLER_4_612 ();
 FILLCELL_X8 FILLER_4_623 ();
 FILLCELL_X16 FILLER_4_632 ();
 FILLCELL_X2 FILLER_4_648 ();
 FILLCELL_X4 FILLER_4_659 ();
 FILLCELL_X8 FILLER_4_666 ();
 FILLCELL_X1 FILLER_4_674 ();
 FILLCELL_X4 FILLER_4_685 ();
 FILLCELL_X1 FILLER_4_689 ();
 FILLCELL_X4 FILLER_4_700 ();
 FILLCELL_X8 FILLER_4_707 ();
 FILLCELL_X2 FILLER_4_715 ();
 FILLCELL_X1 FILLER_4_717 ();
 FILLCELL_X4 FILLER_4_724 ();
 FILLCELL_X8 FILLER_4_731 ();
 FILLCELL_X1 FILLER_4_739 ();
 FILLCELL_X4 FILLER_4_743 ();
 FILLCELL_X4 FILLER_4_751 ();
 FILLCELL_X4 FILLER_4_759 ();
 FILLCELL_X2 FILLER_4_763 ();
 FILLCELL_X1 FILLER_4_765 ();
 FILLCELL_X8 FILLER_4_770 ();
 FILLCELL_X4 FILLER_4_785 ();
 FILLCELL_X8 FILLER_4_792 ();
 FILLCELL_X1 FILLER_4_800 ();
 FILLCELL_X4 FILLER_4_810 ();
 FILLCELL_X2 FILLER_4_814 ();
 FILLCELL_X4 FILLER_4_819 ();
 FILLCELL_X2 FILLER_4_823 ();
 FILLCELL_X1 FILLER_4_825 ();
 FILLCELL_X4 FILLER_4_829 ();
 FILLCELL_X4 FILLER_4_835 ();
 FILLCELL_X8 FILLER_4_849 ();
 FILLCELL_X32 FILLER_4_864 ();
 FILLCELL_X16 FILLER_4_896 ();
 FILLCELL_X8 FILLER_4_912 ();
 FILLCELL_X1 FILLER_4_920 ();
 FILLCELL_X4 FILLER_4_925 ();
 FILLCELL_X4 FILLER_4_938 ();
 FILLCELL_X4 FILLER_4_946 ();
 FILLCELL_X1 FILLER_4_950 ();
 FILLCELL_X4 FILLER_4_954 ();
 FILLCELL_X2 FILLER_4_958 ();
 FILLCELL_X1 FILLER_4_960 ();
 FILLCELL_X4 FILLER_4_963 ();
 FILLCELL_X1 FILLER_4_967 ();
 FILLCELL_X16 FILLER_4_972 ();
 FILLCELL_X4 FILLER_4_992 ();
 FILLCELL_X1 FILLER_4_996 ();
 FILLCELL_X8 FILLER_4_1006 ();
 FILLCELL_X2 FILLER_4_1014 ();
 FILLCELL_X1 FILLER_4_1016 ();
 FILLCELL_X4 FILLER_4_1024 ();
 FILLCELL_X8 FILLER_4_1030 ();
 FILLCELL_X2 FILLER_4_1038 ();
 FILLCELL_X1 FILLER_4_1040 ();
 FILLCELL_X8 FILLER_4_1050 ();
 FILLCELL_X4 FILLER_4_1058 ();
 FILLCELL_X8 FILLER_4_1065 ();
 FILLCELL_X1 FILLER_4_1073 ();
 FILLCELL_X8 FILLER_4_1078 ();
 FILLCELL_X1 FILLER_4_1086 ();
 FILLCELL_X4 FILLER_4_1091 ();
 FILLCELL_X4 FILLER_4_1098 ();
 FILLCELL_X8 FILLER_4_1111 ();
 FILLCELL_X1 FILLER_4_1119 ();
 FILLCELL_X4 FILLER_4_1127 ();
 FILLCELL_X4 FILLER_4_1135 ();
 FILLCELL_X8 FILLER_4_1143 ();
 FILLCELL_X2 FILLER_4_1151 ();
 FILLCELL_X4 FILLER_4_1157 ();
 FILLCELL_X1 FILLER_4_1161 ();
 FILLCELL_X4 FILLER_4_1166 ();
 FILLCELL_X2 FILLER_4_1170 ();
 FILLCELL_X4 FILLER_4_1175 ();
 FILLCELL_X2 FILLER_4_1179 ();
 FILLCELL_X1 FILLER_4_1181 ();
 FILLCELL_X16 FILLER_4_1184 ();
 FILLCELL_X4 FILLER_4_1200 ();
 FILLCELL_X2 FILLER_4_1204 ();
 FILLCELL_X1 FILLER_4_1206 ();
 FILLCELL_X16 FILLER_4_1211 ();
 FILLCELL_X4 FILLER_4_1234 ();
 FILLCELL_X4 FILLER_4_1240 ();
 FILLCELL_X4 FILLER_4_1253 ();
 FILLCELL_X2 FILLER_4_1257 ();
 FILLCELL_X1 FILLER_4_1259 ();
 FILLCELL_X4 FILLER_4_1264 ();
 FILLCELL_X4 FILLER_4_1271 ();
 FILLCELL_X2 FILLER_4_1275 ();
 FILLCELL_X1 FILLER_4_1277 ();
 FILLCELL_X4 FILLER_4_1281 ();
 FILLCELL_X8 FILLER_4_1295 ();
 FILLCELL_X1 FILLER_4_1303 ();
 FILLCELL_X4 FILLER_4_1310 ();
 FILLCELL_X4 FILLER_4_1320 ();
 FILLCELL_X8 FILLER_4_1327 ();
 FILLCELL_X2 FILLER_4_1335 ();
 FILLCELL_X4 FILLER_4_1346 ();
 FILLCELL_X4 FILLER_4_1353 ();
 FILLCELL_X2 FILLER_4_1357 ();
 FILLCELL_X1 FILLER_4_1359 ();
 FILLCELL_X4 FILLER_4_1364 ();
 FILLCELL_X1 FILLER_4_1368 ();
 FILLCELL_X4 FILLER_4_1372 ();
 FILLCELL_X2 FILLER_4_1376 ();
 FILLCELL_X1 FILLER_4_1378 ();
 FILLCELL_X4 FILLER_4_1383 ();
 FILLCELL_X4 FILLER_4_1391 ();
 FILLCELL_X4 FILLER_4_1400 ();
 FILLCELL_X32 FILLER_4_1406 ();
 FILLCELL_X32 FILLER_4_1438 ();
 FILLCELL_X32 FILLER_4_1470 ();
 FILLCELL_X32 FILLER_4_1502 ();
 FILLCELL_X32 FILLER_4_1534 ();
 FILLCELL_X32 FILLER_4_1566 ();
 FILLCELL_X32 FILLER_4_1598 ();
 FILLCELL_X32 FILLER_4_1630 ();
 FILLCELL_X32 FILLER_4_1662 ();
 FILLCELL_X32 FILLER_4_1694 ();
 FILLCELL_X16 FILLER_4_1726 ();
 FILLCELL_X8 FILLER_4_1742 ();
 FILLCELL_X4 FILLER_4_1750 ();
 FILLCELL_X2 FILLER_4_1754 ();
 FILLCELL_X16 FILLER_5_1 ();
 FILLCELL_X8 FILLER_5_17 ();
 FILLCELL_X4 FILLER_5_25 ();
 FILLCELL_X2 FILLER_5_29 ();
 FILLCELL_X4 FILLER_5_35 ();
 FILLCELL_X4 FILLER_5_48 ();
 FILLCELL_X4 FILLER_5_61 ();
 FILLCELL_X2 FILLER_5_65 ();
 FILLCELL_X1 FILLER_5_67 ();
 FILLCELL_X8 FILLER_5_72 ();
 FILLCELL_X8 FILLER_5_90 ();
 FILLCELL_X4 FILLER_5_98 ();
 FILLCELL_X1 FILLER_5_102 ();
 FILLCELL_X4 FILLER_5_113 ();
 FILLCELL_X4 FILLER_5_120 ();
 FILLCELL_X1 FILLER_5_124 ();
 FILLCELL_X16 FILLER_5_128 ();
 FILLCELL_X4 FILLER_5_148 ();
 FILLCELL_X1 FILLER_5_152 ();
 FILLCELL_X4 FILLER_5_156 ();
 FILLCELL_X4 FILLER_5_167 ();
 FILLCELL_X2 FILLER_5_171 ();
 FILLCELL_X8 FILLER_5_183 ();
 FILLCELL_X16 FILLER_5_200 ();
 FILLCELL_X8 FILLER_5_216 ();
 FILLCELL_X4 FILLER_5_224 ();
 FILLCELL_X2 FILLER_5_228 ();
 FILLCELL_X4 FILLER_5_232 ();
 FILLCELL_X8 FILLER_5_239 ();
 FILLCELL_X1 FILLER_5_247 ();
 FILLCELL_X4 FILLER_5_257 ();
 FILLCELL_X8 FILLER_5_264 ();
 FILLCELL_X1 FILLER_5_272 ();
 FILLCELL_X4 FILLER_5_276 ();
 FILLCELL_X4 FILLER_5_283 ();
 FILLCELL_X1 FILLER_5_287 ();
 FILLCELL_X4 FILLER_5_298 ();
 FILLCELL_X4 FILLER_5_321 ();
 FILLCELL_X4 FILLER_5_335 ();
 FILLCELL_X4 FILLER_5_348 ();
 FILLCELL_X8 FILLER_5_355 ();
 FILLCELL_X1 FILLER_5_363 ();
 FILLCELL_X4 FILLER_5_367 ();
 FILLCELL_X8 FILLER_5_380 ();
 FILLCELL_X1 FILLER_5_388 ();
 FILLCELL_X4 FILLER_5_398 ();
 FILLCELL_X4 FILLER_5_406 ();
 FILLCELL_X1 FILLER_5_410 ();
 FILLCELL_X4 FILLER_5_414 ();
 FILLCELL_X4 FILLER_5_425 ();
 FILLCELL_X2 FILLER_5_429 ();
 FILLCELL_X4 FILLER_5_433 ();
 FILLCELL_X8 FILLER_5_447 ();
 FILLCELL_X2 FILLER_5_455 ();
 FILLCELL_X1 FILLER_5_457 ();
 FILLCELL_X4 FILLER_5_467 ();
 FILLCELL_X1 FILLER_5_471 ();
 FILLCELL_X4 FILLER_5_476 ();
 FILLCELL_X8 FILLER_5_490 ();
 FILLCELL_X4 FILLER_5_498 ();
 FILLCELL_X4 FILLER_5_505 ();
 FILLCELL_X4 FILLER_5_512 ();
 FILLCELL_X8 FILLER_5_525 ();
 FILLCELL_X1 FILLER_5_533 ();
 FILLCELL_X4 FILLER_5_543 ();
 FILLCELL_X1 FILLER_5_547 ();
 FILLCELL_X4 FILLER_5_552 ();
 FILLCELL_X8 FILLER_5_566 ();
 FILLCELL_X4 FILLER_5_584 ();
 FILLCELL_X4 FILLER_5_592 ();
 FILLCELL_X2 FILLER_5_596 ();
 FILLCELL_X4 FILLER_5_601 ();
 FILLCELL_X8 FILLER_5_608 ();
 FILLCELL_X2 FILLER_5_616 ();
 FILLCELL_X4 FILLER_5_622 ();
 FILLCELL_X8 FILLER_5_635 ();
 FILLCELL_X4 FILLER_5_643 ();
 FILLCELL_X2 FILLER_5_647 ();
 FILLCELL_X4 FILLER_5_653 ();
 FILLCELL_X8 FILLER_5_661 ();
 FILLCELL_X2 FILLER_5_669 ();
 FILLCELL_X1 FILLER_5_671 ();
 FILLCELL_X4 FILLER_5_681 ();
 FILLCELL_X1 FILLER_5_685 ();
 FILLCELL_X4 FILLER_5_696 ();
 FILLCELL_X8 FILLER_5_710 ();
 FILLCELL_X4 FILLER_5_724 ();
 FILLCELL_X4 FILLER_5_745 ();
 FILLCELL_X2 FILLER_5_749 ();
 FILLCELL_X4 FILLER_5_760 ();
 FILLCELL_X4 FILLER_5_766 ();
 FILLCELL_X4 FILLER_5_774 ();
 FILLCELL_X4 FILLER_5_788 ();
 FILLCELL_X2 FILLER_5_792 ();
 FILLCELL_X8 FILLER_5_798 ();
 FILLCELL_X1 FILLER_5_806 ();
 FILLCELL_X4 FILLER_5_811 ();
 FILLCELL_X2 FILLER_5_815 ();
 FILLCELL_X4 FILLER_5_821 ();
 FILLCELL_X4 FILLER_5_835 ();
 FILLCELL_X2 FILLER_5_839 ();
 FILLCELL_X4 FILLER_5_851 ();
 FILLCELL_X8 FILLER_5_857 ();
 FILLCELL_X1 FILLER_5_865 ();
 FILLCELL_X4 FILLER_5_870 ();
 FILLCELL_X4 FILLER_5_878 ();
 FILLCELL_X4 FILLER_5_886 ();
 FILLCELL_X4 FILLER_5_893 ();
 FILLCELL_X4 FILLER_5_901 ();
 FILLCELL_X8 FILLER_5_912 ();
 FILLCELL_X4 FILLER_5_920 ();
 FILLCELL_X2 FILLER_5_924 ();
 FILLCELL_X1 FILLER_5_926 ();
 FILLCELL_X8 FILLER_5_930 ();
 FILLCELL_X2 FILLER_5_938 ();
 FILLCELL_X4 FILLER_5_949 ();
 FILLCELL_X2 FILLER_5_953 ();
 FILLCELL_X1 FILLER_5_955 ();
 FILLCELL_X4 FILLER_5_966 ();
 FILLCELL_X2 FILLER_5_970 ();
 FILLCELL_X1 FILLER_5_972 ();
 FILLCELL_X4 FILLER_5_977 ();
 FILLCELL_X4 FILLER_5_985 ();
 FILLCELL_X4 FILLER_5_992 ();
 FILLCELL_X16 FILLER_5_1005 ();
 FILLCELL_X8 FILLER_5_1021 ();
 FILLCELL_X4 FILLER_5_1039 ();
 FILLCELL_X4 FILLER_5_1052 ();
 FILLCELL_X1 FILLER_5_1056 ();
 FILLCELL_X4 FILLER_5_1061 ();
 FILLCELL_X4 FILLER_5_1074 ();
 FILLCELL_X4 FILLER_5_1087 ();
 FILLCELL_X8 FILLER_5_1100 ();
 FILLCELL_X8 FILLER_5_1118 ();
 FILLCELL_X4 FILLER_5_1126 ();
 FILLCELL_X2 FILLER_5_1130 ();
 FILLCELL_X4 FILLER_5_1141 ();
 FILLCELL_X4 FILLER_5_1149 ();
 FILLCELL_X4 FILLER_5_1156 ();
 FILLCELL_X1 FILLER_5_1160 ();
 FILLCELL_X4 FILLER_5_1170 ();
 FILLCELL_X8 FILLER_5_1177 ();
 FILLCELL_X1 FILLER_5_1185 ();
 FILLCELL_X4 FILLER_5_1193 ();
 FILLCELL_X4 FILLER_5_1201 ();
 FILLCELL_X1 FILLER_5_1205 ();
 FILLCELL_X4 FILLER_5_1215 ();
 FILLCELL_X4 FILLER_5_1222 ();
 FILLCELL_X4 FILLER_5_1229 ();
 FILLCELL_X2 FILLER_5_1233 ();
 FILLCELL_X1 FILLER_5_1235 ();
 FILLCELL_X4 FILLER_5_1240 ();
 FILLCELL_X4 FILLER_5_1246 ();
 FILLCELL_X1 FILLER_5_1250 ();
 FILLCELL_X8 FILLER_5_1255 ();
 FILLCELL_X4 FILLER_5_1264 ();
 FILLCELL_X4 FILLER_5_1277 ();
 FILLCELL_X4 FILLER_5_1290 ();
 FILLCELL_X8 FILLER_5_1298 ();
 FILLCELL_X4 FILLER_5_1306 ();
 FILLCELL_X2 FILLER_5_1310 ();
 FILLCELL_X8 FILLER_5_1316 ();
 FILLCELL_X4 FILLER_5_1324 ();
 FILLCELL_X2 FILLER_5_1328 ();
 FILLCELL_X1 FILLER_5_1330 ();
 FILLCELL_X8 FILLER_5_1334 ();
 FILLCELL_X4 FILLER_5_1342 ();
 FILLCELL_X2 FILLER_5_1346 ();
 FILLCELL_X4 FILLER_5_1350 ();
 FILLCELL_X2 FILLER_5_1354 ();
 FILLCELL_X8 FILLER_5_1359 ();
 FILLCELL_X4 FILLER_5_1367 ();
 FILLCELL_X4 FILLER_5_1374 ();
 FILLCELL_X4 FILLER_5_1387 ();
 FILLCELL_X2 FILLER_5_1391 ();
 FILLCELL_X1 FILLER_5_1393 ();
 FILLCELL_X4 FILLER_5_1401 ();
 FILLCELL_X32 FILLER_5_1410 ();
 FILLCELL_X32 FILLER_5_1442 ();
 FILLCELL_X32 FILLER_5_1474 ();
 FILLCELL_X32 FILLER_5_1506 ();
 FILLCELL_X32 FILLER_5_1538 ();
 FILLCELL_X32 FILLER_5_1570 ();
 FILLCELL_X32 FILLER_5_1602 ();
 FILLCELL_X32 FILLER_5_1634 ();
 FILLCELL_X32 FILLER_5_1666 ();
 FILLCELL_X32 FILLER_5_1698 ();
 FILLCELL_X16 FILLER_5_1730 ();
 FILLCELL_X8 FILLER_5_1746 ();
 FILLCELL_X2 FILLER_5_1754 ();
 FILLCELL_X4 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_8 ();
 FILLCELL_X4 FILLER_6_40 ();
 FILLCELL_X4 FILLER_6_47 ();
 FILLCELL_X4 FILLER_6_54 ();
 FILLCELL_X1 FILLER_6_58 ();
 FILLCELL_X4 FILLER_6_62 ();
 FILLCELL_X4 FILLER_6_76 ();
 FILLCELL_X8 FILLER_6_82 ();
 FILLCELL_X1 FILLER_6_90 ();
 FILLCELL_X4 FILLER_6_94 ();
 FILLCELL_X1 FILLER_6_98 ();
 FILLCELL_X4 FILLER_6_102 ();
 FILLCELL_X4 FILLER_6_115 ();
 FILLCELL_X4 FILLER_6_122 ();
 FILLCELL_X2 FILLER_6_126 ();
 FILLCELL_X8 FILLER_6_132 ();
 FILLCELL_X4 FILLER_6_143 ();
 FILLCELL_X4 FILLER_6_157 ();
 FILLCELL_X4 FILLER_6_170 ();
 FILLCELL_X4 FILLER_6_176 ();
 FILLCELL_X2 FILLER_6_180 ();
 FILLCELL_X4 FILLER_6_185 ();
 FILLCELL_X4 FILLER_6_192 ();
 FILLCELL_X2 FILLER_6_196 ();
 FILLCELL_X4 FILLER_6_201 ();
 FILLCELL_X8 FILLER_6_215 ();
 FILLCELL_X4 FILLER_6_227 ();
 FILLCELL_X2 FILLER_6_231 ();
 FILLCELL_X1 FILLER_6_233 ();
 FILLCELL_X4 FILLER_6_244 ();
 FILLCELL_X2 FILLER_6_248 ();
 FILLCELL_X1 FILLER_6_250 ();
 FILLCELL_X4 FILLER_6_254 ();
 FILLCELL_X2 FILLER_6_258 ();
 FILLCELL_X1 FILLER_6_260 ();
 FILLCELL_X4 FILLER_6_264 ();
 FILLCELL_X2 FILLER_6_268 ();
 FILLCELL_X1 FILLER_6_270 ();
 FILLCELL_X4 FILLER_6_273 ();
 FILLCELL_X4 FILLER_6_287 ();
 FILLCELL_X8 FILLER_6_300 ();
 FILLCELL_X2 FILLER_6_308 ();
 FILLCELL_X16 FILLER_6_313 ();
 FILLCELL_X1 FILLER_6_329 ();
 FILLCELL_X4 FILLER_6_333 ();
 FILLCELL_X16 FILLER_6_347 ();
 FILLCELL_X2 FILLER_6_363 ();
 FILLCELL_X1 FILLER_6_365 ();
 FILLCELL_X8 FILLER_6_376 ();
 FILLCELL_X2 FILLER_6_384 ();
 FILLCELL_X4 FILLER_6_389 ();
 FILLCELL_X4 FILLER_6_396 ();
 FILLCELL_X8 FILLER_6_409 ();
 FILLCELL_X8 FILLER_6_426 ();
 FILLCELL_X4 FILLER_6_437 ();
 FILLCELL_X4 FILLER_6_450 ();
 FILLCELL_X2 FILLER_6_454 ();
 FILLCELL_X1 FILLER_6_456 ();
 FILLCELL_X8 FILLER_6_460 ();
 FILLCELL_X4 FILLER_6_477 ();
 FILLCELL_X2 FILLER_6_481 ();
 FILLCELL_X4 FILLER_6_490 ();
 FILLCELL_X16 FILLER_6_504 ();
 FILLCELL_X8 FILLER_6_520 ();
 FILLCELL_X2 FILLER_6_528 ();
 FILLCELL_X4 FILLER_6_533 ();
 FILLCELL_X8 FILLER_6_546 ();
 FILLCELL_X4 FILLER_6_554 ();
 FILLCELL_X1 FILLER_6_558 ();
 FILLCELL_X4 FILLER_6_566 ();
 FILLCELL_X8 FILLER_6_572 ();
 FILLCELL_X4 FILLER_6_582 ();
 FILLCELL_X8 FILLER_6_596 ();
 FILLCELL_X4 FILLER_6_608 ();
 FILLCELL_X8 FILLER_6_616 ();
 FILLCELL_X4 FILLER_6_627 ();
 FILLCELL_X4 FILLER_6_632 ();
 FILLCELL_X8 FILLER_6_643 ();
 FILLCELL_X4 FILLER_6_651 ();
 FILLCELL_X1 FILLER_6_655 ();
 FILLCELL_X4 FILLER_6_665 ();
 FILLCELL_X4 FILLER_6_672 ();
 FILLCELL_X4 FILLER_6_679 ();
 FILLCELL_X8 FILLER_6_686 ();
 FILLCELL_X2 FILLER_6_694 ();
 FILLCELL_X1 FILLER_6_696 ();
 FILLCELL_X8 FILLER_6_699 ();
 FILLCELL_X4 FILLER_6_707 ();
 FILLCELL_X4 FILLER_6_715 ();
 FILLCELL_X4 FILLER_6_732 ();
 FILLCELL_X8 FILLER_6_740 ();
 FILLCELL_X4 FILLER_6_752 ();
 FILLCELL_X2 FILLER_6_756 ();
 FILLCELL_X1 FILLER_6_758 ();
 FILLCELL_X4 FILLER_6_762 ();
 FILLCELL_X2 FILLER_6_766 ();
 FILLCELL_X4 FILLER_6_777 ();
 FILLCELL_X2 FILLER_6_781 ();
 FILLCELL_X4 FILLER_6_786 ();
 FILLCELL_X4 FILLER_6_794 ();
 FILLCELL_X4 FILLER_6_807 ();
 FILLCELL_X8 FILLER_6_820 ();
 FILLCELL_X4 FILLER_6_828 ();
 FILLCELL_X8 FILLER_6_839 ();
 FILLCELL_X4 FILLER_6_850 ();
 FILLCELL_X4 FILLER_6_864 ();
 FILLCELL_X4 FILLER_6_877 ();
 FILLCELL_X4 FILLER_6_890 ();
 FILLCELL_X4 FILLER_6_904 ();
 FILLCELL_X16 FILLER_6_918 ();
 FILLCELL_X4 FILLER_6_937 ();
 FILLCELL_X4 FILLER_6_944 ();
 FILLCELL_X4 FILLER_6_955 ();
 FILLCELL_X8 FILLER_6_969 ();
 FILLCELL_X2 FILLER_6_977 ();
 FILLCELL_X4 FILLER_6_988 ();
 FILLCELL_X8 FILLER_6_995 ();
 FILLCELL_X4 FILLER_6_1003 ();
 FILLCELL_X2 FILLER_6_1007 ();
 FILLCELL_X1 FILLER_6_1009 ();
 FILLCELL_X4 FILLER_6_1014 ();
 FILLCELL_X1 FILLER_6_1018 ();
 FILLCELL_X8 FILLER_6_1021 ();
 FILLCELL_X4 FILLER_6_1029 ();
 FILLCELL_X2 FILLER_6_1033 ();
 FILLCELL_X1 FILLER_6_1035 ();
 FILLCELL_X4 FILLER_6_1039 ();
 FILLCELL_X4 FILLER_6_1046 ();
 FILLCELL_X8 FILLER_6_1053 ();
 FILLCELL_X2 FILLER_6_1061 ();
 FILLCELL_X1 FILLER_6_1063 ();
 FILLCELL_X4 FILLER_6_1068 ();
 FILLCELL_X16 FILLER_6_1075 ();
 FILLCELL_X1 FILLER_6_1091 ();
 FILLCELL_X4 FILLER_6_1095 ();
 FILLCELL_X2 FILLER_6_1099 ();
 FILLCELL_X1 FILLER_6_1101 ();
 FILLCELL_X4 FILLER_6_1106 ();
 FILLCELL_X4 FILLER_6_1113 ();
 FILLCELL_X4 FILLER_6_1120 ();
 FILLCELL_X4 FILLER_6_1127 ();
 FILLCELL_X4 FILLER_6_1135 ();
 FILLCELL_X8 FILLER_6_1148 ();
 FILLCELL_X2 FILLER_6_1156 ();
 FILLCELL_X1 FILLER_6_1158 ();
 FILLCELL_X4 FILLER_6_1162 ();
 FILLCELL_X8 FILLER_6_1175 ();
 FILLCELL_X2 FILLER_6_1183 ();
 FILLCELL_X1 FILLER_6_1185 ();
 FILLCELL_X4 FILLER_6_1196 ();
 FILLCELL_X8 FILLER_6_1204 ();
 FILLCELL_X8 FILLER_6_1221 ();
 FILLCELL_X1 FILLER_6_1229 ();
 FILLCELL_X8 FILLER_6_1234 ();
 FILLCELL_X4 FILLER_6_1251 ();
 FILLCELL_X4 FILLER_6_1258 ();
 FILLCELL_X4 FILLER_6_1265 ();
 FILLCELL_X1 FILLER_6_1269 ();
 FILLCELL_X4 FILLER_6_1273 ();
 FILLCELL_X8 FILLER_6_1280 ();
 FILLCELL_X4 FILLER_6_1288 ();
 FILLCELL_X2 FILLER_6_1292 ();
 FILLCELL_X4 FILLER_6_1298 ();
 FILLCELL_X8 FILLER_6_1306 ();
 FILLCELL_X2 FILLER_6_1314 ();
 FILLCELL_X1 FILLER_6_1316 ();
 FILLCELL_X4 FILLER_6_1320 ();
 FILLCELL_X1 FILLER_6_1324 ();
 FILLCELL_X4 FILLER_6_1327 ();
 FILLCELL_X4 FILLER_6_1341 ();
 FILLCELL_X4 FILLER_6_1355 ();
 FILLCELL_X4 FILLER_6_1369 ();
 FILLCELL_X8 FILLER_6_1382 ();
 FILLCELL_X4 FILLER_6_1390 ();
 FILLCELL_X1 FILLER_6_1394 ();
 FILLCELL_X32 FILLER_6_1412 ();
 FILLCELL_X32 FILLER_6_1444 ();
 FILLCELL_X32 FILLER_6_1476 ();
 FILLCELL_X32 FILLER_6_1508 ();
 FILLCELL_X32 FILLER_6_1540 ();
 FILLCELL_X32 FILLER_6_1572 ();
 FILLCELL_X32 FILLER_6_1604 ();
 FILLCELL_X32 FILLER_6_1636 ();
 FILLCELL_X32 FILLER_6_1668 ();
 FILLCELL_X32 FILLER_6_1700 ();
 FILLCELL_X16 FILLER_6_1732 ();
 FILLCELL_X8 FILLER_6_1748 ();
 FILLCELL_X8 FILLER_7_1 ();
 FILLCELL_X4 FILLER_7_9 ();
 FILLCELL_X16 FILLER_7_30 ();
 FILLCELL_X4 FILLER_7_46 ();
 FILLCELL_X2 FILLER_7_50 ();
 FILLCELL_X16 FILLER_7_55 ();
 FILLCELL_X2 FILLER_7_71 ();
 FILLCELL_X1 FILLER_7_73 ();
 FILLCELL_X4 FILLER_7_81 ();
 FILLCELL_X4 FILLER_7_94 ();
 FILLCELL_X8 FILLER_7_108 ();
 FILLCELL_X1 FILLER_7_116 ();
 FILLCELL_X4 FILLER_7_120 ();
 FILLCELL_X4 FILLER_7_128 ();
 FILLCELL_X16 FILLER_7_141 ();
 FILLCELL_X8 FILLER_7_157 ();
 FILLCELL_X2 FILLER_7_165 ();
 FILLCELL_X8 FILLER_7_169 ();
 FILLCELL_X1 FILLER_7_177 ();
 FILLCELL_X8 FILLER_7_180 ();
 FILLCELL_X4 FILLER_7_188 ();
 FILLCELL_X2 FILLER_7_192 ();
 FILLCELL_X1 FILLER_7_194 ();
 FILLCELL_X4 FILLER_7_198 ();
 FILLCELL_X4 FILLER_7_205 ();
 FILLCELL_X4 FILLER_7_218 ();
 FILLCELL_X2 FILLER_7_222 ();
 FILLCELL_X4 FILLER_7_234 ();
 FILLCELL_X1 FILLER_7_238 ();
 FILLCELL_X4 FILLER_7_242 ();
 FILLCELL_X4 FILLER_7_255 ();
 FILLCELL_X4 FILLER_7_269 ();
 FILLCELL_X8 FILLER_7_280 ();
 FILLCELL_X4 FILLER_7_291 ();
 FILLCELL_X2 FILLER_7_295 ();
 FILLCELL_X4 FILLER_7_306 ();
 FILLCELL_X4 FILLER_7_320 ();
 FILLCELL_X2 FILLER_7_324 ();
 FILLCELL_X4 FILLER_7_333 ();
 FILLCELL_X4 FILLER_7_347 ();
 FILLCELL_X2 FILLER_7_351 ();
 FILLCELL_X1 FILLER_7_353 ();
 FILLCELL_X4 FILLER_7_358 ();
 FILLCELL_X4 FILLER_7_372 ();
 FILLCELL_X4 FILLER_7_379 ();
 FILLCELL_X2 FILLER_7_383 ();
 FILLCELL_X16 FILLER_7_388 ();
 FILLCELL_X2 FILLER_7_404 ();
 FILLCELL_X4 FILLER_7_409 ();
 FILLCELL_X4 FILLER_7_416 ();
 FILLCELL_X16 FILLER_7_429 ();
 FILLCELL_X4 FILLER_7_445 ();
 FILLCELL_X1 FILLER_7_449 ();
 FILLCELL_X16 FILLER_7_453 ();
 FILLCELL_X8 FILLER_7_469 ();
 FILLCELL_X4 FILLER_7_477 ();
 FILLCELL_X4 FILLER_7_484 ();
 FILLCELL_X2 FILLER_7_488 ();
 FILLCELL_X1 FILLER_7_490 ();
 FILLCELL_X4 FILLER_7_493 ();
 FILLCELL_X1 FILLER_7_497 ();
 FILLCELL_X4 FILLER_7_501 ();
 FILLCELL_X8 FILLER_7_508 ();
 FILLCELL_X4 FILLER_7_516 ();
 FILLCELL_X1 FILLER_7_520 ();
 FILLCELL_X16 FILLER_7_524 ();
 FILLCELL_X4 FILLER_7_540 ();
 FILLCELL_X4 FILLER_7_547 ();
 FILLCELL_X16 FILLER_7_555 ();
 FILLCELL_X8 FILLER_7_581 ();
 FILLCELL_X4 FILLER_7_593 ();
 FILLCELL_X1 FILLER_7_597 ();
 FILLCELL_X4 FILLER_7_604 ();
 FILLCELL_X4 FILLER_7_621 ();
 FILLCELL_X1 FILLER_7_625 ();
 FILLCELL_X4 FILLER_7_628 ();
 FILLCELL_X1 FILLER_7_632 ();
 FILLCELL_X4 FILLER_7_643 ();
 FILLCELL_X8 FILLER_7_651 ();
 FILLCELL_X2 FILLER_7_659 ();
 FILLCELL_X4 FILLER_7_664 ();
 FILLCELL_X4 FILLER_7_671 ();
 FILLCELL_X1 FILLER_7_675 ();
 FILLCELL_X4 FILLER_7_679 ();
 FILLCELL_X16 FILLER_7_687 ();
 FILLCELL_X8 FILLER_7_703 ();
 FILLCELL_X2 FILLER_7_711 ();
 FILLCELL_X1 FILLER_7_713 ();
 FILLCELL_X32 FILLER_7_717 ();
 FILLCELL_X4 FILLER_7_749 ();
 FILLCELL_X1 FILLER_7_753 ();
 FILLCELL_X32 FILLER_7_757 ();
 FILLCELL_X4 FILLER_7_789 ();
 FILLCELL_X2 FILLER_7_793 ();
 FILLCELL_X4 FILLER_7_798 ();
 FILLCELL_X2 FILLER_7_802 ();
 FILLCELL_X8 FILLER_7_807 ();
 FILLCELL_X4 FILLER_7_815 ();
 FILLCELL_X16 FILLER_7_823 ();
 FILLCELL_X2 FILLER_7_839 ();
 FILLCELL_X8 FILLER_7_844 ();
 FILLCELL_X2 FILLER_7_852 ();
 FILLCELL_X4 FILLER_7_864 ();
 FILLCELL_X2 FILLER_7_868 ();
 FILLCELL_X4 FILLER_7_873 ();
 FILLCELL_X4 FILLER_7_880 ();
 FILLCELL_X1 FILLER_7_884 ();
 FILLCELL_X8 FILLER_7_889 ();
 FILLCELL_X4 FILLER_7_897 ();
 FILLCELL_X2 FILLER_7_901 ();
 FILLCELL_X1 FILLER_7_903 ();
 FILLCELL_X4 FILLER_7_907 ();
 FILLCELL_X8 FILLER_7_913 ();
 FILLCELL_X4 FILLER_7_921 ();
 FILLCELL_X4 FILLER_7_928 ();
 FILLCELL_X32 FILLER_7_942 ();
 FILLCELL_X8 FILLER_7_974 ();
 FILLCELL_X4 FILLER_7_985 ();
 FILLCELL_X8 FILLER_7_992 ();
 FILLCELL_X4 FILLER_7_1003 ();
 FILLCELL_X8 FILLER_7_1017 ();
 FILLCELL_X1 FILLER_7_1025 ();
 FILLCELL_X4 FILLER_7_1029 ();
 FILLCELL_X2 FILLER_7_1033 ();
 FILLCELL_X8 FILLER_7_1045 ();
 FILLCELL_X4 FILLER_7_1053 ();
 FILLCELL_X1 FILLER_7_1057 ();
 FILLCELL_X4 FILLER_7_1062 ();
 FILLCELL_X4 FILLER_7_1069 ();
 FILLCELL_X8 FILLER_7_1076 ();
 FILLCELL_X16 FILLER_7_1087 ();
 FILLCELL_X8 FILLER_7_1103 ();
 FILLCELL_X4 FILLER_7_1111 ();
 FILLCELL_X2 FILLER_7_1115 ();
 FILLCELL_X16 FILLER_7_1119 ();
 FILLCELL_X8 FILLER_7_1138 ();
 FILLCELL_X4 FILLER_7_1146 ();
 FILLCELL_X2 FILLER_7_1150 ();
 FILLCELL_X1 FILLER_7_1152 ();
 FILLCELL_X8 FILLER_7_1156 ();
 FILLCELL_X4 FILLER_7_1164 ();
 FILLCELL_X4 FILLER_7_1175 ();
 FILLCELL_X4 FILLER_7_1182 ();
 FILLCELL_X4 FILLER_7_1188 ();
 FILLCELL_X2 FILLER_7_1192 ();
 FILLCELL_X4 FILLER_7_1198 ();
 FILLCELL_X2 FILLER_7_1202 ();
 FILLCELL_X4 FILLER_7_1207 ();
 FILLCELL_X4 FILLER_7_1214 ();
 FILLCELL_X4 FILLER_7_1222 ();
 FILLCELL_X4 FILLER_7_1236 ();
 FILLCELL_X8 FILLER_7_1243 ();
 FILLCELL_X1 FILLER_7_1251 ();
 FILLCELL_X8 FILLER_7_1255 ();
 FILLCELL_X4 FILLER_7_1264 ();
 FILLCELL_X4 FILLER_7_1272 ();
 FILLCELL_X4 FILLER_7_1278 ();
 FILLCELL_X2 FILLER_7_1282 ();
 FILLCELL_X1 FILLER_7_1284 ();
 FILLCELL_X4 FILLER_7_1291 ();
 FILLCELL_X4 FILLER_7_1302 ();
 FILLCELL_X4 FILLER_7_1312 ();
 FILLCELL_X4 FILLER_7_1323 ();
 FILLCELL_X4 FILLER_7_1330 ();
 FILLCELL_X2 FILLER_7_1334 ();
 FILLCELL_X1 FILLER_7_1336 ();
 FILLCELL_X8 FILLER_7_1344 ();
 FILLCELL_X1 FILLER_7_1352 ();
 FILLCELL_X16 FILLER_7_1357 ();
 FILLCELL_X2 FILLER_7_1373 ();
 FILLCELL_X4 FILLER_7_1378 ();
 FILLCELL_X16 FILLER_7_1385 ();
 FILLCELL_X8 FILLER_7_1401 ();
 FILLCELL_X2 FILLER_7_1409 ();
 FILLCELL_X32 FILLER_7_1430 ();
 FILLCELL_X32 FILLER_7_1462 ();
 FILLCELL_X32 FILLER_7_1494 ();
 FILLCELL_X32 FILLER_7_1526 ();
 FILLCELL_X32 FILLER_7_1558 ();
 FILLCELL_X32 FILLER_7_1590 ();
 FILLCELL_X32 FILLER_7_1622 ();
 FILLCELL_X32 FILLER_7_1654 ();
 FILLCELL_X32 FILLER_7_1686 ();
 FILLCELL_X32 FILLER_7_1718 ();
 FILLCELL_X4 FILLER_7_1750 ();
 FILLCELL_X2 FILLER_7_1754 ();
 FILLCELL_X4 FILLER_8_1 ();
 FILLCELL_X16 FILLER_8_8 ();
 FILLCELL_X4 FILLER_8_24 ();
 FILLCELL_X1 FILLER_8_28 ();
 FILLCELL_X4 FILLER_8_46 ();
 FILLCELL_X2 FILLER_8_50 ();
 FILLCELL_X4 FILLER_8_56 ();
 FILLCELL_X4 FILLER_8_69 ();
 FILLCELL_X8 FILLER_8_77 ();
 FILLCELL_X2 FILLER_8_85 ();
 FILLCELL_X8 FILLER_8_90 ();
 FILLCELL_X4 FILLER_8_98 ();
 FILLCELL_X2 FILLER_8_102 ();
 FILLCELL_X4 FILLER_8_107 ();
 FILLCELL_X8 FILLER_8_120 ();
 FILLCELL_X1 FILLER_8_128 ();
 FILLCELL_X4 FILLER_8_138 ();
 FILLCELL_X8 FILLER_8_145 ();
 FILLCELL_X4 FILLER_8_153 ();
 FILLCELL_X2 FILLER_8_157 ();
 FILLCELL_X4 FILLER_8_162 ();
 FILLCELL_X4 FILLER_8_176 ();
 FILLCELL_X4 FILLER_8_190 ();
 FILLCELL_X2 FILLER_8_194 ();
 FILLCELL_X4 FILLER_8_205 ();
 FILLCELL_X8 FILLER_8_212 ();
 FILLCELL_X4 FILLER_8_222 ();
 FILLCELL_X4 FILLER_8_230 ();
 FILLCELL_X16 FILLER_8_244 ();
 FILLCELL_X8 FILLER_8_260 ();
 FILLCELL_X4 FILLER_8_268 ();
 FILLCELL_X1 FILLER_8_272 ();
 FILLCELL_X4 FILLER_8_276 ();
 FILLCELL_X4 FILLER_8_283 ();
 FILLCELL_X16 FILLER_8_293 ();
 FILLCELL_X16 FILLER_8_316 ();
 FILLCELL_X4 FILLER_8_332 ();
 FILLCELL_X2 FILLER_8_336 ();
 FILLCELL_X8 FILLER_8_341 ();
 FILLCELL_X8 FILLER_8_352 ();
 FILLCELL_X1 FILLER_8_360 ();
 FILLCELL_X4 FILLER_8_368 ();
 FILLCELL_X4 FILLER_8_374 ();
 FILLCELL_X2 FILLER_8_378 ();
 FILLCELL_X1 FILLER_8_380 ();
 FILLCELL_X8 FILLER_8_384 ();
 FILLCELL_X4 FILLER_8_396 ();
 FILLCELL_X16 FILLER_8_402 ();
 FILLCELL_X1 FILLER_8_418 ();
 FILLCELL_X8 FILLER_8_429 ();
 FILLCELL_X1 FILLER_8_437 ();
 FILLCELL_X4 FILLER_8_441 ();
 FILLCELL_X4 FILLER_8_449 ();
 FILLCELL_X1 FILLER_8_453 ();
 FILLCELL_X4 FILLER_8_463 ();
 FILLCELL_X2 FILLER_8_467 ();
 FILLCELL_X1 FILLER_8_469 ();
 FILLCELL_X4 FILLER_8_480 ();
 FILLCELL_X1 FILLER_8_484 ();
 FILLCELL_X8 FILLER_8_487 ();
 FILLCELL_X2 FILLER_8_495 ();
 FILLCELL_X8 FILLER_8_501 ();
 FILLCELL_X2 FILLER_8_509 ();
 FILLCELL_X4 FILLER_8_515 ();
 FILLCELL_X4 FILLER_8_529 ();
 FILLCELL_X8 FILLER_8_540 ();
 FILLCELL_X1 FILLER_8_548 ();
 FILLCELL_X8 FILLER_8_559 ();
 FILLCELL_X4 FILLER_8_567 ();
 FILLCELL_X2 FILLER_8_571 ();
 FILLCELL_X4 FILLER_8_576 ();
 FILLCELL_X4 FILLER_8_583 ();
 FILLCELL_X16 FILLER_8_589 ();
 FILLCELL_X2 FILLER_8_605 ();
 FILLCELL_X4 FILLER_8_617 ();
 FILLCELL_X2 FILLER_8_621 ();
 FILLCELL_X1 FILLER_8_623 ();
 FILLCELL_X4 FILLER_8_627 ();
 FILLCELL_X4 FILLER_8_632 ();
 FILLCELL_X2 FILLER_8_636 ();
 FILLCELL_X8 FILLER_8_641 ();
 FILLCELL_X4 FILLER_8_653 ();
 FILLCELL_X4 FILLER_8_661 ();
 FILLCELL_X8 FILLER_8_674 ();
 FILLCELL_X2 FILLER_8_682 ();
 FILLCELL_X4 FILLER_8_693 ();
 FILLCELL_X8 FILLER_8_701 ();
 FILLCELL_X2 FILLER_8_709 ();
 FILLCELL_X4 FILLER_8_720 ();
 FILLCELL_X2 FILLER_8_724 ();
 FILLCELL_X8 FILLER_8_729 ();
 FILLCELL_X4 FILLER_8_747 ();
 FILLCELL_X4 FILLER_8_755 ();
 FILLCELL_X4 FILLER_8_761 ();
 FILLCELL_X4 FILLER_8_769 ();
 FILLCELL_X4 FILLER_8_776 ();
 FILLCELL_X2 FILLER_8_780 ();
 FILLCELL_X4 FILLER_8_786 ();
 FILLCELL_X2 FILLER_8_790 ();
 FILLCELL_X4 FILLER_8_799 ();
 FILLCELL_X4 FILLER_8_805 ();
 FILLCELL_X4 FILLER_8_812 ();
 FILLCELL_X4 FILLER_8_823 ();
 FILLCELL_X2 FILLER_8_827 ();
 FILLCELL_X1 FILLER_8_829 ();
 FILLCELL_X4 FILLER_8_839 ();
 FILLCELL_X2 FILLER_8_843 ();
 FILLCELL_X1 FILLER_8_845 ();
 FILLCELL_X4 FILLER_8_849 ();
 FILLCELL_X8 FILLER_8_860 ();
 FILLCELL_X4 FILLER_8_872 ();
 FILLCELL_X16 FILLER_8_878 ();
 FILLCELL_X4 FILLER_8_894 ();
 FILLCELL_X4 FILLER_8_907 ();
 FILLCELL_X4 FILLER_8_914 ();
 FILLCELL_X1 FILLER_8_918 ();
 FILLCELL_X4 FILLER_8_921 ();
 FILLCELL_X4 FILLER_8_932 ();
 FILLCELL_X1 FILLER_8_936 ();
 FILLCELL_X4 FILLER_8_946 ();
 FILLCELL_X1 FILLER_8_950 ();
 FILLCELL_X4 FILLER_8_954 ();
 FILLCELL_X4 FILLER_8_967 ();
 FILLCELL_X1 FILLER_8_971 ();
 FILLCELL_X4 FILLER_8_975 ();
 FILLCELL_X4 FILLER_8_983 ();
 FILLCELL_X4 FILLER_8_996 ();
 FILLCELL_X4 FILLER_8_1003 ();
 FILLCELL_X2 FILLER_8_1007 ();
 FILLCELL_X4 FILLER_8_1019 ();
 FILLCELL_X2 FILLER_8_1023 ();
 FILLCELL_X4 FILLER_8_1035 ();
 FILLCELL_X8 FILLER_8_1041 ();
 FILLCELL_X2 FILLER_8_1049 ();
 FILLCELL_X4 FILLER_8_1055 ();
 FILLCELL_X2 FILLER_8_1059 ();
 FILLCELL_X1 FILLER_8_1061 ();
 FILLCELL_X4 FILLER_8_1071 ();
 FILLCELL_X4 FILLER_8_1079 ();
 FILLCELL_X8 FILLER_8_1093 ();
 FILLCELL_X2 FILLER_8_1101 ();
 FILLCELL_X1 FILLER_8_1103 ();
 FILLCELL_X4 FILLER_8_1111 ();
 FILLCELL_X4 FILLER_8_1117 ();
 FILLCELL_X2 FILLER_8_1121 ();
 FILLCELL_X8 FILLER_8_1133 ();
 FILLCELL_X4 FILLER_8_1145 ();
 FILLCELL_X2 FILLER_8_1149 ();
 FILLCELL_X4 FILLER_8_1161 ();
 FILLCELL_X8 FILLER_8_1175 ();
 FILLCELL_X8 FILLER_8_1192 ();
 FILLCELL_X2 FILLER_8_1200 ();
 FILLCELL_X1 FILLER_8_1202 ();
 FILLCELL_X8 FILLER_8_1213 ();
 FILLCELL_X4 FILLER_8_1221 ();
 FILLCELL_X2 FILLER_8_1225 ();
 FILLCELL_X4 FILLER_8_1234 ();
 FILLCELL_X2 FILLER_8_1238 ();
 FILLCELL_X1 FILLER_8_1240 ();
 FILLCELL_X4 FILLER_8_1243 ();
 FILLCELL_X4 FILLER_8_1251 ();
 FILLCELL_X1 FILLER_8_1255 ();
 FILLCELL_X4 FILLER_8_1261 ();
 FILLCELL_X2 FILLER_8_1265 ();
 FILLCELL_X1 FILLER_8_1267 ();
 FILLCELL_X4 FILLER_8_1285 ();
 FILLCELL_X8 FILLER_8_1295 ();
 FILLCELL_X4 FILLER_8_1303 ();
 FILLCELL_X2 FILLER_8_1307 ();
 FILLCELL_X8 FILLER_8_1315 ();
 FILLCELL_X2 FILLER_8_1323 ();
 FILLCELL_X4 FILLER_8_1329 ();
 FILLCELL_X4 FILLER_8_1343 ();
 FILLCELL_X4 FILLER_8_1350 ();
 FILLCELL_X2 FILLER_8_1354 ();
 FILLCELL_X1 FILLER_8_1356 ();
 FILLCELL_X4 FILLER_8_1361 ();
 FILLCELL_X2 FILLER_8_1365 ();
 FILLCELL_X8 FILLER_8_1371 ();
 FILLCELL_X4 FILLER_8_1381 ();
 FILLCELL_X4 FILLER_8_1389 ();
 FILLCELL_X8 FILLER_8_1396 ();
 FILLCELL_X4 FILLER_8_1404 ();
 FILLCELL_X2 FILLER_8_1408 ();
 FILLCELL_X32 FILLER_8_1414 ();
 FILLCELL_X32 FILLER_8_1446 ();
 FILLCELL_X32 FILLER_8_1478 ();
 FILLCELL_X32 FILLER_8_1510 ();
 FILLCELL_X32 FILLER_8_1542 ();
 FILLCELL_X32 FILLER_8_1574 ();
 FILLCELL_X32 FILLER_8_1606 ();
 FILLCELL_X32 FILLER_8_1638 ();
 FILLCELL_X32 FILLER_8_1670 ();
 FILLCELL_X32 FILLER_8_1702 ();
 FILLCELL_X16 FILLER_8_1734 ();
 FILLCELL_X4 FILLER_8_1750 ();
 FILLCELL_X2 FILLER_8_1754 ();
 FILLCELL_X4 FILLER_9_1 ();
 FILLCELL_X4 FILLER_9_8 ();
 FILLCELL_X1 FILLER_9_12 ();
 FILLCELL_X8 FILLER_9_17 ();
 FILLCELL_X2 FILLER_9_25 ();
 FILLCELL_X4 FILLER_9_31 ();
 FILLCELL_X2 FILLER_9_35 ();
 FILLCELL_X4 FILLER_9_41 ();
 FILLCELL_X4 FILLER_9_49 ();
 FILLCELL_X4 FILLER_9_56 ();
 FILLCELL_X4 FILLER_9_64 ();
 FILLCELL_X8 FILLER_9_77 ();
 FILLCELL_X2 FILLER_9_85 ();
 FILLCELL_X4 FILLER_9_96 ();
 FILLCELL_X4 FILLER_9_103 ();
 FILLCELL_X2 FILLER_9_107 ();
 FILLCELL_X8 FILLER_9_116 ();
 FILLCELL_X2 FILLER_9_124 ();
 FILLCELL_X8 FILLER_9_129 ();
 FILLCELL_X2 FILLER_9_137 ();
 FILLCELL_X4 FILLER_9_142 ();
 FILLCELL_X4 FILLER_9_156 ();
 FILLCELL_X4 FILLER_9_170 ();
 FILLCELL_X8 FILLER_9_181 ();
 FILLCELL_X4 FILLER_9_189 ();
 FILLCELL_X2 FILLER_9_193 ();
 FILLCELL_X8 FILLER_9_197 ();
 FILLCELL_X1 FILLER_9_205 ();
 FILLCELL_X4 FILLER_9_210 ();
 FILLCELL_X8 FILLER_9_218 ();
 FILLCELL_X4 FILLER_9_226 ();
 FILLCELL_X1 FILLER_9_230 ();
 FILLCELL_X8 FILLER_9_234 ();
 FILLCELL_X4 FILLER_9_242 ();
 FILLCELL_X2 FILLER_9_246 ();
 FILLCELL_X1 FILLER_9_248 ();
 FILLCELL_X4 FILLER_9_253 ();
 FILLCELL_X4 FILLER_9_264 ();
 FILLCELL_X4 FILLER_9_278 ();
 FILLCELL_X2 FILLER_9_282 ();
 FILLCELL_X1 FILLER_9_284 ();
 FILLCELL_X4 FILLER_9_292 ();
 FILLCELL_X8 FILLER_9_302 ();
 FILLCELL_X2 FILLER_9_310 ();
 FILLCELL_X1 FILLER_9_312 ();
 FILLCELL_X4 FILLER_9_319 ();
 FILLCELL_X4 FILLER_9_325 ();
 FILLCELL_X2 FILLER_9_329 ();
 FILLCELL_X1 FILLER_9_331 ();
 FILLCELL_X4 FILLER_9_335 ();
 FILLCELL_X4 FILLER_9_348 ();
 FILLCELL_X4 FILLER_9_354 ();
 FILLCELL_X1 FILLER_9_358 ();
 FILLCELL_X4 FILLER_9_362 ();
 FILLCELL_X1 FILLER_9_366 ();
 FILLCELL_X8 FILLER_9_376 ();
 FILLCELL_X2 FILLER_9_384 ();
 FILLCELL_X4 FILLER_9_396 ();
 FILLCELL_X8 FILLER_9_410 ();
 FILLCELL_X4 FILLER_9_418 ();
 FILLCELL_X8 FILLER_9_432 ();
 FILLCELL_X2 FILLER_9_440 ();
 FILLCELL_X1 FILLER_9_442 ();
 FILLCELL_X4 FILLER_9_462 ();
 FILLCELL_X4 FILLER_9_469 ();
 FILLCELL_X4 FILLER_9_483 ();
 FILLCELL_X2 FILLER_9_487 ();
 FILLCELL_X4 FILLER_9_493 ();
 FILLCELL_X4 FILLER_9_506 ();
 FILLCELL_X4 FILLER_9_513 ();
 FILLCELL_X4 FILLER_9_520 ();
 FILLCELL_X4 FILLER_9_533 ();
 FILLCELL_X1 FILLER_9_537 ();
 FILLCELL_X4 FILLER_9_548 ();
 FILLCELL_X2 FILLER_9_552 ();
 FILLCELL_X4 FILLER_9_564 ();
 FILLCELL_X4 FILLER_9_577 ();
 FILLCELL_X8 FILLER_9_591 ();
 FILLCELL_X1 FILLER_9_599 ();
 FILLCELL_X8 FILLER_9_606 ();
 FILLCELL_X4 FILLER_9_614 ();
 FILLCELL_X1 FILLER_9_618 ();
 FILLCELL_X4 FILLER_9_622 ();
 FILLCELL_X4 FILLER_9_630 ();
 FILLCELL_X4 FILLER_9_643 ();
 FILLCELL_X4 FILLER_9_651 ();
 FILLCELL_X1 FILLER_9_655 ();
 FILLCELL_X8 FILLER_9_660 ();
 FILLCELL_X4 FILLER_9_668 ();
 FILLCELL_X2 FILLER_9_672 ();
 FILLCELL_X4 FILLER_9_676 ();
 FILLCELL_X4 FILLER_9_690 ();
 FILLCELL_X8 FILLER_9_704 ();
 FILLCELL_X2 FILLER_9_712 ();
 FILLCELL_X1 FILLER_9_714 ();
 FILLCELL_X4 FILLER_9_724 ();
 FILLCELL_X2 FILLER_9_728 ();
 FILLCELL_X4 FILLER_9_734 ();
 FILLCELL_X4 FILLER_9_748 ();
 FILLCELL_X2 FILLER_9_752 ();
 FILLCELL_X1 FILLER_9_754 ();
 FILLCELL_X4 FILLER_9_764 ();
 FILLCELL_X4 FILLER_9_777 ();
 FILLCELL_X2 FILLER_9_781 ();
 FILLCELL_X1 FILLER_9_783 ();
 FILLCELL_X4 FILLER_9_794 ();
 FILLCELL_X1 FILLER_9_798 ();
 FILLCELL_X8 FILLER_9_809 ();
 FILLCELL_X2 FILLER_9_817 ();
 FILLCELL_X4 FILLER_9_829 ();
 FILLCELL_X4 FILLER_9_836 ();
 FILLCELL_X4 FILLER_9_849 ();
 FILLCELL_X2 FILLER_9_853 ();
 FILLCELL_X4 FILLER_9_858 ();
 FILLCELL_X4 FILLER_9_866 ();
 FILLCELL_X8 FILLER_9_879 ();
 FILLCELL_X4 FILLER_9_887 ();
 FILLCELL_X2 FILLER_9_891 ();
 FILLCELL_X4 FILLER_9_896 ();
 FILLCELL_X2 FILLER_9_900 ();
 FILLCELL_X4 FILLER_9_904 ();
 FILLCELL_X2 FILLER_9_908 ();
 FILLCELL_X8 FILLER_9_913 ();
 FILLCELL_X4 FILLER_9_931 ();
 FILLCELL_X4 FILLER_9_938 ();
 FILLCELL_X4 FILLER_9_945 ();
 FILLCELL_X1 FILLER_9_949 ();
 FILLCELL_X4 FILLER_9_952 ();
 FILLCELL_X4 FILLER_9_959 ();
 FILLCELL_X16 FILLER_9_972 ();
 FILLCELL_X4 FILLER_9_995 ();
 FILLCELL_X1 FILLER_9_999 ();
 FILLCELL_X4 FILLER_9_1007 ();
 FILLCELL_X4 FILLER_9_1014 ();
 FILLCELL_X1 FILLER_9_1018 ();
 FILLCELL_X4 FILLER_9_1023 ();
 FILLCELL_X8 FILLER_9_1034 ();
 FILLCELL_X4 FILLER_9_1042 ();
 FILLCELL_X4 FILLER_9_1050 ();
 FILLCELL_X8 FILLER_9_1063 ();
 FILLCELL_X4 FILLER_9_1071 ();
 FILLCELL_X2 FILLER_9_1075 ();
 FILLCELL_X4 FILLER_9_1079 ();
 FILLCELL_X8 FILLER_9_1093 ();
 FILLCELL_X4 FILLER_9_1111 ();
 FILLCELL_X4 FILLER_9_1125 ();
 FILLCELL_X4 FILLER_9_1138 ();
 FILLCELL_X16 FILLER_9_1145 ();
 FILLCELL_X8 FILLER_9_1161 ();
 FILLCELL_X4 FILLER_9_1169 ();
 FILLCELL_X2 FILLER_9_1173 ();
 FILLCELL_X1 FILLER_9_1175 ();
 FILLCELL_X4 FILLER_9_1178 ();
 FILLCELL_X4 FILLER_9_1185 ();
 FILLCELL_X4 FILLER_9_1192 ();
 FILLCELL_X4 FILLER_9_1199 ();
 FILLCELL_X4 FILLER_9_1205 ();
 FILLCELL_X2 FILLER_9_1209 ();
 FILLCELL_X4 FILLER_9_1218 ();
 FILLCELL_X4 FILLER_9_1224 ();
 FILLCELL_X8 FILLER_9_1230 ();
 FILLCELL_X2 FILLER_9_1238 ();
 FILLCELL_X1 FILLER_9_1240 ();
 FILLCELL_X8 FILLER_9_1251 ();
 FILLCELL_X4 FILLER_9_1259 ();
 FILLCELL_X4 FILLER_9_1264 ();
 FILLCELL_X4 FILLER_9_1275 ();
 FILLCELL_X2 FILLER_9_1279 ();
 FILLCELL_X1 FILLER_9_1281 ();
 FILLCELL_X4 FILLER_9_1301 ();
 FILLCELL_X2 FILLER_9_1305 ();
 FILLCELL_X1 FILLER_9_1307 ();
 FILLCELL_X32 FILLER_9_1312 ();
 FILLCELL_X4 FILLER_9_1344 ();
 FILLCELL_X4 FILLER_9_1354 ();
 FILLCELL_X8 FILLER_9_1365 ();
 FILLCELL_X2 FILLER_9_1373 ();
 FILLCELL_X1 FILLER_9_1375 ();
 FILLCELL_X4 FILLER_9_1382 ();
 FILLCELL_X2 FILLER_9_1386 ();
 FILLCELL_X4 FILLER_9_1398 ();
 FILLCELL_X4 FILLER_9_1409 ();
 FILLCELL_X32 FILLER_9_1419 ();
 FILLCELL_X32 FILLER_9_1451 ();
 FILLCELL_X32 FILLER_9_1483 ();
 FILLCELL_X32 FILLER_9_1515 ();
 FILLCELL_X32 FILLER_9_1547 ();
 FILLCELL_X32 FILLER_9_1579 ();
 FILLCELL_X32 FILLER_9_1611 ();
 FILLCELL_X32 FILLER_9_1643 ();
 FILLCELL_X32 FILLER_9_1675 ();
 FILLCELL_X32 FILLER_9_1707 ();
 FILLCELL_X16 FILLER_9_1739 ();
 FILLCELL_X1 FILLER_9_1755 ();
 FILLCELL_X8 FILLER_10_1 ();
 FILLCELL_X1 FILLER_10_9 ();
 FILLCELL_X8 FILLER_10_19 ();
 FILLCELL_X8 FILLER_10_31 ();
 FILLCELL_X1 FILLER_10_39 ();
 FILLCELL_X8 FILLER_10_44 ();
 FILLCELL_X4 FILLER_10_55 ();
 FILLCELL_X16 FILLER_10_66 ();
 FILLCELL_X2 FILLER_10_82 ();
 FILLCELL_X4 FILLER_10_88 ();
 FILLCELL_X4 FILLER_10_95 ();
 FILLCELL_X4 FILLER_10_109 ();
 FILLCELL_X8 FILLER_10_123 ();
 FILLCELL_X8 FILLER_10_141 ();
 FILLCELL_X4 FILLER_10_149 ();
 FILLCELL_X1 FILLER_10_153 ();
 FILLCELL_X4 FILLER_10_163 ();
 FILLCELL_X4 FILLER_10_174 ();
 FILLCELL_X4 FILLER_10_181 ();
 FILLCELL_X4 FILLER_10_195 ();
 FILLCELL_X4 FILLER_10_205 ();
 FILLCELL_X1 FILLER_10_209 ();
 FILLCELL_X4 FILLER_10_216 ();
 FILLCELL_X4 FILLER_10_226 ();
 FILLCELL_X4 FILLER_10_234 ();
 FILLCELL_X4 FILLER_10_247 ();
 FILLCELL_X2 FILLER_10_251 ();
 FILLCELL_X4 FILLER_10_263 ();
 FILLCELL_X8 FILLER_10_269 ();
 FILLCELL_X4 FILLER_10_277 ();
 FILLCELL_X1 FILLER_10_281 ();
 FILLCELL_X4 FILLER_10_285 ();
 FILLCELL_X8 FILLER_10_293 ();
 FILLCELL_X2 FILLER_10_301 ();
 FILLCELL_X8 FILLER_10_307 ();
 FILLCELL_X2 FILLER_10_315 ();
 FILLCELL_X4 FILLER_10_321 ();
 FILLCELL_X4 FILLER_10_329 ();
 FILLCELL_X2 FILLER_10_333 ();
 FILLCELL_X8 FILLER_10_338 ();
 FILLCELL_X4 FILLER_10_346 ();
 FILLCELL_X8 FILLER_10_359 ();
 FILLCELL_X8 FILLER_10_374 ();
 FILLCELL_X1 FILLER_10_382 ();
 FILLCELL_X4 FILLER_10_386 ();
 FILLCELL_X8 FILLER_10_400 ();
 FILLCELL_X4 FILLER_10_408 ();
 FILLCELL_X1 FILLER_10_412 ();
 FILLCELL_X4 FILLER_10_420 ();
 FILLCELL_X4 FILLER_10_427 ();
 FILLCELL_X4 FILLER_10_433 ();
 FILLCELL_X2 FILLER_10_437 ();
 FILLCELL_X1 FILLER_10_439 ();
 FILLCELL_X16 FILLER_10_446 ();
 FILLCELL_X8 FILLER_10_462 ();
 FILLCELL_X2 FILLER_10_470 ();
 FILLCELL_X8 FILLER_10_479 ();
 FILLCELL_X4 FILLER_10_487 ();
 FILLCELL_X2 FILLER_10_491 ();
 FILLCELL_X4 FILLER_10_502 ();
 FILLCELL_X4 FILLER_10_510 ();
 FILLCELL_X2 FILLER_10_514 ();
 FILLCELL_X4 FILLER_10_519 ();
 FILLCELL_X8 FILLER_10_526 ();
 FILLCELL_X1 FILLER_10_534 ();
 FILLCELL_X4 FILLER_10_537 ();
 FILLCELL_X2 FILLER_10_541 ();
 FILLCELL_X1 FILLER_10_543 ();
 FILLCELL_X4 FILLER_10_546 ();
 FILLCELL_X8 FILLER_10_557 ();
 FILLCELL_X4 FILLER_10_565 ();
 FILLCELL_X16 FILLER_10_572 ();
 FILLCELL_X1 FILLER_10_588 ();
 FILLCELL_X8 FILLER_10_596 ();
 FILLCELL_X8 FILLER_10_608 ();
 FILLCELL_X4 FILLER_10_616 ();
 FILLCELL_X2 FILLER_10_620 ();
 FILLCELL_X1 FILLER_10_622 ();
 FILLCELL_X4 FILLER_10_627 ();
 FILLCELL_X8 FILLER_10_632 ();
 FILLCELL_X4 FILLER_10_640 ();
 FILLCELL_X1 FILLER_10_644 ();
 FILLCELL_X8 FILLER_10_654 ();
 FILLCELL_X16 FILLER_10_669 ();
 FILLCELL_X2 FILLER_10_685 ();
 FILLCELL_X4 FILLER_10_694 ();
 FILLCELL_X2 FILLER_10_698 ();
 FILLCELL_X4 FILLER_10_704 ();
 FILLCELL_X4 FILLER_10_713 ();
 FILLCELL_X1 FILLER_10_717 ();
 FILLCELL_X8 FILLER_10_728 ();
 FILLCELL_X1 FILLER_10_736 ();
 FILLCELL_X8 FILLER_10_744 ();
 FILLCELL_X2 FILLER_10_752 ();
 FILLCELL_X4 FILLER_10_757 ();
 FILLCELL_X4 FILLER_10_765 ();
 FILLCELL_X4 FILLER_10_772 ();
 FILLCELL_X2 FILLER_10_776 ();
 FILLCELL_X1 FILLER_10_778 ();
 FILLCELL_X8 FILLER_10_782 ();
 FILLCELL_X1 FILLER_10_790 ();
 FILLCELL_X4 FILLER_10_800 ();
 FILLCELL_X8 FILLER_10_807 ();
 FILLCELL_X4 FILLER_10_825 ();
 FILLCELL_X2 FILLER_10_829 ();
 FILLCELL_X8 FILLER_10_833 ();
 FILLCELL_X2 FILLER_10_841 ();
 FILLCELL_X4 FILLER_10_846 ();
 FILLCELL_X4 FILLER_10_859 ();
 FILLCELL_X4 FILLER_10_866 ();
 FILLCELL_X4 FILLER_10_874 ();
 FILLCELL_X4 FILLER_10_887 ();
 FILLCELL_X4 FILLER_10_900 ();
 FILLCELL_X8 FILLER_10_907 ();
 FILLCELL_X8 FILLER_10_924 ();
 FILLCELL_X4 FILLER_10_941 ();
 FILLCELL_X1 FILLER_10_945 ();
 FILLCELL_X4 FILLER_10_953 ();
 FILLCELL_X2 FILLER_10_957 ();
 FILLCELL_X1 FILLER_10_959 ();
 FILLCELL_X4 FILLER_10_963 ();
 FILLCELL_X2 FILLER_10_967 ();
 FILLCELL_X4 FILLER_10_972 ();
 FILLCELL_X8 FILLER_10_986 ();
 FILLCELL_X2 FILLER_10_994 ();
 FILLCELL_X1 FILLER_10_996 ();
 FILLCELL_X4 FILLER_10_1007 ();
 FILLCELL_X2 FILLER_10_1011 ();
 FILLCELL_X1 FILLER_10_1013 ();
 FILLCELL_X16 FILLER_10_1023 ();
 FILLCELL_X4 FILLER_10_1042 ();
 FILLCELL_X4 FILLER_10_1049 ();
 FILLCELL_X2 FILLER_10_1053 ();
 FILLCELL_X4 FILLER_10_1059 ();
 FILLCELL_X4 FILLER_10_1070 ();
 FILLCELL_X4 FILLER_10_1076 ();
 FILLCELL_X2 FILLER_10_1080 ();
 FILLCELL_X4 FILLER_10_1089 ();
 FILLCELL_X2 FILLER_10_1093 ();
 FILLCELL_X4 FILLER_10_1099 ();
 FILLCELL_X8 FILLER_10_1106 ();
 FILLCELL_X2 FILLER_10_1114 ();
 FILLCELL_X4 FILLER_10_1119 ();
 FILLCELL_X8 FILLER_10_1126 ();
 FILLCELL_X2 FILLER_10_1134 ();
 FILLCELL_X4 FILLER_10_1145 ();
 FILLCELL_X4 FILLER_10_1168 ();
 FILLCELL_X8 FILLER_10_1181 ();
 FILLCELL_X1 FILLER_10_1189 ();
 FILLCELL_X4 FILLER_10_1199 ();
 FILLCELL_X1 FILLER_10_1203 ();
 FILLCELL_X4 FILLER_10_1206 ();
 FILLCELL_X4 FILLER_10_1217 ();
 FILLCELL_X2 FILLER_10_1221 ();
 FILLCELL_X16 FILLER_10_1233 ();
 FILLCELL_X8 FILLER_10_1249 ();
 FILLCELL_X4 FILLER_10_1257 ();
 FILLCELL_X1 FILLER_10_1261 ();
 FILLCELL_X8 FILLER_10_1266 ();
 FILLCELL_X1 FILLER_10_1274 ();
 FILLCELL_X4 FILLER_10_1280 ();
 FILLCELL_X2 FILLER_10_1284 ();
 FILLCELL_X1 FILLER_10_1286 ();
 FILLCELL_X8 FILLER_10_1291 ();
 FILLCELL_X4 FILLER_10_1299 ();
 FILLCELL_X2 FILLER_10_1303 ();
 FILLCELL_X4 FILLER_10_1324 ();
 FILLCELL_X4 FILLER_10_1337 ();
 FILLCELL_X8 FILLER_10_1351 ();
 FILLCELL_X4 FILLER_10_1359 ();
 FILLCELL_X2 FILLER_10_1363 ();
 FILLCELL_X1 FILLER_10_1365 ();
 FILLCELL_X8 FILLER_10_1376 ();
 FILLCELL_X4 FILLER_10_1384 ();
 FILLCELL_X8 FILLER_10_1397 ();
 FILLCELL_X32 FILLER_10_1411 ();
 FILLCELL_X32 FILLER_10_1443 ();
 FILLCELL_X32 FILLER_10_1475 ();
 FILLCELL_X32 FILLER_10_1507 ();
 FILLCELL_X32 FILLER_10_1539 ();
 FILLCELL_X32 FILLER_10_1571 ();
 FILLCELL_X32 FILLER_10_1603 ();
 FILLCELL_X32 FILLER_10_1635 ();
 FILLCELL_X32 FILLER_10_1667 ();
 FILLCELL_X32 FILLER_10_1699 ();
 FILLCELL_X16 FILLER_10_1731 ();
 FILLCELL_X2 FILLER_10_1747 ();
 FILLCELL_X4 FILLER_10_1752 ();
 FILLCELL_X4 FILLER_11_1 ();
 FILLCELL_X1 FILLER_11_5 ();
 FILLCELL_X4 FILLER_11_10 ();
 FILLCELL_X4 FILLER_11_23 ();
 FILLCELL_X2 FILLER_11_27 ();
 FILLCELL_X4 FILLER_11_39 ();
 FILLCELL_X1 FILLER_11_43 ();
 FILLCELL_X4 FILLER_11_54 ();
 FILLCELL_X8 FILLER_11_60 ();
 FILLCELL_X4 FILLER_11_78 ();
 FILLCELL_X2 FILLER_11_82 ();
 FILLCELL_X4 FILLER_11_93 ();
 FILLCELL_X8 FILLER_11_100 ();
 FILLCELL_X4 FILLER_11_108 ();
 FILLCELL_X8 FILLER_11_114 ();
 FILLCELL_X4 FILLER_11_122 ();
 FILLCELL_X4 FILLER_11_135 ();
 FILLCELL_X4 FILLER_11_146 ();
 FILLCELL_X4 FILLER_11_153 ();
 FILLCELL_X2 FILLER_11_157 ();
 FILLCELL_X1 FILLER_11_159 ();
 FILLCELL_X8 FILLER_11_167 ();
 FILLCELL_X4 FILLER_11_175 ();
 FILLCELL_X1 FILLER_11_179 ();
 FILLCELL_X4 FILLER_11_190 ();
 FILLCELL_X8 FILLER_11_201 ();
 FILLCELL_X2 FILLER_11_209 ();
 FILLCELL_X1 FILLER_11_211 ();
 FILLCELL_X8 FILLER_11_219 ();
 FILLCELL_X2 FILLER_11_227 ();
 FILLCELL_X4 FILLER_11_232 ();
 FILLCELL_X8 FILLER_11_245 ();
 FILLCELL_X1 FILLER_11_253 ();
 FILLCELL_X8 FILLER_11_257 ();
 FILLCELL_X4 FILLER_11_272 ();
 FILLCELL_X8 FILLER_11_278 ();
 FILLCELL_X8 FILLER_11_290 ();
 FILLCELL_X2 FILLER_11_298 ();
 FILLCELL_X8 FILLER_11_304 ();
 FILLCELL_X4 FILLER_11_312 ();
 FILLCELL_X2 FILLER_11_316 ();
 FILLCELL_X4 FILLER_11_325 ();
 FILLCELL_X4 FILLER_11_335 ();
 FILLCELL_X2 FILLER_11_339 ();
 FILLCELL_X1 FILLER_11_341 ();
 FILLCELL_X4 FILLER_11_345 ();
 FILLCELL_X4 FILLER_11_359 ();
 FILLCELL_X2 FILLER_11_363 ();
 FILLCELL_X1 FILLER_11_365 ();
 FILLCELL_X4 FILLER_11_376 ();
 FILLCELL_X8 FILLER_11_383 ();
 FILLCELL_X1 FILLER_11_391 ();
 FILLCELL_X4 FILLER_11_396 ();
 FILLCELL_X1 FILLER_11_400 ();
 FILLCELL_X8 FILLER_11_403 ();
 FILLCELL_X2 FILLER_11_411 ();
 FILLCELL_X4 FILLER_11_416 ();
 FILLCELL_X4 FILLER_11_423 ();
 FILLCELL_X4 FILLER_11_436 ();
 FILLCELL_X1 FILLER_11_440 ();
 FILLCELL_X4 FILLER_11_444 ();
 FILLCELL_X8 FILLER_11_454 ();
 FILLCELL_X2 FILLER_11_462 ();
 FILLCELL_X1 FILLER_11_464 ();
 FILLCELL_X8 FILLER_11_468 ();
 FILLCELL_X1 FILLER_11_476 ();
 FILLCELL_X8 FILLER_11_481 ();
 FILLCELL_X1 FILLER_11_489 ();
 FILLCELL_X4 FILLER_11_492 ();
 FILLCELL_X8 FILLER_11_506 ();
 FILLCELL_X4 FILLER_11_517 ();
 FILLCELL_X8 FILLER_11_530 ();
 FILLCELL_X4 FILLER_11_541 ();
 FILLCELL_X4 FILLER_11_548 ();
 FILLCELL_X1 FILLER_11_552 ();
 FILLCELL_X8 FILLER_11_562 ();
 FILLCELL_X2 FILLER_11_570 ();
 FILLCELL_X4 FILLER_11_575 ();
 FILLCELL_X4 FILLER_11_582 ();
 FILLCELL_X8 FILLER_11_596 ();
 FILLCELL_X8 FILLER_11_623 ();
 FILLCELL_X16 FILLER_11_634 ();
 FILLCELL_X2 FILLER_11_650 ();
 FILLCELL_X4 FILLER_11_655 ();
 FILLCELL_X4 FILLER_11_669 ();
 FILLCELL_X4 FILLER_11_683 ();
 FILLCELL_X2 FILLER_11_687 ();
 FILLCELL_X4 FILLER_11_692 ();
 FILLCELL_X4 FILLER_11_700 ();
 FILLCELL_X4 FILLER_11_710 ();
 FILLCELL_X4 FILLER_11_717 ();
 FILLCELL_X4 FILLER_11_731 ();
 FILLCELL_X8 FILLER_11_739 ();
 FILLCELL_X4 FILLER_11_750 ();
 FILLCELL_X8 FILLER_11_757 ();
 FILLCELL_X1 FILLER_11_765 ();
 FILLCELL_X4 FILLER_11_769 ();
 FILLCELL_X2 FILLER_11_773 ();
 FILLCELL_X1 FILLER_11_775 ();
 FILLCELL_X8 FILLER_11_778 ();
 FILLCELL_X4 FILLER_11_786 ();
 FILLCELL_X8 FILLER_11_793 ();
 FILLCELL_X4 FILLER_11_801 ();
 FILLCELL_X16 FILLER_11_808 ();
 FILLCELL_X8 FILLER_11_824 ();
 FILLCELL_X2 FILLER_11_832 ();
 FILLCELL_X1 FILLER_11_834 ();
 FILLCELL_X8 FILLER_11_838 ();
 FILLCELL_X4 FILLER_11_848 ();
 FILLCELL_X4 FILLER_11_855 ();
 FILLCELL_X4 FILLER_11_862 ();
 FILLCELL_X16 FILLER_11_869 ();
 FILLCELL_X8 FILLER_11_885 ();
 FILLCELL_X1 FILLER_11_893 ();
 FILLCELL_X4 FILLER_11_901 ();
 FILLCELL_X1 FILLER_11_905 ();
 FILLCELL_X4 FILLER_11_916 ();
 FILLCELL_X8 FILLER_11_923 ();
 FILLCELL_X1 FILLER_11_931 ();
 FILLCELL_X8 FILLER_11_935 ();
 FILLCELL_X4 FILLER_11_953 ();
 FILLCELL_X16 FILLER_11_967 ();
 FILLCELL_X2 FILLER_11_983 ();
 FILLCELL_X4 FILLER_11_988 ();
 FILLCELL_X1 FILLER_11_992 ();
 FILLCELL_X8 FILLER_11_995 ();
 FILLCELL_X4 FILLER_11_1006 ();
 FILLCELL_X4 FILLER_11_1013 ();
 FILLCELL_X4 FILLER_11_1020 ();
 FILLCELL_X4 FILLER_11_1027 ();
 FILLCELL_X8 FILLER_11_1041 ();
 FILLCELL_X2 FILLER_11_1049 ();
 FILLCELL_X8 FILLER_11_1061 ();
 FILLCELL_X2 FILLER_11_1069 ();
 FILLCELL_X1 FILLER_11_1071 ();
 FILLCELL_X4 FILLER_11_1082 ();
 FILLCELL_X16 FILLER_11_1089 ();
 FILLCELL_X8 FILLER_11_1105 ();
 FILLCELL_X4 FILLER_11_1117 ();
 FILLCELL_X4 FILLER_11_1125 ();
 FILLCELL_X4 FILLER_11_1133 ();
 FILLCELL_X2 FILLER_11_1137 ();
 FILLCELL_X4 FILLER_11_1148 ();
 FILLCELL_X8 FILLER_11_1156 ();
 FILLCELL_X4 FILLER_11_1164 ();
 FILLCELL_X1 FILLER_11_1168 ();
 FILLCELL_X8 FILLER_11_1172 ();
 FILLCELL_X2 FILLER_11_1180 ();
 FILLCELL_X4 FILLER_11_1191 ();
 FILLCELL_X4 FILLER_11_1205 ();
 FILLCELL_X1 FILLER_11_1209 ();
 FILLCELL_X4 FILLER_11_1213 ();
 FILLCELL_X2 FILLER_11_1217 ();
 FILLCELL_X8 FILLER_11_1229 ();
 FILLCELL_X4 FILLER_11_1246 ();
 FILLCELL_X8 FILLER_11_1253 ();
 FILLCELL_X2 FILLER_11_1261 ();
 FILLCELL_X4 FILLER_11_1264 ();
 FILLCELL_X4 FILLER_11_1272 ();
 FILLCELL_X8 FILLER_11_1279 ();
 FILLCELL_X1 FILLER_11_1287 ();
 FILLCELL_X4 FILLER_11_1295 ();
 FILLCELL_X8 FILLER_11_1303 ();
 FILLCELL_X1 FILLER_11_1311 ();
 FILLCELL_X4 FILLER_11_1321 ();
 FILLCELL_X2 FILLER_11_1325 ();
 FILLCELL_X1 FILLER_11_1327 ();
 FILLCELL_X4 FILLER_11_1332 ();
 FILLCELL_X4 FILLER_11_1339 ();
 FILLCELL_X2 FILLER_11_1343 ();
 FILLCELL_X1 FILLER_11_1345 ();
 FILLCELL_X4 FILLER_11_1349 ();
 FILLCELL_X4 FILLER_11_1356 ();
 FILLCELL_X2 FILLER_11_1360 ();
 FILLCELL_X1 FILLER_11_1362 ();
 FILLCELL_X4 FILLER_11_1365 ();
 FILLCELL_X4 FILLER_11_1376 ();
 FILLCELL_X2 FILLER_11_1380 ();
 FILLCELL_X4 FILLER_11_1385 ();
 FILLCELL_X1 FILLER_11_1389 ();
 FILLCELL_X4 FILLER_11_1393 ();
 FILLCELL_X2 FILLER_11_1397 ();
 FILLCELL_X4 FILLER_11_1402 ();
 FILLCELL_X4 FILLER_11_1413 ();
 FILLCELL_X32 FILLER_11_1420 ();
 FILLCELL_X32 FILLER_11_1452 ();
 FILLCELL_X32 FILLER_11_1484 ();
 FILLCELL_X32 FILLER_11_1516 ();
 FILLCELL_X32 FILLER_11_1548 ();
 FILLCELL_X32 FILLER_11_1580 ();
 FILLCELL_X32 FILLER_11_1612 ();
 FILLCELL_X32 FILLER_11_1644 ();
 FILLCELL_X32 FILLER_11_1676 ();
 FILLCELL_X32 FILLER_11_1708 ();
 FILLCELL_X16 FILLER_11_1740 ();
 FILLCELL_X8 FILLER_12_1 ();
 FILLCELL_X2 FILLER_12_9 ();
 FILLCELL_X16 FILLER_12_14 ();
 FILLCELL_X1 FILLER_12_30 ();
 FILLCELL_X8 FILLER_12_34 ();
 FILLCELL_X4 FILLER_12_45 ();
 FILLCELL_X4 FILLER_12_59 ();
 FILLCELL_X2 FILLER_12_63 ();
 FILLCELL_X1 FILLER_12_65 ();
 FILLCELL_X8 FILLER_12_68 ();
 FILLCELL_X4 FILLER_12_76 ();
 FILLCELL_X2 FILLER_12_80 ();
 FILLCELL_X4 FILLER_12_86 ();
 FILLCELL_X1 FILLER_12_90 ();
 FILLCELL_X4 FILLER_12_94 ();
 FILLCELL_X2 FILLER_12_98 ();
 FILLCELL_X8 FILLER_12_109 ();
 FILLCELL_X4 FILLER_12_117 ();
 FILLCELL_X2 FILLER_12_121 ();
 FILLCELL_X4 FILLER_12_126 ();
 FILLCELL_X4 FILLER_12_134 ();
 FILLCELL_X8 FILLER_12_141 ();
 FILLCELL_X2 FILLER_12_149 ();
 FILLCELL_X4 FILLER_12_153 ();
 FILLCELL_X1 FILLER_12_157 ();
 FILLCELL_X4 FILLER_12_168 ();
 FILLCELL_X8 FILLER_12_174 ();
 FILLCELL_X16 FILLER_12_191 ();
 FILLCELL_X2 FILLER_12_207 ();
 FILLCELL_X1 FILLER_12_209 ();
 FILLCELL_X16 FILLER_12_213 ();
 FILLCELL_X4 FILLER_12_229 ();
 FILLCELL_X2 FILLER_12_233 ();
 FILLCELL_X16 FILLER_12_238 ();
 FILLCELL_X4 FILLER_12_254 ();
 FILLCELL_X4 FILLER_12_268 ();
 FILLCELL_X8 FILLER_12_282 ();
 FILLCELL_X2 FILLER_12_290 ();
 FILLCELL_X4 FILLER_12_301 ();
 FILLCELL_X1 FILLER_12_305 ();
 FILLCELL_X8 FILLER_12_315 ();
 FILLCELL_X2 FILLER_12_323 ();
 FILLCELL_X1 FILLER_12_325 ();
 FILLCELL_X8 FILLER_12_332 ();
 FILLCELL_X2 FILLER_12_340 ();
 FILLCELL_X1 FILLER_12_342 ();
 FILLCELL_X4 FILLER_12_350 ();
 FILLCELL_X8 FILLER_12_356 ();
 FILLCELL_X2 FILLER_12_364 ();
 FILLCELL_X8 FILLER_12_370 ();
 FILLCELL_X8 FILLER_12_380 ();
 FILLCELL_X4 FILLER_12_398 ();
 FILLCELL_X4 FILLER_12_405 ();
 FILLCELL_X2 FILLER_12_409 ();
 FILLCELL_X8 FILLER_12_421 ();
 FILLCELL_X2 FILLER_12_429 ();
 FILLCELL_X4 FILLER_12_434 ();
 FILLCELL_X4 FILLER_12_445 ();
 FILLCELL_X4 FILLER_12_458 ();
 FILLCELL_X4 FILLER_12_472 ();
 FILLCELL_X4 FILLER_12_486 ();
 FILLCELL_X4 FILLER_12_492 ();
 FILLCELL_X2 FILLER_12_496 ();
 FILLCELL_X1 FILLER_12_498 ();
 FILLCELL_X8 FILLER_12_509 ();
 FILLCELL_X2 FILLER_12_517 ();
 FILLCELL_X4 FILLER_12_529 ();
 FILLCELL_X4 FILLER_12_543 ();
 FILLCELL_X2 FILLER_12_547 ();
 FILLCELL_X1 FILLER_12_549 ();
 FILLCELL_X4 FILLER_12_553 ();
 FILLCELL_X2 FILLER_12_557 ();
 FILLCELL_X1 FILLER_12_559 ();
 FILLCELL_X8 FILLER_12_569 ();
 FILLCELL_X4 FILLER_12_577 ();
 FILLCELL_X1 FILLER_12_581 ();
 FILLCELL_X16 FILLER_12_591 ();
 FILLCELL_X1 FILLER_12_607 ();
 FILLCELL_X4 FILLER_12_612 ();
 FILLCELL_X4 FILLER_12_625 ();
 FILLCELL_X2 FILLER_12_629 ();
 FILLCELL_X8 FILLER_12_632 ();
 FILLCELL_X4 FILLER_12_640 ();
 FILLCELL_X4 FILLER_12_647 ();
 FILLCELL_X4 FILLER_12_660 ();
 FILLCELL_X2 FILLER_12_664 ();
 FILLCELL_X1 FILLER_12_666 ();
 FILLCELL_X4 FILLER_12_669 ();
 FILLCELL_X4 FILLER_12_676 ();
 FILLCELL_X4 FILLER_12_689 ();
 FILLCELL_X1 FILLER_12_693 ();
 FILLCELL_X4 FILLER_12_698 ();
 FILLCELL_X1 FILLER_12_702 ();
 FILLCELL_X8 FILLER_12_716 ();
 FILLCELL_X4 FILLER_12_724 ();
 FILLCELL_X2 FILLER_12_728 ();
 FILLCELL_X1 FILLER_12_730 ();
 FILLCELL_X4 FILLER_12_741 ();
 FILLCELL_X4 FILLER_12_755 ();
 FILLCELL_X4 FILLER_12_766 ();
 FILLCELL_X1 FILLER_12_770 ();
 FILLCELL_X4 FILLER_12_781 ();
 FILLCELL_X4 FILLER_12_794 ();
 FILLCELL_X4 FILLER_12_803 ();
 FILLCELL_X2 FILLER_12_807 ();
 FILLCELL_X1 FILLER_12_809 ();
 FILLCELL_X4 FILLER_12_819 ();
 FILLCELL_X2 FILLER_12_823 ();
 FILLCELL_X4 FILLER_12_829 ();
 FILLCELL_X4 FILLER_12_843 ();
 FILLCELL_X8 FILLER_12_854 ();
 FILLCELL_X2 FILLER_12_862 ();
 FILLCELL_X4 FILLER_12_873 ();
 FILLCELL_X4 FILLER_12_880 ();
 FILLCELL_X16 FILLER_12_894 ();
 FILLCELL_X4 FILLER_12_913 ();
 FILLCELL_X4 FILLER_12_926 ();
 FILLCELL_X8 FILLER_12_933 ();
 FILLCELL_X4 FILLER_12_945 ();
 FILLCELL_X8 FILLER_12_952 ();
 FILLCELL_X4 FILLER_12_960 ();
 FILLCELL_X2 FILLER_12_964 ();
 FILLCELL_X4 FILLER_12_976 ();
 FILLCELL_X1 FILLER_12_980 ();
 FILLCELL_X4 FILLER_12_990 ();
 FILLCELL_X8 FILLER_12_1003 ();
 FILLCELL_X1 FILLER_12_1011 ();
 FILLCELL_X8 FILLER_12_1021 ();
 FILLCELL_X2 FILLER_12_1029 ();
 FILLCELL_X1 FILLER_12_1031 ();
 FILLCELL_X4 FILLER_12_1042 ();
 FILLCELL_X16 FILLER_12_1048 ();
 FILLCELL_X8 FILLER_12_1064 ();
 FILLCELL_X2 FILLER_12_1072 ();
 FILLCELL_X4 FILLER_12_1077 ();
 FILLCELL_X4 FILLER_12_1090 ();
 FILLCELL_X4 FILLER_12_1113 ();
 FILLCELL_X4 FILLER_12_1121 ();
 FILLCELL_X2 FILLER_12_1125 ();
 FILLCELL_X1 FILLER_12_1127 ();
 FILLCELL_X4 FILLER_12_1137 ();
 FILLCELL_X4 FILLER_12_1144 ();
 FILLCELL_X8 FILLER_12_1151 ();
 FILLCELL_X4 FILLER_12_1159 ();
 FILLCELL_X2 FILLER_12_1163 ();
 FILLCELL_X1 FILLER_12_1165 ();
 FILLCELL_X4 FILLER_12_1173 ();
 FILLCELL_X4 FILLER_12_1180 ();
 FILLCELL_X1 FILLER_12_1184 ();
 FILLCELL_X8 FILLER_12_1187 ();
 FILLCELL_X1 FILLER_12_1195 ();
 FILLCELL_X4 FILLER_12_1201 ();
 FILLCELL_X4 FILLER_12_1208 ();
 FILLCELL_X2 FILLER_12_1212 ();
 FILLCELL_X1 FILLER_12_1214 ();
 FILLCELL_X8 FILLER_12_1224 ();
 FILLCELL_X4 FILLER_12_1235 ();
 FILLCELL_X2 FILLER_12_1239 ();
 FILLCELL_X4 FILLER_12_1244 ();
 FILLCELL_X2 FILLER_12_1248 ();
 FILLCELL_X4 FILLER_12_1259 ();
 FILLCELL_X1 FILLER_12_1263 ();
 FILLCELL_X4 FILLER_12_1269 ();
 FILLCELL_X1 FILLER_12_1273 ();
 FILLCELL_X4 FILLER_12_1283 ();
 FILLCELL_X2 FILLER_12_1287 ();
 FILLCELL_X4 FILLER_12_1299 ();
 FILLCELL_X16 FILLER_12_1307 ();
 FILLCELL_X8 FILLER_12_1326 ();
 FILLCELL_X4 FILLER_12_1334 ();
 FILLCELL_X2 FILLER_12_1338 ();
 FILLCELL_X1 FILLER_12_1340 ();
 FILLCELL_X8 FILLER_12_1345 ();
 FILLCELL_X1 FILLER_12_1353 ();
 FILLCELL_X4 FILLER_12_1358 ();
 FILLCELL_X8 FILLER_12_1372 ();
 FILLCELL_X1 FILLER_12_1380 ();
 FILLCELL_X4 FILLER_12_1390 ();
 FILLCELL_X32 FILLER_12_1397 ();
 FILLCELL_X32 FILLER_12_1429 ();
 FILLCELL_X32 FILLER_12_1461 ();
 FILLCELL_X32 FILLER_12_1493 ();
 FILLCELL_X32 FILLER_12_1525 ();
 FILLCELL_X32 FILLER_12_1557 ();
 FILLCELL_X32 FILLER_12_1589 ();
 FILLCELL_X32 FILLER_12_1621 ();
 FILLCELL_X32 FILLER_12_1653 ();
 FILLCELL_X32 FILLER_12_1685 ();
 FILLCELL_X32 FILLER_12_1717 ();
 FILLCELL_X4 FILLER_12_1749 ();
 FILLCELL_X2 FILLER_12_1753 ();
 FILLCELL_X1 FILLER_12_1755 ();
 FILLCELL_X8 FILLER_13_1 ();
 FILLCELL_X2 FILLER_13_9 ();
 FILLCELL_X4 FILLER_13_14 ();
 FILLCELL_X4 FILLER_13_25 ();
 FILLCELL_X8 FILLER_13_31 ();
 FILLCELL_X4 FILLER_13_39 ();
 FILLCELL_X2 FILLER_13_43 ();
 FILLCELL_X8 FILLER_13_49 ();
 FILLCELL_X1 FILLER_13_57 ();
 FILLCELL_X4 FILLER_13_61 ();
 FILLCELL_X2 FILLER_13_65 ();
 FILLCELL_X1 FILLER_13_67 ();
 FILLCELL_X4 FILLER_13_71 ();
 FILLCELL_X8 FILLER_13_78 ();
 FILLCELL_X4 FILLER_13_86 ();
 FILLCELL_X4 FILLER_13_93 ();
 FILLCELL_X4 FILLER_13_101 ();
 FILLCELL_X4 FILLER_13_109 ();
 FILLCELL_X16 FILLER_13_123 ();
 FILLCELL_X8 FILLER_13_139 ();
 FILLCELL_X1 FILLER_13_147 ();
 FILLCELL_X4 FILLER_13_151 ();
 FILLCELL_X4 FILLER_13_165 ();
 FILLCELL_X2 FILLER_13_169 ();
 FILLCELL_X4 FILLER_13_174 ();
 FILLCELL_X4 FILLER_13_181 ();
 FILLCELL_X4 FILLER_13_191 ();
 FILLCELL_X1 FILLER_13_195 ();
 FILLCELL_X4 FILLER_13_199 ();
 FILLCELL_X8 FILLER_13_207 ();
 FILLCELL_X16 FILLER_13_219 ();
 FILLCELL_X4 FILLER_13_235 ();
 FILLCELL_X1 FILLER_13_239 ();
 FILLCELL_X4 FILLER_13_247 ();
 FILLCELL_X8 FILLER_13_253 ();
 FILLCELL_X4 FILLER_13_264 ();
 FILLCELL_X4 FILLER_13_271 ();
 FILLCELL_X4 FILLER_13_278 ();
 FILLCELL_X1 FILLER_13_282 ();
 FILLCELL_X4 FILLER_13_286 ();
 FILLCELL_X4 FILLER_13_293 ();
 FILLCELL_X32 FILLER_13_300 ();
 FILLCELL_X8 FILLER_13_332 ();
 FILLCELL_X2 FILLER_13_340 ();
 FILLCELL_X4 FILLER_13_345 ();
 FILLCELL_X8 FILLER_13_358 ();
 FILLCELL_X4 FILLER_13_373 ();
 FILLCELL_X4 FILLER_13_381 ();
 FILLCELL_X1 FILLER_13_385 ();
 FILLCELL_X4 FILLER_13_390 ();
 FILLCELL_X8 FILLER_13_404 ();
 FILLCELL_X2 FILLER_13_412 ();
 FILLCELL_X4 FILLER_13_424 ();
 FILLCELL_X4 FILLER_13_435 ();
 FILLCELL_X4 FILLER_13_442 ();
 FILLCELL_X2 FILLER_13_446 ();
 FILLCELL_X16 FILLER_13_458 ();
 FILLCELL_X2 FILLER_13_474 ();
 FILLCELL_X1 FILLER_13_476 ();
 FILLCELL_X8 FILLER_13_480 ();
 FILLCELL_X8 FILLER_13_495 ();
 FILLCELL_X2 FILLER_13_503 ();
 FILLCELL_X1 FILLER_13_505 ();
 FILLCELL_X8 FILLER_13_509 ();
 FILLCELL_X2 FILLER_13_517 ();
 FILLCELL_X1 FILLER_13_519 ();
 FILLCELL_X4 FILLER_13_527 ();
 FILLCELL_X4 FILLER_13_533 ();
 FILLCELL_X1 FILLER_13_537 ();
 FILLCELL_X4 FILLER_13_541 ();
 FILLCELL_X4 FILLER_13_554 ();
 FILLCELL_X2 FILLER_13_558 ();
 FILLCELL_X4 FILLER_13_569 ();
 FILLCELL_X8 FILLER_13_582 ();
 FILLCELL_X2 FILLER_13_590 ();
 FILLCELL_X1 FILLER_13_592 ();
 FILLCELL_X4 FILLER_13_597 ();
 FILLCELL_X4 FILLER_13_610 ();
 FILLCELL_X1 FILLER_13_614 ();
 FILLCELL_X4 FILLER_13_618 ();
 FILLCELL_X4 FILLER_13_632 ();
 FILLCELL_X4 FILLER_13_643 ();
 FILLCELL_X4 FILLER_13_649 ();
 FILLCELL_X4 FILLER_13_656 ();
 FILLCELL_X8 FILLER_13_663 ();
 FILLCELL_X4 FILLER_13_671 ();
 FILLCELL_X4 FILLER_13_678 ();
 FILLCELL_X8 FILLER_13_692 ();
 FILLCELL_X1 FILLER_13_700 ();
 FILLCELL_X8 FILLER_13_705 ();
 FILLCELL_X4 FILLER_13_713 ();
 FILLCELL_X2 FILLER_13_717 ();
 FILLCELL_X4 FILLER_13_722 ();
 FILLCELL_X4 FILLER_13_733 ();
 FILLCELL_X8 FILLER_13_739 ();
 FILLCELL_X1 FILLER_13_747 ();
 FILLCELL_X4 FILLER_13_750 ();
 FILLCELL_X8 FILLER_13_764 ();
 FILLCELL_X4 FILLER_13_772 ();
 FILLCELL_X1 FILLER_13_776 ();
 FILLCELL_X4 FILLER_13_787 ();
 FILLCELL_X2 FILLER_13_791 ();
 FILLCELL_X4 FILLER_13_795 ();
 FILLCELL_X4 FILLER_13_802 ();
 FILLCELL_X4 FILLER_13_816 ();
 FILLCELL_X4 FILLER_13_829 ();
 FILLCELL_X8 FILLER_13_843 ();
 FILLCELL_X4 FILLER_13_851 ();
 FILLCELL_X16 FILLER_13_865 ();
 FILLCELL_X4 FILLER_13_881 ();
 FILLCELL_X1 FILLER_13_885 ();
 FILLCELL_X4 FILLER_13_893 ();
 FILLCELL_X4 FILLER_13_899 ();
 FILLCELL_X1 FILLER_13_903 ();
 FILLCELL_X8 FILLER_13_907 ();
 FILLCELL_X4 FILLER_13_915 ();
 FILLCELL_X8 FILLER_13_928 ();
 FILLCELL_X1 FILLER_13_936 ();
 FILLCELL_X4 FILLER_13_941 ();
 FILLCELL_X4 FILLER_13_947 ();
 FILLCELL_X2 FILLER_13_951 ();
 FILLCELL_X1 FILLER_13_953 ();
 FILLCELL_X4 FILLER_13_961 ();
 FILLCELL_X4 FILLER_13_975 ();
 FILLCELL_X4 FILLER_13_981 ();
 FILLCELL_X8 FILLER_13_988 ();
 FILLCELL_X4 FILLER_13_996 ();
 FILLCELL_X2 FILLER_13_1000 ();
 FILLCELL_X4 FILLER_13_1005 ();
 FILLCELL_X8 FILLER_13_1018 ();
 FILLCELL_X4 FILLER_13_1026 ();
 FILLCELL_X2 FILLER_13_1030 ();
 FILLCELL_X4 FILLER_13_1039 ();
 FILLCELL_X16 FILLER_13_1047 ();
 FILLCELL_X1 FILLER_13_1063 ();
 FILLCELL_X4 FILLER_13_1067 ();
 FILLCELL_X4 FILLER_13_1074 ();
 FILLCELL_X2 FILLER_13_1078 ();
 FILLCELL_X4 FILLER_13_1083 ();
 FILLCELL_X2 FILLER_13_1087 ();
 FILLCELL_X1 FILLER_13_1089 ();
 FILLCELL_X8 FILLER_13_1099 ();
 FILLCELL_X2 FILLER_13_1107 ();
 FILLCELL_X16 FILLER_13_1113 ();
 FILLCELL_X4 FILLER_13_1129 ();
 FILLCELL_X2 FILLER_13_1133 ();
 FILLCELL_X4 FILLER_13_1138 ();
 FILLCELL_X1 FILLER_13_1142 ();
 FILLCELL_X8 FILLER_13_1145 ();
 FILLCELL_X1 FILLER_13_1153 ();
 FILLCELL_X4 FILLER_13_1157 ();
 FILLCELL_X4 FILLER_13_1171 ();
 FILLCELL_X1 FILLER_13_1175 ();
 FILLCELL_X4 FILLER_13_1186 ();
 FILLCELL_X1 FILLER_13_1190 ();
 FILLCELL_X4 FILLER_13_1195 ();
 FILLCELL_X8 FILLER_13_1202 ();
 FILLCELL_X2 FILLER_13_1210 ();
 FILLCELL_X1 FILLER_13_1212 ();
 FILLCELL_X4 FILLER_13_1216 ();
 FILLCELL_X8 FILLER_13_1223 ();
 FILLCELL_X4 FILLER_13_1234 ();
 FILLCELL_X8 FILLER_13_1248 ();
 FILLCELL_X4 FILLER_13_1259 ();
 FILLCELL_X4 FILLER_13_1264 ();
 FILLCELL_X4 FILLER_13_1277 ();
 FILLCELL_X4 FILLER_13_1283 ();
 FILLCELL_X4 FILLER_13_1297 ();
 FILLCELL_X16 FILLER_13_1304 ();
 FILLCELL_X8 FILLER_13_1320 ();
 FILLCELL_X4 FILLER_13_1328 ();
 FILLCELL_X2 FILLER_13_1332 ();
 FILLCELL_X8 FILLER_13_1338 ();
 FILLCELL_X1 FILLER_13_1346 ();
 FILLCELL_X4 FILLER_13_1356 ();
 FILLCELL_X2 FILLER_13_1360 ();
 FILLCELL_X8 FILLER_13_1364 ();
 FILLCELL_X2 FILLER_13_1372 ();
 FILLCELL_X8 FILLER_13_1377 ();
 FILLCELL_X4 FILLER_13_1385 ();
 FILLCELL_X2 FILLER_13_1389 ();
 FILLCELL_X1 FILLER_13_1391 ();
 FILLCELL_X4 FILLER_13_1394 ();
 FILLCELL_X32 FILLER_13_1408 ();
 FILLCELL_X32 FILLER_13_1440 ();
 FILLCELL_X32 FILLER_13_1472 ();
 FILLCELL_X32 FILLER_13_1504 ();
 FILLCELL_X32 FILLER_13_1536 ();
 FILLCELL_X32 FILLER_13_1568 ();
 FILLCELL_X32 FILLER_13_1600 ();
 FILLCELL_X32 FILLER_13_1632 ();
 FILLCELL_X32 FILLER_13_1664 ();
 FILLCELL_X32 FILLER_13_1696 ();
 FILLCELL_X16 FILLER_13_1728 ();
 FILLCELL_X8 FILLER_13_1744 ();
 FILLCELL_X4 FILLER_13_1752 ();
 FILLCELL_X4 FILLER_14_1 ();
 FILLCELL_X2 FILLER_14_5 ();
 FILLCELL_X4 FILLER_14_17 ();
 FILLCELL_X1 FILLER_14_21 ();
 FILLCELL_X4 FILLER_14_32 ();
 FILLCELL_X4 FILLER_14_45 ();
 FILLCELL_X4 FILLER_14_53 ();
 FILLCELL_X4 FILLER_14_66 ();
 FILLCELL_X2 FILLER_14_70 ();
 FILLCELL_X1 FILLER_14_72 ();
 FILLCELL_X16 FILLER_14_92 ();
 FILLCELL_X4 FILLER_14_108 ();
 FILLCELL_X8 FILLER_14_114 ();
 FILLCELL_X2 FILLER_14_122 ();
 FILLCELL_X4 FILLER_14_133 ();
 FILLCELL_X8 FILLER_14_147 ();
 FILLCELL_X4 FILLER_14_155 ();
 FILLCELL_X2 FILLER_14_159 ();
 FILLCELL_X1 FILLER_14_161 ();
 FILLCELL_X4 FILLER_14_166 ();
 FILLCELL_X1 FILLER_14_170 ();
 FILLCELL_X4 FILLER_14_173 ();
 FILLCELL_X4 FILLER_14_180 ();
 FILLCELL_X4 FILLER_14_191 ();
 FILLCELL_X4 FILLER_14_201 ();
 FILLCELL_X2 FILLER_14_205 ();
 FILLCELL_X4 FILLER_14_216 ();
 FILLCELL_X4 FILLER_14_229 ();
 FILLCELL_X2 FILLER_14_233 ();
 FILLCELL_X4 FILLER_14_245 ();
 FILLCELL_X1 FILLER_14_249 ();
 FILLCELL_X4 FILLER_14_260 ();
 FILLCELL_X8 FILLER_14_273 ();
 FILLCELL_X2 FILLER_14_281 ();
 FILLCELL_X8 FILLER_14_287 ();
 FILLCELL_X4 FILLER_14_295 ();
 FILLCELL_X1 FILLER_14_299 ();
 FILLCELL_X8 FILLER_14_304 ();
 FILLCELL_X1 FILLER_14_312 ();
 FILLCELL_X4 FILLER_14_317 ();
 FILLCELL_X2 FILLER_14_321 ();
 FILLCELL_X4 FILLER_14_326 ();
 FILLCELL_X4 FILLER_14_339 ();
 FILLCELL_X8 FILLER_14_353 ();
 FILLCELL_X4 FILLER_14_361 ();
 FILLCELL_X8 FILLER_14_375 ();
 FILLCELL_X4 FILLER_14_393 ();
 FILLCELL_X8 FILLER_14_401 ();
 FILLCELL_X16 FILLER_14_412 ();
 FILLCELL_X8 FILLER_14_428 ();
 FILLCELL_X1 FILLER_14_436 ();
 FILLCELL_X4 FILLER_14_440 ();
 FILLCELL_X8 FILLER_14_446 ();
 FILLCELL_X2 FILLER_14_454 ();
 FILLCELL_X8 FILLER_14_459 ();
 FILLCELL_X2 FILLER_14_467 ();
 FILLCELL_X8 FILLER_14_478 ();
 FILLCELL_X1 FILLER_14_486 ();
 FILLCELL_X4 FILLER_14_489 ();
 FILLCELL_X4 FILLER_14_496 ();
 FILLCELL_X2 FILLER_14_500 ();
 FILLCELL_X1 FILLER_14_502 ();
 FILLCELL_X4 FILLER_14_513 ();
 FILLCELL_X4 FILLER_14_521 ();
 FILLCELL_X1 FILLER_14_525 ();
 FILLCELL_X4 FILLER_14_528 ();
 FILLCELL_X2 FILLER_14_532 ();
 FILLCELL_X1 FILLER_14_534 ();
 FILLCELL_X8 FILLER_14_545 ();
 FILLCELL_X4 FILLER_14_553 ();
 FILLCELL_X2 FILLER_14_557 ();
 FILLCELL_X4 FILLER_14_562 ();
 FILLCELL_X8 FILLER_14_569 ();
 FILLCELL_X4 FILLER_14_577 ();
 FILLCELL_X2 FILLER_14_581 ();
 FILLCELL_X4 FILLER_14_586 ();
 FILLCELL_X4 FILLER_14_592 ();
 FILLCELL_X4 FILLER_14_600 ();
 FILLCELL_X2 FILLER_14_604 ();
 FILLCELL_X1 FILLER_14_606 ();
 FILLCELL_X4 FILLER_14_610 ();
 FILLCELL_X8 FILLER_14_617 ();
 FILLCELL_X4 FILLER_14_625 ();
 FILLCELL_X2 FILLER_14_629 ();
 FILLCELL_X4 FILLER_14_632 ();
 FILLCELL_X4 FILLER_14_639 ();
 FILLCELL_X2 FILLER_14_643 ();
 FILLCELL_X1 FILLER_14_645 ();
 FILLCELL_X8 FILLER_14_655 ();
 FILLCELL_X1 FILLER_14_663 ();
 FILLCELL_X4 FILLER_14_671 ();
 FILLCELL_X16 FILLER_14_678 ();
 FILLCELL_X2 FILLER_14_694 ();
 FILLCELL_X8 FILLER_14_698 ();
 FILLCELL_X4 FILLER_14_706 ();
 FILLCELL_X8 FILLER_14_713 ();
 FILLCELL_X4 FILLER_14_721 ();
 FILLCELL_X2 FILLER_14_725 ();
 FILLCELL_X1 FILLER_14_727 ();
 FILLCELL_X8 FILLER_14_732 ();
 FILLCELL_X2 FILLER_14_740 ();
 FILLCELL_X4 FILLER_14_748 ();
 FILLCELL_X8 FILLER_14_754 ();
 FILLCELL_X4 FILLER_14_762 ();
 FILLCELL_X2 FILLER_14_766 ();
 FILLCELL_X16 FILLER_14_775 ();
 FILLCELL_X8 FILLER_14_791 ();
 FILLCELL_X2 FILLER_14_799 ();
 FILLCELL_X4 FILLER_14_808 ();
 FILLCELL_X16 FILLER_14_815 ();
 FILLCELL_X4 FILLER_14_834 ();
 FILLCELL_X8 FILLER_14_842 ();
 FILLCELL_X1 FILLER_14_850 ();
 FILLCELL_X4 FILLER_14_853 ();
 FILLCELL_X4 FILLER_14_867 ();
 FILLCELL_X1 FILLER_14_871 ();
 FILLCELL_X4 FILLER_14_879 ();
 FILLCELL_X4 FILLER_14_893 ();
 FILLCELL_X4 FILLER_14_907 ();
 FILLCELL_X4 FILLER_14_920 ();
 FILLCELL_X1 FILLER_14_924 ();
 FILLCELL_X8 FILLER_14_935 ();
 FILLCELL_X1 FILLER_14_943 ();
 FILLCELL_X8 FILLER_14_954 ();
 FILLCELL_X4 FILLER_14_962 ();
 FILLCELL_X1 FILLER_14_966 ();
 FILLCELL_X32 FILLER_14_970 ();
 FILLCELL_X8 FILLER_14_1002 ();
 FILLCELL_X4 FILLER_14_1013 ();
 FILLCELL_X2 FILLER_14_1017 ();
 FILLCELL_X1 FILLER_14_1019 ();
 FILLCELL_X4 FILLER_14_1023 ();
 FILLCELL_X4 FILLER_14_1031 ();
 FILLCELL_X2 FILLER_14_1035 ();
 FILLCELL_X4 FILLER_14_1041 ();
 FILLCELL_X8 FILLER_14_1054 ();
 FILLCELL_X2 FILLER_14_1062 ();
 FILLCELL_X4 FILLER_14_1073 ();
 FILLCELL_X8 FILLER_14_1086 ();
 FILLCELL_X8 FILLER_14_1104 ();
 FILLCELL_X4 FILLER_14_1112 ();
 FILLCELL_X2 FILLER_14_1116 ();
 FILLCELL_X1 FILLER_14_1118 ();
 FILLCELL_X4 FILLER_14_1123 ();
 FILLCELL_X2 FILLER_14_1127 ();
 FILLCELL_X1 FILLER_14_1129 ();
 FILLCELL_X4 FILLER_14_1133 ();
 FILLCELL_X4 FILLER_14_1147 ();
 FILLCELL_X4 FILLER_14_1161 ();
 FILLCELL_X2 FILLER_14_1165 ();
 FILLCELL_X4 FILLER_14_1170 ();
 FILLCELL_X4 FILLER_14_1176 ();
 FILLCELL_X2 FILLER_14_1180 ();
 FILLCELL_X4 FILLER_14_1189 ();
 FILLCELL_X4 FILLER_14_1203 ();
 FILLCELL_X8 FILLER_14_1209 ();
 FILLCELL_X2 FILLER_14_1217 ();
 FILLCELL_X4 FILLER_14_1228 ();
 FILLCELL_X4 FILLER_14_1234 ();
 FILLCELL_X1 FILLER_14_1238 ();
 FILLCELL_X4 FILLER_14_1249 ();
 FILLCELL_X1 FILLER_14_1253 ();
 FILLCELL_X8 FILLER_14_1256 ();
 FILLCELL_X4 FILLER_14_1264 ();
 FILLCELL_X4 FILLER_14_1272 ();
 FILLCELL_X8 FILLER_14_1280 ();
 FILLCELL_X4 FILLER_14_1288 ();
 FILLCELL_X2 FILLER_14_1292 ();
 FILLCELL_X1 FILLER_14_1294 ();
 FILLCELL_X8 FILLER_14_1298 ();
 FILLCELL_X16 FILLER_14_1310 ();
 FILLCELL_X4 FILLER_14_1326 ();
 FILLCELL_X4 FILLER_14_1334 ();
 FILLCELL_X4 FILLER_14_1347 ();
 FILLCELL_X4 FILLER_14_1354 ();
 FILLCELL_X4 FILLER_14_1361 ();
 FILLCELL_X2 FILLER_14_1365 ();
 FILLCELL_X4 FILLER_14_1377 ();
 FILLCELL_X4 FILLER_14_1385 ();
 FILLCELL_X4 FILLER_14_1399 ();
 FILLCELL_X32 FILLER_14_1407 ();
 FILLCELL_X32 FILLER_14_1439 ();
 FILLCELL_X32 FILLER_14_1471 ();
 FILLCELL_X32 FILLER_14_1503 ();
 FILLCELL_X32 FILLER_14_1535 ();
 FILLCELL_X32 FILLER_14_1567 ();
 FILLCELL_X32 FILLER_14_1599 ();
 FILLCELL_X32 FILLER_14_1631 ();
 FILLCELL_X32 FILLER_14_1663 ();
 FILLCELL_X32 FILLER_14_1695 ();
 FILLCELL_X16 FILLER_14_1727 ();
 FILLCELL_X8 FILLER_14_1743 ();
 FILLCELL_X4 FILLER_14_1751 ();
 FILLCELL_X1 FILLER_14_1755 ();
 FILLCELL_X4 FILLER_15_1 ();
 FILLCELL_X2 FILLER_15_5 ();
 FILLCELL_X4 FILLER_15_16 ();
 FILLCELL_X4 FILLER_15_24 ();
 FILLCELL_X1 FILLER_15_28 ();
 FILLCELL_X4 FILLER_15_32 ();
 FILLCELL_X4 FILLER_15_39 ();
 FILLCELL_X4 FILLER_15_52 ();
 FILLCELL_X2 FILLER_15_56 ();
 FILLCELL_X16 FILLER_15_60 ();
 FILLCELL_X8 FILLER_15_76 ();
 FILLCELL_X4 FILLER_15_84 ();
 FILLCELL_X8 FILLER_15_97 ();
 FILLCELL_X1 FILLER_15_105 ();
 FILLCELL_X8 FILLER_15_116 ();
 FILLCELL_X4 FILLER_15_124 ();
 FILLCELL_X4 FILLER_15_138 ();
 FILLCELL_X4 FILLER_15_144 ();
 FILLCELL_X2 FILLER_15_148 ();
 FILLCELL_X1 FILLER_15_150 ();
 FILLCELL_X4 FILLER_15_170 ();
 FILLCELL_X8 FILLER_15_177 ();
 FILLCELL_X1 FILLER_15_185 ();
 FILLCELL_X8 FILLER_15_189 ();
 FILLCELL_X4 FILLER_15_197 ();
 FILLCELL_X2 FILLER_15_201 ();
 FILLCELL_X4 FILLER_15_206 ();
 FILLCELL_X4 FILLER_15_214 ();
 FILLCELL_X8 FILLER_15_221 ();
 FILLCELL_X4 FILLER_15_229 ();
 FILLCELL_X2 FILLER_15_233 ();
 FILLCELL_X4 FILLER_15_239 ();
 FILLCELL_X4 FILLER_15_246 ();
 FILLCELL_X8 FILLER_15_252 ();
 FILLCELL_X4 FILLER_15_260 ();
 FILLCELL_X8 FILLER_15_267 ();
 FILLCELL_X2 FILLER_15_275 ();
 FILLCELL_X1 FILLER_15_277 ();
 FILLCELL_X4 FILLER_15_282 ();
 FILLCELL_X4 FILLER_15_295 ();
 FILLCELL_X2 FILLER_15_299 ();
 FILLCELL_X4 FILLER_15_310 ();
 FILLCELL_X8 FILLER_15_324 ();
 FILLCELL_X8 FILLER_15_342 ();
 FILLCELL_X1 FILLER_15_350 ();
 FILLCELL_X8 FILLER_15_354 ();
 FILLCELL_X4 FILLER_15_364 ();
 FILLCELL_X1 FILLER_15_368 ();
 FILLCELL_X4 FILLER_15_372 ();
 FILLCELL_X4 FILLER_15_378 ();
 FILLCELL_X2 FILLER_15_382 ();
 FILLCELL_X1 FILLER_15_384 ();
 FILLCELL_X4 FILLER_15_388 ();
 FILLCELL_X8 FILLER_15_394 ();
 FILLCELL_X4 FILLER_15_402 ();
 FILLCELL_X1 FILLER_15_406 ();
 FILLCELL_X4 FILLER_15_417 ();
 FILLCELL_X1 FILLER_15_421 ();
 FILLCELL_X4 FILLER_15_425 ();
 FILLCELL_X2 FILLER_15_429 ();
 FILLCELL_X8 FILLER_15_435 ();
 FILLCELL_X2 FILLER_15_443 ();
 FILLCELL_X8 FILLER_15_449 ();
 FILLCELL_X2 FILLER_15_457 ();
 FILLCELL_X4 FILLER_15_463 ();
 FILLCELL_X8 FILLER_15_477 ();
 FILLCELL_X4 FILLER_15_485 ();
 FILLCELL_X4 FILLER_15_499 ();
 FILLCELL_X4 FILLER_15_512 ();
 FILLCELL_X2 FILLER_15_516 ();
 FILLCELL_X4 FILLER_15_522 ();
 FILLCELL_X2 FILLER_15_526 ();
 FILLCELL_X1 FILLER_15_528 ();
 FILLCELL_X4 FILLER_15_532 ();
 FILLCELL_X8 FILLER_15_540 ();
 FILLCELL_X2 FILLER_15_548 ();
 FILLCELL_X1 FILLER_15_550 ();
 FILLCELL_X8 FILLER_15_558 ();
 FILLCELL_X4 FILLER_15_566 ();
 FILLCELL_X2 FILLER_15_570 ();
 FILLCELL_X1 FILLER_15_572 ();
 FILLCELL_X8 FILLER_15_580 ();
 FILLCELL_X1 FILLER_15_588 ();
 FILLCELL_X4 FILLER_15_599 ();
 FILLCELL_X8 FILLER_15_606 ();
 FILLCELL_X4 FILLER_15_614 ();
 FILLCELL_X1 FILLER_15_618 ();
 FILLCELL_X4 FILLER_15_626 ();
 FILLCELL_X2 FILLER_15_630 ();
 FILLCELL_X4 FILLER_15_642 ();
 FILLCELL_X4 FILLER_15_656 ();
 FILLCELL_X4 FILLER_15_662 ();
 FILLCELL_X2 FILLER_15_666 ();
 FILLCELL_X4 FILLER_15_678 ();
 FILLCELL_X4 FILLER_15_691 ();
 FILLCELL_X2 FILLER_15_695 ();
 FILLCELL_X1 FILLER_15_697 ();
 FILLCELL_X4 FILLER_15_708 ();
 FILLCELL_X2 FILLER_15_712 ();
 FILLCELL_X1 FILLER_15_714 ();
 FILLCELL_X4 FILLER_15_724 ();
 FILLCELL_X2 FILLER_15_728 ();
 FILLCELL_X1 FILLER_15_730 ();
 FILLCELL_X4 FILLER_15_738 ();
 FILLCELL_X2 FILLER_15_742 ();
 FILLCELL_X1 FILLER_15_744 ();
 FILLCELL_X4 FILLER_15_751 ();
 FILLCELL_X8 FILLER_15_765 ();
 FILLCELL_X4 FILLER_15_773 ();
 FILLCELL_X1 FILLER_15_777 ();
 FILLCELL_X4 FILLER_15_781 ();
 FILLCELL_X8 FILLER_15_794 ();
 FILLCELL_X4 FILLER_15_805 ();
 FILLCELL_X4 FILLER_15_813 ();
 FILLCELL_X4 FILLER_15_821 ();
 FILLCELL_X2 FILLER_15_825 ();
 FILLCELL_X4 FILLER_15_830 ();
 FILLCELL_X4 FILLER_15_838 ();
 FILLCELL_X2 FILLER_15_842 ();
 FILLCELL_X8 FILLER_15_846 ();
 FILLCELL_X2 FILLER_15_854 ();
 FILLCELL_X4 FILLER_15_859 ();
 FILLCELL_X4 FILLER_15_873 ();
 FILLCELL_X1 FILLER_15_877 ();
 FILLCELL_X4 FILLER_15_888 ();
 FILLCELL_X8 FILLER_15_895 ();
 FILLCELL_X2 FILLER_15_903 ();
 FILLCELL_X8 FILLER_15_908 ();
 FILLCELL_X4 FILLER_15_916 ();
 FILLCELL_X4 FILLER_15_923 ();
 FILLCELL_X4 FILLER_15_930 ();
 FILLCELL_X4 FILLER_15_944 ();
 FILLCELL_X2 FILLER_15_948 ();
 FILLCELL_X1 FILLER_15_950 ();
 FILLCELL_X4 FILLER_15_954 ();
 FILLCELL_X2 FILLER_15_958 ();
 FILLCELL_X1 FILLER_15_960 ();
 FILLCELL_X4 FILLER_15_964 ();
 FILLCELL_X8 FILLER_15_977 ();
 FILLCELL_X4 FILLER_15_985 ();
 FILLCELL_X1 FILLER_15_989 ();
 FILLCELL_X4 FILLER_15_993 ();
 FILLCELL_X8 FILLER_15_1006 ();
 FILLCELL_X1 FILLER_15_1014 ();
 FILLCELL_X4 FILLER_15_1025 ();
 FILLCELL_X4 FILLER_15_1031 ();
 FILLCELL_X4 FILLER_15_1045 ();
 FILLCELL_X16 FILLER_15_1052 ();
 FILLCELL_X4 FILLER_15_1068 ();
 FILLCELL_X4 FILLER_15_1075 ();
 FILLCELL_X4 FILLER_15_1081 ();
 FILLCELL_X2 FILLER_15_1085 ();
 FILLCELL_X4 FILLER_15_1090 ();
 FILLCELL_X8 FILLER_15_1104 ();
 FILLCELL_X8 FILLER_15_1116 ();
 FILLCELL_X2 FILLER_15_1124 ();
 FILLCELL_X8 FILLER_15_1135 ();
 FILLCELL_X4 FILLER_15_1150 ();
 FILLCELL_X2 FILLER_15_1154 ();
 FILLCELL_X4 FILLER_15_1159 ();
 FILLCELL_X4 FILLER_15_1172 ();
 FILLCELL_X8 FILLER_15_1185 ();
 FILLCELL_X1 FILLER_15_1193 ();
 FILLCELL_X8 FILLER_15_1204 ();
 FILLCELL_X1 FILLER_15_1212 ();
 FILLCELL_X8 FILLER_15_1215 ();
 FILLCELL_X4 FILLER_15_1233 ();
 FILLCELL_X8 FILLER_15_1244 ();
 FILLCELL_X2 FILLER_15_1252 ();
 FILLCELL_X1 FILLER_15_1254 ();
 FILLCELL_X4 FILLER_15_1259 ();
 FILLCELL_X8 FILLER_15_1264 ();
 FILLCELL_X2 FILLER_15_1272 ();
 FILLCELL_X8 FILLER_15_1278 ();
 FILLCELL_X2 FILLER_15_1286 ();
 FILLCELL_X1 FILLER_15_1288 ();
 FILLCELL_X8 FILLER_15_1293 ();
 FILLCELL_X1 FILLER_15_1301 ();
 FILLCELL_X4 FILLER_15_1321 ();
 FILLCELL_X8 FILLER_15_1330 ();
 FILLCELL_X1 FILLER_15_1338 ();
 FILLCELL_X8 FILLER_15_1342 ();
 FILLCELL_X4 FILLER_15_1350 ();
 FILLCELL_X2 FILLER_15_1354 ();
 FILLCELL_X1 FILLER_15_1356 ();
 FILLCELL_X4 FILLER_15_1367 ();
 FILLCELL_X8 FILLER_15_1378 ();
 FILLCELL_X4 FILLER_15_1386 ();
 FILLCELL_X1 FILLER_15_1390 ();
 FILLCELL_X8 FILLER_15_1394 ();
 FILLCELL_X2 FILLER_15_1402 ();
 FILLCELL_X1 FILLER_15_1404 ();
 FILLCELL_X4 FILLER_15_1409 ();
 FILLCELL_X2 FILLER_15_1413 ();
 FILLCELL_X32 FILLER_15_1421 ();
 FILLCELL_X32 FILLER_15_1453 ();
 FILLCELL_X32 FILLER_15_1485 ();
 FILLCELL_X32 FILLER_15_1517 ();
 FILLCELL_X32 FILLER_15_1549 ();
 FILLCELL_X32 FILLER_15_1581 ();
 FILLCELL_X32 FILLER_15_1613 ();
 FILLCELL_X32 FILLER_15_1645 ();
 FILLCELL_X32 FILLER_15_1677 ();
 FILLCELL_X32 FILLER_15_1709 ();
 FILLCELL_X8 FILLER_15_1741 ();
 FILLCELL_X4 FILLER_15_1749 ();
 FILLCELL_X2 FILLER_15_1753 ();
 FILLCELL_X1 FILLER_15_1755 ();
 FILLCELL_X4 FILLER_16_1 ();
 FILLCELL_X4 FILLER_16_8 ();
 FILLCELL_X4 FILLER_16_15 ();
 FILLCELL_X8 FILLER_16_22 ();
 FILLCELL_X4 FILLER_16_33 ();
 FILLCELL_X2 FILLER_16_37 ();
 FILLCELL_X4 FILLER_16_42 ();
 FILLCELL_X4 FILLER_16_55 ();
 FILLCELL_X1 FILLER_16_59 ();
 FILLCELL_X4 FILLER_16_70 ();
 FILLCELL_X4 FILLER_16_84 ();
 FILLCELL_X1 FILLER_16_88 ();
 FILLCELL_X4 FILLER_16_92 ();
 FILLCELL_X4 FILLER_16_105 ();
 FILLCELL_X4 FILLER_16_112 ();
 FILLCELL_X2 FILLER_16_116 ();
 FILLCELL_X8 FILLER_16_125 ();
 FILLCELL_X2 FILLER_16_133 ();
 FILLCELL_X8 FILLER_16_139 ();
 FILLCELL_X4 FILLER_16_147 ();
 FILLCELL_X4 FILLER_16_154 ();
 FILLCELL_X8 FILLER_16_165 ();
 FILLCELL_X1 FILLER_16_173 ();
 FILLCELL_X8 FILLER_16_183 ();
 FILLCELL_X1 FILLER_16_191 ();
 FILLCELL_X8 FILLER_16_196 ();
 FILLCELL_X2 FILLER_16_204 ();
 FILLCELL_X8 FILLER_16_210 ();
 FILLCELL_X4 FILLER_16_218 ();
 FILLCELL_X2 FILLER_16_222 ();
 FILLCELL_X8 FILLER_16_228 ();
 FILLCELL_X4 FILLER_16_236 ();
 FILLCELL_X2 FILLER_16_240 ();
 FILLCELL_X4 FILLER_16_249 ();
 FILLCELL_X4 FILLER_16_263 ();
 FILLCELL_X4 FILLER_16_276 ();
 FILLCELL_X2 FILLER_16_280 ();
 FILLCELL_X1 FILLER_16_282 ();
 FILLCELL_X4 FILLER_16_286 ();
 FILLCELL_X4 FILLER_16_293 ();
 FILLCELL_X16 FILLER_16_300 ();
 FILLCELL_X4 FILLER_16_319 ();
 FILLCELL_X4 FILLER_16_330 ();
 FILLCELL_X8 FILLER_16_336 ();
 FILLCELL_X2 FILLER_16_344 ();
 FILLCELL_X8 FILLER_16_349 ();
 FILLCELL_X2 FILLER_16_357 ();
 FILLCELL_X1 FILLER_16_359 ();
 FILLCELL_X8 FILLER_16_363 ();
 FILLCELL_X4 FILLER_16_371 ();
 FILLCELL_X2 FILLER_16_375 ();
 FILLCELL_X1 FILLER_16_377 ();
 FILLCELL_X4 FILLER_16_381 ();
 FILLCELL_X1 FILLER_16_385 ();
 FILLCELL_X4 FILLER_16_396 ();
 FILLCELL_X2 FILLER_16_400 ();
 FILLCELL_X4 FILLER_16_406 ();
 FILLCELL_X4 FILLER_16_420 ();
 FILLCELL_X2 FILLER_16_424 ();
 FILLCELL_X4 FILLER_16_430 ();
 FILLCELL_X4 FILLER_16_443 ();
 FILLCELL_X4 FILLER_16_456 ();
 FILLCELL_X4 FILLER_16_465 ();
 FILLCELL_X4 FILLER_16_472 ();
 FILLCELL_X2 FILLER_16_476 ();
 FILLCELL_X1 FILLER_16_478 ();
 FILLCELL_X8 FILLER_16_486 ();
 FILLCELL_X1 FILLER_16_494 ();
 FILLCELL_X4 FILLER_16_498 ();
 FILLCELL_X4 FILLER_16_505 ();
 FILLCELL_X4 FILLER_16_513 ();
 FILLCELL_X4 FILLER_16_526 ();
 FILLCELL_X4 FILLER_16_539 ();
 FILLCELL_X4 FILLER_16_553 ();
 FILLCELL_X4 FILLER_16_567 ();
 FILLCELL_X8 FILLER_16_581 ();
 FILLCELL_X4 FILLER_16_592 ();
 FILLCELL_X4 FILLER_16_599 ();
 FILLCELL_X4 FILLER_16_613 ();
 FILLCELL_X4 FILLER_16_627 ();
 FILLCELL_X8 FILLER_16_632 ();
 FILLCELL_X4 FILLER_16_640 ();
 FILLCELL_X2 FILLER_16_644 ();
 FILLCELL_X4 FILLER_16_649 ();
 FILLCELL_X2 FILLER_16_653 ();
 FILLCELL_X4 FILLER_16_662 ();
 FILLCELL_X2 FILLER_16_666 ();
 FILLCELL_X1 FILLER_16_668 ();
 FILLCELL_X4 FILLER_16_672 ();
 FILLCELL_X4 FILLER_16_679 ();
 FILLCELL_X8 FILLER_16_692 ();
 FILLCELL_X2 FILLER_16_700 ();
 FILLCELL_X4 FILLER_16_705 ();
 FILLCELL_X4 FILLER_16_719 ();
 FILLCELL_X4 FILLER_16_726 ();
 FILLCELL_X4 FILLER_16_740 ();
 FILLCELL_X1 FILLER_16_744 ();
 FILLCELL_X4 FILLER_16_747 ();
 FILLCELL_X4 FILLER_16_761 ();
 FILLCELL_X8 FILLER_16_784 ();
 FILLCELL_X4 FILLER_16_795 ();
 FILLCELL_X4 FILLER_16_809 ();
 FILLCELL_X2 FILLER_16_813 ();
 FILLCELL_X8 FILLER_16_824 ();
 FILLCELL_X4 FILLER_16_842 ();
 FILLCELL_X2 FILLER_16_846 ();
 FILLCELL_X1 FILLER_16_848 ();
 FILLCELL_X16 FILLER_16_859 ();
 FILLCELL_X2 FILLER_16_875 ();
 FILLCELL_X32 FILLER_16_879 ();
 FILLCELL_X16 FILLER_16_911 ();
 FILLCELL_X2 FILLER_16_927 ();
 FILLCELL_X1 FILLER_16_929 ();
 FILLCELL_X4 FILLER_16_932 ();
 FILLCELL_X4 FILLER_16_943 ();
 FILLCELL_X4 FILLER_16_950 ();
 FILLCELL_X2 FILLER_16_954 ();
 FILLCELL_X8 FILLER_16_966 ();
 FILLCELL_X2 FILLER_16_974 ();
 FILLCELL_X4 FILLER_16_986 ();
 FILLCELL_X4 FILLER_16_999 ();
 FILLCELL_X4 FILLER_16_1010 ();
 FILLCELL_X1 FILLER_16_1014 ();
 FILLCELL_X8 FILLER_16_1017 ();
 FILLCELL_X2 FILLER_16_1025 ();
 FILLCELL_X4 FILLER_16_1031 ();
 FILLCELL_X8 FILLER_16_1037 ();
 FILLCELL_X1 FILLER_16_1045 ();
 FILLCELL_X4 FILLER_16_1049 ();
 FILLCELL_X4 FILLER_16_1057 ();
 FILLCELL_X8 FILLER_16_1070 ();
 FILLCELL_X1 FILLER_16_1078 ();
 FILLCELL_X4 FILLER_16_1086 ();
 FILLCELL_X2 FILLER_16_1090 ();
 FILLCELL_X1 FILLER_16_1092 ();
 FILLCELL_X4 FILLER_16_1100 ();
 FILLCELL_X2 FILLER_16_1104 ();
 FILLCELL_X4 FILLER_16_1108 ();
 FILLCELL_X1 FILLER_16_1112 ();
 FILLCELL_X4 FILLER_16_1117 ();
 FILLCELL_X4 FILLER_16_1130 ();
 FILLCELL_X4 FILLER_16_1137 ();
 FILLCELL_X4 FILLER_16_1144 ();
 FILLCELL_X1 FILLER_16_1148 ();
 FILLCELL_X8 FILLER_16_1152 ();
 FILLCELL_X4 FILLER_16_1167 ();
 FILLCELL_X16 FILLER_16_1174 ();
 FILLCELL_X1 FILLER_16_1190 ();
 FILLCELL_X8 FILLER_16_1194 ();
 FILLCELL_X1 FILLER_16_1202 ();
 FILLCELL_X4 FILLER_16_1222 ();
 FILLCELL_X4 FILLER_16_1229 ();
 FILLCELL_X4 FILLER_16_1235 ();
 FILLCELL_X4 FILLER_16_1246 ();
 FILLCELL_X4 FILLER_16_1260 ();
 FILLCELL_X4 FILLER_16_1274 ();
 FILLCELL_X2 FILLER_16_1278 ();
 FILLCELL_X4 FILLER_16_1289 ();
 FILLCELL_X16 FILLER_16_1302 ();
 FILLCELL_X8 FILLER_16_1318 ();
 FILLCELL_X4 FILLER_16_1326 ();
 FILLCELL_X1 FILLER_16_1330 ();
 FILLCELL_X4 FILLER_16_1335 ();
 FILLCELL_X4 FILLER_16_1348 ();
 FILLCELL_X4 FILLER_16_1354 ();
 FILLCELL_X4 FILLER_16_1362 ();
 FILLCELL_X8 FILLER_16_1369 ();
 FILLCELL_X4 FILLER_16_1377 ();
 FILLCELL_X2 FILLER_16_1381 ();
 FILLCELL_X4 FILLER_16_1392 ();
 FILLCELL_X1 FILLER_16_1396 ();
 FILLCELL_X4 FILLER_16_1401 ();
 FILLCELL_X4 FILLER_16_1412 ();
 FILLCELL_X8 FILLER_16_1422 ();
 FILLCELL_X4 FILLER_16_1430 ();
 FILLCELL_X2 FILLER_16_1434 ();
 FILLCELL_X32 FILLER_16_1440 ();
 FILLCELL_X32 FILLER_16_1472 ();
 FILLCELL_X32 FILLER_16_1504 ();
 FILLCELL_X32 FILLER_16_1536 ();
 FILLCELL_X32 FILLER_16_1568 ();
 FILLCELL_X32 FILLER_16_1600 ();
 FILLCELL_X32 FILLER_16_1632 ();
 FILLCELL_X32 FILLER_16_1664 ();
 FILLCELL_X32 FILLER_16_1696 ();
 FILLCELL_X16 FILLER_16_1728 ();
 FILLCELL_X8 FILLER_16_1744 ();
 FILLCELL_X4 FILLER_16_1752 ();
 FILLCELL_X8 FILLER_17_1 ();
 FILLCELL_X2 FILLER_17_9 ();
 FILLCELL_X4 FILLER_17_15 ();
 FILLCELL_X4 FILLER_17_23 ();
 FILLCELL_X8 FILLER_17_31 ();
 FILLCELL_X2 FILLER_17_39 ();
 FILLCELL_X16 FILLER_17_45 ();
 FILLCELL_X1 FILLER_17_61 ();
 FILLCELL_X4 FILLER_17_66 ();
 FILLCELL_X2 FILLER_17_70 ();
 FILLCELL_X16 FILLER_17_74 ();
 FILLCELL_X2 FILLER_17_90 ();
 FILLCELL_X4 FILLER_17_95 ();
 FILLCELL_X1 FILLER_17_99 ();
 FILLCELL_X8 FILLER_17_103 ();
 FILLCELL_X2 FILLER_17_111 ();
 FILLCELL_X4 FILLER_17_116 ();
 FILLCELL_X4 FILLER_17_129 ();
 FILLCELL_X4 FILLER_17_136 ();
 FILLCELL_X1 FILLER_17_140 ();
 FILLCELL_X4 FILLER_17_145 ();
 FILLCELL_X8 FILLER_17_159 ();
 FILLCELL_X2 FILLER_17_167 ();
 FILLCELL_X8 FILLER_17_179 ();
 FILLCELL_X4 FILLER_17_191 ();
 FILLCELL_X8 FILLER_17_204 ();
 FILLCELL_X8 FILLER_17_221 ();
 FILLCELL_X2 FILLER_17_229 ();
 FILLCELL_X1 FILLER_17_231 ();
 FILLCELL_X4 FILLER_17_236 ();
 FILLCELL_X16 FILLER_17_250 ();
 FILLCELL_X4 FILLER_17_266 ();
 FILLCELL_X2 FILLER_17_270 ();
 FILLCELL_X1 FILLER_17_272 ();
 FILLCELL_X4 FILLER_17_280 ();
 FILLCELL_X8 FILLER_17_286 ();
 FILLCELL_X2 FILLER_17_294 ();
 FILLCELL_X1 FILLER_17_296 ();
 FILLCELL_X4 FILLER_17_301 ();
 FILLCELL_X16 FILLER_17_309 ();
 FILLCELL_X2 FILLER_17_325 ();
 FILLCELL_X1 FILLER_17_327 ();
 FILLCELL_X8 FILLER_17_335 ();
 FILLCELL_X2 FILLER_17_343 ();
 FILLCELL_X4 FILLER_17_348 ();
 FILLCELL_X2 FILLER_17_352 ();
 FILLCELL_X4 FILLER_17_364 ();
 FILLCELL_X4 FILLER_17_378 ();
 FILLCELL_X4 FILLER_17_391 ();
 FILLCELL_X4 FILLER_17_398 ();
 FILLCELL_X8 FILLER_17_404 ();
 FILLCELL_X4 FILLER_17_416 ();
 FILLCELL_X4 FILLER_17_423 ();
 FILLCELL_X1 FILLER_17_427 ();
 FILLCELL_X4 FILLER_17_431 ();
 FILLCELL_X4 FILLER_17_438 ();
 FILLCELL_X16 FILLER_17_445 ();
 FILLCELL_X8 FILLER_17_461 ();
 FILLCELL_X4 FILLER_17_469 ();
 FILLCELL_X2 FILLER_17_473 ();
 FILLCELL_X1 FILLER_17_475 ();
 FILLCELL_X4 FILLER_17_483 ();
 FILLCELL_X2 FILLER_17_487 ();
 FILLCELL_X1 FILLER_17_489 ();
 FILLCELL_X4 FILLER_17_499 ();
 FILLCELL_X2 FILLER_17_503 ();
 FILLCELL_X1 FILLER_17_505 ();
 FILLCELL_X8 FILLER_17_510 ();
 FILLCELL_X2 FILLER_17_518 ();
 FILLCELL_X16 FILLER_17_523 ();
 FILLCELL_X8 FILLER_17_539 ();
 FILLCELL_X4 FILLER_17_547 ();
 FILLCELL_X2 FILLER_17_551 ();
 FILLCELL_X4 FILLER_17_556 ();
 FILLCELL_X8 FILLER_17_562 ();
 FILLCELL_X4 FILLER_17_574 ();
 FILLCELL_X2 FILLER_17_578 ();
 FILLCELL_X4 FILLER_17_583 ();
 FILLCELL_X4 FILLER_17_596 ();
 FILLCELL_X8 FILLER_17_609 ();
 FILLCELL_X2 FILLER_17_617 ();
 FILLCELL_X1 FILLER_17_619 ();
 FILLCELL_X8 FILLER_17_622 ();
 FILLCELL_X2 FILLER_17_630 ();
 FILLCELL_X1 FILLER_17_632 ();
 FILLCELL_X8 FILLER_17_642 ();
 FILLCELL_X1 FILLER_17_650 ();
 FILLCELL_X4 FILLER_17_661 ();
 FILLCELL_X2 FILLER_17_665 ();
 FILLCELL_X1 FILLER_17_667 ();
 FILLCELL_X16 FILLER_17_678 ();
 FILLCELL_X2 FILLER_17_694 ();
 FILLCELL_X16 FILLER_17_699 ();
 FILLCELL_X4 FILLER_17_715 ();
 FILLCELL_X2 FILLER_17_719 ();
 FILLCELL_X1 FILLER_17_721 ();
 FILLCELL_X4 FILLER_17_725 ();
 FILLCELL_X8 FILLER_17_734 ();
 FILLCELL_X1 FILLER_17_742 ();
 FILLCELL_X4 FILLER_17_747 ();
 FILLCELL_X4 FILLER_17_754 ();
 FILLCELL_X2 FILLER_17_758 ();
 FILLCELL_X1 FILLER_17_760 ();
 FILLCELL_X4 FILLER_17_765 ();
 FILLCELL_X8 FILLER_17_772 ();
 FILLCELL_X4 FILLER_17_780 ();
 FILLCELL_X2 FILLER_17_784 ();
 FILLCELL_X8 FILLER_17_789 ();
 FILLCELL_X2 FILLER_17_797 ();
 FILLCELL_X1 FILLER_17_799 ();
 FILLCELL_X8 FILLER_17_802 ();
 FILLCELL_X8 FILLER_17_817 ();
 FILLCELL_X4 FILLER_17_825 ();
 FILLCELL_X1 FILLER_17_829 ();
 FILLCELL_X4 FILLER_17_840 ();
 FILLCELL_X2 FILLER_17_844 ();
 FILLCELL_X1 FILLER_17_846 ();
 FILLCELL_X4 FILLER_17_850 ();
 FILLCELL_X4 FILLER_17_861 ();
 FILLCELL_X16 FILLER_17_868 ();
 FILLCELL_X2 FILLER_17_884 ();
 FILLCELL_X8 FILLER_17_889 ();
 FILLCELL_X4 FILLER_17_900 ();
 FILLCELL_X2 FILLER_17_904 ();
 FILLCELL_X4 FILLER_17_915 ();
 FILLCELL_X1 FILLER_17_919 ();
 FILLCELL_X4 FILLER_17_927 ();
 FILLCELL_X2 FILLER_17_931 ();
 FILLCELL_X4 FILLER_17_937 ();
 FILLCELL_X8 FILLER_17_944 ();
 FILLCELL_X1 FILLER_17_952 ();
 FILLCELL_X4 FILLER_17_963 ();
 FILLCELL_X4 FILLER_17_974 ();
 FILLCELL_X4 FILLER_17_980 ();
 FILLCELL_X4 FILLER_17_988 ();
 FILLCELL_X8 FILLER_17_1002 ();
 FILLCELL_X4 FILLER_17_1013 ();
 FILLCELL_X4 FILLER_17_1027 ();
 FILLCELL_X2 FILLER_17_1031 ();
 FILLCELL_X16 FILLER_17_1043 ();
 FILLCELL_X1 FILLER_17_1059 ();
 FILLCELL_X4 FILLER_17_1063 ();
 FILLCELL_X8 FILLER_17_1077 ();
 FILLCELL_X4 FILLER_17_1085 ();
 FILLCELL_X1 FILLER_17_1089 ();
 FILLCELL_X16 FILLER_17_1100 ();
 FILLCELL_X2 FILLER_17_1116 ();
 FILLCELL_X1 FILLER_17_1118 ();
 FILLCELL_X4 FILLER_17_1122 ();
 FILLCELL_X16 FILLER_17_1130 ();
 FILLCELL_X4 FILLER_17_1156 ();
 FILLCELL_X2 FILLER_17_1160 ();
 FILLCELL_X1 FILLER_17_1162 ();
 FILLCELL_X4 FILLER_17_1165 ();
 FILLCELL_X4 FILLER_17_1179 ();
 FILLCELL_X4 FILLER_17_1186 ();
 FILLCELL_X16 FILLER_17_1199 ();
 FILLCELL_X4 FILLER_17_1215 ();
 FILLCELL_X4 FILLER_17_1226 ();
 FILLCELL_X4 FILLER_17_1233 ();
 FILLCELL_X2 FILLER_17_1237 ();
 FILLCELL_X8 FILLER_17_1242 ();
 FILLCELL_X2 FILLER_17_1250 ();
 FILLCELL_X1 FILLER_17_1252 ();
 FILLCELL_X4 FILLER_17_1256 ();
 FILLCELL_X2 FILLER_17_1260 ();
 FILLCELL_X1 FILLER_17_1262 ();
 FILLCELL_X4 FILLER_17_1264 ();
 FILLCELL_X4 FILLER_17_1278 ();
 FILLCELL_X2 FILLER_17_1282 ();
 FILLCELL_X1 FILLER_17_1284 ();
 FILLCELL_X4 FILLER_17_1288 ();
 FILLCELL_X32 FILLER_17_1295 ();
 FILLCELL_X1 FILLER_17_1327 ();
 FILLCELL_X4 FILLER_17_1337 ();
 FILLCELL_X8 FILLER_17_1344 ();
 FILLCELL_X4 FILLER_17_1356 ();
 FILLCELL_X2 FILLER_17_1360 ();
 FILLCELL_X1 FILLER_17_1362 ();
 FILLCELL_X4 FILLER_17_1366 ();
 FILLCELL_X4 FILLER_17_1379 ();
 FILLCELL_X4 FILLER_17_1387 ();
 FILLCELL_X32 FILLER_17_1394 ();
 FILLCELL_X32 FILLER_17_1426 ();
 FILLCELL_X4 FILLER_17_1458 ();
 FILLCELL_X1 FILLER_17_1462 ();
 FILLCELL_X32 FILLER_17_1482 ();
 FILLCELL_X32 FILLER_17_1514 ();
 FILLCELL_X32 FILLER_17_1546 ();
 FILLCELL_X32 FILLER_17_1578 ();
 FILLCELL_X32 FILLER_17_1610 ();
 FILLCELL_X32 FILLER_17_1642 ();
 FILLCELL_X32 FILLER_17_1674 ();
 FILLCELL_X32 FILLER_17_1706 ();
 FILLCELL_X16 FILLER_17_1738 ();
 FILLCELL_X2 FILLER_17_1754 ();
 FILLCELL_X4 FILLER_18_1 ();
 FILLCELL_X2 FILLER_18_5 ();
 FILLCELL_X1 FILLER_18_7 ();
 FILLCELL_X8 FILLER_18_17 ();
 FILLCELL_X4 FILLER_18_34 ();
 FILLCELL_X16 FILLER_18_41 ();
 FILLCELL_X1 FILLER_18_57 ();
 FILLCELL_X4 FILLER_18_68 ();
 FILLCELL_X8 FILLER_18_79 ();
 FILLCELL_X2 FILLER_18_87 ();
 FILLCELL_X8 FILLER_18_99 ();
 FILLCELL_X2 FILLER_18_107 ();
 FILLCELL_X1 FILLER_18_109 ();
 FILLCELL_X4 FILLER_18_113 ();
 FILLCELL_X4 FILLER_18_126 ();
 FILLCELL_X4 FILLER_18_133 ();
 FILLCELL_X1 FILLER_18_137 ();
 FILLCELL_X8 FILLER_18_142 ();
 FILLCELL_X2 FILLER_18_150 ();
 FILLCELL_X16 FILLER_18_156 ();
 FILLCELL_X8 FILLER_18_172 ();
 FILLCELL_X4 FILLER_18_180 ();
 FILLCELL_X4 FILLER_18_187 ();
 FILLCELL_X2 FILLER_18_191 ();
 FILLCELL_X1 FILLER_18_193 ();
 FILLCELL_X4 FILLER_18_197 ();
 FILLCELL_X2 FILLER_18_201 ();
 FILLCELL_X1 FILLER_18_203 ();
 FILLCELL_X4 FILLER_18_210 ();
 FILLCELL_X4 FILLER_18_220 ();
 FILLCELL_X4 FILLER_18_237 ();
 FILLCELL_X16 FILLER_18_244 ();
 FILLCELL_X8 FILLER_18_260 ();
 FILLCELL_X2 FILLER_18_268 ();
 FILLCELL_X1 FILLER_18_270 ();
 FILLCELL_X4 FILLER_18_281 ();
 FILLCELL_X4 FILLER_18_289 ();
 FILLCELL_X4 FILLER_18_302 ();
 FILLCELL_X4 FILLER_18_315 ();
 FILLCELL_X4 FILLER_18_329 ();
 FILLCELL_X4 FILLER_18_343 ();
 FILLCELL_X8 FILLER_18_356 ();
 FILLCELL_X1 FILLER_18_364 ();
 FILLCELL_X8 FILLER_18_368 ();
 FILLCELL_X2 FILLER_18_376 ();
 FILLCELL_X4 FILLER_18_381 ();
 FILLCELL_X1 FILLER_18_385 ();
 FILLCELL_X4 FILLER_18_396 ();
 FILLCELL_X4 FILLER_18_407 ();
 FILLCELL_X4 FILLER_18_418 ();
 FILLCELL_X4 FILLER_18_425 ();
 FILLCELL_X1 FILLER_18_429 ();
 FILLCELL_X4 FILLER_18_434 ();
 FILLCELL_X2 FILLER_18_438 ();
 FILLCELL_X4 FILLER_18_444 ();
 FILLCELL_X4 FILLER_18_451 ();
 FILLCELL_X2 FILLER_18_455 ();
 FILLCELL_X1 FILLER_18_457 ();
 FILLCELL_X4 FILLER_18_461 ();
 FILLCELL_X8 FILLER_18_474 ();
 FILLCELL_X4 FILLER_18_482 ();
 FILLCELL_X4 FILLER_18_496 ();
 FILLCELL_X1 FILLER_18_500 ();
 FILLCELL_X8 FILLER_18_520 ();
 FILLCELL_X4 FILLER_18_528 ();
 FILLCELL_X4 FILLER_18_534 ();
 FILLCELL_X1 FILLER_18_538 ();
 FILLCELL_X16 FILLER_18_548 ();
 FILLCELL_X2 FILLER_18_564 ();
 FILLCELL_X1 FILLER_18_566 ();
 FILLCELL_X4 FILLER_18_571 ();
 FILLCELL_X4 FILLER_18_578 ();
 FILLCELL_X16 FILLER_18_585 ();
 FILLCELL_X4 FILLER_18_601 ();
 FILLCELL_X1 FILLER_18_605 ();
 FILLCELL_X8 FILLER_18_608 ();
 FILLCELL_X4 FILLER_18_625 ();
 FILLCELL_X2 FILLER_18_629 ();
 FILLCELL_X4 FILLER_18_632 ();
 FILLCELL_X1 FILLER_18_636 ();
 FILLCELL_X8 FILLER_18_640 ();
 FILLCELL_X4 FILLER_18_650 ();
 FILLCELL_X4 FILLER_18_658 ();
 FILLCELL_X1 FILLER_18_662 ();
 FILLCELL_X4 FILLER_18_665 ();
 FILLCELL_X2 FILLER_18_669 ();
 FILLCELL_X4 FILLER_18_675 ();
 FILLCELL_X2 FILLER_18_679 ();
 FILLCELL_X1 FILLER_18_681 ();
 FILLCELL_X8 FILLER_18_686 ();
 FILLCELL_X2 FILLER_18_694 ();
 FILLCELL_X4 FILLER_18_699 ();
 FILLCELL_X4 FILLER_18_707 ();
 FILLCELL_X8 FILLER_18_720 ();
 FILLCELL_X1 FILLER_18_728 ();
 FILLCELL_X4 FILLER_18_731 ();
 FILLCELL_X1 FILLER_18_735 ();
 FILLCELL_X4 FILLER_18_739 ();
 FILLCELL_X8 FILLER_18_746 ();
 FILLCELL_X1 FILLER_18_754 ();
 FILLCELL_X4 FILLER_18_764 ();
 FILLCELL_X2 FILLER_18_768 ();
 FILLCELL_X1 FILLER_18_770 ();
 FILLCELL_X4 FILLER_18_774 ();
 FILLCELL_X4 FILLER_18_787 ();
 FILLCELL_X4 FILLER_18_801 ();
 FILLCELL_X8 FILLER_18_812 ();
 FILLCELL_X2 FILLER_18_820 ();
 FILLCELL_X16 FILLER_18_828 ();
 FILLCELL_X4 FILLER_18_844 ();
 FILLCELL_X1 FILLER_18_848 ();
 FILLCELL_X4 FILLER_18_859 ();
 FILLCELL_X8 FILLER_18_872 ();
 FILLCELL_X1 FILLER_18_880 ();
 FILLCELL_X4 FILLER_18_884 ();
 FILLCELL_X8 FILLER_18_897 ();
 FILLCELL_X2 FILLER_18_905 ();
 FILLCELL_X1 FILLER_18_907 ();
 FILLCELL_X4 FILLER_18_918 ();
 FILLCELL_X4 FILLER_18_932 ();
 FILLCELL_X1 FILLER_18_936 ();
 FILLCELL_X8 FILLER_18_946 ();
 FILLCELL_X1 FILLER_18_954 ();
 FILLCELL_X4 FILLER_18_964 ();
 FILLCELL_X8 FILLER_18_971 ();
 FILLCELL_X2 FILLER_18_979 ();
 FILLCELL_X8 FILLER_18_984 ();
 FILLCELL_X1 FILLER_18_992 ();
 FILLCELL_X4 FILLER_18_996 ();
 FILLCELL_X2 FILLER_18_1000 ();
 FILLCELL_X1 FILLER_18_1002 ();
 FILLCELL_X8 FILLER_18_1007 ();
 FILLCELL_X2 FILLER_18_1015 ();
 FILLCELL_X4 FILLER_18_1023 ();
 FILLCELL_X4 FILLER_18_1033 ();
 FILLCELL_X2 FILLER_18_1037 ();
 FILLCELL_X4 FILLER_18_1049 ();
 FILLCELL_X16 FILLER_18_1060 ();
 FILLCELL_X1 FILLER_18_1076 ();
 FILLCELL_X8 FILLER_18_1080 ();
 FILLCELL_X4 FILLER_18_1091 ();
 FILLCELL_X2 FILLER_18_1095 ();
 FILLCELL_X1 FILLER_18_1097 ();
 FILLCELL_X16 FILLER_18_1107 ();
 FILLCELL_X8 FILLER_18_1123 ();
 FILLCELL_X2 FILLER_18_1131 ();
 FILLCELL_X1 FILLER_18_1133 ();
 FILLCELL_X4 FILLER_18_1137 ();
 FILLCELL_X8 FILLER_18_1151 ();
 FILLCELL_X4 FILLER_18_1161 ();
 FILLCELL_X2 FILLER_18_1165 ();
 FILLCELL_X8 FILLER_18_1174 ();
 FILLCELL_X4 FILLER_18_1182 ();
 FILLCELL_X2 FILLER_18_1186 ();
 FILLCELL_X4 FILLER_18_1191 ();
 FILLCELL_X8 FILLER_18_1204 ();
 FILLCELL_X2 FILLER_18_1212 ();
 FILLCELL_X4 FILLER_18_1216 ();
 FILLCELL_X4 FILLER_18_1230 ();
 FILLCELL_X4 FILLER_18_1243 ();
 FILLCELL_X4 FILLER_18_1256 ();
 FILLCELL_X16 FILLER_18_1263 ();
 FILLCELL_X4 FILLER_18_1279 ();
 FILLCELL_X2 FILLER_18_1283 ();
 FILLCELL_X4 FILLER_18_1289 ();
 FILLCELL_X1 FILLER_18_1293 ();
 FILLCELL_X4 FILLER_18_1298 ();
 FILLCELL_X4 FILLER_18_1321 ();
 FILLCELL_X4 FILLER_18_1329 ();
 FILLCELL_X8 FILLER_18_1337 ();
 FILLCELL_X1 FILLER_18_1345 ();
 FILLCELL_X8 FILLER_18_1350 ();
 FILLCELL_X1 FILLER_18_1358 ();
 FILLCELL_X8 FILLER_18_1368 ();
 FILLCELL_X4 FILLER_18_1376 ();
 FILLCELL_X2 FILLER_18_1380 ();
 FILLCELL_X8 FILLER_18_1385 ();
 FILLCELL_X1 FILLER_18_1393 ();
 FILLCELL_X32 FILLER_18_1400 ();
 FILLCELL_X32 FILLER_18_1432 ();
 FILLCELL_X32 FILLER_18_1464 ();
 FILLCELL_X32 FILLER_18_1496 ();
 FILLCELL_X32 FILLER_18_1528 ();
 FILLCELL_X32 FILLER_18_1560 ();
 FILLCELL_X32 FILLER_18_1592 ();
 FILLCELL_X32 FILLER_18_1624 ();
 FILLCELL_X32 FILLER_18_1656 ();
 FILLCELL_X32 FILLER_18_1688 ();
 FILLCELL_X32 FILLER_18_1720 ();
 FILLCELL_X4 FILLER_18_1752 ();
 FILLCELL_X4 FILLER_19_1 ();
 FILLCELL_X4 FILLER_19_7 ();
 FILLCELL_X4 FILLER_19_14 ();
 FILLCELL_X8 FILLER_19_20 ();
 FILLCELL_X4 FILLER_19_31 ();
 FILLCELL_X2 FILLER_19_35 ();
 FILLCELL_X4 FILLER_19_39 ();
 FILLCELL_X4 FILLER_19_53 ();
 FILLCELL_X4 FILLER_19_60 ();
 FILLCELL_X4 FILLER_19_71 ();
 FILLCELL_X4 FILLER_19_85 ();
 FILLCELL_X4 FILLER_19_93 ();
 FILLCELL_X2 FILLER_19_97 ();
 FILLCELL_X1 FILLER_19_99 ();
 FILLCELL_X4 FILLER_19_110 ();
 FILLCELL_X1 FILLER_19_114 ();
 FILLCELL_X4 FILLER_19_125 ();
 FILLCELL_X8 FILLER_19_135 ();
 FILLCELL_X1 FILLER_19_143 ();
 FILLCELL_X4 FILLER_19_150 ();
 FILLCELL_X2 FILLER_19_154 ();
 FILLCELL_X8 FILLER_19_162 ();
 FILLCELL_X4 FILLER_19_170 ();
 FILLCELL_X1 FILLER_19_174 ();
 FILLCELL_X4 FILLER_19_192 ();
 FILLCELL_X4 FILLER_19_202 ();
 FILLCELL_X8 FILLER_19_209 ();
 FILLCELL_X4 FILLER_19_217 ();
 FILLCELL_X2 FILLER_19_221 ();
 FILLCELL_X8 FILLER_19_227 ();
 FILLCELL_X4 FILLER_19_235 ();
 FILLCELL_X1 FILLER_19_239 ();
 FILLCELL_X4 FILLER_19_244 ();
 FILLCELL_X8 FILLER_19_257 ();
 FILLCELL_X4 FILLER_19_268 ();
 FILLCELL_X8 FILLER_19_282 ();
 FILLCELL_X4 FILLER_19_290 ();
 FILLCELL_X4 FILLER_19_297 ();
 FILLCELL_X4 FILLER_19_304 ();
 FILLCELL_X8 FILLER_19_311 ();
 FILLCELL_X4 FILLER_19_319 ();
 FILLCELL_X4 FILLER_19_327 ();
 FILLCELL_X4 FILLER_19_334 ();
 FILLCELL_X4 FILLER_19_340 ();
 FILLCELL_X2 FILLER_19_344 ();
 FILLCELL_X8 FILLER_19_349 ();
 FILLCELL_X4 FILLER_19_366 ();
 FILLCELL_X2 FILLER_19_370 ();
 FILLCELL_X4 FILLER_19_381 ();
 FILLCELL_X2 FILLER_19_385 ();
 FILLCELL_X1 FILLER_19_387 ();
 FILLCELL_X8 FILLER_19_398 ();
 FILLCELL_X2 FILLER_19_406 ();
 FILLCELL_X1 FILLER_19_408 ();
 FILLCELL_X4 FILLER_19_418 ();
 FILLCELL_X4 FILLER_19_427 ();
 FILLCELL_X2 FILLER_19_431 ();
 FILLCELL_X1 FILLER_19_433 ();
 FILLCELL_X4 FILLER_19_443 ();
 FILLCELL_X8 FILLER_19_456 ();
 FILLCELL_X1 FILLER_19_464 ();
 FILLCELL_X4 FILLER_19_475 ();
 FILLCELL_X1 FILLER_19_479 ();
 FILLCELL_X8 FILLER_19_482 ();
 FILLCELL_X16 FILLER_19_493 ();
 FILLCELL_X4 FILLER_19_509 ();
 FILLCELL_X4 FILLER_19_516 ();
 FILLCELL_X4 FILLER_19_523 ();
 FILLCELL_X4 FILLER_19_530 ();
 FILLCELL_X4 FILLER_19_537 ();
 FILLCELL_X4 FILLER_19_551 ();
 FILLCELL_X8 FILLER_19_564 ();
 FILLCELL_X4 FILLER_19_576 ();
 FILLCELL_X8 FILLER_19_589 ();
 FILLCELL_X4 FILLER_19_604 ();
 FILLCELL_X8 FILLER_19_618 ();
 FILLCELL_X2 FILLER_19_626 ();
 FILLCELL_X4 FILLER_19_638 ();
 FILLCELL_X4 FILLER_19_652 ();
 FILLCELL_X4 FILLER_19_659 ();
 FILLCELL_X4 FILLER_19_667 ();
 FILLCELL_X4 FILLER_19_680 ();
 FILLCELL_X8 FILLER_19_693 ();
 FILLCELL_X2 FILLER_19_701 ();
 FILLCELL_X4 FILLER_19_712 ();
 FILLCELL_X4 FILLER_19_720 ();
 FILLCELL_X4 FILLER_19_727 ();
 FILLCELL_X1 FILLER_19_731 ();
 FILLCELL_X4 FILLER_19_736 ();
 FILLCELL_X4 FILLER_19_749 ();
 FILLCELL_X8 FILLER_19_756 ();
 FILLCELL_X8 FILLER_19_773 ();
 FILLCELL_X2 FILLER_19_781 ();
 FILLCELL_X4 FILLER_19_793 ();
 FILLCELL_X2 FILLER_19_797 ();
 FILLCELL_X1 FILLER_19_799 ();
 FILLCELL_X4 FILLER_19_803 ();
 FILLCELL_X4 FILLER_19_811 ();
 FILLCELL_X2 FILLER_19_815 ();
 FILLCELL_X1 FILLER_19_817 ();
 FILLCELL_X4 FILLER_19_821 ();
 FILLCELL_X4 FILLER_19_829 ();
 FILLCELL_X16 FILLER_19_842 ();
 FILLCELL_X4 FILLER_19_858 ();
 FILLCELL_X1 FILLER_19_862 ();
 FILLCELL_X4 FILLER_19_870 ();
 FILLCELL_X4 FILLER_19_884 ();
 FILLCELL_X4 FILLER_19_898 ();
 FILLCELL_X4 FILLER_19_906 ();
 FILLCELL_X1 FILLER_19_910 ();
 FILLCELL_X8 FILLER_19_914 ();
 FILLCELL_X8 FILLER_19_924 ();
 FILLCELL_X2 FILLER_19_932 ();
 FILLCELL_X8 FILLER_19_938 ();
 FILLCELL_X4 FILLER_19_949 ();
 FILLCELL_X8 FILLER_19_957 ();
 FILLCELL_X4 FILLER_19_965 ();
 FILLCELL_X4 FILLER_19_972 ();
 FILLCELL_X4 FILLER_19_983 ();
 FILLCELL_X4 FILLER_19_989 ();
 FILLCELL_X1 FILLER_19_993 ();
 FILLCELL_X4 FILLER_19_998 ();
 FILLCELL_X8 FILLER_19_1015 ();
 FILLCELL_X2 FILLER_19_1023 ();
 FILLCELL_X1 FILLER_19_1025 ();
 FILLCELL_X4 FILLER_19_1036 ();
 FILLCELL_X4 FILLER_19_1043 ();
 FILLCELL_X2 FILLER_19_1047 ();
 FILLCELL_X1 FILLER_19_1049 ();
 FILLCELL_X8 FILLER_19_1060 ();
 FILLCELL_X4 FILLER_19_1072 ();
 FILLCELL_X4 FILLER_19_1086 ();
 FILLCELL_X4 FILLER_19_1097 ();
 FILLCELL_X4 FILLER_19_1104 ();
 FILLCELL_X8 FILLER_19_1110 ();
 FILLCELL_X1 FILLER_19_1118 ();
 FILLCELL_X4 FILLER_19_1122 ();
 FILLCELL_X2 FILLER_19_1126 ();
 FILLCELL_X8 FILLER_19_1137 ();
 FILLCELL_X2 FILLER_19_1145 ();
 FILLCELL_X1 FILLER_19_1147 ();
 FILLCELL_X4 FILLER_19_1152 ();
 FILLCELL_X2 FILLER_19_1156 ();
 FILLCELL_X4 FILLER_19_1161 ();
 FILLCELL_X4 FILLER_19_1175 ();
 FILLCELL_X2 FILLER_19_1179 ();
 FILLCELL_X1 FILLER_19_1181 ();
 FILLCELL_X8 FILLER_19_1192 ();
 FILLCELL_X4 FILLER_19_1203 ();
 FILLCELL_X16 FILLER_19_1209 ();
 FILLCELL_X8 FILLER_19_1225 ();
 FILLCELL_X4 FILLER_19_1233 ();
 FILLCELL_X2 FILLER_19_1237 ();
 FILLCELL_X1 FILLER_19_1239 ();
 FILLCELL_X8 FILLER_19_1243 ();
 FILLCELL_X1 FILLER_19_1251 ();
 FILLCELL_X4 FILLER_19_1259 ();
 FILLCELL_X4 FILLER_19_1264 ();
 FILLCELL_X2 FILLER_19_1268 ();
 FILLCELL_X1 FILLER_19_1270 ();
 FILLCELL_X4 FILLER_19_1274 ();
 FILLCELL_X4 FILLER_19_1285 ();
 FILLCELL_X16 FILLER_19_1291 ();
 FILLCELL_X4 FILLER_19_1307 ();
 FILLCELL_X1 FILLER_19_1311 ();
 FILLCELL_X16 FILLER_19_1315 ();
 FILLCELL_X8 FILLER_19_1331 ();
 FILLCELL_X1 FILLER_19_1339 ();
 FILLCELL_X4 FILLER_19_1344 ();
 FILLCELL_X4 FILLER_19_1351 ();
 FILLCELL_X4 FILLER_19_1360 ();
 FILLCELL_X8 FILLER_19_1369 ();
 FILLCELL_X4 FILLER_19_1377 ();
 FILLCELL_X4 FILLER_19_1383 ();
 FILLCELL_X32 FILLER_19_1406 ();
 FILLCELL_X32 FILLER_19_1438 ();
 FILLCELL_X32 FILLER_19_1470 ();
 FILLCELL_X32 FILLER_19_1502 ();
 FILLCELL_X32 FILLER_19_1534 ();
 FILLCELL_X32 FILLER_19_1566 ();
 FILLCELL_X32 FILLER_19_1598 ();
 FILLCELL_X32 FILLER_19_1630 ();
 FILLCELL_X32 FILLER_19_1662 ();
 FILLCELL_X32 FILLER_19_1694 ();
 FILLCELL_X16 FILLER_19_1726 ();
 FILLCELL_X8 FILLER_19_1742 ();
 FILLCELL_X4 FILLER_19_1750 ();
 FILLCELL_X2 FILLER_19_1754 ();
 FILLCELL_X4 FILLER_20_1 ();
 FILLCELL_X8 FILLER_20_9 ();
 FILLCELL_X4 FILLER_20_22 ();
 FILLCELL_X8 FILLER_20_30 ();
 FILLCELL_X4 FILLER_20_38 ();
 FILLCELL_X2 FILLER_20_42 ();
 FILLCELL_X1 FILLER_20_44 ();
 FILLCELL_X8 FILLER_20_52 ();
 FILLCELL_X4 FILLER_20_60 ();
 FILLCELL_X2 FILLER_20_64 ();
 FILLCELL_X4 FILLER_20_75 ();
 FILLCELL_X4 FILLER_20_82 ();
 FILLCELL_X2 FILLER_20_86 ();
 FILLCELL_X1 FILLER_20_88 ();
 FILLCELL_X8 FILLER_20_91 ();
 FILLCELL_X8 FILLER_20_101 ();
 FILLCELL_X4 FILLER_20_109 ();
 FILLCELL_X2 FILLER_20_113 ();
 FILLCELL_X8 FILLER_20_117 ();
 FILLCELL_X2 FILLER_20_125 ();
 FILLCELL_X16 FILLER_20_129 ();
 FILLCELL_X2 FILLER_20_145 ();
 FILLCELL_X8 FILLER_20_154 ();
 FILLCELL_X4 FILLER_20_169 ();
 FILLCELL_X4 FILLER_20_182 ();
 FILLCELL_X8 FILLER_20_193 ();
 FILLCELL_X4 FILLER_20_208 ();
 FILLCELL_X4 FILLER_20_215 ();
 FILLCELL_X2 FILLER_20_219 ();
 FILLCELL_X8 FILLER_20_225 ();
 FILLCELL_X4 FILLER_20_233 ();
 FILLCELL_X1 FILLER_20_237 ();
 FILLCELL_X4 FILLER_20_242 ();
 FILLCELL_X4 FILLER_20_255 ();
 FILLCELL_X4 FILLER_20_262 ();
 FILLCELL_X4 FILLER_20_275 ();
 FILLCELL_X8 FILLER_20_283 ();
 FILLCELL_X4 FILLER_20_291 ();
 FILLCELL_X1 FILLER_20_295 ();
 FILLCELL_X4 FILLER_20_300 ();
 FILLCELL_X1 FILLER_20_304 ();
 FILLCELL_X16 FILLER_20_309 ();
 FILLCELL_X4 FILLER_20_325 ();
 FILLCELL_X2 FILLER_20_329 ();
 FILLCELL_X1 FILLER_20_331 ();
 FILLCELL_X16 FILLER_20_335 ();
 FILLCELL_X2 FILLER_20_351 ();
 FILLCELL_X8 FILLER_20_355 ();
 FILLCELL_X2 FILLER_20_363 ();
 FILLCELL_X16 FILLER_20_375 ();
 FILLCELL_X4 FILLER_20_391 ();
 FILLCELL_X1 FILLER_20_395 ();
 FILLCELL_X8 FILLER_20_398 ();
 FILLCELL_X4 FILLER_20_406 ();
 FILLCELL_X1 FILLER_20_410 ();
 FILLCELL_X4 FILLER_20_420 ();
 FILLCELL_X8 FILLER_20_428 ();
 FILLCELL_X4 FILLER_20_440 ();
 FILLCELL_X8 FILLER_20_447 ();
 FILLCELL_X4 FILLER_20_455 ();
 FILLCELL_X8 FILLER_20_463 ();
 FILLCELL_X1 FILLER_20_471 ();
 FILLCELL_X4 FILLER_20_479 ();
 FILLCELL_X4 FILLER_20_486 ();
 FILLCELL_X1 FILLER_20_490 ();
 FILLCELL_X4 FILLER_20_494 ();
 FILLCELL_X8 FILLER_20_501 ();
 FILLCELL_X4 FILLER_20_513 ();
 FILLCELL_X4 FILLER_20_527 ();
 FILLCELL_X8 FILLER_20_538 ();
 FILLCELL_X1 FILLER_20_546 ();
 FILLCELL_X4 FILLER_20_550 ();
 FILLCELL_X4 FILLER_20_557 ();
 FILLCELL_X4 FILLER_20_565 ();
 FILLCELL_X4 FILLER_20_578 ();
 FILLCELL_X2 FILLER_20_582 ();
 FILLCELL_X1 FILLER_20_584 ();
 FILLCELL_X4 FILLER_20_589 ();
 FILLCELL_X4 FILLER_20_603 ();
 FILLCELL_X2 FILLER_20_607 ();
 FILLCELL_X4 FILLER_20_612 ();
 FILLCELL_X4 FILLER_20_619 ();
 FILLCELL_X4 FILLER_20_627 ();
 FILLCELL_X4 FILLER_20_632 ();
 FILLCELL_X8 FILLER_20_639 ();
 FILLCELL_X4 FILLER_20_647 ();
 FILLCELL_X2 FILLER_20_651 ();
 FILLCELL_X1 FILLER_20_653 ();
 FILLCELL_X4 FILLER_20_658 ();
 FILLCELL_X4 FILLER_20_665 ();
 FILLCELL_X2 FILLER_20_669 ();
 FILLCELL_X1 FILLER_20_671 ();
 FILLCELL_X4 FILLER_20_675 ();
 FILLCELL_X16 FILLER_20_682 ();
 FILLCELL_X2 FILLER_20_698 ();
 FILLCELL_X1 FILLER_20_700 ();
 FILLCELL_X8 FILLER_20_705 ();
 FILLCELL_X2 FILLER_20_713 ();
 FILLCELL_X4 FILLER_20_718 ();
 FILLCELL_X4 FILLER_20_731 ();
 FILLCELL_X16 FILLER_20_744 ();
 FILLCELL_X2 FILLER_20_760 ();
 FILLCELL_X16 FILLER_20_765 ();
 FILLCELL_X8 FILLER_20_785 ();
 FILLCELL_X2 FILLER_20_793 ();
 FILLCELL_X4 FILLER_20_798 ();
 FILLCELL_X4 FILLER_20_806 ();
 FILLCELL_X16 FILLER_20_819 ();
 FILLCELL_X8 FILLER_20_839 ();
 FILLCELL_X2 FILLER_20_847 ();
 FILLCELL_X1 FILLER_20_849 ();
 FILLCELL_X4 FILLER_20_853 ();
 FILLCELL_X4 FILLER_20_867 ();
 FILLCELL_X4 FILLER_20_873 ();
 FILLCELL_X2 FILLER_20_877 ();
 FILLCELL_X4 FILLER_20_882 ();
 FILLCELL_X4 FILLER_20_893 ();
 FILLCELL_X8 FILLER_20_899 ();
 FILLCELL_X4 FILLER_20_907 ();
 FILLCELL_X4 FILLER_20_915 ();
 FILLCELL_X1 FILLER_20_919 ();
 FILLCELL_X32 FILLER_20_924 ();
 FILLCELL_X2 FILLER_20_956 ();
 FILLCELL_X1 FILLER_20_958 ();
 FILLCELL_X4 FILLER_20_969 ();
 FILLCELL_X2 FILLER_20_973 ();
 FILLCELL_X1 FILLER_20_975 ();
 FILLCELL_X4 FILLER_20_986 ();
 FILLCELL_X16 FILLER_20_999 ();
 FILLCELL_X4 FILLER_20_1015 ();
 FILLCELL_X1 FILLER_20_1019 ();
 FILLCELL_X4 FILLER_20_1022 ();
 FILLCELL_X4 FILLER_20_1033 ();
 FILLCELL_X2 FILLER_20_1037 ();
 FILLCELL_X1 FILLER_20_1039 ();
 FILLCELL_X4 FILLER_20_1043 ();
 FILLCELL_X4 FILLER_20_1050 ();
 FILLCELL_X4 FILLER_20_1057 ();
 FILLCELL_X4 FILLER_20_1064 ();
 FILLCELL_X2 FILLER_20_1068 ();
 FILLCELL_X4 FILLER_20_1079 ();
 FILLCELL_X2 FILLER_20_1083 ();
 FILLCELL_X1 FILLER_20_1085 ();
 FILLCELL_X4 FILLER_20_1090 ();
 FILLCELL_X1 FILLER_20_1094 ();
 FILLCELL_X4 FILLER_20_1114 ();
 FILLCELL_X8 FILLER_20_1128 ();
 FILLCELL_X4 FILLER_20_1146 ();
 FILLCELL_X32 FILLER_20_1152 ();
 FILLCELL_X8 FILLER_20_1184 ();
 FILLCELL_X1 FILLER_20_1192 ();
 FILLCELL_X4 FILLER_20_1203 ();
 FILLCELL_X4 FILLER_20_1216 ();
 FILLCELL_X4 FILLER_20_1223 ();
 FILLCELL_X4 FILLER_20_1230 ();
 FILLCELL_X4 FILLER_20_1237 ();
 FILLCELL_X1 FILLER_20_1241 ();
 FILLCELL_X4 FILLER_20_1245 ();
 FILLCELL_X4 FILLER_20_1259 ();
 FILLCELL_X4 FILLER_20_1273 ();
 FILLCELL_X4 FILLER_20_1287 ();
 FILLCELL_X1 FILLER_20_1291 ();
 FILLCELL_X4 FILLER_20_1302 ();
 FILLCELL_X1 FILLER_20_1306 ();
 FILLCELL_X4 FILLER_20_1310 ();
 FILLCELL_X4 FILLER_20_1320 ();
 FILLCELL_X4 FILLER_20_1330 ();
 FILLCELL_X8 FILLER_20_1338 ();
 FILLCELL_X4 FILLER_20_1346 ();
 FILLCELL_X2 FILLER_20_1350 ();
 FILLCELL_X1 FILLER_20_1352 ();
 FILLCELL_X4 FILLER_20_1357 ();
 FILLCELL_X2 FILLER_20_1361 ();
 FILLCELL_X1 FILLER_20_1363 ();
 FILLCELL_X8 FILLER_20_1367 ();
 FILLCELL_X2 FILLER_20_1375 ();
 FILLCELL_X4 FILLER_20_1381 ();
 FILLCELL_X32 FILLER_20_1395 ();
 FILLCELL_X32 FILLER_20_1427 ();
 FILLCELL_X32 FILLER_20_1459 ();
 FILLCELL_X32 FILLER_20_1491 ();
 FILLCELL_X32 FILLER_20_1523 ();
 FILLCELL_X32 FILLER_20_1555 ();
 FILLCELL_X32 FILLER_20_1587 ();
 FILLCELL_X32 FILLER_20_1619 ();
 FILLCELL_X32 FILLER_20_1651 ();
 FILLCELL_X32 FILLER_20_1683 ();
 FILLCELL_X32 FILLER_20_1715 ();
 FILLCELL_X2 FILLER_20_1747 ();
 FILLCELL_X4 FILLER_20_1752 ();
 FILLCELL_X4 FILLER_21_1 ();
 FILLCELL_X2 FILLER_21_5 ();
 FILLCELL_X4 FILLER_21_14 ();
 FILLCELL_X4 FILLER_21_35 ();
 FILLCELL_X1 FILLER_21_39 ();
 FILLCELL_X4 FILLER_21_50 ();
 FILLCELL_X8 FILLER_21_58 ();
 FILLCELL_X8 FILLER_21_75 ();
 FILLCELL_X2 FILLER_21_83 ();
 FILLCELL_X4 FILLER_21_88 ();
 FILLCELL_X4 FILLER_21_102 ();
 FILLCELL_X4 FILLER_21_113 ();
 FILLCELL_X4 FILLER_21_121 ();
 FILLCELL_X2 FILLER_21_125 ();
 FILLCELL_X1 FILLER_21_127 ();
 FILLCELL_X4 FILLER_21_135 ();
 FILLCELL_X2 FILLER_21_139 ();
 FILLCELL_X1 FILLER_21_141 ();
 FILLCELL_X16 FILLER_21_145 ();
 FILLCELL_X1 FILLER_21_161 ();
 FILLCELL_X4 FILLER_21_167 ();
 FILLCELL_X4 FILLER_21_180 ();
 FILLCELL_X8 FILLER_21_186 ();
 FILLCELL_X8 FILLER_21_200 ();
 FILLCELL_X2 FILLER_21_208 ();
 FILLCELL_X4 FILLER_21_220 ();
 FILLCELL_X4 FILLER_21_234 ();
 FILLCELL_X4 FILLER_21_241 ();
 FILLCELL_X2 FILLER_21_245 ();
 FILLCELL_X4 FILLER_21_252 ();
 FILLCELL_X8 FILLER_21_259 ();
 FILLCELL_X16 FILLER_21_271 ();
 FILLCELL_X4 FILLER_21_290 ();
 FILLCELL_X4 FILLER_21_303 ();
 FILLCELL_X4 FILLER_21_310 ();
 FILLCELL_X4 FILLER_21_318 ();
 FILLCELL_X4 FILLER_21_326 ();
 FILLCELL_X4 FILLER_21_334 ();
 FILLCELL_X4 FILLER_21_343 ();
 FILLCELL_X8 FILLER_21_364 ();
 FILLCELL_X1 FILLER_21_372 ();
 FILLCELL_X4 FILLER_21_383 ();
 FILLCELL_X16 FILLER_21_390 ();
 FILLCELL_X8 FILLER_21_406 ();
 FILLCELL_X2 FILLER_21_414 ();
 FILLCELL_X8 FILLER_21_419 ();
 FILLCELL_X4 FILLER_21_427 ();
 FILLCELL_X4 FILLER_21_434 ();
 FILLCELL_X4 FILLER_21_441 ();
 FILLCELL_X8 FILLER_21_449 ();
 FILLCELL_X1 FILLER_21_457 ();
 FILLCELL_X4 FILLER_21_461 ();
 FILLCELL_X4 FILLER_21_475 ();
 FILLCELL_X4 FILLER_21_489 ();
 FILLCELL_X4 FILLER_21_497 ();
 FILLCELL_X2 FILLER_21_501 ();
 FILLCELL_X16 FILLER_21_512 ();
 FILLCELL_X8 FILLER_21_528 ();
 FILLCELL_X2 FILLER_21_536 ();
 FILLCELL_X1 FILLER_21_538 ();
 FILLCELL_X4 FILLER_21_542 ();
 FILLCELL_X8 FILLER_21_555 ();
 FILLCELL_X4 FILLER_21_563 ();
 FILLCELL_X1 FILLER_21_567 ();
 FILLCELL_X16 FILLER_21_571 ();
 FILLCELL_X2 FILLER_21_587 ();
 FILLCELL_X4 FILLER_21_592 ();
 FILLCELL_X8 FILLER_21_599 ();
 FILLCELL_X1 FILLER_21_607 ();
 FILLCELL_X4 FILLER_21_612 ();
 FILLCELL_X16 FILLER_21_619 ();
 FILLCELL_X4 FILLER_21_635 ();
 FILLCELL_X1 FILLER_21_639 ();
 FILLCELL_X4 FILLER_21_643 ();
 FILLCELL_X4 FILLER_21_651 ();
 FILLCELL_X8 FILLER_21_664 ();
 FILLCELL_X8 FILLER_21_676 ();
 FILLCELL_X4 FILLER_21_684 ();
 FILLCELL_X2 FILLER_21_688 ();
 FILLCELL_X1 FILLER_21_690 ();
 FILLCELL_X8 FILLER_21_695 ();
 FILLCELL_X4 FILLER_21_703 ();
 FILLCELL_X4 FILLER_21_710 ();
 FILLCELL_X1 FILLER_21_714 ();
 FILLCELL_X4 FILLER_21_719 ();
 FILLCELL_X4 FILLER_21_727 ();
 FILLCELL_X2 FILLER_21_731 ();
 FILLCELL_X1 FILLER_21_733 ();
 FILLCELL_X4 FILLER_21_737 ();
 FILLCELL_X4 FILLER_21_743 ();
 FILLCELL_X2 FILLER_21_747 ();
 FILLCELL_X4 FILLER_21_756 ();
 FILLCELL_X4 FILLER_21_770 ();
 FILLCELL_X2 FILLER_21_774 ();
 FILLCELL_X1 FILLER_21_776 ();
 FILLCELL_X4 FILLER_21_780 ();
 FILLCELL_X4 FILLER_21_787 ();
 FILLCELL_X4 FILLER_21_795 ();
 FILLCELL_X2 FILLER_21_799 ();
 FILLCELL_X4 FILLER_21_804 ();
 FILLCELL_X8 FILLER_21_812 ();
 FILLCELL_X1 FILLER_21_820 ();
 FILLCELL_X4 FILLER_21_827 ();
 FILLCELL_X2 FILLER_21_831 ();
 FILLCELL_X4 FILLER_21_842 ();
 FILLCELL_X4 FILLER_21_850 ();
 FILLCELL_X2 FILLER_21_854 ();
 FILLCELL_X1 FILLER_21_856 ();
 FILLCELL_X8 FILLER_21_861 ();
 FILLCELL_X1 FILLER_21_869 ();
 FILLCELL_X4 FILLER_21_874 ();
 FILLCELL_X8 FILLER_21_888 ();
 FILLCELL_X2 FILLER_21_896 ();
 FILLCELL_X4 FILLER_21_901 ();
 FILLCELL_X4 FILLER_21_909 ();
 FILLCELL_X4 FILLER_21_922 ();
 FILLCELL_X4 FILLER_21_935 ();
 FILLCELL_X4 FILLER_21_943 ();
 FILLCELL_X8 FILLER_21_950 ();
 FILLCELL_X8 FILLER_21_962 ();
 FILLCELL_X4 FILLER_21_970 ();
 FILLCELL_X1 FILLER_21_974 ();
 FILLCELL_X4 FILLER_21_978 ();
 FILLCELL_X8 FILLER_21_985 ();
 FILLCELL_X4 FILLER_21_993 ();
 FILLCELL_X4 FILLER_21_1001 ();
 FILLCELL_X8 FILLER_21_1008 ();
 FILLCELL_X4 FILLER_21_1016 ();
 FILLCELL_X4 FILLER_21_1023 ();
 FILLCELL_X4 FILLER_21_1036 ();
 FILLCELL_X4 FILLER_21_1043 ();
 FILLCELL_X2 FILLER_21_1047 ();
 FILLCELL_X4 FILLER_21_1058 ();
 FILLCELL_X2 FILLER_21_1062 ();
 FILLCELL_X1 FILLER_21_1064 ();
 FILLCELL_X4 FILLER_21_1069 ();
 FILLCELL_X4 FILLER_21_1076 ();
 FILLCELL_X2 FILLER_21_1080 ();
 FILLCELL_X8 FILLER_21_1086 ();
 FILLCELL_X2 FILLER_21_1094 ();
 FILLCELL_X1 FILLER_21_1096 ();
 FILLCELL_X4 FILLER_21_1101 ();
 FILLCELL_X16 FILLER_21_1108 ();
 FILLCELL_X4 FILLER_21_1124 ();
 FILLCELL_X2 FILLER_21_1128 ();
 FILLCELL_X1 FILLER_21_1130 ();
 FILLCELL_X4 FILLER_21_1134 ();
 FILLCELL_X1 FILLER_21_1138 ();
 FILLCELL_X4 FILLER_21_1146 ();
 FILLCELL_X2 FILLER_21_1150 ();
 FILLCELL_X1 FILLER_21_1152 ();
 FILLCELL_X4 FILLER_21_1160 ();
 FILLCELL_X8 FILLER_21_1170 ();
 FILLCELL_X8 FILLER_21_1188 ();
 FILLCELL_X4 FILLER_21_1196 ();
 FILLCELL_X1 FILLER_21_1200 ();
 FILLCELL_X8 FILLER_21_1204 ();
 FILLCELL_X2 FILLER_21_1212 ();
 FILLCELL_X4 FILLER_21_1223 ();
 FILLCELL_X4 FILLER_21_1236 ();
 FILLCELL_X4 FILLER_21_1249 ();
 FILLCELL_X4 FILLER_21_1256 ();
 FILLCELL_X2 FILLER_21_1260 ();
 FILLCELL_X1 FILLER_21_1262 ();
 FILLCELL_X8 FILLER_21_1264 ();
 FILLCELL_X4 FILLER_21_1281 ();
 FILLCELL_X4 FILLER_21_1288 ();
 FILLCELL_X8 FILLER_21_1295 ();
 FILLCELL_X2 FILLER_21_1303 ();
 FILLCELL_X4 FILLER_21_1308 ();
 FILLCELL_X1 FILLER_21_1312 ();
 FILLCELL_X4 FILLER_21_1326 ();
 FILLCELL_X1 FILLER_21_1330 ();
 FILLCELL_X4 FILLER_21_1350 ();
 FILLCELL_X4 FILLER_21_1358 ();
 FILLCELL_X4 FILLER_21_1371 ();
 FILLCELL_X4 FILLER_21_1384 ();
 FILLCELL_X2 FILLER_21_1388 ();
 FILLCELL_X1 FILLER_21_1390 ();
 FILLCELL_X4 FILLER_21_1398 ();
 FILLCELL_X32 FILLER_21_1405 ();
 FILLCELL_X32 FILLER_21_1437 ();
 FILLCELL_X32 FILLER_21_1469 ();
 FILLCELL_X32 FILLER_21_1501 ();
 FILLCELL_X32 FILLER_21_1533 ();
 FILLCELL_X32 FILLER_21_1565 ();
 FILLCELL_X32 FILLER_21_1597 ();
 FILLCELL_X32 FILLER_21_1629 ();
 FILLCELL_X32 FILLER_21_1661 ();
 FILLCELL_X32 FILLER_21_1693 ();
 FILLCELL_X16 FILLER_21_1725 ();
 FILLCELL_X8 FILLER_21_1741 ();
 FILLCELL_X4 FILLER_21_1749 ();
 FILLCELL_X2 FILLER_21_1753 ();
 FILLCELL_X1 FILLER_21_1755 ();
 FILLCELL_X4 FILLER_22_1 ();
 FILLCELL_X8 FILLER_22_8 ();
 FILLCELL_X4 FILLER_22_21 ();
 FILLCELL_X16 FILLER_22_29 ();
 FILLCELL_X4 FILLER_22_49 ();
 FILLCELL_X4 FILLER_22_56 ();
 FILLCELL_X1 FILLER_22_60 ();
 FILLCELL_X4 FILLER_22_64 ();
 FILLCELL_X4 FILLER_22_71 ();
 FILLCELL_X8 FILLER_22_78 ();
 FILLCELL_X1 FILLER_22_86 ();
 FILLCELL_X4 FILLER_22_94 ();
 FILLCELL_X4 FILLER_22_101 ();
 FILLCELL_X2 FILLER_22_105 ();
 FILLCELL_X1 FILLER_22_107 ();
 FILLCELL_X4 FILLER_22_117 ();
 FILLCELL_X4 FILLER_22_131 ();
 FILLCELL_X1 FILLER_22_135 ();
 FILLCELL_X4 FILLER_22_139 ();
 FILLCELL_X4 FILLER_22_153 ();
 FILLCELL_X4 FILLER_22_164 ();
 FILLCELL_X16 FILLER_22_173 ();
 FILLCELL_X2 FILLER_22_189 ();
 FILLCELL_X4 FILLER_22_195 ();
 FILLCELL_X16 FILLER_22_203 ();
 FILLCELL_X16 FILLER_22_221 ();
 FILLCELL_X4 FILLER_22_239 ();
 FILLCELL_X16 FILLER_22_246 ();
 FILLCELL_X8 FILLER_22_262 ();
 FILLCELL_X8 FILLER_22_274 ();
 FILLCELL_X2 FILLER_22_282 ();
 FILLCELL_X4 FILLER_22_293 ();
 FILLCELL_X8 FILLER_22_301 ();
 FILLCELL_X2 FILLER_22_309 ();
 FILLCELL_X4 FILLER_22_314 ();
 FILLCELL_X8 FILLER_22_327 ();
 FILLCELL_X2 FILLER_22_335 ();
 FILLCELL_X4 FILLER_22_342 ();
 FILLCELL_X8 FILLER_22_353 ();
 FILLCELL_X4 FILLER_22_363 ();
 FILLCELL_X4 FILLER_22_371 ();
 FILLCELL_X8 FILLER_22_382 ();
 FILLCELL_X4 FILLER_22_390 ();
 FILLCELL_X1 FILLER_22_394 ();
 FILLCELL_X4 FILLER_22_399 ();
 FILLCELL_X1 FILLER_22_403 ();
 FILLCELL_X8 FILLER_22_413 ();
 FILLCELL_X4 FILLER_22_421 ();
 FILLCELL_X2 FILLER_22_425 ();
 FILLCELL_X4 FILLER_22_430 ();
 FILLCELL_X8 FILLER_22_443 ();
 FILLCELL_X8 FILLER_22_460 ();
 FILLCELL_X1 FILLER_22_468 ();
 FILLCELL_X4 FILLER_22_473 ();
 FILLCELL_X8 FILLER_22_479 ();
 FILLCELL_X4 FILLER_22_491 ();
 FILLCELL_X4 FILLER_22_504 ();
 FILLCELL_X8 FILLER_22_512 ();
 FILLCELL_X4 FILLER_22_520 ();
 FILLCELL_X2 FILLER_22_524 ();
 FILLCELL_X4 FILLER_22_529 ();
 FILLCELL_X16 FILLER_22_542 ();
 FILLCELL_X4 FILLER_22_561 ();
 FILLCELL_X8 FILLER_22_568 ();
 FILLCELL_X8 FILLER_22_585 ();
 FILLCELL_X2 FILLER_22_593 ();
 FILLCELL_X8 FILLER_22_605 ();
 FILLCELL_X1 FILLER_22_613 ();
 FILLCELL_X8 FILLER_22_623 ();
 FILLCELL_X4 FILLER_22_632 ();
 FILLCELL_X4 FILLER_22_642 ();
 FILLCELL_X1 FILLER_22_646 ();
 FILLCELL_X8 FILLER_22_651 ();
 FILLCELL_X4 FILLER_22_668 ();
 FILLCELL_X2 FILLER_22_672 ();
 FILLCELL_X1 FILLER_22_674 ();
 FILLCELL_X8 FILLER_22_679 ();
 FILLCELL_X1 FILLER_22_687 ();
 FILLCELL_X4 FILLER_22_693 ();
 FILLCELL_X2 FILLER_22_697 ();
 FILLCELL_X1 FILLER_22_699 ();
 FILLCELL_X4 FILLER_22_704 ();
 FILLCELL_X2 FILLER_22_708 ();
 FILLCELL_X1 FILLER_22_710 ();
 FILLCELL_X8 FILLER_22_715 ();
 FILLCELL_X4 FILLER_22_723 ();
 FILLCELL_X2 FILLER_22_727 ();
 FILLCELL_X4 FILLER_22_732 ();
 FILLCELL_X2 FILLER_22_736 ();
 FILLCELL_X4 FILLER_22_741 ();
 FILLCELL_X4 FILLER_22_748 ();
 FILLCELL_X4 FILLER_22_762 ();
 FILLCELL_X4 FILLER_22_768 ();
 FILLCELL_X4 FILLER_22_775 ();
 FILLCELL_X8 FILLER_22_788 ();
 FILLCELL_X1 FILLER_22_796 ();
 FILLCELL_X4 FILLER_22_806 ();
 FILLCELL_X4 FILLER_22_814 ();
 FILLCELL_X4 FILLER_22_827 ();
 FILLCELL_X8 FILLER_22_840 ();
 FILLCELL_X1 FILLER_22_848 ();
 FILLCELL_X4 FILLER_22_853 ();
 FILLCELL_X4 FILLER_22_861 ();
 FILLCELL_X16 FILLER_22_869 ();
 FILLCELL_X4 FILLER_22_885 ();
 FILLCELL_X2 FILLER_22_889 ();
 FILLCELL_X4 FILLER_22_895 ();
 FILLCELL_X8 FILLER_22_903 ();
 FILLCELL_X4 FILLER_22_914 ();
 FILLCELL_X8 FILLER_22_921 ();
 FILLCELL_X2 FILLER_22_929 ();
 FILLCELL_X4 FILLER_22_935 ();
 FILLCELL_X4 FILLER_22_948 ();
 FILLCELL_X16 FILLER_22_956 ();
 FILLCELL_X2 FILLER_22_972 ();
 FILLCELL_X1 FILLER_22_974 ();
 FILLCELL_X4 FILLER_22_978 ();
 FILLCELL_X2 FILLER_22_982 ();
 FILLCELL_X4 FILLER_22_987 ();
 FILLCELL_X4 FILLER_22_995 ();
 FILLCELL_X4 FILLER_22_1008 ();
 FILLCELL_X8 FILLER_22_1015 ();
 FILLCELL_X1 FILLER_22_1023 ();
 FILLCELL_X4 FILLER_22_1034 ();
 FILLCELL_X2 FILLER_22_1038 ();
 FILLCELL_X4 FILLER_22_1047 ();
 FILLCELL_X4 FILLER_22_1054 ();
 FILLCELL_X1 FILLER_22_1058 ();
 FILLCELL_X8 FILLER_22_1063 ();
 FILLCELL_X1 FILLER_22_1071 ();
 FILLCELL_X4 FILLER_22_1081 ();
 FILLCELL_X1 FILLER_22_1085 ();
 FILLCELL_X8 FILLER_22_1095 ();
 FILLCELL_X8 FILLER_22_1113 ();
 FILLCELL_X1 FILLER_22_1121 ();
 FILLCELL_X4 FILLER_22_1131 ();
 FILLCELL_X4 FILLER_22_1145 ();
 FILLCELL_X1 FILLER_22_1149 ();
 FILLCELL_X4 FILLER_22_1152 ();
 FILLCELL_X4 FILLER_22_1166 ();
 FILLCELL_X2 FILLER_22_1170 ();
 FILLCELL_X4 FILLER_22_1178 ();
 FILLCELL_X8 FILLER_22_1195 ();
 FILLCELL_X2 FILLER_22_1203 ();
 FILLCELL_X1 FILLER_22_1205 ();
 FILLCELL_X4 FILLER_22_1209 ();
 FILLCELL_X4 FILLER_22_1216 ();
 FILLCELL_X2 FILLER_22_1220 ();
 FILLCELL_X1 FILLER_22_1222 ();
 FILLCELL_X8 FILLER_22_1226 ();
 FILLCELL_X4 FILLER_22_1244 ();
 FILLCELL_X4 FILLER_22_1250 ();
 FILLCELL_X4 FILLER_22_1264 ();
 FILLCELL_X4 FILLER_22_1271 ();
 FILLCELL_X4 FILLER_22_1277 ();
 FILLCELL_X4 FILLER_22_1283 ();
 FILLCELL_X2 FILLER_22_1287 ();
 FILLCELL_X4 FILLER_22_1298 ();
 FILLCELL_X1 FILLER_22_1302 ();
 FILLCELL_X4 FILLER_22_1309 ();
 FILLCELL_X32 FILLER_22_1317 ();
 FILLCELL_X8 FILLER_22_1349 ();
 FILLCELL_X2 FILLER_22_1357 ();
 FILLCELL_X1 FILLER_22_1359 ();
 FILLCELL_X4 FILLER_22_1364 ();
 FILLCELL_X4 FILLER_22_1371 ();
 FILLCELL_X4 FILLER_22_1378 ();
 FILLCELL_X4 FILLER_22_1385 ();
 FILLCELL_X2 FILLER_22_1389 ();
 FILLCELL_X32 FILLER_22_1400 ();
 FILLCELL_X32 FILLER_22_1432 ();
 FILLCELL_X32 FILLER_22_1464 ();
 FILLCELL_X32 FILLER_22_1496 ();
 FILLCELL_X32 FILLER_22_1528 ();
 FILLCELL_X32 FILLER_22_1560 ();
 FILLCELL_X32 FILLER_22_1592 ();
 FILLCELL_X32 FILLER_22_1624 ();
 FILLCELL_X32 FILLER_22_1656 ();
 FILLCELL_X32 FILLER_22_1688 ();
 FILLCELL_X32 FILLER_22_1720 ();
 FILLCELL_X4 FILLER_22_1752 ();
 FILLCELL_X4 FILLER_23_1 ();
 FILLCELL_X2 FILLER_23_5 ();
 FILLCELL_X8 FILLER_23_17 ();
 FILLCELL_X8 FILLER_23_28 ();
 FILLCELL_X1 FILLER_23_36 ();
 FILLCELL_X8 FILLER_23_56 ();
 FILLCELL_X4 FILLER_23_64 ();
 FILLCELL_X1 FILLER_23_68 ();
 FILLCELL_X8 FILLER_23_73 ();
 FILLCELL_X2 FILLER_23_81 ();
 FILLCELL_X4 FILLER_23_87 ();
 FILLCELL_X8 FILLER_23_101 ();
 FILLCELL_X2 FILLER_23_109 ();
 FILLCELL_X8 FILLER_23_121 ();
 FILLCELL_X2 FILLER_23_129 ();
 FILLCELL_X1 FILLER_23_131 ();
 FILLCELL_X4 FILLER_23_135 ();
 FILLCELL_X8 FILLER_23_148 ();
 FILLCELL_X1 FILLER_23_156 ();
 FILLCELL_X4 FILLER_23_163 ();
 FILLCELL_X4 FILLER_23_174 ();
 FILLCELL_X2 FILLER_23_178 ();
 FILLCELL_X4 FILLER_23_197 ();
 FILLCELL_X8 FILLER_23_218 ();
 FILLCELL_X4 FILLER_23_226 ();
 FILLCELL_X1 FILLER_23_230 ();
 FILLCELL_X4 FILLER_23_238 ();
 FILLCELL_X8 FILLER_23_252 ();
 FILLCELL_X1 FILLER_23_260 ();
 FILLCELL_X4 FILLER_23_264 ();
 FILLCELL_X4 FILLER_23_278 ();
 FILLCELL_X8 FILLER_23_285 ();
 FILLCELL_X4 FILLER_23_293 ();
 FILLCELL_X1 FILLER_23_297 ();
 FILLCELL_X4 FILLER_23_301 ();
 FILLCELL_X4 FILLER_23_314 ();
 FILLCELL_X4 FILLER_23_322 ();
 FILLCELL_X8 FILLER_23_329 ();
 FILLCELL_X4 FILLER_23_341 ();
 FILLCELL_X16 FILLER_23_349 ();
 FILLCELL_X8 FILLER_23_365 ();
 FILLCELL_X4 FILLER_23_373 ();
 FILLCELL_X2 FILLER_23_377 ();
 FILLCELL_X1 FILLER_23_379 ();
 FILLCELL_X4 FILLER_23_384 ();
 FILLCELL_X4 FILLER_23_392 ();
 FILLCELL_X4 FILLER_23_400 ();
 FILLCELL_X4 FILLER_23_413 ();
 FILLCELL_X4 FILLER_23_423 ();
 FILLCELL_X1 FILLER_23_427 ();
 FILLCELL_X4 FILLER_23_432 ();
 FILLCELL_X8 FILLER_23_440 ();
 FILLCELL_X4 FILLER_23_448 ();
 FILLCELL_X4 FILLER_23_456 ();
 FILLCELL_X8 FILLER_23_464 ();
 FILLCELL_X2 FILLER_23_472 ();
 FILLCELL_X1 FILLER_23_474 ();
 FILLCELL_X4 FILLER_23_477 ();
 FILLCELL_X4 FILLER_23_484 ();
 FILLCELL_X4 FILLER_23_493 ();
 FILLCELL_X4 FILLER_23_500 ();
 FILLCELL_X2 FILLER_23_504 ();
 FILLCELL_X1 FILLER_23_506 ();
 FILLCELL_X4 FILLER_23_532 ();
 FILLCELL_X1 FILLER_23_536 ();
 FILLCELL_X4 FILLER_23_547 ();
 FILLCELL_X2 FILLER_23_551 ();
 FILLCELL_X4 FILLER_23_556 ();
 FILLCELL_X8 FILLER_23_569 ();
 FILLCELL_X2 FILLER_23_577 ();
 FILLCELL_X1 FILLER_23_579 ();
 FILLCELL_X4 FILLER_23_584 ();
 FILLCELL_X4 FILLER_23_598 ();
 FILLCELL_X4 FILLER_23_604 ();
 FILLCELL_X2 FILLER_23_608 ();
 FILLCELL_X8 FILLER_23_614 ();
 FILLCELL_X1 FILLER_23_622 ();
 FILLCELL_X4 FILLER_23_632 ();
 FILLCELL_X8 FILLER_23_645 ();
 FILLCELL_X1 FILLER_23_653 ();
 FILLCELL_X4 FILLER_23_660 ();
 FILLCELL_X4 FILLER_23_673 ();
 FILLCELL_X4 FILLER_23_683 ();
 FILLCELL_X4 FILLER_23_696 ();
 FILLCELL_X8 FILLER_23_709 ();
 FILLCELL_X1 FILLER_23_717 ();
 FILLCELL_X4 FILLER_23_722 ();
 FILLCELL_X4 FILLER_23_731 ();
 FILLCELL_X4 FILLER_23_752 ();
 FILLCELL_X8 FILLER_23_760 ();
 FILLCELL_X4 FILLER_23_768 ();
 FILLCELL_X2 FILLER_23_772 ();
 FILLCELL_X4 FILLER_23_778 ();
 FILLCELL_X16 FILLER_23_786 ();
 FILLCELL_X8 FILLER_23_802 ();
 FILLCELL_X2 FILLER_23_810 ();
 FILLCELL_X8 FILLER_23_815 ();
 FILLCELL_X4 FILLER_23_823 ();
 FILLCELL_X4 FILLER_23_831 ();
 FILLCELL_X4 FILLER_23_840 ();
 FILLCELL_X8 FILLER_23_847 ();
 FILLCELL_X2 FILLER_23_855 ();
 FILLCELL_X16 FILLER_23_861 ();
 FILLCELL_X8 FILLER_23_881 ();
 FILLCELL_X4 FILLER_23_889 ();
 FILLCELL_X2 FILLER_23_893 ();
 FILLCELL_X4 FILLER_23_904 ();
 FILLCELL_X1 FILLER_23_908 ();
 FILLCELL_X8 FILLER_23_912 ();
 FILLCELL_X8 FILLER_23_924 ();
 FILLCELL_X4 FILLER_23_932 ();
 FILLCELL_X2 FILLER_23_936 ();
 FILLCELL_X8 FILLER_23_941 ();
 FILLCELL_X2 FILLER_23_949 ();
 FILLCELL_X4 FILLER_23_960 ();
 FILLCELL_X4 FILLER_23_971 ();
 FILLCELL_X8 FILLER_23_984 ();
 FILLCELL_X4 FILLER_23_992 ();
 FILLCELL_X2 FILLER_23_996 ();
 FILLCELL_X1 FILLER_23_998 ();
 FILLCELL_X4 FILLER_23_1003 ();
 FILLCELL_X4 FILLER_23_1016 ();
 FILLCELL_X4 FILLER_23_1023 ();
 FILLCELL_X4 FILLER_23_1037 ();
 FILLCELL_X2 FILLER_23_1041 ();
 FILLCELL_X4 FILLER_23_1045 ();
 FILLCELL_X4 FILLER_23_1059 ();
 FILLCELL_X4 FILLER_23_1066 ();
 FILLCELL_X4 FILLER_23_1073 ();
 FILLCELL_X2 FILLER_23_1077 ();
 FILLCELL_X8 FILLER_23_1082 ();
 FILLCELL_X1 FILLER_23_1090 ();
 FILLCELL_X8 FILLER_23_1094 ();
 FILLCELL_X2 FILLER_23_1102 ();
 FILLCELL_X1 FILLER_23_1104 ();
 FILLCELL_X4 FILLER_23_1107 ();
 FILLCELL_X4 FILLER_23_1121 ();
 FILLCELL_X4 FILLER_23_1128 ();
 FILLCELL_X4 FILLER_23_1135 ();
 FILLCELL_X8 FILLER_23_1142 ();
 FILLCELL_X16 FILLER_23_1153 ();
 FILLCELL_X8 FILLER_23_1169 ();
 FILLCELL_X4 FILLER_23_1177 ();
 FILLCELL_X1 FILLER_23_1181 ();
 FILLCELL_X4 FILLER_23_1186 ();
 FILLCELL_X8 FILLER_23_1194 ();
 FILLCELL_X4 FILLER_23_1202 ();
 FILLCELL_X4 FILLER_23_1213 ();
 FILLCELL_X2 FILLER_23_1217 ();
 FILLCELL_X4 FILLER_23_1222 ();
 FILLCELL_X2 FILLER_23_1226 ();
 FILLCELL_X4 FILLER_23_1232 ();
 FILLCELL_X4 FILLER_23_1243 ();
 FILLCELL_X4 FILLER_23_1249 ();
 FILLCELL_X4 FILLER_23_1256 ();
 FILLCELL_X2 FILLER_23_1260 ();
 FILLCELL_X1 FILLER_23_1262 ();
 FILLCELL_X4 FILLER_23_1264 ();
 FILLCELL_X8 FILLER_23_1271 ();
 FILLCELL_X4 FILLER_23_1286 ();
 FILLCELL_X4 FILLER_23_1293 ();
 FILLCELL_X8 FILLER_23_1299 ();
 FILLCELL_X4 FILLER_23_1307 ();
 FILLCELL_X1 FILLER_23_1311 ();
 FILLCELL_X4 FILLER_23_1314 ();
 FILLCELL_X8 FILLER_23_1324 ();
 FILLCELL_X2 FILLER_23_1332 ();
 FILLCELL_X32 FILLER_23_1340 ();
 FILLCELL_X8 FILLER_23_1376 ();
 FILLCELL_X1 FILLER_23_1384 ();
 FILLCELL_X4 FILLER_23_1389 ();
 FILLCELL_X32 FILLER_23_1403 ();
 FILLCELL_X32 FILLER_23_1435 ();
 FILLCELL_X32 FILLER_23_1467 ();
 FILLCELL_X32 FILLER_23_1499 ();
 FILLCELL_X32 FILLER_23_1531 ();
 FILLCELL_X32 FILLER_23_1563 ();
 FILLCELL_X32 FILLER_23_1595 ();
 FILLCELL_X32 FILLER_23_1627 ();
 FILLCELL_X32 FILLER_23_1659 ();
 FILLCELL_X32 FILLER_23_1691 ();
 FILLCELL_X32 FILLER_23_1723 ();
 FILLCELL_X1 FILLER_23_1755 ();
 FILLCELL_X4 FILLER_24_1 ();
 FILLCELL_X2 FILLER_24_5 ();
 FILLCELL_X4 FILLER_24_14 ();
 FILLCELL_X4 FILLER_24_27 ();
 FILLCELL_X8 FILLER_24_40 ();
 FILLCELL_X4 FILLER_24_57 ();
 FILLCELL_X16 FILLER_24_80 ();
 FILLCELL_X4 FILLER_24_100 ();
 FILLCELL_X2 FILLER_24_104 ();
 FILLCELL_X8 FILLER_24_109 ();
 FILLCELL_X2 FILLER_24_117 ();
 FILLCELL_X1 FILLER_24_119 ();
 FILLCELL_X8 FILLER_24_123 ();
 FILLCELL_X16 FILLER_24_134 ();
 FILLCELL_X4 FILLER_24_150 ();
 FILLCELL_X4 FILLER_24_158 ();
 FILLCELL_X4 FILLER_24_168 ();
 FILLCELL_X32 FILLER_24_176 ();
 FILLCELL_X8 FILLER_24_208 ();
 FILLCELL_X1 FILLER_24_216 ();
 FILLCELL_X4 FILLER_24_220 ();
 FILLCELL_X4 FILLER_24_227 ();
 FILLCELL_X1 FILLER_24_231 ();
 FILLCELL_X4 FILLER_24_242 ();
 FILLCELL_X4 FILLER_24_253 ();
 FILLCELL_X4 FILLER_24_259 ();
 FILLCELL_X1 FILLER_24_263 ();
 FILLCELL_X8 FILLER_24_271 ();
 FILLCELL_X1 FILLER_24_279 ();
 FILLCELL_X8 FILLER_24_283 ();
 FILLCELL_X2 FILLER_24_291 ();
 FILLCELL_X8 FILLER_24_296 ();
 FILLCELL_X4 FILLER_24_308 ();
 FILLCELL_X1 FILLER_24_312 ();
 FILLCELL_X4 FILLER_24_317 ();
 FILLCELL_X8 FILLER_24_325 ();
 FILLCELL_X4 FILLER_24_333 ();
 FILLCELL_X2 FILLER_24_337 ();
 FILLCELL_X4 FILLER_24_343 ();
 FILLCELL_X16 FILLER_24_351 ();
 FILLCELL_X4 FILLER_24_373 ();
 FILLCELL_X8 FILLER_24_380 ();
 FILLCELL_X4 FILLER_24_388 ();
 FILLCELL_X2 FILLER_24_392 ();
 FILLCELL_X4 FILLER_24_399 ();
 FILLCELL_X1 FILLER_24_403 ();
 FILLCELL_X4 FILLER_24_413 ();
 FILLCELL_X2 FILLER_24_417 ();
 FILLCELL_X8 FILLER_24_424 ();
 FILLCELL_X2 FILLER_24_432 ();
 FILLCELL_X8 FILLER_24_437 ();
 FILLCELL_X1 FILLER_24_445 ();
 FILLCELL_X4 FILLER_24_450 ();
 FILLCELL_X4 FILLER_24_463 ();
 FILLCELL_X2 FILLER_24_467 ();
 FILLCELL_X1 FILLER_24_469 ();
 FILLCELL_X4 FILLER_24_475 ();
 FILLCELL_X2 FILLER_24_479 ();
 FILLCELL_X1 FILLER_24_481 ();
 FILLCELL_X4 FILLER_24_486 ();
 FILLCELL_X1 FILLER_24_490 ();
 FILLCELL_X4 FILLER_24_494 ();
 FILLCELL_X4 FILLER_24_502 ();
 FILLCELL_X2 FILLER_24_506 ();
 FILLCELL_X8 FILLER_24_512 ();
 FILLCELL_X4 FILLER_24_520 ();
 FILLCELL_X2 FILLER_24_524 ();
 FILLCELL_X1 FILLER_24_526 ();
 FILLCELL_X4 FILLER_24_534 ();
 FILLCELL_X16 FILLER_24_540 ();
 FILLCELL_X1 FILLER_24_556 ();
 FILLCELL_X4 FILLER_24_561 ();
 FILLCELL_X4 FILLER_24_569 ();
 FILLCELL_X8 FILLER_24_577 ();
 FILLCELL_X4 FILLER_24_585 ();
 FILLCELL_X4 FILLER_24_596 ();
 FILLCELL_X2 FILLER_24_600 ();
 FILLCELL_X4 FILLER_24_606 ();
 FILLCELL_X4 FILLER_24_619 ();
 FILLCELL_X4 FILLER_24_626 ();
 FILLCELL_X1 FILLER_24_630 ();
 FILLCELL_X8 FILLER_24_632 ();
 FILLCELL_X2 FILLER_24_640 ();
 FILLCELL_X8 FILLER_24_647 ();
 FILLCELL_X1 FILLER_24_655 ();
 FILLCELL_X4 FILLER_24_659 ();
 FILLCELL_X4 FILLER_24_668 ();
 FILLCELL_X8 FILLER_24_676 ();
 FILLCELL_X1 FILLER_24_684 ();
 FILLCELL_X4 FILLER_24_688 ();
 FILLCELL_X8 FILLER_24_701 ();
 FILLCELL_X2 FILLER_24_709 ();
 FILLCELL_X1 FILLER_24_711 ();
 FILLCELL_X4 FILLER_24_716 ();
 FILLCELL_X4 FILLER_24_724 ();
 FILLCELL_X4 FILLER_24_735 ();
 FILLCELL_X8 FILLER_24_744 ();
 FILLCELL_X16 FILLER_24_761 ();
 FILLCELL_X2 FILLER_24_777 ();
 FILLCELL_X1 FILLER_24_779 ();
 FILLCELL_X4 FILLER_24_786 ();
 FILLCELL_X4 FILLER_24_793 ();
 FILLCELL_X32 FILLER_24_806 ();
 FILLCELL_X8 FILLER_24_838 ();
 FILLCELL_X2 FILLER_24_846 ();
 FILLCELL_X1 FILLER_24_848 ();
 FILLCELL_X4 FILLER_24_854 ();
 FILLCELL_X8 FILLER_24_867 ();
 FILLCELL_X1 FILLER_24_875 ();
 FILLCELL_X4 FILLER_24_880 ();
 FILLCELL_X4 FILLER_24_893 ();
 FILLCELL_X4 FILLER_24_903 ();
 FILLCELL_X4 FILLER_24_911 ();
 FILLCELL_X1 FILLER_24_915 ();
 FILLCELL_X4 FILLER_24_920 ();
 FILLCELL_X8 FILLER_24_929 ();
 FILLCELL_X4 FILLER_24_937 ();
 FILLCELL_X4 FILLER_24_945 ();
 FILLCELL_X8 FILLER_24_952 ();
 FILLCELL_X4 FILLER_24_970 ();
 FILLCELL_X2 FILLER_24_974 ();
 FILLCELL_X4 FILLER_24_986 ();
 FILLCELL_X4 FILLER_24_992 ();
 FILLCELL_X1 FILLER_24_996 ();
 FILLCELL_X4 FILLER_24_1000 ();
 FILLCELL_X16 FILLER_24_1008 ();
 FILLCELL_X16 FILLER_24_1028 ();
 FILLCELL_X8 FILLER_24_1044 ();
 FILLCELL_X4 FILLER_24_1052 ();
 FILLCELL_X4 FILLER_24_1065 ();
 FILLCELL_X8 FILLER_24_1073 ();
 FILLCELL_X4 FILLER_24_1081 ();
 FILLCELL_X4 FILLER_24_1089 ();
 FILLCELL_X8 FILLER_24_1102 ();
 FILLCELL_X1 FILLER_24_1110 ();
 FILLCELL_X8 FILLER_24_1118 ();
 FILLCELL_X4 FILLER_24_1126 ();
 FILLCELL_X1 FILLER_24_1130 ();
 FILLCELL_X8 FILLER_24_1135 ();
 FILLCELL_X4 FILLER_24_1143 ();
 FILLCELL_X4 FILLER_24_1156 ();
 FILLCELL_X4 FILLER_24_1164 ();
 FILLCELL_X16 FILLER_24_1172 ();
 FILLCELL_X2 FILLER_24_1188 ();
 FILLCELL_X1 FILLER_24_1190 ();
 FILLCELL_X4 FILLER_24_1194 ();
 FILLCELL_X4 FILLER_24_1208 ();
 FILLCELL_X4 FILLER_24_1222 ();
 FILLCELL_X4 FILLER_24_1236 ();
 FILLCELL_X8 FILLER_24_1250 ();
 FILLCELL_X4 FILLER_24_1267 ();
 FILLCELL_X4 FILLER_24_1278 ();
 FILLCELL_X2 FILLER_24_1282 ();
 FILLCELL_X4 FILLER_24_1294 ();
 FILLCELL_X4 FILLER_24_1302 ();
 FILLCELL_X16 FILLER_24_1309 ();
 FILLCELL_X4 FILLER_24_1329 ();
 FILLCELL_X16 FILLER_24_1346 ();
 FILLCELL_X2 FILLER_24_1362 ();
 FILLCELL_X1 FILLER_24_1364 ();
 FILLCELL_X8 FILLER_24_1369 ();
 FILLCELL_X1 FILLER_24_1377 ();
 FILLCELL_X4 FILLER_24_1383 ();
 FILLCELL_X2 FILLER_24_1387 ();
 FILLCELL_X4 FILLER_24_1393 ();
 FILLCELL_X2 FILLER_24_1397 ();
 FILLCELL_X1 FILLER_24_1399 ();
 FILLCELL_X32 FILLER_24_1419 ();
 FILLCELL_X32 FILLER_24_1451 ();
 FILLCELL_X32 FILLER_24_1483 ();
 FILLCELL_X32 FILLER_24_1515 ();
 FILLCELL_X32 FILLER_24_1547 ();
 FILLCELL_X32 FILLER_24_1579 ();
 FILLCELL_X32 FILLER_24_1611 ();
 FILLCELL_X32 FILLER_24_1643 ();
 FILLCELL_X32 FILLER_24_1675 ();
 FILLCELL_X32 FILLER_24_1707 ();
 FILLCELL_X16 FILLER_24_1739 ();
 FILLCELL_X1 FILLER_24_1755 ();
 FILLCELL_X4 FILLER_25_1 ();
 FILLCELL_X2 FILLER_25_5 ();
 FILLCELL_X4 FILLER_25_17 ();
 FILLCELL_X4 FILLER_25_24 ();
 FILLCELL_X4 FILLER_25_31 ();
 FILLCELL_X2 FILLER_25_35 ();
 FILLCELL_X1 FILLER_25_37 ();
 FILLCELL_X4 FILLER_25_48 ();
 FILLCELL_X2 FILLER_25_52 ();
 FILLCELL_X1 FILLER_25_54 ();
 FILLCELL_X16 FILLER_25_59 ();
 FILLCELL_X4 FILLER_25_77 ();
 FILLCELL_X4 FILLER_25_91 ();
 FILLCELL_X1 FILLER_25_95 ();
 FILLCELL_X4 FILLER_25_105 ();
 FILLCELL_X4 FILLER_25_113 ();
 FILLCELL_X2 FILLER_25_117 ();
 FILLCELL_X1 FILLER_25_119 ();
 FILLCELL_X4 FILLER_25_129 ();
 FILLCELL_X2 FILLER_25_133 ();
 FILLCELL_X1 FILLER_25_135 ();
 FILLCELL_X4 FILLER_25_146 ();
 FILLCELL_X2 FILLER_25_150 ();
 FILLCELL_X1 FILLER_25_152 ();
 FILLCELL_X4 FILLER_25_158 ();
 FILLCELL_X4 FILLER_25_165 ();
 FILLCELL_X1 FILLER_25_169 ();
 FILLCELL_X4 FILLER_25_176 ();
 FILLCELL_X4 FILLER_25_182 ();
 FILLCELL_X8 FILLER_25_193 ();
 FILLCELL_X4 FILLER_25_201 ();
 FILLCELL_X2 FILLER_25_205 ();
 FILLCELL_X4 FILLER_25_216 ();
 FILLCELL_X8 FILLER_25_230 ();
 FILLCELL_X1 FILLER_25_238 ();
 FILLCELL_X4 FILLER_25_243 ();
 FILLCELL_X4 FILLER_25_257 ();
 FILLCELL_X2 FILLER_25_261 ();
 FILLCELL_X1 FILLER_25_263 ();
 FILLCELL_X4 FILLER_25_273 ();
 FILLCELL_X4 FILLER_25_280 ();
 FILLCELL_X4 FILLER_25_288 ();
 FILLCELL_X8 FILLER_25_302 ();
 FILLCELL_X8 FILLER_25_319 ();
 FILLCELL_X4 FILLER_25_331 ();
 FILLCELL_X2 FILLER_25_335 ();
 FILLCELL_X4 FILLER_25_346 ();
 FILLCELL_X4 FILLER_25_359 ();
 FILLCELL_X4 FILLER_25_372 ();
 FILLCELL_X16 FILLER_25_385 ();
 FILLCELL_X8 FILLER_25_405 ();
 FILLCELL_X1 FILLER_25_413 ();
 FILLCELL_X4 FILLER_25_417 ();
 FILLCELL_X4 FILLER_25_426 ();
 FILLCELL_X4 FILLER_25_434 ();
 FILLCELL_X1 FILLER_25_438 ();
 FILLCELL_X4 FILLER_25_443 ();
 FILLCELL_X2 FILLER_25_447 ();
 FILLCELL_X1 FILLER_25_449 ();
 FILLCELL_X4 FILLER_25_455 ();
 FILLCELL_X8 FILLER_25_468 ();
 FILLCELL_X4 FILLER_25_480 ();
 FILLCELL_X4 FILLER_25_493 ();
 FILLCELL_X4 FILLER_25_506 ();
 FILLCELL_X16 FILLER_25_520 ();
 FILLCELL_X2 FILLER_25_536 ();
 FILLCELL_X4 FILLER_25_543 ();
 FILLCELL_X4 FILLER_25_551 ();
 FILLCELL_X4 FILLER_25_557 ();
 FILLCELL_X1 FILLER_25_561 ();
 FILLCELL_X4 FILLER_25_565 ();
 FILLCELL_X4 FILLER_25_572 ();
 FILLCELL_X4 FILLER_25_579 ();
 FILLCELL_X16 FILLER_25_592 ();
 FILLCELL_X2 FILLER_25_608 ();
 FILLCELL_X1 FILLER_25_610 ();
 FILLCELL_X8 FILLER_25_614 ();
 FILLCELL_X4 FILLER_25_622 ();
 FILLCELL_X2 FILLER_25_626 ();
 FILLCELL_X4 FILLER_25_631 ();
 FILLCELL_X16 FILLER_25_640 ();
 FILLCELL_X4 FILLER_25_656 ();
 FILLCELL_X2 FILLER_25_660 ();
 FILLCELL_X16 FILLER_25_666 ();
 FILLCELL_X4 FILLER_25_682 ();
 FILLCELL_X8 FILLER_25_691 ();
 FILLCELL_X4 FILLER_25_699 ();
 FILLCELL_X4 FILLER_25_707 ();
 FILLCELL_X4 FILLER_25_715 ();
 FILLCELL_X16 FILLER_25_723 ();
 FILLCELL_X4 FILLER_25_739 ();
 FILLCELL_X1 FILLER_25_743 ();
 FILLCELL_X4 FILLER_25_748 ();
 FILLCELL_X4 FILLER_25_756 ();
 FILLCELL_X16 FILLER_25_764 ();
 FILLCELL_X4 FILLER_25_789 ();
 FILLCELL_X4 FILLER_25_798 ();
 FILLCELL_X4 FILLER_25_806 ();
 FILLCELL_X8 FILLER_25_813 ();
 FILLCELL_X2 FILLER_25_821 ();
 FILLCELL_X8 FILLER_25_829 ();
 FILLCELL_X4 FILLER_25_837 ();
 FILLCELL_X1 FILLER_25_841 ();
 FILLCELL_X4 FILLER_25_848 ();
 FILLCELL_X4 FILLER_25_861 ();
 FILLCELL_X8 FILLER_25_870 ();
 FILLCELL_X4 FILLER_25_878 ();
 FILLCELL_X1 FILLER_25_882 ();
 FILLCELL_X4 FILLER_25_886 ();
 FILLCELL_X4 FILLER_25_895 ();
 FILLCELL_X2 FILLER_25_899 ();
 FILLCELL_X1 FILLER_25_901 ();
 FILLCELL_X4 FILLER_25_905 ();
 FILLCELL_X4 FILLER_25_915 ();
 FILLCELL_X8 FILLER_25_928 ();
 FILLCELL_X4 FILLER_25_945 ();
 FILLCELL_X4 FILLER_25_953 ();
 FILLCELL_X4 FILLER_25_961 ();
 FILLCELL_X16 FILLER_25_968 ();
 FILLCELL_X4 FILLER_25_984 ();
 FILLCELL_X4 FILLER_25_992 ();
 FILLCELL_X4 FILLER_25_1000 ();
 FILLCELL_X2 FILLER_25_1004 ();
 FILLCELL_X4 FILLER_25_1015 ();
 FILLCELL_X4 FILLER_25_1023 ();
 FILLCELL_X4 FILLER_25_1030 ();
 FILLCELL_X4 FILLER_25_1041 ();
 FILLCELL_X4 FILLER_25_1048 ();
 FILLCELL_X4 FILLER_25_1055 ();
 FILLCELL_X4 FILLER_25_1062 ();
 FILLCELL_X1 FILLER_25_1066 ();
 FILLCELL_X4 FILLER_25_1071 ();
 FILLCELL_X2 FILLER_25_1075 ();
 FILLCELL_X4 FILLER_25_1086 ();
 FILLCELL_X4 FILLER_25_1093 ();
 FILLCELL_X8 FILLER_25_1100 ();
 FILLCELL_X2 FILLER_25_1108 ();
 FILLCELL_X1 FILLER_25_1110 ();
 FILLCELL_X4 FILLER_25_1114 ();
 FILLCELL_X4 FILLER_25_1127 ();
 FILLCELL_X4 FILLER_25_1133 ();
 FILLCELL_X2 FILLER_25_1137 ();
 FILLCELL_X4 FILLER_25_1142 ();
 FILLCELL_X4 FILLER_25_1155 ();
 FILLCELL_X4 FILLER_25_1168 ();
 FILLCELL_X4 FILLER_25_1175 ();
 FILLCELL_X4 FILLER_25_1189 ();
 FILLCELL_X4 FILLER_25_1197 ();
 FILLCELL_X4 FILLER_25_1203 ();
 FILLCELL_X8 FILLER_25_1209 ();
 FILLCELL_X4 FILLER_25_1217 ();
 FILLCELL_X4 FILLER_25_1223 ();
 FILLCELL_X8 FILLER_25_1229 ();
 FILLCELL_X1 FILLER_25_1237 ();
 FILLCELL_X4 FILLER_25_1248 ();
 FILLCELL_X8 FILLER_25_1254 ();
 FILLCELL_X1 FILLER_25_1262 ();
 FILLCELL_X4 FILLER_25_1264 ();
 FILLCELL_X4 FILLER_25_1278 ();
 FILLCELL_X2 FILLER_25_1282 ();
 FILLCELL_X1 FILLER_25_1284 ();
 FILLCELL_X4 FILLER_25_1295 ();
 FILLCELL_X4 FILLER_25_1309 ();
 FILLCELL_X8 FILLER_25_1322 ();
 FILLCELL_X2 FILLER_25_1330 ();
 FILLCELL_X4 FILLER_25_1336 ();
 FILLCELL_X8 FILLER_25_1346 ();
 FILLCELL_X4 FILLER_25_1358 ();
 FILLCELL_X4 FILLER_25_1367 ();
 FILLCELL_X4 FILLER_25_1378 ();
 FILLCELL_X4 FILLER_25_1399 ();
 FILLCELL_X32 FILLER_25_1407 ();
 FILLCELL_X32 FILLER_25_1439 ();
 FILLCELL_X32 FILLER_25_1471 ();
 FILLCELL_X32 FILLER_25_1503 ();
 FILLCELL_X32 FILLER_25_1535 ();
 FILLCELL_X32 FILLER_25_1567 ();
 FILLCELL_X32 FILLER_25_1599 ();
 FILLCELL_X32 FILLER_25_1631 ();
 FILLCELL_X32 FILLER_25_1663 ();
 FILLCELL_X32 FILLER_25_1695 ();
 FILLCELL_X16 FILLER_25_1727 ();
 FILLCELL_X8 FILLER_25_1743 ();
 FILLCELL_X4 FILLER_25_1751 ();
 FILLCELL_X1 FILLER_25_1755 ();
 FILLCELL_X8 FILLER_26_1 ();
 FILLCELL_X1 FILLER_26_9 ();
 FILLCELL_X4 FILLER_26_14 ();
 FILLCELL_X8 FILLER_26_21 ();
 FILLCELL_X4 FILLER_26_29 ();
 FILLCELL_X2 FILLER_26_33 ();
 FILLCELL_X8 FILLER_26_37 ();
 FILLCELL_X2 FILLER_26_45 ();
 FILLCELL_X4 FILLER_26_51 ();
 FILLCELL_X4 FILLER_26_59 ();
 FILLCELL_X8 FILLER_26_66 ();
 FILLCELL_X2 FILLER_26_74 ();
 FILLCELL_X1 FILLER_26_76 ();
 FILLCELL_X4 FILLER_26_87 ();
 FILLCELL_X4 FILLER_26_98 ();
 FILLCELL_X2 FILLER_26_102 ();
 FILLCELL_X4 FILLER_26_113 ();
 FILLCELL_X8 FILLER_26_121 ();
 FILLCELL_X2 FILLER_26_129 ();
 FILLCELL_X4 FILLER_26_134 ();
 FILLCELL_X4 FILLER_26_148 ();
 FILLCELL_X4 FILLER_26_156 ();
 FILLCELL_X4 FILLER_26_169 ();
 FILLCELL_X4 FILLER_26_176 ();
 FILLCELL_X4 FILLER_26_183 ();
 FILLCELL_X4 FILLER_26_197 ();
 FILLCELL_X2 FILLER_26_201 ();
 FILLCELL_X4 FILLER_26_206 ();
 FILLCELL_X2 FILLER_26_210 ();
 FILLCELL_X16 FILLER_26_215 ();
 FILLCELL_X1 FILLER_26_231 ();
 FILLCELL_X4 FILLER_26_234 ();
 FILLCELL_X16 FILLER_26_241 ();
 FILLCELL_X2 FILLER_26_257 ();
 FILLCELL_X4 FILLER_26_262 ();
 FILLCELL_X4 FILLER_26_269 ();
 FILLCELL_X4 FILLER_26_282 ();
 FILLCELL_X8 FILLER_26_293 ();
 FILLCELL_X4 FILLER_26_305 ();
 FILLCELL_X4 FILLER_26_318 ();
 FILLCELL_X4 FILLER_26_331 ();
 FILLCELL_X8 FILLER_26_340 ();
 FILLCELL_X1 FILLER_26_348 ();
 FILLCELL_X4 FILLER_26_353 ();
 FILLCELL_X4 FILLER_26_361 ();
 FILLCELL_X1 FILLER_26_365 ();
 FILLCELL_X8 FILLER_26_371 ();
 FILLCELL_X8 FILLER_26_384 ();
 FILLCELL_X1 FILLER_26_392 ();
 FILLCELL_X4 FILLER_26_399 ();
 FILLCELL_X8 FILLER_26_406 ();
 FILLCELL_X4 FILLER_26_414 ();
 FILLCELL_X4 FILLER_26_424 ();
 FILLCELL_X8 FILLER_26_437 ();
 FILLCELL_X2 FILLER_26_445 ();
 FILLCELL_X4 FILLER_26_453 ();
 FILLCELL_X4 FILLER_26_466 ();
 FILLCELL_X8 FILLER_26_473 ();
 FILLCELL_X2 FILLER_26_481 ();
 FILLCELL_X1 FILLER_26_483 ();
 FILLCELL_X16 FILLER_26_487 ();
 FILLCELL_X8 FILLER_26_503 ();
 FILLCELL_X1 FILLER_26_511 ();
 FILLCELL_X16 FILLER_26_515 ();
 FILLCELL_X4 FILLER_26_538 ();
 FILLCELL_X8 FILLER_26_559 ();
 FILLCELL_X8 FILLER_26_576 ();
 FILLCELL_X1 FILLER_26_584 ();
 FILLCELL_X4 FILLER_26_589 ();
 FILLCELL_X16 FILLER_26_597 ();
 FILLCELL_X4 FILLER_26_616 ();
 FILLCELL_X4 FILLER_26_626 ();
 FILLCELL_X1 FILLER_26_630 ();
 FILLCELL_X4 FILLER_26_632 ();
 FILLCELL_X4 FILLER_26_641 ();
 FILLCELL_X2 FILLER_26_645 ();
 FILLCELL_X1 FILLER_26_647 ();
 FILLCELL_X4 FILLER_26_652 ();
 FILLCELL_X4 FILLER_26_662 ();
 FILLCELL_X2 FILLER_26_666 ();
 FILLCELL_X8 FILLER_26_677 ();
 FILLCELL_X2 FILLER_26_685 ();
 FILLCELL_X1 FILLER_26_687 ();
 FILLCELL_X4 FILLER_26_692 ();
 FILLCELL_X4 FILLER_26_700 ();
 FILLCELL_X2 FILLER_26_704 ();
 FILLCELL_X1 FILLER_26_706 ();
 FILLCELL_X4 FILLER_26_712 ();
 FILLCELL_X1 FILLER_26_716 ();
 FILLCELL_X4 FILLER_26_722 ();
 FILLCELL_X2 FILLER_26_726 ();
 FILLCELL_X4 FILLER_26_734 ();
 FILLCELL_X2 FILLER_26_738 ();
 FILLCELL_X1 FILLER_26_740 ();
 FILLCELL_X16 FILLER_26_745 ();
 FILLCELL_X8 FILLER_26_761 ();
 FILLCELL_X8 FILLER_26_773 ();
 FILLCELL_X8 FILLER_26_786 ();
 FILLCELL_X4 FILLER_26_797 ();
 FILLCELL_X2 FILLER_26_801 ();
 FILLCELL_X4 FILLER_26_807 ();
 FILLCELL_X4 FILLER_26_820 ();
 FILLCELL_X4 FILLER_26_833 ();
 FILLCELL_X8 FILLER_26_840 ();
 FILLCELL_X2 FILLER_26_848 ();
 FILLCELL_X1 FILLER_26_850 ();
 FILLCELL_X4 FILLER_26_855 ();
 FILLCELL_X2 FILLER_26_859 ();
 FILLCELL_X1 FILLER_26_861 ();
 FILLCELL_X8 FILLER_26_865 ();
 FILLCELL_X1 FILLER_26_873 ();
 FILLCELL_X8 FILLER_26_883 ();
 FILLCELL_X4 FILLER_26_891 ();
 FILLCELL_X2 FILLER_26_895 ();
 FILLCELL_X1 FILLER_26_897 ();
 FILLCELL_X16 FILLER_26_901 ();
 FILLCELL_X1 FILLER_26_917 ();
 FILLCELL_X4 FILLER_26_923 ();
 FILLCELL_X2 FILLER_26_927 ();
 FILLCELL_X1 FILLER_26_929 ();
 FILLCELL_X16 FILLER_26_934 ();
 FILLCELL_X4 FILLER_26_950 ();
 FILLCELL_X1 FILLER_26_954 ();
 FILLCELL_X4 FILLER_26_964 ();
 FILLCELL_X8 FILLER_26_985 ();
 FILLCELL_X1 FILLER_26_993 ();
 FILLCELL_X4 FILLER_26_1003 ();
 FILLCELL_X4 FILLER_26_1010 ();
 FILLCELL_X2 FILLER_26_1014 ();
 FILLCELL_X1 FILLER_26_1016 ();
 FILLCELL_X4 FILLER_26_1027 ();
 FILLCELL_X4 FILLER_26_1033 ();
 FILLCELL_X4 FILLER_26_1047 ();
 FILLCELL_X4 FILLER_26_1060 ();
 FILLCELL_X4 FILLER_26_1067 ();
 FILLCELL_X8 FILLER_26_1074 ();
 FILLCELL_X4 FILLER_26_1082 ();
 FILLCELL_X1 FILLER_26_1086 ();
 FILLCELL_X8 FILLER_26_1090 ();
 FILLCELL_X1 FILLER_26_1098 ();
 FILLCELL_X4 FILLER_26_1106 ();
 FILLCELL_X2 FILLER_26_1110 ();
 FILLCELL_X1 FILLER_26_1112 ();
 FILLCELL_X4 FILLER_26_1117 ();
 FILLCELL_X4 FILLER_26_1128 ();
 FILLCELL_X4 FILLER_26_1142 ();
 FILLCELL_X1 FILLER_26_1146 ();
 FILLCELL_X4 FILLER_26_1150 ();
 FILLCELL_X4 FILLER_26_1158 ();
 FILLCELL_X2 FILLER_26_1162 ();
 FILLCELL_X4 FILLER_26_1167 ();
 FILLCELL_X4 FILLER_26_1174 ();
 FILLCELL_X1 FILLER_26_1178 ();
 FILLCELL_X32 FILLER_26_1188 ();
 FILLCELL_X4 FILLER_26_1220 ();
 FILLCELL_X1 FILLER_26_1224 ();
 FILLCELL_X4 FILLER_26_1227 ();
 FILLCELL_X4 FILLER_26_1234 ();
 FILLCELL_X8 FILLER_26_1241 ();
 FILLCELL_X1 FILLER_26_1249 ();
 FILLCELL_X4 FILLER_26_1253 ();
 FILLCELL_X2 FILLER_26_1257 ();
 FILLCELL_X1 FILLER_26_1259 ();
 FILLCELL_X4 FILLER_26_1267 ();
 FILLCELL_X2 FILLER_26_1271 ();
 FILLCELL_X1 FILLER_26_1273 ();
 FILLCELL_X4 FILLER_26_1284 ();
 FILLCELL_X4 FILLER_26_1291 ();
 FILLCELL_X4 FILLER_26_1297 ();
 FILLCELL_X4 FILLER_26_1303 ();
 FILLCELL_X4 FILLER_26_1310 ();
 FILLCELL_X4 FILLER_26_1323 ();
 FILLCELL_X4 FILLER_26_1330 ();
 FILLCELL_X8 FILLER_26_1336 ();
 FILLCELL_X4 FILLER_26_1344 ();
 FILLCELL_X1 FILLER_26_1348 ();
 FILLCELL_X16 FILLER_26_1353 ();
 FILLCELL_X8 FILLER_26_1369 ();
 FILLCELL_X2 FILLER_26_1377 ();
 FILLCELL_X1 FILLER_26_1379 ();
 FILLCELL_X8 FILLER_26_1382 ();
 FILLCELL_X4 FILLER_26_1390 ();
 FILLCELL_X1 FILLER_26_1394 ();
 FILLCELL_X32 FILLER_26_1398 ();
 FILLCELL_X32 FILLER_26_1430 ();
 FILLCELL_X32 FILLER_26_1462 ();
 FILLCELL_X32 FILLER_26_1494 ();
 FILLCELL_X32 FILLER_26_1526 ();
 FILLCELL_X32 FILLER_26_1558 ();
 FILLCELL_X32 FILLER_26_1590 ();
 FILLCELL_X32 FILLER_26_1622 ();
 FILLCELL_X32 FILLER_26_1654 ();
 FILLCELL_X32 FILLER_26_1686 ();
 FILLCELL_X32 FILLER_26_1718 ();
 FILLCELL_X4 FILLER_26_1750 ();
 FILLCELL_X2 FILLER_26_1754 ();
 FILLCELL_X4 FILLER_27_1 ();
 FILLCELL_X8 FILLER_27_8 ();
 FILLCELL_X2 FILLER_27_16 ();
 FILLCELL_X1 FILLER_27_18 ();
 FILLCELL_X8 FILLER_27_23 ();
 FILLCELL_X4 FILLER_27_31 ();
 FILLCELL_X2 FILLER_27_35 ();
 FILLCELL_X8 FILLER_27_44 ();
 FILLCELL_X1 FILLER_27_52 ();
 FILLCELL_X4 FILLER_27_62 ();
 FILLCELL_X8 FILLER_27_69 ();
 FILLCELL_X2 FILLER_27_77 ();
 FILLCELL_X1 FILLER_27_79 ();
 FILLCELL_X8 FILLER_27_83 ();
 FILLCELL_X4 FILLER_27_91 ();
 FILLCELL_X2 FILLER_27_95 ();
 FILLCELL_X1 FILLER_27_97 ();
 FILLCELL_X4 FILLER_27_101 ();
 FILLCELL_X4 FILLER_27_108 ();
 FILLCELL_X8 FILLER_27_115 ();
 FILLCELL_X1 FILLER_27_123 ();
 FILLCELL_X8 FILLER_27_127 ();
 FILLCELL_X2 FILLER_27_135 ();
 FILLCELL_X4 FILLER_27_139 ();
 FILLCELL_X8 FILLER_27_152 ();
 FILLCELL_X2 FILLER_27_160 ();
 FILLCELL_X4 FILLER_27_165 ();
 FILLCELL_X4 FILLER_27_179 ();
 FILLCELL_X4 FILLER_27_185 ();
 FILLCELL_X1 FILLER_27_189 ();
 FILLCELL_X4 FILLER_27_199 ();
 FILLCELL_X4 FILLER_27_213 ();
 FILLCELL_X8 FILLER_27_227 ();
 FILLCELL_X4 FILLER_27_244 ();
 FILLCELL_X8 FILLER_27_251 ();
 FILLCELL_X1 FILLER_27_259 ();
 FILLCELL_X4 FILLER_27_264 ();
 FILLCELL_X2 FILLER_27_268 ();
 FILLCELL_X1 FILLER_27_270 ();
 FILLCELL_X4 FILLER_27_281 ();
 FILLCELL_X32 FILLER_27_287 ();
 FILLCELL_X2 FILLER_27_319 ();
 FILLCELL_X4 FILLER_27_327 ();
 FILLCELL_X8 FILLER_27_334 ();
 FILLCELL_X2 FILLER_27_342 ();
 FILLCELL_X4 FILLER_27_348 ();
 FILLCELL_X4 FILLER_27_356 ();
 FILLCELL_X2 FILLER_27_360 ();
 FILLCELL_X4 FILLER_27_365 ();
 FILLCELL_X4 FILLER_27_373 ();
 FILLCELL_X4 FILLER_27_386 ();
 FILLCELL_X4 FILLER_27_399 ();
 FILLCELL_X4 FILLER_27_412 ();
 FILLCELL_X8 FILLER_27_421 ();
 FILLCELL_X1 FILLER_27_429 ();
 FILLCELL_X4 FILLER_27_439 ();
 FILLCELL_X8 FILLER_27_448 ();
 FILLCELL_X4 FILLER_27_460 ();
 FILLCELL_X1 FILLER_27_464 ();
 FILLCELL_X8 FILLER_27_469 ();
 FILLCELL_X2 FILLER_27_477 ();
 FILLCELL_X1 FILLER_27_479 ();
 FILLCELL_X32 FILLER_27_484 ();
 FILLCELL_X8 FILLER_27_516 ();
 FILLCELL_X4 FILLER_27_524 ();
 FILLCELL_X1 FILLER_27_528 ();
 FILLCELL_X4 FILLER_27_533 ();
 FILLCELL_X4 FILLER_27_542 ();
 FILLCELL_X8 FILLER_27_550 ();
 FILLCELL_X4 FILLER_27_558 ();
 FILLCELL_X4 FILLER_27_566 ();
 FILLCELL_X8 FILLER_27_574 ();
 FILLCELL_X2 FILLER_27_582 ();
 FILLCELL_X4 FILLER_27_603 ();
 FILLCELL_X4 FILLER_27_613 ();
 FILLCELL_X2 FILLER_27_617 ();
 FILLCELL_X1 FILLER_27_619 ();
 FILLCELL_X4 FILLER_27_629 ();
 FILLCELL_X2 FILLER_27_633 ();
 FILLCELL_X1 FILLER_27_635 ();
 FILLCELL_X8 FILLER_27_645 ();
 FILLCELL_X4 FILLER_27_662 ();
 FILLCELL_X4 FILLER_27_675 ();
 FILLCELL_X8 FILLER_27_684 ();
 FILLCELL_X4 FILLER_27_696 ();
 FILLCELL_X8 FILLER_27_709 ();
 FILLCELL_X8 FILLER_27_726 ();
 FILLCELL_X2 FILLER_27_734 ();
 FILLCELL_X4 FILLER_27_745 ();
 FILLCELL_X4 FILLER_27_758 ();
 FILLCELL_X4 FILLER_27_771 ();
 FILLCELL_X4 FILLER_27_779 ();
 FILLCELL_X4 FILLER_27_787 ();
 FILLCELL_X2 FILLER_27_791 ();
 FILLCELL_X4 FILLER_27_797 ();
 FILLCELL_X4 FILLER_27_805 ();
 FILLCELL_X4 FILLER_27_813 ();
 FILLCELL_X1 FILLER_27_817 ();
 FILLCELL_X4 FILLER_27_823 ();
 FILLCELL_X4 FILLER_27_831 ();
 FILLCELL_X8 FILLER_27_838 ();
 FILLCELL_X4 FILLER_27_846 ();
 FILLCELL_X4 FILLER_27_855 ();
 FILLCELL_X4 FILLER_27_862 ();
 FILLCELL_X4 FILLER_27_870 ();
 FILLCELL_X4 FILLER_27_883 ();
 FILLCELL_X2 FILLER_27_887 ();
 FILLCELL_X1 FILLER_27_889 ();
 FILLCELL_X4 FILLER_27_899 ();
 FILLCELL_X16 FILLER_27_907 ();
 FILLCELL_X2 FILLER_27_923 ();
 FILLCELL_X4 FILLER_27_928 ();
 FILLCELL_X1 FILLER_27_932 ();
 FILLCELL_X8 FILLER_27_936 ();
 FILLCELL_X4 FILLER_27_944 ();
 FILLCELL_X8 FILLER_27_952 ();
 FILLCELL_X4 FILLER_27_960 ();
 FILLCELL_X2 FILLER_27_964 ();
 FILLCELL_X1 FILLER_27_966 ();
 FILLCELL_X4 FILLER_27_974 ();
 FILLCELL_X8 FILLER_27_980 ();
 FILLCELL_X1 FILLER_27_988 ();
 FILLCELL_X4 FILLER_27_992 ();
 FILLCELL_X4 FILLER_27_999 ();
 FILLCELL_X2 FILLER_27_1003 ();
 FILLCELL_X1 FILLER_27_1005 ();
 FILLCELL_X4 FILLER_27_1010 ();
 FILLCELL_X8 FILLER_27_1018 ();
 FILLCELL_X4 FILLER_27_1026 ();
 FILLCELL_X1 FILLER_27_1030 ();
 FILLCELL_X8 FILLER_27_1033 ();
 FILLCELL_X2 FILLER_27_1041 ();
 FILLCELL_X1 FILLER_27_1043 ();
 FILLCELL_X4 FILLER_27_1047 ();
 FILLCELL_X4 FILLER_27_1054 ();
 FILLCELL_X2 FILLER_27_1058 ();
 FILLCELL_X1 FILLER_27_1060 ();
 FILLCELL_X4 FILLER_27_1065 ();
 FILLCELL_X2 FILLER_27_1069 ();
 FILLCELL_X4 FILLER_27_1075 ();
 FILLCELL_X8 FILLER_27_1082 ();
 FILLCELL_X2 FILLER_27_1090 ();
 FILLCELL_X4 FILLER_27_1102 ();
 FILLCELL_X4 FILLER_27_1116 ();
 FILLCELL_X1 FILLER_27_1120 ();
 FILLCELL_X4 FILLER_27_1131 ();
 FILLCELL_X2 FILLER_27_1135 ();
 FILLCELL_X4 FILLER_27_1141 ();
 FILLCELL_X8 FILLER_27_1148 ();
 FILLCELL_X4 FILLER_27_1156 ();
 FILLCELL_X4 FILLER_27_1162 ();
 FILLCELL_X4 FILLER_27_1169 ();
 FILLCELL_X2 FILLER_27_1173 ();
 FILLCELL_X1 FILLER_27_1175 ();
 FILLCELL_X8 FILLER_27_1185 ();
 FILLCELL_X4 FILLER_27_1193 ();
 FILLCELL_X2 FILLER_27_1197 ();
 FILLCELL_X4 FILLER_27_1204 ();
 FILLCELL_X4 FILLER_27_1210 ();
 FILLCELL_X2 FILLER_27_1214 ();
 FILLCELL_X4 FILLER_27_1219 ();
 FILLCELL_X4 FILLER_27_1232 ();
 FILLCELL_X4 FILLER_27_1245 ();
 FILLCELL_X4 FILLER_27_1259 ();
 FILLCELL_X8 FILLER_27_1264 ();
 FILLCELL_X1 FILLER_27_1272 ();
 FILLCELL_X4 FILLER_27_1283 ();
 FILLCELL_X1 FILLER_27_1287 ();
 FILLCELL_X8 FILLER_27_1291 ();
 FILLCELL_X2 FILLER_27_1299 ();
 FILLCELL_X1 FILLER_27_1301 ();
 FILLCELL_X4 FILLER_27_1305 ();
 FILLCELL_X2 FILLER_27_1309 ();
 FILLCELL_X1 FILLER_27_1311 ();
 FILLCELL_X4 FILLER_27_1314 ();
 FILLCELL_X1 FILLER_27_1318 ();
 FILLCELL_X4 FILLER_27_1322 ();
 FILLCELL_X4 FILLER_27_1336 ();
 FILLCELL_X4 FILLER_27_1344 ();
 FILLCELL_X2 FILLER_27_1348 ();
 FILLCELL_X1 FILLER_27_1350 ();
 FILLCELL_X8 FILLER_27_1370 ();
 FILLCELL_X4 FILLER_27_1378 ();
 FILLCELL_X2 FILLER_27_1382 ();
 FILLCELL_X1 FILLER_27_1384 ();
 FILLCELL_X4 FILLER_27_1389 ();
 FILLCELL_X32 FILLER_27_1397 ();
 FILLCELL_X32 FILLER_27_1429 ();
 FILLCELL_X32 FILLER_27_1461 ();
 FILLCELL_X32 FILLER_27_1493 ();
 FILLCELL_X32 FILLER_27_1525 ();
 FILLCELL_X32 FILLER_27_1557 ();
 FILLCELL_X32 FILLER_27_1589 ();
 FILLCELL_X32 FILLER_27_1621 ();
 FILLCELL_X32 FILLER_27_1653 ();
 FILLCELL_X32 FILLER_27_1685 ();
 FILLCELL_X32 FILLER_27_1717 ();
 FILLCELL_X4 FILLER_27_1749 ();
 FILLCELL_X2 FILLER_27_1753 ();
 FILLCELL_X1 FILLER_27_1755 ();
 FILLCELL_X4 FILLER_28_1 ();
 FILLCELL_X2 FILLER_28_5 ();
 FILLCELL_X1 FILLER_28_7 ();
 FILLCELL_X4 FILLER_28_17 ();
 FILLCELL_X2 FILLER_28_21 ();
 FILLCELL_X1 FILLER_28_23 ();
 FILLCELL_X4 FILLER_28_28 ();
 FILLCELL_X4 FILLER_28_42 ();
 FILLCELL_X8 FILLER_28_49 ();
 FILLCELL_X8 FILLER_28_60 ();
 FILLCELL_X4 FILLER_28_68 ();
 FILLCELL_X2 FILLER_28_72 ();
 FILLCELL_X1 FILLER_28_74 ();
 FILLCELL_X4 FILLER_28_77 ();
 FILLCELL_X16 FILLER_28_91 ();
 FILLCELL_X2 FILLER_28_107 ();
 FILLCELL_X16 FILLER_28_118 ();
 FILLCELL_X1 FILLER_28_134 ();
 FILLCELL_X16 FILLER_28_137 ();
 FILLCELL_X2 FILLER_28_153 ();
 FILLCELL_X1 FILLER_28_155 ();
 FILLCELL_X16 FILLER_28_166 ();
 FILLCELL_X4 FILLER_28_182 ();
 FILLCELL_X1 FILLER_28_186 ();
 FILLCELL_X32 FILLER_28_191 ();
 FILLCELL_X8 FILLER_28_223 ();
 FILLCELL_X4 FILLER_28_231 ();
 FILLCELL_X2 FILLER_28_235 ();
 FILLCELL_X4 FILLER_28_246 ();
 FILLCELL_X4 FILLER_28_253 ();
 FILLCELL_X4 FILLER_28_266 ();
 FILLCELL_X8 FILLER_28_274 ();
 FILLCELL_X4 FILLER_28_282 ();
 FILLCELL_X2 FILLER_28_286 ();
 FILLCELL_X4 FILLER_28_292 ();
 FILLCELL_X4 FILLER_28_300 ();
 FILLCELL_X8 FILLER_28_309 ();
 FILLCELL_X4 FILLER_28_317 ();
 FILLCELL_X2 FILLER_28_321 ();
 FILLCELL_X4 FILLER_28_326 ();
 FILLCELL_X2 FILLER_28_330 ();
 FILLCELL_X4 FILLER_28_336 ();
 FILLCELL_X1 FILLER_28_340 ();
 FILLCELL_X4 FILLER_28_350 ();
 FILLCELL_X4 FILLER_28_363 ();
 FILLCELL_X8 FILLER_28_372 ();
 FILLCELL_X2 FILLER_28_380 ();
 FILLCELL_X1 FILLER_28_382 ();
 FILLCELL_X4 FILLER_28_387 ();
 FILLCELL_X4 FILLER_28_394 ();
 FILLCELL_X16 FILLER_28_402 ();
 FILLCELL_X8 FILLER_28_418 ();
 FILLCELL_X1 FILLER_28_426 ();
 FILLCELL_X16 FILLER_28_436 ();
 FILLCELL_X8 FILLER_28_452 ();
 FILLCELL_X4 FILLER_28_460 ();
 FILLCELL_X2 FILLER_28_464 ();
 FILLCELL_X1 FILLER_28_466 ();
 FILLCELL_X4 FILLER_28_470 ();
 FILLCELL_X4 FILLER_28_478 ();
 FILLCELL_X4 FILLER_28_491 ();
 FILLCELL_X8 FILLER_28_500 ();
 FILLCELL_X16 FILLER_28_533 ();
 FILLCELL_X8 FILLER_28_549 ();
 FILLCELL_X1 FILLER_28_557 ();
 FILLCELL_X16 FILLER_28_562 ();
 FILLCELL_X4 FILLER_28_578 ();
 FILLCELL_X2 FILLER_28_582 ();
 FILLCELL_X8 FILLER_28_588 ();
 FILLCELL_X2 FILLER_28_596 ();
 FILLCELL_X4 FILLER_28_604 ();
 FILLCELL_X8 FILLER_28_615 ();
 FILLCELL_X1 FILLER_28_623 ();
 FILLCELL_X4 FILLER_28_627 ();
 FILLCELL_X4 FILLER_28_632 ();
 FILLCELL_X4 FILLER_28_640 ();
 FILLCELL_X2 FILLER_28_644 ();
 FILLCELL_X1 FILLER_28_646 ();
 FILLCELL_X4 FILLER_28_650 ();
 FILLCELL_X8 FILLER_28_658 ();
 FILLCELL_X2 FILLER_28_666 ();
 FILLCELL_X8 FILLER_28_671 ();
 FILLCELL_X2 FILLER_28_679 ();
 FILLCELL_X8 FILLER_28_685 ();
 FILLCELL_X2 FILLER_28_693 ();
 FILLCELL_X1 FILLER_28_695 ();
 FILLCELL_X4 FILLER_28_699 ();
 FILLCELL_X1 FILLER_28_703 ();
 FILLCELL_X4 FILLER_28_707 ();
 FILLCELL_X4 FILLER_28_715 ();
 FILLCELL_X4 FILLER_28_722 ();
 FILLCELL_X1 FILLER_28_726 ();
 FILLCELL_X4 FILLER_28_732 ();
 FILLCELL_X2 FILLER_28_736 ();
 FILLCELL_X4 FILLER_28_742 ();
 FILLCELL_X4 FILLER_28_751 ();
 FILLCELL_X2 FILLER_28_755 ();
 FILLCELL_X1 FILLER_28_757 ();
 FILLCELL_X4 FILLER_28_764 ();
 FILLCELL_X8 FILLER_28_773 ();
 FILLCELL_X16 FILLER_28_800 ();
 FILLCELL_X8 FILLER_28_816 ();
 FILLCELL_X4 FILLER_28_824 ();
 FILLCELL_X2 FILLER_28_828 ();
 FILLCELL_X1 FILLER_28_830 ();
 FILLCELL_X4 FILLER_28_835 ();
 FILLCELL_X8 FILLER_28_848 ();
 FILLCELL_X2 FILLER_28_856 ();
 FILLCELL_X4 FILLER_28_863 ();
 FILLCELL_X4 FILLER_28_873 ();
 FILLCELL_X1 FILLER_28_877 ();
 FILLCELL_X4 FILLER_28_883 ();
 FILLCELL_X1 FILLER_28_887 ();
 FILLCELL_X4 FILLER_28_892 ();
 FILLCELL_X4 FILLER_28_900 ();
 FILLCELL_X8 FILLER_28_913 ();
 FILLCELL_X4 FILLER_28_921 ();
 FILLCELL_X1 FILLER_28_925 ();
 FILLCELL_X4 FILLER_28_929 ();
 FILLCELL_X4 FILLER_28_939 ();
 FILLCELL_X8 FILLER_28_948 ();
 FILLCELL_X2 FILLER_28_956 ();
 FILLCELL_X4 FILLER_28_963 ();
 FILLCELL_X4 FILLER_28_976 ();
 FILLCELL_X4 FILLER_28_987 ();
 FILLCELL_X8 FILLER_28_995 ();
 FILLCELL_X1 FILLER_28_1003 ();
 FILLCELL_X8 FILLER_28_1013 ();
 FILLCELL_X4 FILLER_28_1028 ();
 FILLCELL_X4 FILLER_28_1042 ();
 FILLCELL_X4 FILLER_28_1050 ();
 FILLCELL_X1 FILLER_28_1054 ();
 FILLCELL_X8 FILLER_28_1059 ();
 FILLCELL_X4 FILLER_28_1076 ();
 FILLCELL_X4 FILLER_28_1089 ();
 FILLCELL_X4 FILLER_28_1097 ();
 FILLCELL_X4 FILLER_28_1103 ();
 FILLCELL_X1 FILLER_28_1107 ();
 FILLCELL_X4 FILLER_28_1111 ();
 FILLCELL_X4 FILLER_28_1118 ();
 FILLCELL_X8 FILLER_28_1125 ();
 FILLCELL_X2 FILLER_28_1133 ();
 FILLCELL_X8 FILLER_28_1139 ();
 FILLCELL_X2 FILLER_28_1147 ();
 FILLCELL_X8 FILLER_28_1159 ();
 FILLCELL_X2 FILLER_28_1167 ();
 FILLCELL_X1 FILLER_28_1169 ();
 FILLCELL_X8 FILLER_28_1177 ();
 FILLCELL_X1 FILLER_28_1185 ();
 FILLCELL_X4 FILLER_28_1190 ();
 FILLCELL_X4 FILLER_28_1199 ();
 FILLCELL_X4 FILLER_28_1212 ();
 FILLCELL_X4 FILLER_28_1226 ();
 FILLCELL_X4 FILLER_28_1240 ();
 FILLCELL_X8 FILLER_28_1246 ();
 FILLCELL_X4 FILLER_28_1254 ();
 FILLCELL_X1 FILLER_28_1258 ();
 FILLCELL_X4 FILLER_28_1261 ();
 FILLCELL_X1 FILLER_28_1265 ();
 FILLCELL_X4 FILLER_28_1268 ();
 FILLCELL_X2 FILLER_28_1272 ();
 FILLCELL_X4 FILLER_28_1276 ();
 FILLCELL_X4 FILLER_28_1283 ();
 FILLCELL_X4 FILLER_28_1296 ();
 FILLCELL_X4 FILLER_28_1310 ();
 FILLCELL_X4 FILLER_28_1321 ();
 FILLCELL_X2 FILLER_28_1325 ();
 FILLCELL_X1 FILLER_28_1327 ();
 FILLCELL_X4 FILLER_28_1330 ();
 FILLCELL_X32 FILLER_28_1344 ();
 FILLCELL_X1 FILLER_28_1376 ();
 FILLCELL_X4 FILLER_28_1381 ();
 FILLCELL_X4 FILLER_28_1391 ();
 FILLCELL_X4 FILLER_28_1401 ();
 FILLCELL_X32 FILLER_28_1409 ();
 FILLCELL_X32 FILLER_28_1441 ();
 FILLCELL_X32 FILLER_28_1473 ();
 FILLCELL_X32 FILLER_28_1505 ();
 FILLCELL_X32 FILLER_28_1537 ();
 FILLCELL_X32 FILLER_28_1569 ();
 FILLCELL_X32 FILLER_28_1601 ();
 FILLCELL_X32 FILLER_28_1633 ();
 FILLCELL_X32 FILLER_28_1665 ();
 FILLCELL_X32 FILLER_28_1697 ();
 FILLCELL_X16 FILLER_28_1729 ();
 FILLCELL_X8 FILLER_28_1745 ();
 FILLCELL_X2 FILLER_28_1753 ();
 FILLCELL_X1 FILLER_28_1755 ();
 FILLCELL_X8 FILLER_29_1 ();
 FILLCELL_X4 FILLER_29_18 ();
 FILLCELL_X4 FILLER_29_26 ();
 FILLCELL_X8 FILLER_29_32 ();
 FILLCELL_X4 FILLER_29_40 ();
 FILLCELL_X2 FILLER_29_44 ();
 FILLCELL_X1 FILLER_29_46 ();
 FILLCELL_X4 FILLER_29_49 ();
 FILLCELL_X2 FILLER_29_53 ();
 FILLCELL_X1 FILLER_29_55 ();
 FILLCELL_X8 FILLER_29_66 ();
 FILLCELL_X4 FILLER_29_74 ();
 FILLCELL_X2 FILLER_29_78 ();
 FILLCELL_X4 FILLER_29_87 ();
 FILLCELL_X8 FILLER_29_100 ();
 FILLCELL_X4 FILLER_29_108 ();
 FILLCELL_X4 FILLER_29_115 ();
 FILLCELL_X4 FILLER_29_122 ();
 FILLCELL_X4 FILLER_29_129 ();
 FILLCELL_X4 FILLER_29_143 ();
 FILLCELL_X4 FILLER_29_154 ();
 FILLCELL_X1 FILLER_29_158 ();
 FILLCELL_X4 FILLER_29_169 ();
 FILLCELL_X4 FILLER_29_180 ();
 FILLCELL_X4 FILLER_29_188 ();
 FILLCELL_X2 FILLER_29_192 ();
 FILLCELL_X4 FILLER_29_198 ();
 FILLCELL_X8 FILLER_29_221 ();
 FILLCELL_X1 FILLER_29_229 ();
 FILLCELL_X16 FILLER_29_235 ();
 FILLCELL_X2 FILLER_29_251 ();
 FILLCELL_X1 FILLER_29_253 ();
 FILLCELL_X4 FILLER_29_257 ();
 FILLCELL_X2 FILLER_29_261 ();
 FILLCELL_X4 FILLER_29_266 ();
 FILLCELL_X2 FILLER_29_270 ();
 FILLCELL_X1 FILLER_29_272 ();
 FILLCELL_X4 FILLER_29_280 ();
 FILLCELL_X4 FILLER_29_293 ();
 FILLCELL_X4 FILLER_29_306 ();
 FILLCELL_X8 FILLER_29_314 ();
 FILLCELL_X8 FILLER_29_327 ();
 FILLCELL_X1 FILLER_29_335 ();
 FILLCELL_X4 FILLER_29_340 ();
 FILLCELL_X4 FILLER_29_353 ();
 FILLCELL_X1 FILLER_29_357 ();
 FILLCELL_X8 FILLER_29_364 ();
 FILLCELL_X4 FILLER_29_372 ();
 FILLCELL_X2 FILLER_29_376 ();
 FILLCELL_X1 FILLER_29_378 ();
 FILLCELL_X16 FILLER_29_392 ();
 FILLCELL_X2 FILLER_29_408 ();
 FILLCELL_X1 FILLER_29_410 ();
 FILLCELL_X8 FILLER_29_415 ();
 FILLCELL_X2 FILLER_29_423 ();
 FILLCELL_X4 FILLER_29_429 ();
 FILLCELL_X4 FILLER_29_437 ();
 FILLCELL_X2 FILLER_29_441 ();
 FILLCELL_X1 FILLER_29_443 ();
 FILLCELL_X4 FILLER_29_448 ();
 FILLCELL_X4 FILLER_29_456 ();
 FILLCELL_X2 FILLER_29_460 ();
 FILLCELL_X1 FILLER_29_462 ();
 FILLCELL_X8 FILLER_29_469 ();
 FILLCELL_X1 FILLER_29_477 ();
 FILLCELL_X4 FILLER_29_484 ();
 FILLCELL_X4 FILLER_29_497 ();
 FILLCELL_X4 FILLER_29_510 ();
 FILLCELL_X16 FILLER_29_518 ();
 FILLCELL_X2 FILLER_29_534 ();
 FILLCELL_X1 FILLER_29_536 ();
 FILLCELL_X4 FILLER_29_541 ();
 FILLCELL_X4 FILLER_29_549 ();
 FILLCELL_X1 FILLER_29_553 ();
 FILLCELL_X4 FILLER_29_558 ();
 FILLCELL_X8 FILLER_29_568 ();
 FILLCELL_X4 FILLER_29_576 ();
 FILLCELL_X4 FILLER_29_589 ();
 FILLCELL_X8 FILLER_29_597 ();
 FILLCELL_X2 FILLER_29_605 ();
 FILLCELL_X4 FILLER_29_610 ();
 FILLCELL_X8 FILLER_29_618 ();
 FILLCELL_X4 FILLER_29_630 ();
 FILLCELL_X4 FILLER_29_640 ();
 FILLCELL_X8 FILLER_29_647 ();
 FILLCELL_X2 FILLER_29_655 ();
 FILLCELL_X4 FILLER_29_661 ();
 FILLCELL_X8 FILLER_29_669 ();
 FILLCELL_X2 FILLER_29_677 ();
 FILLCELL_X1 FILLER_29_679 ();
 FILLCELL_X4 FILLER_29_686 ();
 FILLCELL_X8 FILLER_29_695 ();
 FILLCELL_X4 FILLER_29_712 ();
 FILLCELL_X8 FILLER_29_720 ();
 FILLCELL_X4 FILLER_29_728 ();
 FILLCELL_X16 FILLER_29_736 ();
 FILLCELL_X1 FILLER_29_752 ();
 FILLCELL_X4 FILLER_29_756 ();
 FILLCELL_X2 FILLER_29_760 ();
 FILLCELL_X32 FILLER_29_766 ();
 FILLCELL_X2 FILLER_29_798 ();
 FILLCELL_X4 FILLER_29_809 ();
 FILLCELL_X4 FILLER_29_818 ();
 FILLCELL_X2 FILLER_29_822 ();
 FILLCELL_X4 FILLER_29_827 ();
 FILLCELL_X4 FILLER_29_837 ();
 FILLCELL_X4 FILLER_29_850 ();
 FILLCELL_X16 FILLER_29_857 ();
 FILLCELL_X1 FILLER_29_873 ();
 FILLCELL_X8 FILLER_29_877 ();
 FILLCELL_X8 FILLER_29_888 ();
 FILLCELL_X4 FILLER_29_901 ();
 FILLCELL_X4 FILLER_29_914 ();
 FILLCELL_X2 FILLER_29_918 ();
 FILLCELL_X1 FILLER_29_920 ();
 FILLCELL_X4 FILLER_29_925 ();
 FILLCELL_X4 FILLER_29_938 ();
 FILLCELL_X4 FILLER_29_951 ();
 FILLCELL_X8 FILLER_29_959 ();
 FILLCELL_X8 FILLER_29_972 ();
 FILLCELL_X4 FILLER_29_980 ();
 FILLCELL_X4 FILLER_29_989 ();
 FILLCELL_X8 FILLER_29_1002 ();
 FILLCELL_X4 FILLER_29_1010 ();
 FILLCELL_X1 FILLER_29_1014 ();
 FILLCELL_X8 FILLER_29_1025 ();
 FILLCELL_X2 FILLER_29_1033 ();
 FILLCELL_X4 FILLER_29_1039 ();
 FILLCELL_X4 FILLER_29_1046 ();
 FILLCELL_X16 FILLER_29_1059 ();
 FILLCELL_X8 FILLER_29_1075 ();
 FILLCELL_X4 FILLER_29_1083 ();
 FILLCELL_X1 FILLER_29_1087 ();
 FILLCELL_X8 FILLER_29_1091 ();
 FILLCELL_X4 FILLER_29_1099 ();
 FILLCELL_X2 FILLER_29_1103 ();
 FILLCELL_X4 FILLER_29_1109 ();
 FILLCELL_X4 FILLER_29_1122 ();
 FILLCELL_X8 FILLER_29_1135 ();
 FILLCELL_X1 FILLER_29_1143 ();
 FILLCELL_X4 FILLER_29_1154 ();
 FILLCELL_X8 FILLER_29_1160 ();
 FILLCELL_X1 FILLER_29_1168 ();
 FILLCELL_X4 FILLER_29_1176 ();
 FILLCELL_X4 FILLER_29_1182 ();
 FILLCELL_X4 FILLER_29_1188 ();
 FILLCELL_X1 FILLER_29_1192 ();
 FILLCELL_X4 FILLER_29_1197 ();
 FILLCELL_X16 FILLER_29_1205 ();
 FILLCELL_X4 FILLER_29_1221 ();
 FILLCELL_X2 FILLER_29_1225 ();
 FILLCELL_X8 FILLER_29_1229 ();
 FILLCELL_X4 FILLER_29_1237 ();
 FILLCELL_X2 FILLER_29_1241 ();
 FILLCELL_X4 FILLER_29_1246 ();
 FILLCELL_X4 FILLER_29_1259 ();
 FILLCELL_X4 FILLER_29_1264 ();
 FILLCELL_X4 FILLER_29_1270 ();
 FILLCELL_X2 FILLER_29_1274 ();
 FILLCELL_X1 FILLER_29_1276 ();
 FILLCELL_X4 FILLER_29_1279 ();
 FILLCELL_X4 FILLER_29_1286 ();
 FILLCELL_X4 FILLER_29_1293 ();
 FILLCELL_X8 FILLER_29_1299 ();
 FILLCELL_X4 FILLER_29_1309 ();
 FILLCELL_X8 FILLER_29_1323 ();
 FILLCELL_X4 FILLER_29_1331 ();
 FILLCELL_X4 FILLER_29_1338 ();
 FILLCELL_X4 FILLER_29_1349 ();
 FILLCELL_X4 FILLER_29_1356 ();
 FILLCELL_X16 FILLER_29_1362 ();
 FILLCELL_X8 FILLER_29_1378 ();
 FILLCELL_X2 FILLER_29_1386 ();
 FILLCELL_X8 FILLER_29_1392 ();
 FILLCELL_X2 FILLER_29_1400 ();
 FILLCELL_X1 FILLER_29_1402 ();
 FILLCELL_X32 FILLER_29_1422 ();
 FILLCELL_X32 FILLER_29_1454 ();
 FILLCELL_X32 FILLER_29_1486 ();
 FILLCELL_X32 FILLER_29_1518 ();
 FILLCELL_X32 FILLER_29_1550 ();
 FILLCELL_X32 FILLER_29_1582 ();
 FILLCELL_X32 FILLER_29_1614 ();
 FILLCELL_X32 FILLER_29_1646 ();
 FILLCELL_X32 FILLER_29_1678 ();
 FILLCELL_X32 FILLER_29_1710 ();
 FILLCELL_X8 FILLER_29_1742 ();
 FILLCELL_X4 FILLER_29_1750 ();
 FILLCELL_X2 FILLER_29_1754 ();
 FILLCELL_X4 FILLER_30_1 ();
 FILLCELL_X4 FILLER_30_8 ();
 FILLCELL_X8 FILLER_30_16 ();
 FILLCELL_X2 FILLER_30_24 ();
 FILLCELL_X4 FILLER_30_30 ();
 FILLCELL_X8 FILLER_30_43 ();
 FILLCELL_X4 FILLER_30_55 ();
 FILLCELL_X4 FILLER_30_69 ();
 FILLCELL_X4 FILLER_30_77 ();
 FILLCELL_X4 FILLER_30_91 ();
 FILLCELL_X4 FILLER_30_98 ();
 FILLCELL_X4 FILLER_30_105 ();
 FILLCELL_X4 FILLER_30_119 ();
 FILLCELL_X4 FILLER_30_132 ();
 FILLCELL_X8 FILLER_30_146 ();
 FILLCELL_X1 FILLER_30_154 ();
 FILLCELL_X4 FILLER_30_157 ();
 FILLCELL_X2 FILLER_30_161 ();
 FILLCELL_X4 FILLER_30_166 ();
 FILLCELL_X1 FILLER_30_170 ();
 FILLCELL_X4 FILLER_30_178 ();
 FILLCELL_X4 FILLER_30_192 ();
 FILLCELL_X4 FILLER_30_205 ();
 FILLCELL_X4 FILLER_30_212 ();
 FILLCELL_X4 FILLER_30_220 ();
 FILLCELL_X4 FILLER_30_229 ();
 FILLCELL_X4 FILLER_30_242 ();
 FILLCELL_X8 FILLER_30_255 ();
 FILLCELL_X2 FILLER_30_263 ();
 FILLCELL_X1 FILLER_30_265 ();
 FILLCELL_X4 FILLER_30_270 ();
 FILLCELL_X8 FILLER_30_284 ();
 FILLCELL_X2 FILLER_30_292 ();
 FILLCELL_X4 FILLER_30_297 ();
 FILLCELL_X4 FILLER_30_304 ();
 FILLCELL_X4 FILLER_30_312 ();
 FILLCELL_X4 FILLER_30_325 ();
 FILLCELL_X16 FILLER_30_338 ();
 FILLCELL_X2 FILLER_30_354 ();
 FILLCELL_X4 FILLER_30_359 ();
 FILLCELL_X2 FILLER_30_363 ();
 FILLCELL_X1 FILLER_30_365 ();
 FILLCELL_X4 FILLER_30_370 ();
 FILLCELL_X8 FILLER_30_380 ();
 FILLCELL_X1 FILLER_30_388 ();
 FILLCELL_X8 FILLER_30_393 ();
 FILLCELL_X2 FILLER_30_401 ();
 FILLCELL_X1 FILLER_30_403 ();
 FILLCELL_X16 FILLER_30_421 ();
 FILLCELL_X8 FILLER_30_437 ();
 FILLCELL_X4 FILLER_30_445 ();
 FILLCELL_X4 FILLER_30_458 ();
 FILLCELL_X4 FILLER_30_471 ();
 FILLCELL_X4 FILLER_30_480 ();
 FILLCELL_X1 FILLER_30_484 ();
 FILLCELL_X4 FILLER_30_490 ();
 FILLCELL_X8 FILLER_30_498 ();
 FILLCELL_X1 FILLER_30_506 ();
 FILLCELL_X8 FILLER_30_511 ();
 FILLCELL_X2 FILLER_30_519 ();
 FILLCELL_X4 FILLER_30_525 ();
 FILLCELL_X4 FILLER_30_533 ();
 FILLCELL_X8 FILLER_30_546 ();
 FILLCELL_X1 FILLER_30_554 ();
 FILLCELL_X4 FILLER_30_564 ();
 FILLCELL_X4 FILLER_30_577 ();
 FILLCELL_X8 FILLER_30_584 ();
 FILLCELL_X4 FILLER_30_592 ();
 FILLCELL_X2 FILLER_30_596 ();
 FILLCELL_X4 FILLER_30_601 ();
 FILLCELL_X4 FILLER_30_609 ();
 FILLCELL_X8 FILLER_30_622 ();
 FILLCELL_X1 FILLER_30_630 ();
 FILLCELL_X8 FILLER_30_632 ();
 FILLCELL_X2 FILLER_30_640 ();
 FILLCELL_X8 FILLER_30_648 ();
 FILLCELL_X2 FILLER_30_656 ();
 FILLCELL_X1 FILLER_30_658 ();
 FILLCELL_X4 FILLER_30_668 ();
 FILLCELL_X4 FILLER_30_681 ();
 FILLCELL_X8 FILLER_30_694 ();
 FILLCELL_X2 FILLER_30_702 ();
 FILLCELL_X8 FILLER_30_713 ();
 FILLCELL_X4 FILLER_30_725 ();
 FILLCELL_X4 FILLER_30_738 ();
 FILLCELL_X4 FILLER_30_748 ();
 FILLCELL_X4 FILLER_30_756 ();
 FILLCELL_X1 FILLER_30_760 ();
 FILLCELL_X4 FILLER_30_765 ();
 FILLCELL_X2 FILLER_30_769 ();
 FILLCELL_X1 FILLER_30_771 ();
 FILLCELL_X4 FILLER_30_781 ();
 FILLCELL_X1 FILLER_30_785 ();
 FILLCELL_X4 FILLER_30_791 ();
 FILLCELL_X2 FILLER_30_795 ();
 FILLCELL_X4 FILLER_30_800 ();
 FILLCELL_X4 FILLER_30_810 ();
 FILLCELL_X4 FILLER_30_823 ();
 FILLCELL_X8 FILLER_30_830 ();
 FILLCELL_X2 FILLER_30_838 ();
 FILLCELL_X4 FILLER_30_844 ();
 FILLCELL_X16 FILLER_30_851 ();
 FILLCELL_X4 FILLER_30_867 ();
 FILLCELL_X1 FILLER_30_871 ();
 FILLCELL_X4 FILLER_30_878 ();
 FILLCELL_X4 FILLER_30_886 ();
 FILLCELL_X2 FILLER_30_890 ();
 FILLCELL_X1 FILLER_30_892 ();
 FILLCELL_X4 FILLER_30_896 ();
 FILLCELL_X4 FILLER_30_906 ();
 FILLCELL_X4 FILLER_30_914 ();
 FILLCELL_X4 FILLER_30_921 ();
 FILLCELL_X1 FILLER_30_925 ();
 FILLCELL_X4 FILLER_30_930 ();
 FILLCELL_X4 FILLER_30_939 ();
 FILLCELL_X8 FILLER_30_947 ();
 FILLCELL_X4 FILLER_30_955 ();
 FILLCELL_X2 FILLER_30_959 ();
 FILLCELL_X1 FILLER_30_961 ();
 FILLCELL_X4 FILLER_30_966 ();
 FILLCELL_X1 FILLER_30_970 ();
 FILLCELL_X8 FILLER_30_975 ();
 FILLCELL_X4 FILLER_30_987 ();
 FILLCELL_X4 FILLER_30_995 ();
 FILLCELL_X1 FILLER_30_999 ();
 FILLCELL_X16 FILLER_30_1003 ();
 FILLCELL_X8 FILLER_30_1019 ();
 FILLCELL_X2 FILLER_30_1027 ();
 FILLCELL_X1 FILLER_30_1029 ();
 FILLCELL_X4 FILLER_30_1034 ();
 FILLCELL_X16 FILLER_30_1047 ();
 FILLCELL_X2 FILLER_30_1063 ();
 FILLCELL_X1 FILLER_30_1065 ();
 FILLCELL_X4 FILLER_30_1070 ();
 FILLCELL_X1 FILLER_30_1074 ();
 FILLCELL_X4 FILLER_30_1078 ();
 FILLCELL_X4 FILLER_30_1085 ();
 FILLCELL_X4 FILLER_30_1098 ();
 FILLCELL_X4 FILLER_30_1106 ();
 FILLCELL_X8 FILLER_30_1114 ();
 FILLCELL_X16 FILLER_30_1125 ();
 FILLCELL_X4 FILLER_30_1141 ();
 FILLCELL_X8 FILLER_30_1148 ();
 FILLCELL_X1 FILLER_30_1156 ();
 FILLCELL_X4 FILLER_30_1161 ();
 FILLCELL_X4 FILLER_30_1167 ();
 FILLCELL_X16 FILLER_30_1174 ();
 FILLCELL_X4 FILLER_30_1190 ();
 FILLCELL_X1 FILLER_30_1194 ();
 FILLCELL_X4 FILLER_30_1199 ();
 FILLCELL_X4 FILLER_30_1207 ();
 FILLCELL_X2 FILLER_30_1211 ();
 FILLCELL_X4 FILLER_30_1216 ();
 FILLCELL_X4 FILLER_30_1223 ();
 FILLCELL_X2 FILLER_30_1227 ();
 FILLCELL_X4 FILLER_30_1232 ();
 FILLCELL_X4 FILLER_30_1246 ();
 FILLCELL_X4 FILLER_30_1257 ();
 FILLCELL_X4 FILLER_30_1263 ();
 FILLCELL_X4 FILLER_30_1277 ();
 FILLCELL_X8 FILLER_30_1290 ();
 FILLCELL_X2 FILLER_30_1298 ();
 FILLCELL_X1 FILLER_30_1300 ();
 FILLCELL_X4 FILLER_30_1308 ();
 FILLCELL_X8 FILLER_30_1314 ();
 FILLCELL_X2 FILLER_30_1322 ();
 FILLCELL_X1 FILLER_30_1324 ();
 FILLCELL_X4 FILLER_30_1328 ();
 FILLCELL_X4 FILLER_30_1335 ();
 FILLCELL_X1 FILLER_30_1339 ();
 FILLCELL_X4 FILLER_30_1346 ();
 FILLCELL_X4 FILLER_30_1352 ();
 FILLCELL_X2 FILLER_30_1356 ();
 FILLCELL_X4 FILLER_30_1377 ();
 FILLCELL_X32 FILLER_30_1383 ();
 FILLCELL_X32 FILLER_30_1415 ();
 FILLCELL_X32 FILLER_30_1447 ();
 FILLCELL_X32 FILLER_30_1479 ();
 FILLCELL_X32 FILLER_30_1511 ();
 FILLCELL_X32 FILLER_30_1543 ();
 FILLCELL_X32 FILLER_30_1575 ();
 FILLCELL_X32 FILLER_30_1607 ();
 FILLCELL_X32 FILLER_30_1639 ();
 FILLCELL_X32 FILLER_30_1671 ();
 FILLCELL_X32 FILLER_30_1703 ();
 FILLCELL_X8 FILLER_30_1735 ();
 FILLCELL_X4 FILLER_30_1743 ();
 FILLCELL_X2 FILLER_30_1747 ();
 FILLCELL_X4 FILLER_30_1752 ();
 FILLCELL_X4 FILLER_31_1 ();
 FILLCELL_X2 FILLER_31_5 ();
 FILLCELL_X8 FILLER_31_10 ();
 FILLCELL_X4 FILLER_31_28 ();
 FILLCELL_X2 FILLER_31_32 ();
 FILLCELL_X1 FILLER_31_34 ();
 FILLCELL_X4 FILLER_31_38 ();
 FILLCELL_X8 FILLER_31_45 ();
 FILLCELL_X4 FILLER_31_56 ();
 FILLCELL_X16 FILLER_31_67 ();
 FILLCELL_X2 FILLER_31_83 ();
 FILLCELL_X1 FILLER_31_85 ();
 FILLCELL_X4 FILLER_31_89 ();
 FILLCELL_X8 FILLER_31_96 ();
 FILLCELL_X4 FILLER_31_104 ();
 FILLCELL_X2 FILLER_31_108 ();
 FILLCELL_X16 FILLER_31_112 ();
 FILLCELL_X4 FILLER_31_128 ();
 FILLCELL_X2 FILLER_31_132 ();
 FILLCELL_X1 FILLER_31_134 ();
 FILLCELL_X4 FILLER_31_138 ();
 FILLCELL_X8 FILLER_31_145 ();
 FILLCELL_X1 FILLER_31_153 ();
 FILLCELL_X4 FILLER_31_156 ();
 FILLCELL_X4 FILLER_31_170 ();
 FILLCELL_X8 FILLER_31_177 ();
 FILLCELL_X4 FILLER_31_188 ();
 FILLCELL_X1 FILLER_31_192 ();
 FILLCELL_X4 FILLER_31_196 ();
 FILLCELL_X8 FILLER_31_202 ();
 FILLCELL_X2 FILLER_31_210 ();
 FILLCELL_X1 FILLER_31_212 ();
 FILLCELL_X4 FILLER_31_217 ();
 FILLCELL_X4 FILLER_31_225 ();
 FILLCELL_X4 FILLER_31_233 ();
 FILLCELL_X4 FILLER_31_239 ();
 FILLCELL_X2 FILLER_31_243 ();
 FILLCELL_X1 FILLER_31_245 ();
 FILLCELL_X8 FILLER_31_250 ();
 FILLCELL_X4 FILLER_31_258 ();
 FILLCELL_X2 FILLER_31_262 ();
 FILLCELL_X4 FILLER_31_274 ();
 FILLCELL_X4 FILLER_31_280 ();
 FILLCELL_X2 FILLER_31_284 ();
 FILLCELL_X16 FILLER_31_289 ();
 FILLCELL_X2 FILLER_31_305 ();
 FILLCELL_X4 FILLER_31_310 ();
 FILLCELL_X2 FILLER_31_314 ();
 FILLCELL_X4 FILLER_31_319 ();
 FILLCELL_X4 FILLER_31_327 ();
 FILLCELL_X4 FILLER_31_336 ();
 FILLCELL_X4 FILLER_31_343 ();
 FILLCELL_X1 FILLER_31_347 ();
 FILLCELL_X4 FILLER_31_354 ();
 FILLCELL_X4 FILLER_31_362 ();
 FILLCELL_X4 FILLER_31_369 ();
 FILLCELL_X2 FILLER_31_373 ();
 FILLCELL_X4 FILLER_31_381 ();
 FILLCELL_X2 FILLER_31_385 ();
 FILLCELL_X8 FILLER_31_406 ();
 FILLCELL_X1 FILLER_31_414 ();
 FILLCELL_X8 FILLER_31_421 ();
 FILLCELL_X1 FILLER_31_429 ();
 FILLCELL_X4 FILLER_31_443 ();
 FILLCELL_X4 FILLER_31_451 ();
 FILLCELL_X4 FILLER_31_464 ();
 FILLCELL_X4 FILLER_31_472 ();
 FILLCELL_X8 FILLER_31_481 ();
 FILLCELL_X2 FILLER_31_489 ();
 FILLCELL_X4 FILLER_31_494 ();
 FILLCELL_X4 FILLER_31_507 ();
 FILLCELL_X2 FILLER_31_511 ();
 FILLCELL_X8 FILLER_31_522 ();
 FILLCELL_X4 FILLER_31_539 ();
 FILLCELL_X8 FILLER_31_552 ();
 FILLCELL_X2 FILLER_31_560 ();
 FILLCELL_X8 FILLER_31_567 ();
 FILLCELL_X2 FILLER_31_575 ();
 FILLCELL_X4 FILLER_31_582 ();
 FILLCELL_X8 FILLER_31_595 ();
 FILLCELL_X4 FILLER_31_603 ();
 FILLCELL_X8 FILLER_31_612 ();
 FILLCELL_X4 FILLER_31_624 ();
 FILLCELL_X4 FILLER_31_641 ();
 FILLCELL_X8 FILLER_31_664 ();
 FILLCELL_X4 FILLER_31_672 ();
 FILLCELL_X1 FILLER_31_676 ();
 FILLCELL_X4 FILLER_31_681 ();
 FILLCELL_X4 FILLER_31_690 ();
 FILLCELL_X1 FILLER_31_694 ();
 FILLCELL_X4 FILLER_31_700 ();
 FILLCELL_X4 FILLER_31_713 ();
 FILLCELL_X4 FILLER_31_723 ();
 FILLCELL_X1 FILLER_31_727 ();
 FILLCELL_X4 FILLER_31_737 ();
 FILLCELL_X4 FILLER_31_750 ();
 FILLCELL_X8 FILLER_31_759 ();
 FILLCELL_X4 FILLER_31_776 ();
 FILLCELL_X2 FILLER_31_780 ();
 FILLCELL_X1 FILLER_31_782 ();
 FILLCELL_X4 FILLER_31_789 ();
 FILLCELL_X8 FILLER_31_798 ();
 FILLCELL_X4 FILLER_31_806 ();
 FILLCELL_X4 FILLER_31_814 ();
 FILLCELL_X16 FILLER_31_821 ();
 FILLCELL_X8 FILLER_31_837 ();
 FILLCELL_X2 FILLER_31_845 ();
 FILLCELL_X1 FILLER_31_847 ();
 FILLCELL_X8 FILLER_31_857 ();
 FILLCELL_X4 FILLER_31_874 ();
 FILLCELL_X16 FILLER_31_887 ();
 FILLCELL_X2 FILLER_31_903 ();
 FILLCELL_X16 FILLER_31_908 ();
 FILLCELL_X4 FILLER_31_924 ();
 FILLCELL_X1 FILLER_31_928 ();
 FILLCELL_X32 FILLER_31_932 ();
 FILLCELL_X2 FILLER_31_964 ();
 FILLCELL_X4 FILLER_31_975 ();
 FILLCELL_X4 FILLER_31_988 ();
 FILLCELL_X4 FILLER_31_996 ();
 FILLCELL_X2 FILLER_31_1000 ();
 FILLCELL_X4 FILLER_31_1006 ();
 FILLCELL_X8 FILLER_31_1013 ();
 FILLCELL_X4 FILLER_31_1025 ();
 FILLCELL_X4 FILLER_31_1033 ();
 FILLCELL_X1 FILLER_31_1037 ();
 FILLCELL_X16 FILLER_31_1041 ();
 FILLCELL_X2 FILLER_31_1057 ();
 FILLCELL_X1 FILLER_31_1059 ();
 FILLCELL_X8 FILLER_31_1064 ();
 FILLCELL_X1 FILLER_31_1072 ();
 FILLCELL_X4 FILLER_31_1082 ();
 FILLCELL_X32 FILLER_31_1090 ();
 FILLCELL_X4 FILLER_31_1122 ();
 FILLCELL_X4 FILLER_31_1129 ();
 FILLCELL_X8 FILLER_31_1136 ();
 FILLCELL_X1 FILLER_31_1144 ();
 FILLCELL_X4 FILLER_31_1149 ();
 FILLCELL_X4 FILLER_31_1157 ();
 FILLCELL_X2 FILLER_31_1161 ();
 FILLCELL_X4 FILLER_31_1172 ();
 FILLCELL_X4 FILLER_31_1182 ();
 FILLCELL_X16 FILLER_31_1189 ();
 FILLCELL_X2 FILLER_31_1205 ();
 FILLCELL_X1 FILLER_31_1207 ();
 FILLCELL_X4 FILLER_31_1211 ();
 FILLCELL_X4 FILLER_31_1224 ();
 FILLCELL_X4 FILLER_31_1237 ();
 FILLCELL_X8 FILLER_31_1243 ();
 FILLCELL_X1 FILLER_31_1251 ();
 FILLCELL_X4 FILLER_31_1259 ();
 FILLCELL_X4 FILLER_31_1264 ();
 FILLCELL_X1 FILLER_31_1268 ();
 FILLCELL_X8 FILLER_31_1279 ();
 FILLCELL_X1 FILLER_31_1287 ();
 FILLCELL_X8 FILLER_31_1298 ();
 FILLCELL_X1 FILLER_31_1306 ();
 FILLCELL_X4 FILLER_31_1317 ();
 FILLCELL_X2 FILLER_31_1321 ();
 FILLCELL_X4 FILLER_31_1332 ();
 FILLCELL_X8 FILLER_31_1339 ();
 FILLCELL_X1 FILLER_31_1347 ();
 FILLCELL_X4 FILLER_31_1354 ();
 FILLCELL_X4 FILLER_31_1362 ();
 FILLCELL_X4 FILLER_31_1385 ();
 FILLCELL_X4 FILLER_31_1395 ();
 FILLCELL_X4 FILLER_31_1403 ();
 FILLCELL_X4 FILLER_31_1411 ();
 FILLCELL_X1 FILLER_31_1415 ();
 FILLCELL_X32 FILLER_31_1418 ();
 FILLCELL_X32 FILLER_31_1450 ();
 FILLCELL_X32 FILLER_31_1482 ();
 FILLCELL_X32 FILLER_31_1514 ();
 FILLCELL_X32 FILLER_31_1546 ();
 FILLCELL_X32 FILLER_31_1578 ();
 FILLCELL_X32 FILLER_31_1610 ();
 FILLCELL_X32 FILLER_31_1642 ();
 FILLCELL_X32 FILLER_31_1674 ();
 FILLCELL_X32 FILLER_31_1706 ();
 FILLCELL_X16 FILLER_31_1738 ();
 FILLCELL_X2 FILLER_31_1754 ();
 FILLCELL_X16 FILLER_32_1 ();
 FILLCELL_X4 FILLER_32_17 ();
 FILLCELL_X2 FILLER_32_21 ();
 FILLCELL_X1 FILLER_32_23 ();
 FILLCELL_X4 FILLER_32_31 ();
 FILLCELL_X4 FILLER_32_44 ();
 FILLCELL_X8 FILLER_32_51 ();
 FILLCELL_X8 FILLER_32_62 ();
 FILLCELL_X4 FILLER_32_70 ();
 FILLCELL_X1 FILLER_32_74 ();
 FILLCELL_X4 FILLER_32_79 ();
 FILLCELL_X4 FILLER_32_92 ();
 FILLCELL_X4 FILLER_32_99 ();
 FILLCELL_X2 FILLER_32_103 ();
 FILLCELL_X4 FILLER_32_108 ();
 FILLCELL_X8 FILLER_32_119 ();
 FILLCELL_X4 FILLER_32_127 ();
 FILLCELL_X8 FILLER_32_140 ();
 FILLCELL_X2 FILLER_32_148 ();
 FILLCELL_X8 FILLER_32_159 ();
 FILLCELL_X1 FILLER_32_167 ();
 FILLCELL_X4 FILLER_32_171 ();
 FILLCELL_X4 FILLER_32_178 ();
 FILLCELL_X4 FILLER_32_185 ();
 FILLCELL_X2 FILLER_32_189 ();
 FILLCELL_X1 FILLER_32_191 ();
 FILLCELL_X4 FILLER_32_201 ();
 FILLCELL_X4 FILLER_32_208 ();
 FILLCELL_X1 FILLER_32_212 ();
 FILLCELL_X4 FILLER_32_217 ();
 FILLCELL_X8 FILLER_32_224 ();
 FILLCELL_X4 FILLER_32_235 ();
 FILLCELL_X4 FILLER_32_242 ();
 FILLCELL_X2 FILLER_32_246 ();
 FILLCELL_X4 FILLER_32_251 ();
 FILLCELL_X4 FILLER_32_258 ();
 FILLCELL_X4 FILLER_32_266 ();
 FILLCELL_X2 FILLER_32_270 ();
 FILLCELL_X8 FILLER_32_276 ();
 FILLCELL_X2 FILLER_32_284 ();
 FILLCELL_X4 FILLER_32_290 ();
 FILLCELL_X4 FILLER_32_299 ();
 FILLCELL_X4 FILLER_32_307 ();
 FILLCELL_X2 FILLER_32_311 ();
 FILLCELL_X1 FILLER_32_313 ();
 FILLCELL_X4 FILLER_32_317 ();
 FILLCELL_X2 FILLER_32_321 ();
 FILLCELL_X8 FILLER_32_329 ();
 FILLCELL_X2 FILLER_32_337 ();
 FILLCELL_X1 FILLER_32_339 ();
 FILLCELL_X4 FILLER_32_349 ();
 FILLCELL_X4 FILLER_32_362 ();
 FILLCELL_X32 FILLER_32_369 ();
 FILLCELL_X16 FILLER_32_401 ();
 FILLCELL_X4 FILLER_32_417 ();
 FILLCELL_X8 FILLER_32_427 ();
 FILLCELL_X4 FILLER_32_439 ();
 FILLCELL_X4 FILLER_32_447 ();
 FILLCELL_X16 FILLER_32_455 ();
 FILLCELL_X4 FILLER_32_471 ();
 FILLCELL_X2 FILLER_32_475 ();
 FILLCELL_X4 FILLER_32_486 ();
 FILLCELL_X2 FILLER_32_490 ();
 FILLCELL_X4 FILLER_32_495 ();
 FILLCELL_X4 FILLER_32_516 ();
 FILLCELL_X4 FILLER_32_530 ();
 FILLCELL_X2 FILLER_32_534 ();
 FILLCELL_X4 FILLER_32_540 ();
 FILLCELL_X2 FILLER_32_544 ();
 FILLCELL_X16 FILLER_32_551 ();
 FILLCELL_X2 FILLER_32_567 ();
 FILLCELL_X8 FILLER_32_573 ();
 FILLCELL_X2 FILLER_32_581 ();
 FILLCELL_X1 FILLER_32_583 ();
 FILLCELL_X4 FILLER_32_593 ();
 FILLCELL_X4 FILLER_32_606 ();
 FILLCELL_X4 FILLER_32_616 ();
 FILLCELL_X4 FILLER_32_625 ();
 FILLCELL_X2 FILLER_32_629 ();
 FILLCELL_X8 FILLER_32_632 ();
 FILLCELL_X4 FILLER_32_640 ();
 FILLCELL_X2 FILLER_32_644 ();
 FILLCELL_X1 FILLER_32_646 ();
 FILLCELL_X32 FILLER_32_651 ();
 FILLCELL_X16 FILLER_32_683 ();
 FILLCELL_X4 FILLER_32_699 ();
 FILLCELL_X1 FILLER_32_703 ();
 FILLCELL_X8 FILLER_32_707 ();
 FILLCELL_X1 FILLER_32_715 ();
 FILLCELL_X4 FILLER_32_721 ();
 FILLCELL_X4 FILLER_32_730 ();
 FILLCELL_X8 FILLER_32_737 ();
 FILLCELL_X1 FILLER_32_745 ();
 FILLCELL_X4 FILLER_32_750 ();
 FILLCELL_X4 FILLER_32_758 ();
 FILLCELL_X2 FILLER_32_762 ();
 FILLCELL_X1 FILLER_32_764 ();
 FILLCELL_X4 FILLER_32_774 ();
 FILLCELL_X32 FILLER_32_781 ();
 FILLCELL_X1 FILLER_32_813 ();
 FILLCELL_X4 FILLER_32_823 ();
 FILLCELL_X4 FILLER_32_830 ();
 FILLCELL_X4 FILLER_32_837 ();
 FILLCELL_X4 FILLER_32_846 ();
 FILLCELL_X8 FILLER_32_860 ();
 FILLCELL_X1 FILLER_32_868 ();
 FILLCELL_X4 FILLER_32_872 ();
 FILLCELL_X4 FILLER_32_881 ();
 FILLCELL_X8 FILLER_32_888 ();
 FILLCELL_X4 FILLER_32_896 ();
 FILLCELL_X2 FILLER_32_900 ();
 FILLCELL_X8 FILLER_32_907 ();
 FILLCELL_X4 FILLER_32_915 ();
 FILLCELL_X2 FILLER_32_919 ();
 FILLCELL_X4 FILLER_32_924 ();
 FILLCELL_X4 FILLER_32_934 ();
 FILLCELL_X8 FILLER_32_943 ();
 FILLCELL_X4 FILLER_32_955 ();
 FILLCELL_X4 FILLER_32_968 ();
 FILLCELL_X4 FILLER_32_975 ();
 FILLCELL_X16 FILLER_32_982 ();
 FILLCELL_X2 FILLER_32_998 ();
 FILLCELL_X4 FILLER_32_1005 ();
 FILLCELL_X2 FILLER_32_1009 ();
 FILLCELL_X1 FILLER_32_1011 ();
 FILLCELL_X4 FILLER_32_1021 ();
 FILLCELL_X8 FILLER_32_1029 ();
 FILLCELL_X1 FILLER_32_1037 ();
 FILLCELL_X4 FILLER_32_1047 ();
 FILLCELL_X2 FILLER_32_1051 ();
 FILLCELL_X1 FILLER_32_1053 ();
 FILLCELL_X4 FILLER_32_1057 ();
 FILLCELL_X2 FILLER_32_1061 ();
 FILLCELL_X8 FILLER_32_1068 ();
 FILLCELL_X4 FILLER_32_1076 ();
 FILLCELL_X1 FILLER_32_1080 ();
 FILLCELL_X8 FILLER_32_1086 ();
 FILLCELL_X4 FILLER_32_1097 ();
 FILLCELL_X4 FILLER_32_1104 ();
 FILLCELL_X1 FILLER_32_1108 ();
 FILLCELL_X4 FILLER_32_1113 ();
 FILLCELL_X2 FILLER_32_1117 ();
 FILLCELL_X1 FILLER_32_1119 ();
 FILLCELL_X4 FILLER_32_1125 ();
 FILLCELL_X4 FILLER_32_1133 ();
 FILLCELL_X2 FILLER_32_1137 ();
 FILLCELL_X8 FILLER_32_1143 ();
 FILLCELL_X2 FILLER_32_1151 ();
 FILLCELL_X4 FILLER_32_1162 ();
 FILLCELL_X4 FILLER_32_1171 ();
 FILLCELL_X4 FILLER_32_1178 ();
 FILLCELL_X8 FILLER_32_1188 ();
 FILLCELL_X4 FILLER_32_1196 ();
 FILLCELL_X4 FILLER_32_1209 ();
 FILLCELL_X4 FILLER_32_1216 ();
 FILLCELL_X4 FILLER_32_1223 ();
 FILLCELL_X1 FILLER_32_1227 ();
 FILLCELL_X4 FILLER_32_1232 ();
 FILLCELL_X8 FILLER_32_1240 ();
 FILLCELL_X4 FILLER_32_1248 ();
 FILLCELL_X1 FILLER_32_1252 ();
 FILLCELL_X4 FILLER_32_1256 ();
 FILLCELL_X4 FILLER_32_1270 ();
 FILLCELL_X8 FILLER_32_1277 ();
 FILLCELL_X4 FILLER_32_1289 ();
 FILLCELL_X4 FILLER_32_1297 ();
 FILLCELL_X2 FILLER_32_1301 ();
 FILLCELL_X1 FILLER_32_1303 ();
 FILLCELL_X4 FILLER_32_1307 ();
 FILLCELL_X4 FILLER_32_1314 ();
 FILLCELL_X8 FILLER_32_1320 ();
 FILLCELL_X4 FILLER_32_1337 ();
 FILLCELL_X8 FILLER_32_1343 ();
 FILLCELL_X1 FILLER_32_1351 ();
 FILLCELL_X4 FILLER_32_1356 ();
 FILLCELL_X4 FILLER_32_1364 ();
 FILLCELL_X8 FILLER_32_1370 ();
 FILLCELL_X1 FILLER_32_1378 ();
 FILLCELL_X4 FILLER_32_1382 ();
 FILLCELL_X4 FILLER_32_1392 ();
 FILLCELL_X1 FILLER_32_1396 ();
 FILLCELL_X4 FILLER_32_1416 ();
 FILLCELL_X4 FILLER_32_1422 ();
 FILLCELL_X32 FILLER_32_1428 ();
 FILLCELL_X32 FILLER_32_1460 ();
 FILLCELL_X32 FILLER_32_1492 ();
 FILLCELL_X32 FILLER_32_1524 ();
 FILLCELL_X32 FILLER_32_1556 ();
 FILLCELL_X32 FILLER_32_1588 ();
 FILLCELL_X32 FILLER_32_1620 ();
 FILLCELL_X32 FILLER_32_1652 ();
 FILLCELL_X32 FILLER_32_1684 ();
 FILLCELL_X32 FILLER_32_1716 ();
 FILLCELL_X8 FILLER_32_1748 ();
 FILLCELL_X4 FILLER_33_1 ();
 FILLCELL_X16 FILLER_33_8 ();
 FILLCELL_X1 FILLER_33_24 ();
 FILLCELL_X8 FILLER_33_29 ();
 FILLCELL_X2 FILLER_33_37 ();
 FILLCELL_X1 FILLER_33_39 ();
 FILLCELL_X4 FILLER_33_44 ();
 FILLCELL_X4 FILLER_33_52 ();
 FILLCELL_X4 FILLER_33_65 ();
 FILLCELL_X4 FILLER_33_74 ();
 FILLCELL_X4 FILLER_33_87 ();
 FILLCELL_X4 FILLER_33_94 ();
 FILLCELL_X2 FILLER_33_98 ();
 FILLCELL_X4 FILLER_33_109 ();
 FILLCELL_X4 FILLER_33_123 ();
 FILLCELL_X4 FILLER_33_131 ();
 FILLCELL_X4 FILLER_33_144 ();
 FILLCELL_X2 FILLER_33_148 ();
 FILLCELL_X1 FILLER_33_150 ();
 FILLCELL_X4 FILLER_33_154 ();
 FILLCELL_X2 FILLER_33_158 ();
 FILLCELL_X4 FILLER_33_169 ();
 FILLCELL_X2 FILLER_33_173 ();
 FILLCELL_X1 FILLER_33_175 ();
 FILLCELL_X8 FILLER_33_186 ();
 FILLCELL_X1 FILLER_33_194 ();
 FILLCELL_X8 FILLER_33_202 ();
 FILLCELL_X1 FILLER_33_210 ();
 FILLCELL_X4 FILLER_33_220 ();
 FILLCELL_X2 FILLER_33_224 ();
 FILLCELL_X4 FILLER_33_230 ();
 FILLCELL_X2 FILLER_33_234 ();
 FILLCELL_X4 FILLER_33_240 ();
 FILLCELL_X4 FILLER_33_253 ();
 FILLCELL_X8 FILLER_33_266 ();
 FILLCELL_X2 FILLER_33_274 ();
 FILLCELL_X4 FILLER_33_280 ();
 FILLCELL_X4 FILLER_33_293 ();
 FILLCELL_X4 FILLER_33_306 ();
 FILLCELL_X4 FILLER_33_314 ();
 FILLCELL_X16 FILLER_33_321 ();
 FILLCELL_X8 FILLER_33_337 ();
 FILLCELL_X4 FILLER_33_345 ();
 FILLCELL_X1 FILLER_33_349 ();
 FILLCELL_X4 FILLER_33_355 ();
 FILLCELL_X4 FILLER_33_362 ();
 FILLCELL_X2 FILLER_33_366 ();
 FILLCELL_X1 FILLER_33_368 ();
 FILLCELL_X4 FILLER_33_373 ();
 FILLCELL_X4 FILLER_33_381 ();
 FILLCELL_X2 FILLER_33_385 ();
 FILLCELL_X1 FILLER_33_387 ();
 FILLCELL_X4 FILLER_33_392 ();
 FILLCELL_X4 FILLER_33_400 ();
 FILLCELL_X4 FILLER_33_408 ();
 FILLCELL_X4 FILLER_33_416 ();
 FILLCELL_X2 FILLER_33_420 ();
 FILLCELL_X1 FILLER_33_422 ();
 FILLCELL_X4 FILLER_33_427 ();
 FILLCELL_X4 FILLER_33_435 ();
 FILLCELL_X4 FILLER_33_445 ();
 FILLCELL_X1 FILLER_33_449 ();
 FILLCELL_X4 FILLER_33_454 ();
 FILLCELL_X4 FILLER_33_462 ();
 FILLCELL_X4 FILLER_33_472 ();
 FILLCELL_X4 FILLER_33_485 ();
 FILLCELL_X8 FILLER_33_493 ();
 FILLCELL_X8 FILLER_33_510 ();
 FILLCELL_X1 FILLER_33_518 ();
 FILLCELL_X4 FILLER_33_528 ();
 FILLCELL_X1 FILLER_33_532 ();
 FILLCELL_X4 FILLER_33_539 ();
 FILLCELL_X8 FILLER_33_546 ();
 FILLCELL_X1 FILLER_33_554 ();
 FILLCELL_X4 FILLER_33_559 ();
 FILLCELL_X4 FILLER_33_567 ();
 FILLCELL_X4 FILLER_33_574 ();
 FILLCELL_X8 FILLER_33_581 ();
 FILLCELL_X8 FILLER_33_593 ();
 FILLCELL_X2 FILLER_33_601 ();
 FILLCELL_X1 FILLER_33_603 ();
 FILLCELL_X8 FILLER_33_607 ();
 FILLCELL_X8 FILLER_33_620 ();
 FILLCELL_X1 FILLER_33_628 ();
 FILLCELL_X4 FILLER_33_648 ();
 FILLCELL_X1 FILLER_33_652 ();
 FILLCELL_X4 FILLER_33_657 ();
 FILLCELL_X4 FILLER_33_680 ();
 FILLCELL_X4 FILLER_33_703 ();
 FILLCELL_X8 FILLER_33_726 ();
 FILLCELL_X2 FILLER_33_734 ();
 FILLCELL_X1 FILLER_33_736 ();
 FILLCELL_X16 FILLER_33_742 ();
 FILLCELL_X8 FILLER_33_758 ();
 FILLCELL_X2 FILLER_33_766 ();
 FILLCELL_X1 FILLER_33_768 ();
 FILLCELL_X8 FILLER_33_788 ();
 FILLCELL_X8 FILLER_33_815 ();
 FILLCELL_X4 FILLER_33_832 ();
 FILLCELL_X8 FILLER_33_842 ();
 FILLCELL_X2 FILLER_33_850 ();
 FILLCELL_X4 FILLER_33_859 ();
 FILLCELL_X8 FILLER_33_866 ();
 FILLCELL_X4 FILLER_33_874 ();
 FILLCELL_X1 FILLER_33_878 ();
 FILLCELL_X16 FILLER_33_882 ();
 FILLCELL_X2 FILLER_33_898 ();
 FILLCELL_X4 FILLER_33_909 ();
 FILLCELL_X8 FILLER_33_922 ();
 FILLCELL_X4 FILLER_33_939 ();
 FILLCELL_X8 FILLER_33_952 ();
 FILLCELL_X4 FILLER_33_966 ();
 FILLCELL_X16 FILLER_33_975 ();
 FILLCELL_X2 FILLER_33_991 ();
 FILLCELL_X1 FILLER_33_993 ();
 FILLCELL_X4 FILLER_33_1000 ();
 FILLCELL_X4 FILLER_33_1013 ();
 FILLCELL_X4 FILLER_33_1026 ();
 FILLCELL_X2 FILLER_33_1030 ();
 FILLCELL_X1 FILLER_33_1032 ();
 FILLCELL_X4 FILLER_33_1037 ();
 FILLCELL_X4 FILLER_33_1051 ();
 FILLCELL_X4 FILLER_33_1064 ();
 FILLCELL_X8 FILLER_33_1077 ();
 FILLCELL_X2 FILLER_33_1085 ();
 FILLCELL_X1 FILLER_33_1087 ();
 FILLCELL_X4 FILLER_33_1094 ();
 FILLCELL_X4 FILLER_33_1102 ();
 FILLCELL_X4 FILLER_33_1110 ();
 FILLCELL_X2 FILLER_33_1114 ();
 FILLCELL_X4 FILLER_33_1125 ();
 FILLCELL_X4 FILLER_33_1138 ();
 FILLCELL_X4 FILLER_33_1148 ();
 FILLCELL_X8 FILLER_33_1157 ();
 FILLCELL_X4 FILLER_33_1165 ();
 FILLCELL_X2 FILLER_33_1169 ();
 FILLCELL_X4 FILLER_33_1175 ();
 FILLCELL_X2 FILLER_33_1179 ();
 FILLCELL_X1 FILLER_33_1181 ();
 FILLCELL_X4 FILLER_33_1191 ();
 FILLCELL_X4 FILLER_33_1198 ();
 FILLCELL_X16 FILLER_33_1205 ();
 FILLCELL_X8 FILLER_33_1221 ();
 FILLCELL_X1 FILLER_33_1229 ();
 FILLCELL_X8 FILLER_33_1234 ();
 FILLCELL_X2 FILLER_33_1242 ();
 FILLCELL_X1 FILLER_33_1244 ();
 FILLCELL_X8 FILLER_33_1254 ();
 FILLCELL_X1 FILLER_33_1262 ();
 FILLCELL_X4 FILLER_33_1264 ();
 FILLCELL_X4 FILLER_33_1271 ();
 FILLCELL_X2 FILLER_33_1275 ();
 FILLCELL_X1 FILLER_33_1277 ();
 FILLCELL_X4 FILLER_33_1280 ();
 FILLCELL_X2 FILLER_33_1284 ();
 FILLCELL_X4 FILLER_33_1290 ();
 FILLCELL_X1 FILLER_33_1294 ();
 FILLCELL_X4 FILLER_33_1298 ();
 FILLCELL_X4 FILLER_33_1308 ();
 FILLCELL_X4 FILLER_33_1319 ();
 FILLCELL_X8 FILLER_33_1329 ();
 FILLCELL_X4 FILLER_33_1347 ();
 FILLCELL_X4 FILLER_33_1358 ();
 FILLCELL_X4 FILLER_33_1366 ();
 FILLCELL_X4 FILLER_33_1374 ();
 FILLCELL_X8 FILLER_33_1380 ();
 FILLCELL_X32 FILLER_33_1391 ();
 FILLCELL_X32 FILLER_33_1423 ();
 FILLCELL_X32 FILLER_33_1455 ();
 FILLCELL_X32 FILLER_33_1487 ();
 FILLCELL_X32 FILLER_33_1519 ();
 FILLCELL_X32 FILLER_33_1551 ();
 FILLCELL_X32 FILLER_33_1583 ();
 FILLCELL_X32 FILLER_33_1615 ();
 FILLCELL_X32 FILLER_33_1647 ();
 FILLCELL_X32 FILLER_33_1679 ();
 FILLCELL_X32 FILLER_33_1711 ();
 FILLCELL_X8 FILLER_33_1743 ();
 FILLCELL_X4 FILLER_33_1751 ();
 FILLCELL_X1 FILLER_33_1755 ();
 FILLCELL_X4 FILLER_34_1 ();
 FILLCELL_X4 FILLER_34_24 ();
 FILLCELL_X4 FILLER_34_38 ();
 FILLCELL_X4 FILLER_34_45 ();
 FILLCELL_X2 FILLER_34_49 ();
 FILLCELL_X1 FILLER_34_51 ();
 FILLCELL_X4 FILLER_34_61 ();
 FILLCELL_X4 FILLER_34_68 ();
 FILLCELL_X4 FILLER_34_76 ();
 FILLCELL_X4 FILLER_34_84 ();
 FILLCELL_X4 FILLER_34_97 ();
 FILLCELL_X4 FILLER_34_105 ();
 FILLCELL_X2 FILLER_34_109 ();
 FILLCELL_X1 FILLER_34_111 ();
 FILLCELL_X4 FILLER_34_116 ();
 FILLCELL_X8 FILLER_34_123 ();
 FILLCELL_X2 FILLER_34_131 ();
 FILLCELL_X4 FILLER_34_137 ();
 FILLCELL_X4 FILLER_34_145 ();
 FILLCELL_X8 FILLER_34_152 ();
 FILLCELL_X2 FILLER_34_160 ();
 FILLCELL_X1 FILLER_34_162 ();
 FILLCELL_X4 FILLER_34_173 ();
 FILLCELL_X2 FILLER_34_177 ();
 FILLCELL_X1 FILLER_34_179 ();
 FILLCELL_X8 FILLER_34_190 ();
 FILLCELL_X1 FILLER_34_198 ();
 FILLCELL_X8 FILLER_34_209 ();
 FILLCELL_X4 FILLER_34_217 ();
 FILLCELL_X2 FILLER_34_221 ();
 FILLCELL_X4 FILLER_34_232 ();
 FILLCELL_X16 FILLER_34_240 ();
 FILLCELL_X4 FILLER_34_256 ();
 FILLCELL_X1 FILLER_34_260 ();
 FILLCELL_X4 FILLER_34_265 ();
 FILLCELL_X16 FILLER_34_272 ();
 FILLCELL_X8 FILLER_34_288 ();
 FILLCELL_X2 FILLER_34_296 ();
 FILLCELL_X4 FILLER_34_304 ();
 FILLCELL_X8 FILLER_34_313 ();
 FILLCELL_X1 FILLER_34_321 ();
 FILLCELL_X4 FILLER_34_331 ();
 FILLCELL_X16 FILLER_34_338 ();
 FILLCELL_X1 FILLER_34_354 ();
 FILLCELL_X4 FILLER_34_358 ();
 FILLCELL_X4 FILLER_34_366 ();
 FILLCELL_X8 FILLER_34_379 ();
 FILLCELL_X1 FILLER_34_387 ();
 FILLCELL_X4 FILLER_34_397 ();
 FILLCELL_X8 FILLER_34_410 ();
 FILLCELL_X4 FILLER_34_422 ();
 FILLCELL_X8 FILLER_34_435 ();
 FILLCELL_X4 FILLER_34_443 ();
 FILLCELL_X8 FILLER_34_456 ();
 FILLCELL_X2 FILLER_34_464 ();
 FILLCELL_X1 FILLER_34_466 ();
 FILLCELL_X4 FILLER_34_472 ();
 FILLCELL_X8 FILLER_34_485 ();
 FILLCELL_X8 FILLER_34_496 ();
 FILLCELL_X1 FILLER_34_504 ();
 FILLCELL_X4 FILLER_34_508 ();
 FILLCELL_X16 FILLER_34_516 ();
 FILLCELL_X2 FILLER_34_532 ();
 FILLCELL_X8 FILLER_34_539 ();
 FILLCELL_X2 FILLER_34_547 ();
 FILLCELL_X4 FILLER_34_555 ();
 FILLCELL_X4 FILLER_34_568 ();
 FILLCELL_X1 FILLER_34_572 ();
 FILLCELL_X4 FILLER_34_577 ();
 FILLCELL_X4 FILLER_34_585 ();
 FILLCELL_X8 FILLER_34_593 ();
 FILLCELL_X4 FILLER_34_601 ();
 FILLCELL_X2 FILLER_34_605 ();
 FILLCELL_X1 FILLER_34_607 ();
 FILLCELL_X16 FILLER_34_612 ();
 FILLCELL_X2 FILLER_34_628 ();
 FILLCELL_X1 FILLER_34_630 ();
 FILLCELL_X4 FILLER_34_632 ();
 FILLCELL_X8 FILLER_34_640 ();
 FILLCELL_X4 FILLER_34_648 ();
 FILLCELL_X4 FILLER_34_671 ();
 FILLCELL_X8 FILLER_34_679 ();
 FILLCELL_X4 FILLER_34_687 ();
 FILLCELL_X8 FILLER_34_695 ();
 FILLCELL_X4 FILLER_34_703 ();
 FILLCELL_X2 FILLER_34_707 ();
 FILLCELL_X1 FILLER_34_709 ();
 FILLCELL_X4 FILLER_34_729 ();
 FILLCELL_X4 FILLER_34_752 ();
 FILLCELL_X8 FILLER_34_775 ();
 FILLCELL_X2 FILLER_34_783 ();
 FILLCELL_X1 FILLER_34_785 ();
 FILLCELL_X4 FILLER_34_805 ();
 FILLCELL_X2 FILLER_34_809 ();
 FILLCELL_X1 FILLER_34_811 ();
 FILLCELL_X4 FILLER_34_816 ();
 FILLCELL_X4 FILLER_34_825 ();
 FILLCELL_X8 FILLER_34_832 ();
 FILLCELL_X2 FILLER_34_840 ();
 FILLCELL_X1 FILLER_34_842 ();
 FILLCELL_X8 FILLER_34_862 ();
 FILLCELL_X4 FILLER_34_879 ();
 FILLCELL_X2 FILLER_34_883 ();
 FILLCELL_X4 FILLER_34_888 ();
 FILLCELL_X4 FILLER_34_895 ();
 FILLCELL_X4 FILLER_34_905 ();
 FILLCELL_X4 FILLER_34_913 ();
 FILLCELL_X4 FILLER_34_920 ();
 FILLCELL_X4 FILLER_34_928 ();
 FILLCELL_X8 FILLER_34_937 ();
 FILLCELL_X2 FILLER_34_945 ();
 FILLCELL_X1 FILLER_34_947 ();
 FILLCELL_X4 FILLER_34_953 ();
 FILLCELL_X4 FILLER_34_961 ();
 FILLCELL_X2 FILLER_34_965 ();
 FILLCELL_X1 FILLER_34_967 ();
 FILLCELL_X4 FILLER_34_971 ();
 FILLCELL_X4 FILLER_34_981 ();
 FILLCELL_X8 FILLER_34_990 ();
 FILLCELL_X4 FILLER_34_998 ();
 FILLCELL_X4 FILLER_34_1007 ();
 FILLCELL_X1 FILLER_34_1011 ();
 FILLCELL_X16 FILLER_34_1016 ();
 FILLCELL_X4 FILLER_34_1035 ();
 FILLCELL_X32 FILLER_34_1048 ();
 FILLCELL_X4 FILLER_34_1080 ();
 FILLCELL_X4 FILLER_34_1093 ();
 FILLCELL_X8 FILLER_34_1106 ();
 FILLCELL_X1 FILLER_34_1114 ();
 FILLCELL_X4 FILLER_34_1119 ();
 FILLCELL_X16 FILLER_34_1127 ();
 FILLCELL_X4 FILLER_34_1143 ();
 FILLCELL_X2 FILLER_34_1147 ();
 FILLCELL_X1 FILLER_34_1149 ();
 FILLCELL_X16 FILLER_34_1155 ();
 FILLCELL_X2 FILLER_34_1171 ();
 FILLCELL_X4 FILLER_34_1178 ();
 FILLCELL_X2 FILLER_34_1182 ();
 FILLCELL_X1 FILLER_34_1184 ();
 FILLCELL_X8 FILLER_34_1190 ();
 FILLCELL_X2 FILLER_34_1198 ();
 FILLCELL_X1 FILLER_34_1200 ();
 FILLCELL_X4 FILLER_34_1204 ();
 FILLCELL_X4 FILLER_34_1217 ();
 FILLCELL_X2 FILLER_34_1221 ();
 FILLCELL_X1 FILLER_34_1223 ();
 FILLCELL_X4 FILLER_34_1229 ();
 FILLCELL_X4 FILLER_34_1242 ();
 FILLCELL_X4 FILLER_34_1252 ();
 FILLCELL_X4 FILLER_34_1261 ();
 FILLCELL_X8 FILLER_34_1269 ();
 FILLCELL_X4 FILLER_34_1277 ();
 FILLCELL_X2 FILLER_34_1281 ();
 FILLCELL_X1 FILLER_34_1283 ();
 FILLCELL_X4 FILLER_34_1288 ();
 FILLCELL_X4 FILLER_34_1296 ();
 FILLCELL_X2 FILLER_34_1300 ();
 FILLCELL_X1 FILLER_34_1302 ();
 FILLCELL_X4 FILLER_34_1309 ();
 FILLCELL_X8 FILLER_34_1317 ();
 FILLCELL_X1 FILLER_34_1325 ();
 FILLCELL_X4 FILLER_34_1329 ();
 FILLCELL_X4 FILLER_34_1343 ();
 FILLCELL_X4 FILLER_34_1349 ();
 FILLCELL_X4 FILLER_34_1355 ();
 FILLCELL_X2 FILLER_34_1359 ();
 FILLCELL_X4 FILLER_34_1367 ();
 FILLCELL_X2 FILLER_34_1371 ();
 FILLCELL_X4 FILLER_34_1379 ();
 FILLCELL_X32 FILLER_34_1385 ();
 FILLCELL_X32 FILLER_34_1417 ();
 FILLCELL_X32 FILLER_34_1449 ();
 FILLCELL_X32 FILLER_34_1481 ();
 FILLCELL_X32 FILLER_34_1513 ();
 FILLCELL_X32 FILLER_34_1545 ();
 FILLCELL_X32 FILLER_34_1577 ();
 FILLCELL_X32 FILLER_34_1609 ();
 FILLCELL_X32 FILLER_34_1641 ();
 FILLCELL_X32 FILLER_34_1673 ();
 FILLCELL_X32 FILLER_34_1705 ();
 FILLCELL_X16 FILLER_34_1737 ();
 FILLCELL_X2 FILLER_34_1753 ();
 FILLCELL_X1 FILLER_34_1755 ();
 FILLCELL_X4 FILLER_35_1 ();
 FILLCELL_X2 FILLER_35_5 ();
 FILLCELL_X1 FILLER_35_7 ();
 FILLCELL_X32 FILLER_35_12 ();
 FILLCELL_X8 FILLER_35_44 ();
 FILLCELL_X32 FILLER_35_57 ();
 FILLCELL_X4 FILLER_35_89 ();
 FILLCELL_X1 FILLER_35_93 ();
 FILLCELL_X4 FILLER_35_97 ();
 FILLCELL_X4 FILLER_35_104 ();
 FILLCELL_X2 FILLER_35_108 ();
 FILLCELL_X4 FILLER_35_112 ();
 FILLCELL_X32 FILLER_35_123 ();
 FILLCELL_X2 FILLER_35_155 ();
 FILLCELL_X4 FILLER_35_160 ();
 FILLCELL_X2 FILLER_35_164 ();
 FILLCELL_X4 FILLER_35_168 ();
 FILLCELL_X4 FILLER_35_176 ();
 FILLCELL_X4 FILLER_35_187 ();
 FILLCELL_X2 FILLER_35_191 ();
 FILLCELL_X1 FILLER_35_193 ();
 FILLCELL_X4 FILLER_35_197 ();
 FILLCELL_X32 FILLER_35_205 ();
 FILLCELL_X4 FILLER_35_237 ();
 FILLCELL_X1 FILLER_35_241 ();
 FILLCELL_X16 FILLER_35_246 ();
 FILLCELL_X2 FILLER_35_262 ();
 FILLCELL_X1 FILLER_35_264 ();
 FILLCELL_X4 FILLER_35_269 ();
 FILLCELL_X4 FILLER_35_277 ();
 FILLCELL_X16 FILLER_35_285 ();
 FILLCELL_X8 FILLER_35_301 ();
 FILLCELL_X4 FILLER_35_309 ();
 FILLCELL_X4 FILLER_35_319 ();
 FILLCELL_X2 FILLER_35_323 ();
 FILLCELL_X4 FILLER_35_329 ();
 FILLCELL_X8 FILLER_35_336 ();
 FILLCELL_X4 FILLER_35_353 ();
 FILLCELL_X2 FILLER_35_357 ();
 FILLCELL_X4 FILLER_35_363 ();
 FILLCELL_X4 FILLER_35_372 ();
 FILLCELL_X4 FILLER_35_380 ();
 FILLCELL_X8 FILLER_35_388 ();
 FILLCELL_X4 FILLER_35_405 ();
 FILLCELL_X4 FILLER_35_415 ();
 FILLCELL_X1 FILLER_35_419 ();
 FILLCELL_X8 FILLER_35_423 ();
 FILLCELL_X4 FILLER_35_440 ();
 FILLCELL_X1 FILLER_35_444 ();
 FILLCELL_X16 FILLER_35_450 ();
 FILLCELL_X4 FILLER_35_466 ();
 FILLCELL_X8 FILLER_35_475 ();
 FILLCELL_X2 FILLER_35_483 ();
 FILLCELL_X4 FILLER_35_490 ();
 FILLCELL_X4 FILLER_35_499 ();
 FILLCELL_X4 FILLER_35_509 ();
 FILLCELL_X8 FILLER_35_518 ();
 FILLCELL_X4 FILLER_35_526 ();
 FILLCELL_X1 FILLER_35_530 ();
 FILLCELL_X8 FILLER_35_540 ();
 FILLCELL_X2 FILLER_35_548 ();
 FILLCELL_X1 FILLER_35_550 ();
 FILLCELL_X4 FILLER_35_556 ();
 FILLCELL_X4 FILLER_35_565 ();
 FILLCELL_X4 FILLER_35_573 ();
 FILLCELL_X2 FILLER_35_577 ();
 FILLCELL_X1 FILLER_35_579 ();
 FILLCELL_X8 FILLER_35_589 ();
 FILLCELL_X4 FILLER_35_597 ();
 FILLCELL_X2 FILLER_35_601 ();
 FILLCELL_X1 FILLER_35_603 ();
 FILLCELL_X32 FILLER_35_623 ();
 FILLCELL_X16 FILLER_35_655 ();
 FILLCELL_X8 FILLER_35_671 ();
 FILLCELL_X2 FILLER_35_679 ();
 FILLCELL_X1 FILLER_35_681 ();
 FILLCELL_X32 FILLER_35_701 ();
 FILLCELL_X4 FILLER_35_733 ();
 FILLCELL_X4 FILLER_35_742 ();
 FILLCELL_X4 FILLER_35_750 ();
 FILLCELL_X1 FILLER_35_754 ();
 FILLCELL_X16 FILLER_35_759 ();
 FILLCELL_X2 FILLER_35_775 ();
 FILLCELL_X4 FILLER_35_781 ();
 FILLCELL_X16 FILLER_35_789 ();
 FILLCELL_X2 FILLER_35_805 ();
 FILLCELL_X32 FILLER_35_811 ();
 FILLCELL_X2 FILLER_35_843 ();
 FILLCELL_X1 FILLER_35_845 ();
 FILLCELL_X8 FILLER_35_850 ();
 FILLCELL_X4 FILLER_35_858 ();
 FILLCELL_X4 FILLER_35_869 ();
 FILLCELL_X4 FILLER_35_883 ();
 FILLCELL_X4 FILLER_35_891 ();
 FILLCELL_X1 FILLER_35_895 ();
 FILLCELL_X4 FILLER_35_899 ();
 FILLCELL_X8 FILLER_35_907 ();
 FILLCELL_X4 FILLER_35_915 ();
 FILLCELL_X2 FILLER_35_919 ();
 FILLCELL_X1 FILLER_35_921 ();
 FILLCELL_X4 FILLER_35_926 ();
 FILLCELL_X8 FILLER_35_935 ();
 FILLCELL_X4 FILLER_35_948 ();
 FILLCELL_X8 FILLER_35_961 ();
 FILLCELL_X2 FILLER_35_969 ();
 FILLCELL_X4 FILLER_35_975 ();
 FILLCELL_X4 FILLER_35_988 ();
 FILLCELL_X4 FILLER_35_996 ();
 FILLCELL_X4 FILLER_35_1004 ();
 FILLCELL_X2 FILLER_35_1008 ();
 FILLCELL_X8 FILLER_35_1013 ();
 FILLCELL_X4 FILLER_35_1021 ();
 FILLCELL_X8 FILLER_35_1029 ();
 FILLCELL_X2 FILLER_35_1037 ();
 FILLCELL_X4 FILLER_35_1043 ();
 FILLCELL_X4 FILLER_35_1051 ();
 FILLCELL_X4 FILLER_35_1064 ();
 FILLCELL_X4 FILLER_35_1074 ();
 FILLCELL_X8 FILLER_35_1081 ();
 FILLCELL_X2 FILLER_35_1089 ();
 FILLCELL_X4 FILLER_35_1096 ();
 FILLCELL_X4 FILLER_35_1103 ();
 FILLCELL_X2 FILLER_35_1107 ();
 FILLCELL_X4 FILLER_35_1113 ();
 FILLCELL_X8 FILLER_35_1120 ();
 FILLCELL_X4 FILLER_35_1128 ();
 FILLCELL_X1 FILLER_35_1132 ();
 FILLCELL_X4 FILLER_35_1136 ();
 FILLCELL_X2 FILLER_35_1140 ();
 FILLCELL_X4 FILLER_35_1145 ();
 FILLCELL_X4 FILLER_35_1158 ();
 FILLCELL_X4 FILLER_35_1166 ();
 FILLCELL_X8 FILLER_35_1174 ();
 FILLCELL_X2 FILLER_35_1182 ();
 FILLCELL_X1 FILLER_35_1184 ();
 FILLCELL_X4 FILLER_35_1194 ();
 FILLCELL_X4 FILLER_35_1201 ();
 FILLCELL_X4 FILLER_35_1208 ();
 FILLCELL_X4 FILLER_35_1215 ();
 FILLCELL_X8 FILLER_35_1222 ();
 FILLCELL_X1 FILLER_35_1230 ();
 FILLCELL_X4 FILLER_35_1235 ();
 FILLCELL_X8 FILLER_35_1244 ();
 FILLCELL_X2 FILLER_35_1252 ();
 FILLCELL_X1 FILLER_35_1254 ();
 FILLCELL_X4 FILLER_35_1259 ();
 FILLCELL_X4 FILLER_35_1264 ();
 FILLCELL_X4 FILLER_35_1285 ();
 FILLCELL_X8 FILLER_35_1298 ();
 FILLCELL_X4 FILLER_35_1306 ();
 FILLCELL_X1 FILLER_35_1310 ();
 FILLCELL_X4 FILLER_35_1318 ();
 FILLCELL_X4 FILLER_35_1328 ();
 FILLCELL_X2 FILLER_35_1332 ();
 FILLCELL_X32 FILLER_35_1338 ();
 FILLCELL_X4 FILLER_35_1370 ();
 FILLCELL_X1 FILLER_35_1374 ();
 FILLCELL_X4 FILLER_35_1379 ();
 FILLCELL_X32 FILLER_35_1402 ();
 FILLCELL_X32 FILLER_35_1434 ();
 FILLCELL_X32 FILLER_35_1466 ();
 FILLCELL_X32 FILLER_35_1498 ();
 FILLCELL_X32 FILLER_35_1530 ();
 FILLCELL_X32 FILLER_35_1562 ();
 FILLCELL_X32 FILLER_35_1594 ();
 FILLCELL_X32 FILLER_35_1626 ();
 FILLCELL_X32 FILLER_35_1658 ();
 FILLCELL_X32 FILLER_35_1690 ();
 FILLCELL_X32 FILLER_35_1722 ();
 FILLCELL_X2 FILLER_35_1754 ();
 FILLCELL_X8 FILLER_36_1 ();
 FILLCELL_X4 FILLER_36_9 ();
 FILLCELL_X2 FILLER_36_13 ();
 FILLCELL_X4 FILLER_36_19 ();
 FILLCELL_X8 FILLER_36_32 ();
 FILLCELL_X2 FILLER_36_40 ();
 FILLCELL_X1 FILLER_36_42 ();
 FILLCELL_X4 FILLER_36_60 ();
 FILLCELL_X4 FILLER_36_69 ();
 FILLCELL_X4 FILLER_36_77 ();
 FILLCELL_X2 FILLER_36_81 ();
 FILLCELL_X4 FILLER_36_87 ();
 FILLCELL_X1 FILLER_36_91 ();
 FILLCELL_X4 FILLER_36_101 ();
 FILLCELL_X4 FILLER_36_108 ();
 FILLCELL_X2 FILLER_36_112 ();
 FILLCELL_X16 FILLER_36_124 ();
 FILLCELL_X4 FILLER_36_144 ();
 FILLCELL_X2 FILLER_36_148 ();
 FILLCELL_X1 FILLER_36_150 ();
 FILLCELL_X4 FILLER_36_155 ();
 FILLCELL_X4 FILLER_36_162 ();
 FILLCELL_X8 FILLER_36_169 ();
 FILLCELL_X4 FILLER_36_177 ();
 FILLCELL_X4 FILLER_36_185 ();
 FILLCELL_X8 FILLER_36_193 ();
 FILLCELL_X4 FILLER_36_201 ();
 FILLCELL_X2 FILLER_36_205 ();
 FILLCELL_X4 FILLER_36_211 ();
 FILLCELL_X8 FILLER_36_219 ();
 FILLCELL_X4 FILLER_36_231 ();
 FILLCELL_X2 FILLER_36_235 ();
 FILLCELL_X4 FILLER_36_241 ();
 FILLCELL_X2 FILLER_36_245 ();
 FILLCELL_X8 FILLER_36_256 ();
 FILLCELL_X2 FILLER_36_264 ();
 FILLCELL_X1 FILLER_36_266 ();
 FILLCELL_X4 FILLER_36_271 ();
 FILLCELL_X2 FILLER_36_275 ();
 FILLCELL_X1 FILLER_36_277 ();
 FILLCELL_X8 FILLER_36_287 ();
 FILLCELL_X4 FILLER_36_295 ();
 FILLCELL_X1 FILLER_36_299 ();
 FILLCELL_X4 FILLER_36_303 ();
 FILLCELL_X4 FILLER_36_316 ();
 FILLCELL_X8 FILLER_36_325 ();
 FILLCELL_X1 FILLER_36_333 ();
 FILLCELL_X4 FILLER_36_340 ();
 FILLCELL_X4 FILLER_36_353 ();
 FILLCELL_X1 FILLER_36_357 ();
 FILLCELL_X4 FILLER_36_361 ();
 FILLCELL_X16 FILLER_36_374 ();
 FILLCELL_X4 FILLER_36_390 ();
 FILLCELL_X4 FILLER_36_399 ();
 FILLCELL_X8 FILLER_36_406 ();
 FILLCELL_X2 FILLER_36_414 ();
 FILLCELL_X1 FILLER_36_416 ();
 FILLCELL_X4 FILLER_36_422 ();
 FILLCELL_X1 FILLER_36_426 ();
 FILLCELL_X4 FILLER_36_432 ();
 FILLCELL_X4 FILLER_36_439 ();
 FILLCELL_X2 FILLER_36_443 ();
 FILLCELL_X8 FILLER_36_449 ();
 FILLCELL_X1 FILLER_36_457 ();
 FILLCELL_X4 FILLER_36_461 ();
 FILLCELL_X8 FILLER_36_469 ();
 FILLCELL_X4 FILLER_36_483 ();
 FILLCELL_X8 FILLER_36_490 ();
 FILLCELL_X1 FILLER_36_498 ();
 FILLCELL_X4 FILLER_36_503 ();
 FILLCELL_X8 FILLER_36_516 ();
 FILLCELL_X4 FILLER_36_529 ();
 FILLCELL_X4 FILLER_36_542 ();
 FILLCELL_X4 FILLER_36_550 ();
 FILLCELL_X2 FILLER_36_554 ();
 FILLCELL_X1 FILLER_36_556 ();
 FILLCELL_X16 FILLER_36_566 ();
 FILLCELL_X2 FILLER_36_582 ();
 FILLCELL_X1 FILLER_36_584 ();
 FILLCELL_X4 FILLER_36_604 ();
 FILLCELL_X4 FILLER_36_627 ();
 FILLCELL_X4 FILLER_36_632 ();
 FILLCELL_X4 FILLER_36_655 ();
 FILLCELL_X4 FILLER_36_678 ();
 FILLCELL_X4 FILLER_36_687 ();
 FILLCELL_X8 FILLER_36_695 ();
 FILLCELL_X4 FILLER_36_703 ();
 FILLCELL_X1 FILLER_36_707 ();
 FILLCELL_X8 FILLER_36_712 ();
 FILLCELL_X1 FILLER_36_720 ();
 FILLCELL_X8 FILLER_36_725 ();
 FILLCELL_X4 FILLER_36_733 ();
 FILLCELL_X4 FILLER_36_756 ();
 FILLCELL_X16 FILLER_36_779 ();
 FILLCELL_X8 FILLER_36_795 ();
 FILLCELL_X4 FILLER_36_803 ();
 FILLCELL_X2 FILLER_36_807 ();
 FILLCELL_X4 FILLER_36_828 ();
 FILLCELL_X1 FILLER_36_832 ();
 FILLCELL_X4 FILLER_36_837 ();
 FILLCELL_X4 FILLER_36_847 ();
 FILLCELL_X1 FILLER_36_851 ();
 FILLCELL_X8 FILLER_36_858 ();
 FILLCELL_X1 FILLER_36_866 ();
 FILLCELL_X4 FILLER_36_870 ();
 FILLCELL_X4 FILLER_36_877 ();
 FILLCELL_X4 FILLER_36_888 ();
 FILLCELL_X4 FILLER_36_898 ();
 FILLCELL_X8 FILLER_36_906 ();
 FILLCELL_X4 FILLER_36_920 ();
 FILLCELL_X4 FILLER_36_933 ();
 FILLCELL_X1 FILLER_36_937 ();
 FILLCELL_X4 FILLER_36_944 ();
 FILLCELL_X4 FILLER_36_957 ();
 FILLCELL_X4 FILLER_36_970 ();
 FILLCELL_X4 FILLER_36_979 ();
 FILLCELL_X1 FILLER_36_983 ();
 FILLCELL_X4 FILLER_36_988 ();
 FILLCELL_X8 FILLER_36_995 ();
 FILLCELL_X4 FILLER_36_1003 ();
 FILLCELL_X1 FILLER_36_1007 ();
 FILLCELL_X4 FILLER_36_1012 ();
 FILLCELL_X4 FILLER_36_1020 ();
 FILLCELL_X1 FILLER_36_1024 ();
 FILLCELL_X4 FILLER_36_1034 ();
 FILLCELL_X4 FILLER_36_1044 ();
 FILLCELL_X4 FILLER_36_1051 ();
 FILLCELL_X4 FILLER_36_1060 ();
 FILLCELL_X4 FILLER_36_1073 ();
 FILLCELL_X4 FILLER_36_1081 ();
 FILLCELL_X8 FILLER_36_1088 ();
 FILLCELL_X4 FILLER_36_1096 ();
 FILLCELL_X2 FILLER_36_1100 ();
 FILLCELL_X8 FILLER_36_1106 ();
 FILLCELL_X2 FILLER_36_1114 ();
 FILLCELL_X1 FILLER_36_1116 ();
 FILLCELL_X4 FILLER_36_1123 ();
 FILLCELL_X8 FILLER_36_1130 ();
 FILLCELL_X2 FILLER_36_1138 ();
 FILLCELL_X4 FILLER_36_1149 ();
 FILLCELL_X2 FILLER_36_1153 ();
 FILLCELL_X1 FILLER_36_1155 ();
 FILLCELL_X4 FILLER_36_1160 ();
 FILLCELL_X2 FILLER_36_1164 ();
 FILLCELL_X4 FILLER_36_1171 ();
 FILLCELL_X4 FILLER_36_1179 ();
 FILLCELL_X4 FILLER_36_1187 ();
 FILLCELL_X4 FILLER_36_1194 ();
 FILLCELL_X4 FILLER_36_1201 ();
 FILLCELL_X1 FILLER_36_1205 ();
 FILLCELL_X4 FILLER_36_1212 ();
 FILLCELL_X4 FILLER_36_1220 ();
 FILLCELL_X16 FILLER_36_1228 ();
 FILLCELL_X1 FILLER_36_1244 ();
 FILLCELL_X8 FILLER_36_1254 ();
 FILLCELL_X1 FILLER_36_1262 ();
 FILLCELL_X4 FILLER_36_1268 ();
 FILLCELL_X4 FILLER_36_1276 ();
 FILLCELL_X2 FILLER_36_1280 ();
 FILLCELL_X1 FILLER_36_1282 ();
 FILLCELL_X4 FILLER_36_1287 ();
 FILLCELL_X8 FILLER_36_1295 ();
 FILLCELL_X4 FILLER_36_1303 ();
 FILLCELL_X8 FILLER_36_1311 ();
 FILLCELL_X4 FILLER_36_1319 ();
 FILLCELL_X1 FILLER_36_1323 ();
 FILLCELL_X8 FILLER_36_1326 ();
 FILLCELL_X1 FILLER_36_1334 ();
 FILLCELL_X4 FILLER_36_1340 ();
 FILLCELL_X1 FILLER_36_1344 ();
 FILLCELL_X4 FILLER_36_1349 ();
 FILLCELL_X2 FILLER_36_1353 ();
 FILLCELL_X1 FILLER_36_1355 ();
 FILLCELL_X16 FILLER_36_1375 ();
 FILLCELL_X2 FILLER_36_1391 ();
 FILLCELL_X4 FILLER_36_1397 ();
 FILLCELL_X32 FILLER_36_1420 ();
 FILLCELL_X32 FILLER_36_1452 ();
 FILLCELL_X32 FILLER_36_1484 ();
 FILLCELL_X32 FILLER_36_1520 ();
 FILLCELL_X32 FILLER_36_1552 ();
 FILLCELL_X32 FILLER_36_1584 ();
 FILLCELL_X32 FILLER_36_1616 ();
 FILLCELL_X32 FILLER_36_1648 ();
 FILLCELL_X32 FILLER_36_1680 ();
 FILLCELL_X32 FILLER_36_1712 ();
 FILLCELL_X8 FILLER_36_1744 ();
 FILLCELL_X4 FILLER_36_1752 ();
 FILLCELL_X16 FILLER_37_1 ();
 FILLCELL_X4 FILLER_37_17 ();
 FILLCELL_X2 FILLER_37_21 ();
 FILLCELL_X4 FILLER_37_26 ();
 FILLCELL_X4 FILLER_37_33 ();
 FILLCELL_X2 FILLER_37_37 ();
 FILLCELL_X1 FILLER_37_39 ();
 FILLCELL_X4 FILLER_37_42 ();
 FILLCELL_X8 FILLER_37_53 ();
 FILLCELL_X2 FILLER_37_61 ();
 FILLCELL_X4 FILLER_37_69 ();
 FILLCELL_X16 FILLER_37_77 ();
 FILLCELL_X4 FILLER_37_97 ();
 FILLCELL_X4 FILLER_37_105 ();
 FILLCELL_X2 FILLER_37_109 ();
 FILLCELL_X1 FILLER_37_111 ();
 FILLCELL_X4 FILLER_37_116 ();
 FILLCELL_X4 FILLER_37_130 ();
 FILLCELL_X2 FILLER_37_134 ();
 FILLCELL_X4 FILLER_37_145 ();
 FILLCELL_X4 FILLER_37_158 ();
 FILLCELL_X8 FILLER_37_166 ();
 FILLCELL_X4 FILLER_37_187 ();
 FILLCELL_X2 FILLER_37_191 ();
 FILLCELL_X4 FILLER_37_202 ();
 FILLCELL_X8 FILLER_37_215 ();
 FILLCELL_X4 FILLER_37_227 ();
 FILLCELL_X8 FILLER_37_240 ();
 FILLCELL_X2 FILLER_37_248 ();
 FILLCELL_X4 FILLER_37_256 ();
 FILLCELL_X4 FILLER_37_265 ();
 FILLCELL_X4 FILLER_37_273 ();
 FILLCELL_X4 FILLER_37_286 ();
 FILLCELL_X8 FILLER_37_299 ();
 FILLCELL_X2 FILLER_37_307 ();
 FILLCELL_X8 FILLER_37_314 ();
 FILLCELL_X4 FILLER_37_322 ();
 FILLCELL_X4 FILLER_37_335 ();
 FILLCELL_X4 FILLER_37_356 ();
 FILLCELL_X2 FILLER_37_360 ();
 FILLCELL_X1 FILLER_37_362 ();
 FILLCELL_X4 FILLER_37_366 ();
 FILLCELL_X4 FILLER_37_376 ();
 FILLCELL_X8 FILLER_37_385 ();
 FILLCELL_X1 FILLER_37_393 ();
 FILLCELL_X4 FILLER_37_403 ();
 FILLCELL_X2 FILLER_37_407 ();
 FILLCELL_X4 FILLER_37_413 ();
 FILLCELL_X2 FILLER_37_417 ();
 FILLCELL_X1 FILLER_37_419 ();
 FILLCELL_X8 FILLER_37_426 ();
 FILLCELL_X8 FILLER_37_443 ();
 FILLCELL_X2 FILLER_37_451 ();
 FILLCELL_X4 FILLER_37_458 ();
 FILLCELL_X4 FILLER_37_471 ();
 FILLCELL_X4 FILLER_37_484 ();
 FILLCELL_X8 FILLER_37_492 ();
 FILLCELL_X4 FILLER_37_500 ();
 FILLCELL_X2 FILLER_37_504 ();
 FILLCELL_X1 FILLER_37_506 ();
 FILLCELL_X8 FILLER_37_516 ();
 FILLCELL_X2 FILLER_37_524 ();
 FILLCELL_X1 FILLER_37_526 ();
 FILLCELL_X4 FILLER_37_530 ();
 FILLCELL_X8 FILLER_37_543 ();
 FILLCELL_X4 FILLER_37_555 ();
 FILLCELL_X16 FILLER_37_563 ();
 FILLCELL_X2 FILLER_37_579 ();
 FILLCELL_X8 FILLER_37_585 ();
 FILLCELL_X8 FILLER_37_597 ();
 FILLCELL_X2 FILLER_37_605 ();
 FILLCELL_X4 FILLER_37_611 ();
 FILLCELL_X4 FILLER_37_634 ();
 FILLCELL_X4 FILLER_37_657 ();
 FILLCELL_X4 FILLER_37_680 ();
 FILLCELL_X4 FILLER_37_703 ();
 FILLCELL_X4 FILLER_37_726 ();
 FILLCELL_X4 FILLER_37_749 ();
 FILLCELL_X8 FILLER_37_757 ();
 FILLCELL_X1 FILLER_37_765 ();
 FILLCELL_X4 FILLER_37_785 ();
 FILLCELL_X8 FILLER_37_808 ();
 FILLCELL_X8 FILLER_37_835 ();
 FILLCELL_X1 FILLER_37_843 ();
 FILLCELL_X4 FILLER_37_857 ();
 FILLCELL_X2 FILLER_37_861 ();
 FILLCELL_X8 FILLER_37_882 ();
 FILLCELL_X2 FILLER_37_890 ();
 FILLCELL_X8 FILLER_37_898 ();
 FILLCELL_X2 FILLER_37_906 ();
 FILLCELL_X4 FILLER_37_917 ();
 FILLCELL_X4 FILLER_37_930 ();
 FILLCELL_X4 FILLER_37_938 ();
 FILLCELL_X4 FILLER_37_945 ();
 FILLCELL_X1 FILLER_37_949 ();
 FILLCELL_X8 FILLER_37_953 ();
 FILLCELL_X2 FILLER_37_961 ();
 FILLCELL_X1 FILLER_37_963 ();
 FILLCELL_X4 FILLER_37_968 ();
 FILLCELL_X8 FILLER_37_981 ();
 FILLCELL_X1 FILLER_37_989 ();
 FILLCELL_X4 FILLER_37_1009 ();
 FILLCELL_X4 FILLER_37_1017 ();
 FILLCELL_X4 FILLER_37_1030 ();
 FILLCELL_X16 FILLER_37_1037 ();
 FILLCELL_X1 FILLER_37_1053 ();
 FILLCELL_X4 FILLER_37_1058 ();
 FILLCELL_X8 FILLER_37_1066 ();
 FILLCELL_X2 FILLER_37_1074 ();
 FILLCELL_X4 FILLER_37_1095 ();
 FILLCELL_X2 FILLER_37_1099 ();
 FILLCELL_X1 FILLER_37_1101 ();
 FILLCELL_X4 FILLER_37_1106 ();
 FILLCELL_X2 FILLER_37_1110 ();
 FILLCELL_X1 FILLER_37_1112 ();
 FILLCELL_X4 FILLER_37_1122 ();
 FILLCELL_X4 FILLER_37_1135 ();
 FILLCELL_X4 FILLER_37_1143 ();
 FILLCELL_X2 FILLER_37_1147 ();
 FILLCELL_X1 FILLER_37_1149 ();
 FILLCELL_X8 FILLER_37_1154 ();
 FILLCELL_X4 FILLER_37_1171 ();
 FILLCELL_X4 FILLER_37_1184 ();
 FILLCELL_X4 FILLER_37_1194 ();
 FILLCELL_X1 FILLER_37_1198 ();
 FILLCELL_X4 FILLER_37_1208 ();
 FILLCELL_X2 FILLER_37_1212 ();
 FILLCELL_X8 FILLER_37_1223 ();
 FILLCELL_X2 FILLER_37_1231 ();
 FILLCELL_X4 FILLER_37_1238 ();
 FILLCELL_X4 FILLER_37_1259 ();
 FILLCELL_X4 FILLER_37_1264 ();
 FILLCELL_X8 FILLER_37_1277 ();
 FILLCELL_X4 FILLER_37_1285 ();
 FILLCELL_X4 FILLER_37_1292 ();
 FILLCELL_X4 FILLER_37_1302 ();
 FILLCELL_X1 FILLER_37_1306 ();
 FILLCELL_X4 FILLER_37_1313 ();
 FILLCELL_X2 FILLER_37_1317 ();
 FILLCELL_X1 FILLER_37_1319 ();
 FILLCELL_X16 FILLER_37_1324 ();
 FILLCELL_X2 FILLER_37_1340 ();
 FILLCELL_X1 FILLER_37_1342 ();
 FILLCELL_X32 FILLER_37_1362 ();
 FILLCELL_X32 FILLER_37_1394 ();
 FILLCELL_X32 FILLER_37_1426 ();
 FILLCELL_X32 FILLER_37_1458 ();
 FILLCELL_X16 FILLER_37_1490 ();
 FILLCELL_X4 FILLER_37_1506 ();
 FILLCELL_X2 FILLER_37_1510 ();
 FILLCELL_X32 FILLER_37_1531 ();
 FILLCELL_X32 FILLER_37_1563 ();
 FILLCELL_X32 FILLER_37_1595 ();
 FILLCELL_X32 FILLER_37_1627 ();
 FILLCELL_X32 FILLER_37_1659 ();
 FILLCELL_X32 FILLER_37_1691 ();
 FILLCELL_X32 FILLER_37_1723 ();
 FILLCELL_X1 FILLER_37_1755 ();
 FILLCELL_X16 FILLER_38_1 ();
 FILLCELL_X1 FILLER_38_17 ();
 FILLCELL_X4 FILLER_38_27 ();
 FILLCELL_X8 FILLER_38_34 ();
 FILLCELL_X4 FILLER_38_42 ();
 FILLCELL_X2 FILLER_38_46 ();
 FILLCELL_X1 FILLER_38_48 ();
 FILLCELL_X4 FILLER_38_53 ();
 FILLCELL_X4 FILLER_38_66 ();
 FILLCELL_X4 FILLER_38_79 ();
 FILLCELL_X1 FILLER_38_83 ();
 FILLCELL_X4 FILLER_38_88 ();
 FILLCELL_X16 FILLER_38_96 ();
 FILLCELL_X8 FILLER_38_112 ();
 FILLCELL_X2 FILLER_38_120 ();
 FILLCELL_X16 FILLER_38_125 ();
 FILLCELL_X4 FILLER_38_141 ();
 FILLCELL_X2 FILLER_38_145 ();
 FILLCELL_X4 FILLER_38_151 ();
 FILLCELL_X8 FILLER_38_159 ();
 FILLCELL_X4 FILLER_38_167 ();
 FILLCELL_X2 FILLER_38_171 ();
 FILLCELL_X4 FILLER_38_176 ();
 FILLCELL_X8 FILLER_38_183 ();
 FILLCELL_X2 FILLER_38_191 ();
 FILLCELL_X4 FILLER_38_202 ();
 FILLCELL_X4 FILLER_38_212 ();
 FILLCELL_X4 FILLER_38_221 ();
 FILLCELL_X4 FILLER_38_228 ();
 FILLCELL_X2 FILLER_38_232 ();
 FILLCELL_X1 FILLER_38_234 ();
 FILLCELL_X4 FILLER_38_238 ();
 FILLCELL_X4 FILLER_38_247 ();
 FILLCELL_X4 FILLER_38_255 ();
 FILLCELL_X8 FILLER_38_262 ();
 FILLCELL_X2 FILLER_38_270 ();
 FILLCELL_X4 FILLER_38_277 ();
 FILLCELL_X4 FILLER_38_287 ();
 FILLCELL_X4 FILLER_38_294 ();
 FILLCELL_X2 FILLER_38_298 ();
 FILLCELL_X1 FILLER_38_300 ();
 FILLCELL_X4 FILLER_38_304 ();
 FILLCELL_X4 FILLER_38_317 ();
 FILLCELL_X16 FILLER_38_324 ();
 FILLCELL_X1 FILLER_38_340 ();
 FILLCELL_X4 FILLER_38_345 ();
 FILLCELL_X8 FILLER_38_352 ();
 FILLCELL_X8 FILLER_38_369 ();
 FILLCELL_X1 FILLER_38_377 ();
 FILLCELL_X4 FILLER_38_382 ();
 FILLCELL_X4 FILLER_38_390 ();
 FILLCELL_X1 FILLER_38_394 ();
 FILLCELL_X4 FILLER_38_404 ();
 FILLCELL_X1 FILLER_38_408 ();
 FILLCELL_X8 FILLER_38_418 ();
 FILLCELL_X2 FILLER_38_426 ();
 FILLCELL_X4 FILLER_38_437 ();
 FILLCELL_X4 FILLER_38_450 ();
 FILLCELL_X4 FILLER_38_460 ();
 FILLCELL_X1 FILLER_38_464 ();
 FILLCELL_X8 FILLER_38_469 ();
 FILLCELL_X4 FILLER_38_477 ();
 FILLCELL_X4 FILLER_38_490 ();
 FILLCELL_X2 FILLER_38_494 ();
 FILLCELL_X4 FILLER_38_500 ();
 FILLCELL_X8 FILLER_38_513 ();
 FILLCELL_X1 FILLER_38_521 ();
 FILLCELL_X4 FILLER_38_526 ();
 FILLCELL_X2 FILLER_38_530 ();
 FILLCELL_X8 FILLER_38_538 ();
 FILLCELL_X4 FILLER_38_546 ();
 FILLCELL_X4 FILLER_38_569 ();
 FILLCELL_X4 FILLER_38_592 ();
 FILLCELL_X1 FILLER_38_596 ();
 FILLCELL_X4 FILLER_38_616 ();
 FILLCELL_X2 FILLER_38_620 ();
 FILLCELL_X1 FILLER_38_622 ();
 FILLCELL_X4 FILLER_38_627 ();
 FILLCELL_X4 FILLER_38_632 ();
 FILLCELL_X2 FILLER_38_636 ();
 FILLCELL_X1 FILLER_38_638 ();
 FILLCELL_X4 FILLER_38_643 ();
 FILLCELL_X1 FILLER_38_647 ();
 FILLCELL_X8 FILLER_38_652 ();
 FILLCELL_X1 FILLER_38_660 ();
 FILLCELL_X8 FILLER_38_665 ();
 FILLCELL_X2 FILLER_38_673 ();
 FILLCELL_X8 FILLER_38_679 ();
 FILLCELL_X1 FILLER_38_687 ();
 FILLCELL_X4 FILLER_38_690 ();
 FILLCELL_X4 FILLER_38_699 ();
 FILLCELL_X4 FILLER_38_707 ();
 FILLCELL_X2 FILLER_38_711 ();
 FILLCELL_X8 FILLER_38_717 ();
 FILLCELL_X4 FILLER_38_725 ();
 FILLCELL_X2 FILLER_38_729 ();
 FILLCELL_X4 FILLER_38_735 ();
 FILLCELL_X1 FILLER_38_739 ();
 FILLCELL_X16 FILLER_38_743 ();
 FILLCELL_X1 FILLER_38_759 ();
 FILLCELL_X4 FILLER_38_764 ();
 FILLCELL_X2 FILLER_38_768 ();
 FILLCELL_X16 FILLER_38_774 ();
 FILLCELL_X1 FILLER_38_790 ();
 FILLCELL_X8 FILLER_38_795 ();
 FILLCELL_X1 FILLER_38_803 ();
 FILLCELL_X4 FILLER_38_808 ();
 FILLCELL_X16 FILLER_38_816 ();
 FILLCELL_X8 FILLER_38_832 ();
 FILLCELL_X1 FILLER_38_840 ();
 FILLCELL_X8 FILLER_38_845 ();
 FILLCELL_X2 FILLER_38_853 ();
 FILLCELL_X1 FILLER_38_855 ();
 FILLCELL_X16 FILLER_38_860 ();
 FILLCELL_X8 FILLER_38_876 ();
 FILLCELL_X2 FILLER_38_884 ();
 FILLCELL_X32 FILLER_38_890 ();
 FILLCELL_X4 FILLER_38_922 ();
 FILLCELL_X2 FILLER_38_926 ();
 FILLCELL_X1 FILLER_38_928 ();
 FILLCELL_X32 FILLER_38_933 ();
 FILLCELL_X4 FILLER_38_965 ();
 FILLCELL_X2 FILLER_38_969 ();
 FILLCELL_X32 FILLER_38_975 ();
 FILLCELL_X4 FILLER_38_1007 ();
 FILLCELL_X2 FILLER_38_1011 ();
 FILLCELL_X4 FILLER_38_1017 ();
 FILLCELL_X1 FILLER_38_1021 ();
 FILLCELL_X32 FILLER_38_1027 ();
 FILLCELL_X8 FILLER_38_1059 ();
 FILLCELL_X2 FILLER_38_1067 ();
 FILLCELL_X1 FILLER_38_1069 ();
 FILLCELL_X16 FILLER_38_1074 ();
 FILLCELL_X8 FILLER_38_1090 ();
 FILLCELL_X4 FILLER_38_1098 ();
 FILLCELL_X2 FILLER_38_1102 ();
 FILLCELL_X8 FILLER_38_1108 ();
 FILLCELL_X2 FILLER_38_1116 ();
 FILLCELL_X1 FILLER_38_1118 ();
 FILLCELL_X16 FILLER_38_1124 ();
 FILLCELL_X8 FILLER_38_1140 ();
 FILLCELL_X2 FILLER_38_1148 ();
 FILLCELL_X1 FILLER_38_1150 ();
 FILLCELL_X32 FILLER_38_1154 ();
 FILLCELL_X8 FILLER_38_1186 ();
 FILLCELL_X8 FILLER_38_1198 ();
 FILLCELL_X1 FILLER_38_1206 ();
 FILLCELL_X4 FILLER_38_1212 ();
 FILLCELL_X8 FILLER_38_1220 ();
 FILLCELL_X2 FILLER_38_1228 ();
 FILLCELL_X1 FILLER_38_1230 ();
 FILLCELL_X4 FILLER_38_1235 ();
 FILLCELL_X2 FILLER_38_1239 ();
 FILLCELL_X4 FILLER_38_1250 ();
 FILLCELL_X2 FILLER_38_1254 ();
 FILLCELL_X1 FILLER_38_1256 ();
 FILLCELL_X4 FILLER_38_1260 ();
 FILLCELL_X2 FILLER_38_1264 ();
 FILLCELL_X1 FILLER_38_1266 ();
 FILLCELL_X4 FILLER_38_1273 ();
 FILLCELL_X4 FILLER_38_1282 ();
 FILLCELL_X4 FILLER_38_1289 ();
 FILLCELL_X2 FILLER_38_1293 ();
 FILLCELL_X8 FILLER_38_1308 ();
 FILLCELL_X1 FILLER_38_1316 ();
 FILLCELL_X4 FILLER_38_1336 ();
 FILLCELL_X32 FILLER_38_1359 ();
 FILLCELL_X32 FILLER_38_1391 ();
 FILLCELL_X32 FILLER_38_1423 ();
 FILLCELL_X32 FILLER_38_1455 ();
 FILLCELL_X32 FILLER_38_1487 ();
 FILLCELL_X32 FILLER_38_1519 ();
 FILLCELL_X32 FILLER_38_1551 ();
 FILLCELL_X32 FILLER_38_1583 ();
 FILLCELL_X32 FILLER_38_1615 ();
 FILLCELL_X32 FILLER_38_1647 ();
 FILLCELL_X32 FILLER_38_1679 ();
 FILLCELL_X32 FILLER_38_1711 ();
 FILLCELL_X8 FILLER_38_1743 ();
 FILLCELL_X4 FILLER_38_1751 ();
 FILLCELL_X1 FILLER_38_1755 ();
 FILLCELL_X4 FILLER_39_1 ();
 FILLCELL_X1 FILLER_39_5 ();
 FILLCELL_X4 FILLER_39_10 ();
 FILLCELL_X4 FILLER_39_18 ();
 FILLCELL_X8 FILLER_39_26 ();
 FILLCELL_X8 FILLER_39_38 ();
 FILLCELL_X2 FILLER_39_46 ();
 FILLCELL_X1 FILLER_39_48 ();
 FILLCELL_X4 FILLER_39_53 ();
 FILLCELL_X1 FILLER_39_57 ();
 FILLCELL_X4 FILLER_39_61 ();
 FILLCELL_X4 FILLER_39_69 ();
 FILLCELL_X8 FILLER_39_82 ();
 FILLCELL_X4 FILLER_39_94 ();
 FILLCELL_X16 FILLER_39_102 ();
 FILLCELL_X4 FILLER_39_118 ();
 FILLCELL_X2 FILLER_39_122 ();
 FILLCELL_X4 FILLER_39_133 ();
 FILLCELL_X1 FILLER_39_137 ();
 FILLCELL_X4 FILLER_39_141 ();
 FILLCELL_X4 FILLER_39_150 ();
 FILLCELL_X4 FILLER_39_158 ();
 FILLCELL_X8 FILLER_39_165 ();
 FILLCELL_X1 FILLER_39_173 ();
 FILLCELL_X16 FILLER_39_180 ();
 FILLCELL_X4 FILLER_39_196 ();
 FILLCELL_X2 FILLER_39_200 ();
 FILLCELL_X4 FILLER_39_207 ();
 FILLCELL_X16 FILLER_39_215 ();
 FILLCELL_X8 FILLER_39_231 ();
 FILLCELL_X1 FILLER_39_239 ();
 FILLCELL_X8 FILLER_39_244 ();
 FILLCELL_X4 FILLER_39_261 ();
 FILLCELL_X16 FILLER_39_270 ();
 FILLCELL_X1 FILLER_39_286 ();
 FILLCELL_X4 FILLER_39_292 ();
 FILLCELL_X4 FILLER_39_302 ();
 FILLCELL_X4 FILLER_39_315 ();
 FILLCELL_X8 FILLER_39_323 ();
 FILLCELL_X4 FILLER_39_331 ();
 FILLCELL_X4 FILLER_39_339 ();
 FILLCELL_X1 FILLER_39_343 ();
 FILLCELL_X8 FILLER_39_347 ();
 FILLCELL_X4 FILLER_39_358 ();
 FILLCELL_X4 FILLER_39_371 ();
 FILLCELL_X8 FILLER_39_379 ();
 FILLCELL_X2 FILLER_39_387 ();
 FILLCELL_X1 FILLER_39_389 ();
 FILLCELL_X4 FILLER_39_395 ();
 FILLCELL_X2 FILLER_39_399 ();
 FILLCELL_X4 FILLER_39_404 ();
 FILLCELL_X16 FILLER_39_413 ();
 FILLCELL_X4 FILLER_39_429 ();
 FILLCELL_X2 FILLER_39_433 ();
 FILLCELL_X1 FILLER_39_435 ();
 FILLCELL_X4 FILLER_39_441 ();
 FILLCELL_X16 FILLER_39_448 ();
 FILLCELL_X8 FILLER_39_464 ();
 FILLCELL_X4 FILLER_39_472 ();
 FILLCELL_X2 FILLER_39_476 ();
 FILLCELL_X4 FILLER_39_482 ();
 FILLCELL_X8 FILLER_39_490 ();
 FILLCELL_X2 FILLER_39_498 ();
 FILLCELL_X4 FILLER_39_504 ();
 FILLCELL_X4 FILLER_39_513 ();
 FILLCELL_X16 FILLER_39_521 ();
 FILLCELL_X2 FILLER_39_537 ();
 FILLCELL_X1 FILLER_39_539 ();
 FILLCELL_X16 FILLER_39_545 ();
 FILLCELL_X4 FILLER_39_561 ();
 FILLCELL_X16 FILLER_39_569 ();
 FILLCELL_X8 FILLER_39_585 ();
 FILLCELL_X4 FILLER_39_593 ();
 FILLCELL_X2 FILLER_39_597 ();
 FILLCELL_X1 FILLER_39_599 ();
 FILLCELL_X16 FILLER_39_604 ();
 FILLCELL_X8 FILLER_39_620 ();
 FILLCELL_X2 FILLER_39_628 ();
 FILLCELL_X1 FILLER_39_630 ();
 FILLCELL_X32 FILLER_39_632 ();
 FILLCELL_X32 FILLER_39_664 ();
 FILLCELL_X4 FILLER_39_696 ();
 FILLCELL_X2 FILLER_39_700 ();
 FILLCELL_X4 FILLER_39_707 ();
 FILLCELL_X32 FILLER_39_714 ();
 FILLCELL_X16 FILLER_39_746 ();
 FILLCELL_X8 FILLER_39_762 ();
 FILLCELL_X4 FILLER_39_770 ();
 FILLCELL_X1 FILLER_39_774 ();
 FILLCELL_X32 FILLER_39_780 ();
 FILLCELL_X16 FILLER_39_812 ();
 FILLCELL_X8 FILLER_39_828 ();
 FILLCELL_X4 FILLER_39_836 ();
 FILLCELL_X4 FILLER_39_845 ();
 FILLCELL_X32 FILLER_39_854 ();
 FILLCELL_X32 FILLER_39_886 ();
 FILLCELL_X32 FILLER_39_918 ();
 FILLCELL_X32 FILLER_39_950 ();
 FILLCELL_X32 FILLER_39_982 ();
 FILLCELL_X32 FILLER_39_1014 ();
 FILLCELL_X32 FILLER_39_1046 ();
 FILLCELL_X32 FILLER_39_1078 ();
 FILLCELL_X16 FILLER_39_1110 ();
 FILLCELL_X8 FILLER_39_1126 ();
 FILLCELL_X4 FILLER_39_1134 ();
 FILLCELL_X2 FILLER_39_1138 ();
 FILLCELL_X32 FILLER_39_1145 ();
 FILLCELL_X16 FILLER_39_1177 ();
 FILLCELL_X4 FILLER_39_1193 ();
 FILLCELL_X2 FILLER_39_1197 ();
 FILLCELL_X1 FILLER_39_1199 ();
 FILLCELL_X32 FILLER_39_1204 ();
 FILLCELL_X16 FILLER_39_1236 ();
 FILLCELL_X8 FILLER_39_1252 ();
 FILLCELL_X2 FILLER_39_1260 ();
 FILLCELL_X4 FILLER_39_1263 ();
 FILLCELL_X2 FILLER_39_1267 ();
 FILLCELL_X16 FILLER_39_1274 ();
 FILLCELL_X4 FILLER_39_1290 ();
 FILLCELL_X8 FILLER_39_1297 ();
 FILLCELL_X4 FILLER_39_1305 ();
 FILLCELL_X2 FILLER_39_1309 ();
 FILLCELL_X32 FILLER_39_1315 ();
 FILLCELL_X32 FILLER_39_1347 ();
 FILLCELL_X2 FILLER_39_1379 ();
 FILLCELL_X4 FILLER_39_1386 ();
 FILLCELL_X32 FILLER_39_1393 ();
 FILLCELL_X8 FILLER_39_1425 ();
 FILLCELL_X4 FILLER_39_1433 ();
 FILLCELL_X2 FILLER_39_1437 ();
 FILLCELL_X1 FILLER_39_1439 ();
 FILLCELL_X32 FILLER_39_1443 ();
 FILLCELL_X32 FILLER_39_1475 ();
 FILLCELL_X32 FILLER_39_1507 ();
 FILLCELL_X32 FILLER_39_1539 ();
 FILLCELL_X32 FILLER_39_1571 ();
 FILLCELL_X32 FILLER_39_1603 ();
 FILLCELL_X32 FILLER_39_1635 ();
 FILLCELL_X32 FILLER_39_1667 ();
 FILLCELL_X32 FILLER_39_1699 ();
 FILLCELL_X16 FILLER_39_1731 ();
 FILLCELL_X8 FILLER_39_1747 ();
 FILLCELL_X1 FILLER_39_1755 ();
 FILLCELL_X4 FILLER_40_1 ();
 FILLCELL_X4 FILLER_40_24 ();
 FILLCELL_X1 FILLER_40_28 ();
 FILLCELL_X4 FILLER_40_33 ();
 FILLCELL_X8 FILLER_40_46 ();
 FILLCELL_X4 FILLER_40_58 ();
 FILLCELL_X4 FILLER_40_67 ();
 FILLCELL_X4 FILLER_40_76 ();
 FILLCELL_X4 FILLER_40_84 ();
 FILLCELL_X1 FILLER_40_88 ();
 FILLCELL_X4 FILLER_40_93 ();
 FILLCELL_X1 FILLER_40_97 ();
 FILLCELL_X4 FILLER_40_102 ();
 FILLCELL_X4 FILLER_40_110 ();
 FILLCELL_X4 FILLER_40_120 ();
 FILLCELL_X4 FILLER_40_133 ();
 FILLCELL_X4 FILLER_40_142 ();
 FILLCELL_X1 FILLER_40_146 ();
 FILLCELL_X4 FILLER_40_166 ();
 FILLCELL_X2 FILLER_40_170 ();
 FILLCELL_X1 FILLER_40_172 ();
 FILLCELL_X4 FILLER_40_179 ();
 FILLCELL_X16 FILLER_40_187 ();
 FILLCELL_X8 FILLER_40_203 ();
 FILLCELL_X2 FILLER_40_211 ();
 FILLCELL_X4 FILLER_40_217 ();
 FILLCELL_X4 FILLER_40_225 ();
 FILLCELL_X4 FILLER_40_238 ();
 FILLCELL_X2 FILLER_40_242 ();
 FILLCELL_X1 FILLER_40_244 ();
 FILLCELL_X4 FILLER_40_249 ();
 FILLCELL_X4 FILLER_40_262 ();
 FILLCELL_X4 FILLER_40_272 ();
 FILLCELL_X4 FILLER_40_281 ();
 FILLCELL_X1 FILLER_40_285 ();
 FILLCELL_X16 FILLER_40_290 ();
 FILLCELL_X8 FILLER_40_311 ();
 FILLCELL_X4 FILLER_40_319 ();
 FILLCELL_X2 FILLER_40_323 ();
 FILLCELL_X4 FILLER_40_329 ();
 FILLCELL_X8 FILLER_40_342 ();
 FILLCELL_X2 FILLER_40_350 ();
 FILLCELL_X4 FILLER_40_358 ();
 FILLCELL_X8 FILLER_40_371 ();
 FILLCELL_X1 FILLER_40_379 ();
 FILLCELL_X32 FILLER_40_1518 ();
 FILLCELL_X32 FILLER_40_1550 ();
 FILLCELL_X32 FILLER_40_1582 ();
 FILLCELL_X32 FILLER_40_1614 ();
 FILLCELL_X32 FILLER_40_1646 ();
 FILLCELL_X32 FILLER_40_1678 ();
 FILLCELL_X32 FILLER_40_1710 ();
 FILLCELL_X8 FILLER_40_1742 ();
 FILLCELL_X4 FILLER_40_1750 ();
 FILLCELL_X2 FILLER_40_1754 ();
 FILLCELL_X4 FILLER_41_1 ();
 FILLCELL_X16 FILLER_41_8 ();
 FILLCELL_X1 FILLER_41_24 ();
 FILLCELL_X4 FILLER_41_34 ();
 FILLCELL_X4 FILLER_41_47 ();
 FILLCELL_X8 FILLER_41_55 ();
 FILLCELL_X2 FILLER_41_63 ();
 FILLCELL_X1 FILLER_41_65 ();
 FILLCELL_X4 FILLER_41_75 ();
 FILLCELL_X8 FILLER_41_84 ();
 FILLCELL_X2 FILLER_41_92 ();
 FILLCELL_X1 FILLER_41_94 ();
 FILLCELL_X8 FILLER_41_104 ();
 FILLCELL_X4 FILLER_41_112 ();
 FILLCELL_X2 FILLER_41_116 ();
 FILLCELL_X1 FILLER_41_118 ();
 FILLCELL_X4 FILLER_41_124 ();
 FILLCELL_X4 FILLER_41_132 ();
 FILLCELL_X4 FILLER_41_139 ();
 FILLCELL_X1 FILLER_41_143 ();
 FILLCELL_X4 FILLER_41_148 ();
 FILLCELL_X8 FILLER_41_156 ();
 FILLCELL_X4 FILLER_41_164 ();
 FILLCELL_X2 FILLER_41_168 ();
 FILLCELL_X4 FILLER_41_187 ();
 FILLCELL_X1 FILLER_41_191 ();
 FILLCELL_X4 FILLER_41_196 ();
 FILLCELL_X4 FILLER_41_204 ();
 FILLCELL_X4 FILLER_41_213 ();
 FILLCELL_X4 FILLER_41_226 ();
 FILLCELL_X4 FILLER_41_239 ();
 FILLCELL_X4 FILLER_41_248 ();
 FILLCELL_X1 FILLER_41_252 ();
 FILLCELL_X8 FILLER_41_262 ();
 FILLCELL_X1 FILLER_41_270 ();
 FILLCELL_X4 FILLER_41_288 ();
 FILLCELL_X8 FILLER_41_301 ();
 FILLCELL_X1 FILLER_41_309 ();
 FILLCELL_X4 FILLER_41_313 ();
 FILLCELL_X16 FILLER_41_320 ();
 FILLCELL_X4 FILLER_41_342 ();
 FILLCELL_X4 FILLER_41_351 ();
 FILLCELL_X2 FILLER_41_355 ();
 FILLCELL_X8 FILLER_41_362 ();
 FILLCELL_X1 FILLER_41_370 ();
 FILLCELL_X4 FILLER_41_376 ();
 FILLCELL_X32 FILLER_41_1518 ();
 FILLCELL_X32 FILLER_41_1550 ();
 FILLCELL_X32 FILLER_41_1582 ();
 FILLCELL_X32 FILLER_41_1614 ();
 FILLCELL_X32 FILLER_41_1646 ();
 FILLCELL_X32 FILLER_41_1678 ();
 FILLCELL_X32 FILLER_41_1710 ();
 FILLCELL_X8 FILLER_41_1742 ();
 FILLCELL_X4 FILLER_41_1750 ();
 FILLCELL_X2 FILLER_41_1754 ();
 FILLCELL_X4 FILLER_42_1 ();
 FILLCELL_X16 FILLER_42_9 ();
 FILLCELL_X8 FILLER_42_25 ();
 FILLCELL_X2 FILLER_42_33 ();
 FILLCELL_X1 FILLER_42_35 ();
 FILLCELL_X4 FILLER_42_42 ();
 FILLCELL_X4 FILLER_42_49 ();
 FILLCELL_X2 FILLER_42_53 ();
 FILLCELL_X4 FILLER_42_64 ();
 FILLCELL_X4 FILLER_42_77 ();
 FILLCELL_X2 FILLER_42_81 ();
 FILLCELL_X1 FILLER_42_83 ();
 FILLCELL_X4 FILLER_42_90 ();
 FILLCELL_X4 FILLER_42_103 ();
 FILLCELL_X8 FILLER_42_112 ();
 FILLCELL_X2 FILLER_42_120 ();
 FILLCELL_X1 FILLER_42_122 ();
 FILLCELL_X4 FILLER_42_127 ();
 FILLCELL_X1 FILLER_42_131 ();
 FILLCELL_X32 FILLER_42_135 ();
 FILLCELL_X1 FILLER_42_167 ();
 FILLCELL_X4 FILLER_42_173 ();
 FILLCELL_X8 FILLER_42_180 ();
 FILLCELL_X4 FILLER_42_194 ();
 FILLCELL_X4 FILLER_42_207 ();
 FILLCELL_X8 FILLER_42_214 ();
 FILLCELL_X4 FILLER_42_228 ();
 FILLCELL_X4 FILLER_42_236 ();
 FILLCELL_X16 FILLER_42_243 ();
 FILLCELL_X1 FILLER_42_259 ();
 FILLCELL_X4 FILLER_42_265 ();
 FILLCELL_X8 FILLER_42_273 ();
 FILLCELL_X4 FILLER_42_281 ();
 FILLCELL_X2 FILLER_42_285 ();
 FILLCELL_X4 FILLER_42_296 ();
 FILLCELL_X4 FILLER_42_309 ();
 FILLCELL_X4 FILLER_42_319 ();
 FILLCELL_X4 FILLER_42_328 ();
 FILLCELL_X2 FILLER_42_332 ();
 FILLCELL_X1 FILLER_42_334 ();
 FILLCELL_X4 FILLER_42_344 ();
 FILLCELL_X4 FILLER_42_352 ();
 FILLCELL_X2 FILLER_42_356 ();
 FILLCELL_X4 FILLER_42_361 ();
 FILLCELL_X8 FILLER_42_371 ();
 FILLCELL_X1 FILLER_42_379 ();
 FILLCELL_X32 FILLER_42_1518 ();
 FILLCELL_X32 FILLER_42_1550 ();
 FILLCELL_X32 FILLER_42_1582 ();
 FILLCELL_X32 FILLER_42_1614 ();
 FILLCELL_X32 FILLER_42_1646 ();
 FILLCELL_X32 FILLER_42_1678 ();
 FILLCELL_X32 FILLER_42_1710 ();
 FILLCELL_X8 FILLER_42_1742 ();
 FILLCELL_X4 FILLER_42_1750 ();
 FILLCELL_X2 FILLER_42_1754 ();
 FILLCELL_X4 FILLER_43_1 ();
 FILLCELL_X1 FILLER_43_5 ();
 FILLCELL_X4 FILLER_43_10 ();
 FILLCELL_X2 FILLER_43_14 ();
 FILLCELL_X16 FILLER_43_20 ();
 FILLCELL_X4 FILLER_43_39 ();
 FILLCELL_X8 FILLER_43_48 ();
 FILLCELL_X4 FILLER_43_56 ();
 FILLCELL_X4 FILLER_43_66 ();
 FILLCELL_X1 FILLER_43_70 ();
 FILLCELL_X4 FILLER_43_76 ();
 FILLCELL_X8 FILLER_43_83 ();
 FILLCELL_X1 FILLER_43_91 ();
 FILLCELL_X4 FILLER_43_95 ();
 FILLCELL_X8 FILLER_43_103 ();
 FILLCELL_X4 FILLER_43_111 ();
 FILLCELL_X2 FILLER_43_115 ();
 FILLCELL_X4 FILLER_43_121 ();
 FILLCELL_X8 FILLER_43_130 ();
 FILLCELL_X4 FILLER_43_141 ();
 FILLCELL_X4 FILLER_43_151 ();
 FILLCELL_X4 FILLER_43_164 ();
 FILLCELL_X2 FILLER_43_168 ();
 FILLCELL_X1 FILLER_43_170 ();
 FILLCELL_X4 FILLER_43_180 ();
 FILLCELL_X1 FILLER_43_184 ();
 FILLCELL_X4 FILLER_43_194 ();
 FILLCELL_X4 FILLER_43_207 ();
 FILLCELL_X16 FILLER_43_216 ();
 FILLCELL_X8 FILLER_43_232 ();
 FILLCELL_X4 FILLER_43_240 ();
 FILLCELL_X2 FILLER_43_244 ();
 FILLCELL_X4 FILLER_43_249 ();
 FILLCELL_X4 FILLER_43_262 ();
 FILLCELL_X4 FILLER_43_269 ();
 FILLCELL_X2 FILLER_43_273 ();
 FILLCELL_X16 FILLER_43_279 ();
 FILLCELL_X4 FILLER_43_295 ();
 FILLCELL_X16 FILLER_43_303 ();
 FILLCELL_X8 FILLER_43_319 ();
 FILLCELL_X4 FILLER_43_331 ();
 FILLCELL_X4 FILLER_43_339 ();
 FILLCELL_X4 FILLER_43_346 ();
 FILLCELL_X2 FILLER_43_350 ();
 FILLCELL_X1 FILLER_43_352 ();
 FILLCELL_X4 FILLER_43_362 ();
 FILLCELL_X4 FILLER_43_375 ();
 FILLCELL_X1 FILLER_43_379 ();
 FILLCELL_X32 FILLER_43_1518 ();
 FILLCELL_X32 FILLER_43_1550 ();
 FILLCELL_X32 FILLER_43_1582 ();
 FILLCELL_X32 FILLER_43_1614 ();
 FILLCELL_X32 FILLER_43_1646 ();
 FILLCELL_X32 FILLER_43_1678 ();
 FILLCELL_X32 FILLER_43_1710 ();
 FILLCELL_X8 FILLER_43_1742 ();
 FILLCELL_X4 FILLER_43_1750 ();
 FILLCELL_X2 FILLER_43_1754 ();
 FILLCELL_X8 FILLER_44_1 ();
 FILLCELL_X2 FILLER_44_9 ();
 FILLCELL_X4 FILLER_44_20 ();
 FILLCELL_X4 FILLER_44_28 ();
 FILLCELL_X16 FILLER_44_35 ();
 FILLCELL_X8 FILLER_44_51 ();
 FILLCELL_X4 FILLER_44_59 ();
 FILLCELL_X4 FILLER_44_66 ();
 FILLCELL_X8 FILLER_44_79 ();
 FILLCELL_X2 FILLER_44_87 ();
 FILLCELL_X1 FILLER_44_89 ();
 FILLCELL_X8 FILLER_44_93 ();
 FILLCELL_X4 FILLER_44_101 ();
 FILLCELL_X2 FILLER_44_105 ();
 FILLCELL_X1 FILLER_44_107 ();
 FILLCELL_X4 FILLER_44_114 ();
 FILLCELL_X4 FILLER_44_127 ();
 FILLCELL_X8 FILLER_44_140 ();
 FILLCELL_X1 FILLER_44_148 ();
 FILLCELL_X4 FILLER_44_152 ();
 FILLCELL_X4 FILLER_44_159 ();
 FILLCELL_X4 FILLER_44_166 ();
 FILLCELL_X16 FILLER_44_174 ();
 FILLCELL_X2 FILLER_44_190 ();
 FILLCELL_X4 FILLER_44_197 ();
 FILLCELL_X2 FILLER_44_201 ();
 FILLCELL_X1 FILLER_44_203 ();
 FILLCELL_X4 FILLER_44_209 ();
 FILLCELL_X8 FILLER_44_222 ();
 FILLCELL_X1 FILLER_44_230 ();
 FILLCELL_X4 FILLER_44_236 ();
 FILLCELL_X4 FILLER_44_245 ();
 FILLCELL_X4 FILLER_44_258 ();
 FILLCELL_X8 FILLER_44_271 ();
 FILLCELL_X2 FILLER_44_279 ();
 FILLCELL_X4 FILLER_44_287 ();
 FILLCELL_X8 FILLER_44_296 ();
 FILLCELL_X1 FILLER_44_304 ();
 FILLCELL_X4 FILLER_44_310 ();
 FILLCELL_X8 FILLER_44_319 ();
 FILLCELL_X4 FILLER_44_327 ();
 FILLCELL_X2 FILLER_44_331 ();
 FILLCELL_X16 FILLER_44_337 ();
 FILLCELL_X4 FILLER_44_353 ();
 FILLCELL_X1 FILLER_44_357 ();
 FILLCELL_X4 FILLER_44_361 ();
 FILLCELL_X8 FILLER_44_370 ();
 FILLCELL_X2 FILLER_44_378 ();
 FILLCELL_X32 FILLER_44_1518 ();
 FILLCELL_X32 FILLER_44_1550 ();
 FILLCELL_X32 FILLER_44_1582 ();
 FILLCELL_X32 FILLER_44_1614 ();
 FILLCELL_X32 FILLER_44_1646 ();
 FILLCELL_X32 FILLER_44_1678 ();
 FILLCELL_X32 FILLER_44_1710 ();
 FILLCELL_X8 FILLER_44_1742 ();
 FILLCELL_X4 FILLER_44_1750 ();
 FILLCELL_X2 FILLER_44_1754 ();
 FILLCELL_X8 FILLER_45_1 ();
 FILLCELL_X1 FILLER_45_9 ();
 FILLCELL_X4 FILLER_45_19 ();
 FILLCELL_X4 FILLER_45_32 ();
 FILLCELL_X1 FILLER_45_36 ();
 FILLCELL_X16 FILLER_45_42 ();
 FILLCELL_X1 FILLER_45_58 ();
 FILLCELL_X4 FILLER_45_68 ();
 FILLCELL_X4 FILLER_45_81 ();
 FILLCELL_X16 FILLER_45_90 ();
 FILLCELL_X2 FILLER_45_106 ();
 FILLCELL_X1 FILLER_45_108 ();
 FILLCELL_X4 FILLER_45_113 ();
 FILLCELL_X4 FILLER_45_122 ();
 FILLCELL_X8 FILLER_45_130 ();
 FILLCELL_X4 FILLER_45_138 ();
 FILLCELL_X2 FILLER_45_142 ();
 FILLCELL_X1 FILLER_45_144 ();
 FILLCELL_X8 FILLER_45_154 ();
 FILLCELL_X1 FILLER_45_162 ();
 FILLCELL_X4 FILLER_45_167 ();
 FILLCELL_X4 FILLER_45_175 ();
 FILLCELL_X8 FILLER_45_183 ();
 FILLCELL_X4 FILLER_45_191 ();
 FILLCELL_X2 FILLER_45_195 ();
 FILLCELL_X4 FILLER_45_201 ();
 FILLCELL_X4 FILLER_45_209 ();
 FILLCELL_X4 FILLER_45_222 ();
 FILLCELL_X4 FILLER_45_235 ();
 FILLCELL_X4 FILLER_45_242 ();
 FILLCELL_X4 FILLER_45_249 ();
 FILLCELL_X4 FILLER_45_259 ();
 FILLCELL_X4 FILLER_45_267 ();
 FILLCELL_X1 FILLER_45_271 ();
 FILLCELL_X4 FILLER_45_277 ();
 FILLCELL_X8 FILLER_45_290 ();
 FILLCELL_X2 FILLER_45_298 ();
 FILLCELL_X4 FILLER_45_306 ();
 FILLCELL_X4 FILLER_45_319 ();
 FILLCELL_X8 FILLER_45_326 ();
 FILLCELL_X8 FILLER_45_353 ();
 FILLCELL_X2 FILLER_45_361 ();
 FILLCELL_X4 FILLER_45_366 ();
 FILLCELL_X2 FILLER_45_370 ();
 FILLCELL_X4 FILLER_45_376 ();
 FILLCELL_X32 FILLER_45_1518 ();
 FILLCELL_X32 FILLER_45_1550 ();
 FILLCELL_X32 FILLER_45_1582 ();
 FILLCELL_X32 FILLER_45_1614 ();
 FILLCELL_X32 FILLER_45_1646 ();
 FILLCELL_X32 FILLER_45_1678 ();
 FILLCELL_X32 FILLER_45_1710 ();
 FILLCELL_X8 FILLER_45_1742 ();
 FILLCELL_X4 FILLER_45_1750 ();
 FILLCELL_X2 FILLER_45_1754 ();
 FILLCELL_X8 FILLER_46_1 ();
 FILLCELL_X2 FILLER_46_9 ();
 FILLCELL_X8 FILLER_46_15 ();
 FILLCELL_X2 FILLER_46_23 ();
 FILLCELL_X1 FILLER_46_25 ();
 FILLCELL_X8 FILLER_46_32 ();
 FILLCELL_X4 FILLER_46_40 ();
 FILLCELL_X4 FILLER_46_48 ();
 FILLCELL_X8 FILLER_46_56 ();
 FILLCELL_X2 FILLER_46_64 ();
 FILLCELL_X1 FILLER_46_66 ();
 FILLCELL_X4 FILLER_46_71 ();
 FILLCELL_X8 FILLER_46_81 ();
 FILLCELL_X1 FILLER_46_89 ();
 FILLCELL_X32 FILLER_46_107 ();
 FILLCELL_X8 FILLER_46_139 ();
 FILLCELL_X4 FILLER_46_152 ();
 FILLCELL_X8 FILLER_46_159 ();
 FILLCELL_X2 FILLER_46_167 ();
 FILLCELL_X1 FILLER_46_169 ();
 FILLCELL_X16 FILLER_46_179 ();
 FILLCELL_X2 FILLER_46_195 ();
 FILLCELL_X8 FILLER_46_201 ();
 FILLCELL_X2 FILLER_46_209 ();
 FILLCELL_X4 FILLER_46_214 ();
 FILLCELL_X2 FILLER_46_218 ();
 FILLCELL_X1 FILLER_46_220 ();
 FILLCELL_X8 FILLER_46_227 ();
 FILLCELL_X4 FILLER_46_235 ();
 FILLCELL_X2 FILLER_46_239 ();
 FILLCELL_X1 FILLER_46_241 ();
 FILLCELL_X8 FILLER_46_247 ();
 FILLCELL_X2 FILLER_46_255 ();
 FILLCELL_X4 FILLER_46_262 ();
 FILLCELL_X1 FILLER_46_266 ();
 FILLCELL_X8 FILLER_46_270 ();
 FILLCELL_X4 FILLER_46_278 ();
 FILLCELL_X1 FILLER_46_282 ();
 FILLCELL_X4 FILLER_46_292 ();
 FILLCELL_X8 FILLER_46_299 ();
 FILLCELL_X2 FILLER_46_307 ();
 FILLCELL_X4 FILLER_46_313 ();
 FILLCELL_X8 FILLER_46_321 ();
 FILLCELL_X4 FILLER_46_329 ();
 FILLCELL_X2 FILLER_46_333 ();
 FILLCELL_X4 FILLER_46_344 ();
 FILLCELL_X2 FILLER_46_348 ();
 FILLCELL_X4 FILLER_46_353 ();
 FILLCELL_X4 FILLER_46_360 ();
 FILLCELL_X8 FILLER_46_371 ();
 FILLCELL_X1 FILLER_46_379 ();
 FILLCELL_X32 FILLER_46_1518 ();
 FILLCELL_X32 FILLER_46_1550 ();
 FILLCELL_X32 FILLER_46_1582 ();
 FILLCELL_X32 FILLER_46_1614 ();
 FILLCELL_X32 FILLER_46_1646 ();
 FILLCELL_X32 FILLER_46_1678 ();
 FILLCELL_X32 FILLER_46_1710 ();
 FILLCELL_X8 FILLER_46_1742 ();
 FILLCELL_X4 FILLER_46_1750 ();
 FILLCELL_X2 FILLER_46_1754 ();
 FILLCELL_X16 FILLER_47_1 ();
 FILLCELL_X8 FILLER_47_17 ();
 FILLCELL_X4 FILLER_47_25 ();
 FILLCELL_X8 FILLER_47_34 ();
 FILLCELL_X2 FILLER_47_42 ();
 FILLCELL_X4 FILLER_47_53 ();
 FILLCELL_X8 FILLER_47_60 ();
 FILLCELL_X4 FILLER_47_68 ();
 FILLCELL_X2 FILLER_47_72 ();
 FILLCELL_X1 FILLER_47_74 ();
 FILLCELL_X4 FILLER_47_79 ();
 FILLCELL_X8 FILLER_47_88 ();
 FILLCELL_X2 FILLER_47_96 ();
 FILLCELL_X1 FILLER_47_98 ();
 FILLCELL_X8 FILLER_47_103 ();
 FILLCELL_X1 FILLER_47_111 ();
 FILLCELL_X4 FILLER_47_118 ();
 FILLCELL_X2 FILLER_47_122 ();
 FILLCELL_X8 FILLER_47_128 ();
 FILLCELL_X2 FILLER_47_136 ();
 FILLCELL_X4 FILLER_47_144 ();
 FILLCELL_X8 FILLER_47_157 ();
 FILLCELL_X4 FILLER_47_165 ();
 FILLCELL_X2 FILLER_47_169 ();
 FILLCELL_X1 FILLER_47_171 ();
 FILLCELL_X4 FILLER_47_175 ();
 FILLCELL_X4 FILLER_47_188 ();
 FILLCELL_X4 FILLER_47_195 ();
 FILLCELL_X1 FILLER_47_199 ();
 FILLCELL_X4 FILLER_47_209 ();
 FILLCELL_X2 FILLER_47_213 ();
 FILLCELL_X4 FILLER_47_218 ();
 FILLCELL_X16 FILLER_47_226 ();
 FILLCELL_X2 FILLER_47_242 ();
 FILLCELL_X1 FILLER_47_244 ();
 FILLCELL_X4 FILLER_47_251 ();
 FILLCELL_X1 FILLER_47_255 ();
 FILLCELL_X8 FILLER_47_265 ();
 FILLCELL_X1 FILLER_47_273 ();
 FILLCELL_X4 FILLER_47_278 ();
 FILLCELL_X8 FILLER_47_291 ();
 FILLCELL_X4 FILLER_47_299 ();
 FILLCELL_X2 FILLER_47_303 ();
 FILLCELL_X4 FILLER_47_314 ();
 FILLCELL_X8 FILLER_47_327 ();
 FILLCELL_X2 FILLER_47_335 ();
 FILLCELL_X4 FILLER_47_340 ();
 FILLCELL_X4 FILLER_47_347 ();
 FILLCELL_X1 FILLER_47_351 ();
 FILLCELL_X4 FILLER_47_358 ();
 FILLCELL_X8 FILLER_47_368 ();
 FILLCELL_X4 FILLER_47_376 ();
 FILLCELL_X32 FILLER_47_1518 ();
 FILLCELL_X32 FILLER_47_1550 ();
 FILLCELL_X32 FILLER_47_1582 ();
 FILLCELL_X32 FILLER_47_1614 ();
 FILLCELL_X32 FILLER_47_1646 ();
 FILLCELL_X32 FILLER_47_1678 ();
 FILLCELL_X32 FILLER_47_1710 ();
 FILLCELL_X8 FILLER_47_1742 ();
 FILLCELL_X4 FILLER_47_1750 ();
 FILLCELL_X2 FILLER_47_1754 ();
 FILLCELL_X16 FILLER_48_1 ();
 FILLCELL_X8 FILLER_48_17 ();
 FILLCELL_X2 FILLER_48_25 ();
 FILLCELL_X8 FILLER_48_31 ();
 FILLCELL_X2 FILLER_48_39 ();
 FILLCELL_X1 FILLER_48_41 ();
 FILLCELL_X4 FILLER_48_45 ();
 FILLCELL_X4 FILLER_48_58 ();
 FILLCELL_X4 FILLER_48_67 ();
 FILLCELL_X4 FILLER_48_75 ();
 FILLCELL_X4 FILLER_48_82 ();
 FILLCELL_X4 FILLER_48_90 ();
 FILLCELL_X8 FILLER_48_98 ();
 FILLCELL_X4 FILLER_48_106 ();
 FILLCELL_X2 FILLER_48_110 ();
 FILLCELL_X1 FILLER_48_112 ();
 FILLCELL_X4 FILLER_48_119 ();
 FILLCELL_X8 FILLER_48_136 ();
 FILLCELL_X1 FILLER_48_144 ();
 FILLCELL_X4 FILLER_48_149 ();
 FILLCELL_X1 FILLER_48_153 ();
 FILLCELL_X8 FILLER_48_157 ();
 FILLCELL_X2 FILLER_48_165 ();
 FILLCELL_X4 FILLER_48_170 ();
 FILLCELL_X4 FILLER_48_179 ();
 FILLCELL_X4 FILLER_48_188 ();
 FILLCELL_X2 FILLER_48_192 ();
 FILLCELL_X4 FILLER_48_198 ();
 FILLCELL_X4 FILLER_48_208 ();
 FILLCELL_X8 FILLER_48_217 ();
 FILLCELL_X1 FILLER_48_225 ();
 FILLCELL_X4 FILLER_48_230 ();
 FILLCELL_X4 FILLER_48_238 ();
 FILLCELL_X4 FILLER_48_251 ();
 FILLCELL_X4 FILLER_48_264 ();
 FILLCELL_X2 FILLER_48_268 ();
 FILLCELL_X1 FILLER_48_270 ();
 FILLCELL_X4 FILLER_48_275 ();
 FILLCELL_X4 FILLER_48_283 ();
 FILLCELL_X4 FILLER_48_291 ();
 FILLCELL_X4 FILLER_48_299 ();
 FILLCELL_X4 FILLER_48_307 ();
 FILLCELL_X8 FILLER_48_315 ();
 FILLCELL_X2 FILLER_48_323 ();
 FILLCELL_X1 FILLER_48_325 ();
 FILLCELL_X4 FILLER_48_331 ();
 FILLCELL_X4 FILLER_48_341 ();
 FILLCELL_X4 FILLER_48_349 ();
 FILLCELL_X8 FILLER_48_356 ();
 FILLCELL_X4 FILLER_48_364 ();
 FILLCELL_X8 FILLER_48_372 ();
 FILLCELL_X32 FILLER_48_1518 ();
 FILLCELL_X32 FILLER_48_1550 ();
 FILLCELL_X32 FILLER_48_1582 ();
 FILLCELL_X32 FILLER_48_1614 ();
 FILLCELL_X32 FILLER_48_1646 ();
 FILLCELL_X32 FILLER_48_1678 ();
 FILLCELL_X32 FILLER_48_1710 ();
 FILLCELL_X8 FILLER_48_1742 ();
 FILLCELL_X4 FILLER_48_1750 ();
 FILLCELL_X2 FILLER_48_1754 ();
 FILLCELL_X16 FILLER_49_1 ();
 FILLCELL_X2 FILLER_49_17 ();
 FILLCELL_X4 FILLER_49_36 ();
 FILLCELL_X2 FILLER_49_40 ();
 FILLCELL_X1 FILLER_49_42 ();
 FILLCELL_X4 FILLER_49_49 ();
 FILLCELL_X2 FILLER_49_53 ();
 FILLCELL_X1 FILLER_49_55 ();
 FILLCELL_X8 FILLER_49_60 ();
 FILLCELL_X4 FILLER_49_68 ();
 FILLCELL_X2 FILLER_49_72 ();
 FILLCELL_X1 FILLER_49_74 ();
 FILLCELL_X8 FILLER_49_84 ();
 FILLCELL_X4 FILLER_49_96 ();
 FILLCELL_X2 FILLER_49_100 ();
 FILLCELL_X1 FILLER_49_102 ();
 FILLCELL_X4 FILLER_49_112 ();
 FILLCELL_X4 FILLER_49_119 ();
 FILLCELL_X1 FILLER_49_123 ();
 FILLCELL_X8 FILLER_49_128 ();
 FILLCELL_X4 FILLER_49_139 ();
 FILLCELL_X4 FILLER_49_146 ();
 FILLCELL_X4 FILLER_49_159 ();
 FILLCELL_X4 FILLER_49_168 ();
 FILLCELL_X4 FILLER_49_178 ();
 FILLCELL_X8 FILLER_49_191 ();
 FILLCELL_X4 FILLER_49_199 ();
 FILLCELL_X1 FILLER_49_203 ();
 FILLCELL_X4 FILLER_49_213 ();
 FILLCELL_X4 FILLER_49_220 ();
 FILLCELL_X1 FILLER_49_224 ();
 FILLCELL_X4 FILLER_49_234 ();
 FILLCELL_X4 FILLER_49_242 ();
 FILLCELL_X2 FILLER_49_246 ();
 FILLCELL_X1 FILLER_49_248 ();
 FILLCELL_X4 FILLER_49_253 ();
 FILLCELL_X4 FILLER_49_261 ();
 FILLCELL_X4 FILLER_49_269 ();
 FILLCELL_X32 FILLER_49_277 ();
 FILLCELL_X8 FILLER_49_309 ();
 FILLCELL_X2 FILLER_49_317 ();
 FILLCELL_X1 FILLER_49_319 ();
 FILLCELL_X4 FILLER_49_323 ();
 FILLCELL_X2 FILLER_49_327 ();
 FILLCELL_X8 FILLER_49_338 ();
 FILLCELL_X2 FILLER_49_346 ();
 FILLCELL_X4 FILLER_49_352 ();
 FILLCELL_X1 FILLER_49_356 ();
 FILLCELL_X4 FILLER_49_376 ();
 FILLCELL_X32 FILLER_49_1518 ();
 FILLCELL_X32 FILLER_49_1550 ();
 FILLCELL_X32 FILLER_49_1582 ();
 FILLCELL_X32 FILLER_49_1614 ();
 FILLCELL_X32 FILLER_49_1646 ();
 FILLCELL_X32 FILLER_49_1678 ();
 FILLCELL_X32 FILLER_49_1710 ();
 FILLCELL_X4 FILLER_49_1742 ();
 FILLCELL_X2 FILLER_49_1746 ();
 FILLCELL_X1 FILLER_49_1748 ();
 FILLCELL_X4 FILLER_49_1752 ();
 FILLCELL_X16 FILLER_50_1 ();
 FILLCELL_X2 FILLER_50_17 ();
 FILLCELL_X1 FILLER_50_19 ();
 FILLCELL_X16 FILLER_50_24 ();
 FILLCELL_X4 FILLER_50_40 ();
 FILLCELL_X1 FILLER_50_44 ();
 FILLCELL_X4 FILLER_50_50 ();
 FILLCELL_X16 FILLER_50_58 ();
 FILLCELL_X4 FILLER_50_83 ();
 FILLCELL_X8 FILLER_50_92 ();
 FILLCELL_X4 FILLER_50_104 ();
 FILLCELL_X8 FILLER_50_113 ();
 FILLCELL_X4 FILLER_50_124 ();
 FILLCELL_X2 FILLER_50_128 ();
 FILLCELL_X1 FILLER_50_130 ();
 FILLCELL_X4 FILLER_50_135 ();
 FILLCELL_X8 FILLER_50_142 ();
 FILLCELL_X1 FILLER_50_150 ();
 FILLCELL_X4 FILLER_50_157 ();
 FILLCELL_X16 FILLER_50_165 ();
 FILLCELL_X2 FILLER_50_181 ();
 FILLCELL_X16 FILLER_50_187 ();
 FILLCELL_X8 FILLER_50_203 ();
 FILLCELL_X4 FILLER_50_211 ();
 FILLCELL_X1 FILLER_50_215 ();
 FILLCELL_X4 FILLER_50_219 ();
 FILLCELL_X2 FILLER_50_223 ();
 FILLCELL_X8 FILLER_50_230 ();
 FILLCELL_X16 FILLER_50_242 ();
 FILLCELL_X4 FILLER_50_258 ();
 FILLCELL_X1 FILLER_50_262 ();
 FILLCELL_X16 FILLER_50_267 ();
 FILLCELL_X2 FILLER_50_283 ();
 FILLCELL_X4 FILLER_50_289 ();
 FILLCELL_X4 FILLER_50_297 ();
 FILLCELL_X4 FILLER_50_310 ();
 FILLCELL_X4 FILLER_50_319 ();
 FILLCELL_X2 FILLER_50_323 ();
 FILLCELL_X8 FILLER_50_328 ();
 FILLCELL_X4 FILLER_50_342 ();
 FILLCELL_X4 FILLER_50_353 ();
 FILLCELL_X8 FILLER_50_367 ();
 FILLCELL_X4 FILLER_50_375 ();
 FILLCELL_X1 FILLER_50_379 ();
 FILLCELL_X32 FILLER_50_1518 ();
 FILLCELL_X32 FILLER_50_1550 ();
 FILLCELL_X32 FILLER_50_1582 ();
 FILLCELL_X32 FILLER_50_1614 ();
 FILLCELL_X32 FILLER_50_1646 ();
 FILLCELL_X32 FILLER_50_1678 ();
 FILLCELL_X32 FILLER_50_1710 ();
 FILLCELL_X8 FILLER_50_1742 ();
 FILLCELL_X4 FILLER_50_1750 ();
 FILLCELL_X2 FILLER_50_1754 ();
 FILLCELL_X4 FILLER_51_1 ();
 FILLCELL_X4 FILLER_51_8 ();
 FILLCELL_X4 FILLER_51_16 ();
 FILLCELL_X8 FILLER_51_25 ();
 FILLCELL_X2 FILLER_51_33 ();
 FILLCELL_X1 FILLER_51_35 ();
 FILLCELL_X4 FILLER_51_45 ();
 FILLCELL_X16 FILLER_51_53 ();
 FILLCELL_X4 FILLER_51_75 ();
 FILLCELL_X4 FILLER_51_83 ();
 FILLCELL_X4 FILLER_51_90 ();
 FILLCELL_X2 FILLER_51_94 ();
 FILLCELL_X4 FILLER_51_102 ();
 FILLCELL_X8 FILLER_51_115 ();
 FILLCELL_X1 FILLER_51_123 ();
 FILLCELL_X4 FILLER_51_129 ();
 FILLCELL_X4 FILLER_51_142 ();
 FILLCELL_X2 FILLER_51_146 ();
 FILLCELL_X4 FILLER_51_153 ();
 FILLCELL_X4 FILLER_51_166 ();
 FILLCELL_X1 FILLER_51_170 ();
 FILLCELL_X4 FILLER_51_174 ();
 FILLCELL_X4 FILLER_51_182 ();
 FILLCELL_X4 FILLER_51_192 ();
 FILLCELL_X8 FILLER_51_199 ();
 FILLCELL_X4 FILLER_51_207 ();
 FILLCELL_X4 FILLER_51_217 ();
 FILLCELL_X2 FILLER_51_221 ();
 FILLCELL_X4 FILLER_51_232 ();
 FILLCELL_X1 FILLER_51_236 ();
 FILLCELL_X4 FILLER_51_243 ();
 FILLCELL_X8 FILLER_51_253 ();
 FILLCELL_X4 FILLER_51_280 ();
 FILLCELL_X4 FILLER_51_288 ();
 FILLCELL_X4 FILLER_51_296 ();
 FILLCELL_X2 FILLER_51_300 ();
 FILLCELL_X1 FILLER_51_302 ();
 FILLCELL_X4 FILLER_51_307 ();
 FILLCELL_X4 FILLER_51_320 ();
 FILLCELL_X4 FILLER_51_330 ();
 FILLCELL_X8 FILLER_51_337 ();
 FILLCELL_X2 FILLER_51_345 ();
 FILLCELL_X1 FILLER_51_347 ();
 FILLCELL_X4 FILLER_51_352 ();
 FILLCELL_X2 FILLER_51_356 ();
 FILLCELL_X1 FILLER_51_358 ();
 FILLCELL_X4 FILLER_51_365 ();
 FILLCELL_X8 FILLER_51_372 ();
 FILLCELL_X32 FILLER_51_1518 ();
 FILLCELL_X32 FILLER_51_1550 ();
 FILLCELL_X32 FILLER_51_1582 ();
 FILLCELL_X32 FILLER_51_1614 ();
 FILLCELL_X32 FILLER_51_1646 ();
 FILLCELL_X32 FILLER_51_1678 ();
 FILLCELL_X32 FILLER_51_1710 ();
 FILLCELL_X8 FILLER_51_1742 ();
 FILLCELL_X4 FILLER_51_1750 ();
 FILLCELL_X2 FILLER_51_1754 ();
 FILLCELL_X8 FILLER_52_1 ();
 FILLCELL_X8 FILLER_52_18 ();
 FILLCELL_X4 FILLER_52_35 ();
 FILLCELL_X4 FILLER_52_48 ();
 FILLCELL_X4 FILLER_52_58 ();
 FILLCELL_X4 FILLER_52_65 ();
 FILLCELL_X2 FILLER_52_69 ();
 FILLCELL_X4 FILLER_52_74 ();
 FILLCELL_X2 FILLER_52_78 ();
 FILLCELL_X16 FILLER_52_83 ();
 FILLCELL_X2 FILLER_52_99 ();
 FILLCELL_X1 FILLER_52_101 ();
 FILLCELL_X4 FILLER_52_107 ();
 FILLCELL_X2 FILLER_52_111 ();
 FILLCELL_X8 FILLER_52_116 ();
 FILLCELL_X4 FILLER_52_133 ();
 FILLCELL_X16 FILLER_52_143 ();
 FILLCELL_X4 FILLER_52_159 ();
 FILLCELL_X2 FILLER_52_163 ();
 FILLCELL_X1 FILLER_52_165 ();
 FILLCELL_X4 FILLER_52_170 ();
 FILLCELL_X4 FILLER_52_183 ();
 FILLCELL_X4 FILLER_52_196 ();
 FILLCELL_X4 FILLER_52_205 ();
 FILLCELL_X2 FILLER_52_209 ();
 FILLCELL_X8 FILLER_52_216 ();
 FILLCELL_X4 FILLER_52_228 ();
 FILLCELL_X8 FILLER_52_237 ();
 FILLCELL_X2 FILLER_52_245 ();
 FILLCELL_X4 FILLER_52_251 ();
 FILLCELL_X8 FILLER_52_262 ();
 FILLCELL_X2 FILLER_52_270 ();
 FILLCELL_X1 FILLER_52_272 ();
 FILLCELL_X4 FILLER_52_277 ();
 FILLCELL_X4 FILLER_52_290 ();
 FILLCELL_X16 FILLER_52_299 ();
 FILLCELL_X4 FILLER_52_315 ();
 FILLCELL_X1 FILLER_52_319 ();
 FILLCELL_X4 FILLER_52_323 ();
 FILLCELL_X4 FILLER_52_330 ();
 FILLCELL_X8 FILLER_52_339 ();
 FILLCELL_X4 FILLER_52_347 ();
 FILLCELL_X4 FILLER_52_364 ();
 FILLCELL_X4 FILLER_52_374 ();
 FILLCELL_X2 FILLER_52_378 ();
 FILLCELL_X32 FILLER_52_1518 ();
 FILLCELL_X32 FILLER_52_1550 ();
 FILLCELL_X32 FILLER_52_1582 ();
 FILLCELL_X32 FILLER_52_1614 ();
 FILLCELL_X32 FILLER_52_1646 ();
 FILLCELL_X32 FILLER_52_1678 ();
 FILLCELL_X32 FILLER_52_1710 ();
 FILLCELL_X8 FILLER_52_1742 ();
 FILLCELL_X4 FILLER_52_1750 ();
 FILLCELL_X2 FILLER_52_1754 ();
 FILLCELL_X8 FILLER_53_1 ();
 FILLCELL_X1 FILLER_53_9 ();
 FILLCELL_X4 FILLER_53_19 ();
 FILLCELL_X8 FILLER_53_26 ();
 FILLCELL_X4 FILLER_53_34 ();
 FILLCELL_X1 FILLER_53_38 ();
 FILLCELL_X4 FILLER_53_42 ();
 FILLCELL_X8 FILLER_53_51 ();
 FILLCELL_X1 FILLER_53_59 ();
 FILLCELL_X16 FILLER_53_69 ();
 FILLCELL_X2 FILLER_53_85 ();
 FILLCELL_X1 FILLER_53_87 ();
 FILLCELL_X4 FILLER_53_93 ();
 FILLCELL_X2 FILLER_53_97 ();
 FILLCELL_X4 FILLER_53_103 ();
 FILLCELL_X4 FILLER_53_110 ();
 FILLCELL_X8 FILLER_53_117 ();
 FILLCELL_X2 FILLER_53_125 ();
 FILLCELL_X1 FILLER_53_127 ();
 FILLCELL_X8 FILLER_53_131 ();
 FILLCELL_X2 FILLER_53_139 ();
 FILLCELL_X1 FILLER_53_141 ();
 FILLCELL_X4 FILLER_53_145 ();
 FILLCELL_X4 FILLER_53_154 ();
 FILLCELL_X4 FILLER_53_162 ();
 FILLCELL_X4 FILLER_53_170 ();
 FILLCELL_X4 FILLER_53_178 ();
 FILLCELL_X4 FILLER_53_191 ();
 FILLCELL_X4 FILLER_53_200 ();
 FILLCELL_X4 FILLER_53_210 ();
 FILLCELL_X4 FILLER_53_219 ();
 FILLCELL_X4 FILLER_53_226 ();
 FILLCELL_X1 FILLER_53_230 ();
 FILLCELL_X4 FILLER_53_237 ();
 FILLCELL_X8 FILLER_53_244 ();
 FILLCELL_X1 FILLER_53_252 ();
 FILLCELL_X16 FILLER_53_257 ();
 FILLCELL_X8 FILLER_53_273 ();
 FILLCELL_X2 FILLER_53_281 ();
 FILLCELL_X1 FILLER_53_283 ();
 FILLCELL_X8 FILLER_53_290 ();
 FILLCELL_X2 FILLER_53_298 ();
 FILLCELL_X1 FILLER_53_300 ();
 FILLCELL_X4 FILLER_53_305 ();
 FILLCELL_X2 FILLER_53_309 ();
 FILLCELL_X1 FILLER_53_311 ();
 FILLCELL_X8 FILLER_53_317 ();
 FILLCELL_X2 FILLER_53_325 ();
 FILLCELL_X8 FILLER_53_333 ();
 FILLCELL_X1 FILLER_53_341 ();
 FILLCELL_X4 FILLER_53_345 ();
 FILLCELL_X4 FILLER_53_352 ();
 FILLCELL_X8 FILLER_53_359 ();
 FILLCELL_X1 FILLER_53_367 ();
 FILLCELL_X8 FILLER_53_372 ();
 FILLCELL_X32 FILLER_53_1518 ();
 FILLCELL_X32 FILLER_53_1550 ();
 FILLCELL_X32 FILLER_53_1582 ();
 FILLCELL_X32 FILLER_53_1614 ();
 FILLCELL_X32 FILLER_53_1646 ();
 FILLCELL_X32 FILLER_53_1678 ();
 FILLCELL_X32 FILLER_53_1710 ();
 FILLCELL_X8 FILLER_53_1742 ();
 FILLCELL_X4 FILLER_53_1750 ();
 FILLCELL_X2 FILLER_53_1754 ();
 FILLCELL_X8 FILLER_54_1 ();
 FILLCELL_X4 FILLER_54_15 ();
 FILLCELL_X2 FILLER_54_19 ();
 FILLCELL_X4 FILLER_54_25 ();
 FILLCELL_X16 FILLER_54_33 ();
 FILLCELL_X4 FILLER_54_49 ();
 FILLCELL_X4 FILLER_54_58 ();
 FILLCELL_X4 FILLER_54_71 ();
 FILLCELL_X4 FILLER_54_84 ();
 FILLCELL_X8 FILLER_54_97 ();
 FILLCELL_X1 FILLER_54_105 ();
 FILLCELL_X4 FILLER_54_113 ();
 FILLCELL_X8 FILLER_54_127 ();
 FILLCELL_X1 FILLER_54_135 ();
 FILLCELL_X4 FILLER_54_139 ();
 FILLCELL_X4 FILLER_54_149 ();
 FILLCELL_X2 FILLER_54_153 ();
 FILLCELL_X8 FILLER_54_164 ();
 FILLCELL_X4 FILLER_54_172 ();
 FILLCELL_X2 FILLER_54_176 ();
 FILLCELL_X1 FILLER_54_178 ();
 FILLCELL_X16 FILLER_54_183 ();
 FILLCELL_X2 FILLER_54_199 ();
 FILLCELL_X1 FILLER_54_201 ();
 FILLCELL_X8 FILLER_54_211 ();
 FILLCELL_X4 FILLER_54_219 ();
 FILLCELL_X1 FILLER_54_223 ();
 FILLCELL_X8 FILLER_54_229 ();
 FILLCELL_X4 FILLER_54_246 ();
 FILLCELL_X4 FILLER_54_254 ();
 FILLCELL_X1 FILLER_54_258 ();
 FILLCELL_X4 FILLER_54_265 ();
 FILLCELL_X2 FILLER_54_269 ();
 FILLCELL_X1 FILLER_54_271 ();
 FILLCELL_X4 FILLER_54_275 ();
 FILLCELL_X4 FILLER_54_288 ();
 FILLCELL_X2 FILLER_54_292 ();
 FILLCELL_X1 FILLER_54_294 ();
 FILLCELL_X4 FILLER_54_299 ();
 FILLCELL_X4 FILLER_54_312 ();
 FILLCELL_X4 FILLER_54_325 ();
 FILLCELL_X2 FILLER_54_329 ();
 FILLCELL_X4 FILLER_54_334 ();
 FILLCELL_X8 FILLER_54_347 ();
 FILLCELL_X2 FILLER_54_355 ();
 FILLCELL_X4 FILLER_54_376 ();
 FILLCELL_X32 FILLER_54_1518 ();
 FILLCELL_X32 FILLER_54_1550 ();
 FILLCELL_X32 FILLER_54_1582 ();
 FILLCELL_X32 FILLER_54_1614 ();
 FILLCELL_X32 FILLER_54_1646 ();
 FILLCELL_X32 FILLER_54_1678 ();
 FILLCELL_X32 FILLER_54_1710 ();
 FILLCELL_X8 FILLER_54_1742 ();
 FILLCELL_X4 FILLER_54_1750 ();
 FILLCELL_X2 FILLER_54_1754 ();
 FILLCELL_X4 FILLER_55_1 ();
 FILLCELL_X1 FILLER_55_5 ();
 FILLCELL_X4 FILLER_55_10 ();
 FILLCELL_X8 FILLER_55_19 ();
 FILLCELL_X1 FILLER_55_27 ();
 FILLCELL_X4 FILLER_55_32 ();
 FILLCELL_X4 FILLER_55_40 ();
 FILLCELL_X4 FILLER_55_48 ();
 FILLCELL_X4 FILLER_55_57 ();
 FILLCELL_X4 FILLER_55_67 ();
 FILLCELL_X8 FILLER_55_75 ();
 FILLCELL_X4 FILLER_55_86 ();
 FILLCELL_X4 FILLER_55_96 ();
 FILLCELL_X4 FILLER_55_103 ();
 FILLCELL_X1 FILLER_55_107 ();
 FILLCELL_X4 FILLER_55_111 ();
 FILLCELL_X8 FILLER_55_124 ();
 FILLCELL_X4 FILLER_55_132 ();
 FILLCELL_X2 FILLER_55_136 ();
 FILLCELL_X4 FILLER_55_147 ();
 FILLCELL_X8 FILLER_55_160 ();
 FILLCELL_X4 FILLER_55_168 ();
 FILLCELL_X1 FILLER_55_172 ();
 FILLCELL_X4 FILLER_55_179 ();
 FILLCELL_X4 FILLER_55_186 ();
 FILLCELL_X2 FILLER_55_190 ();
 FILLCELL_X4 FILLER_55_201 ();
 FILLCELL_X4 FILLER_55_214 ();
 FILLCELL_X4 FILLER_55_227 ();
 FILLCELL_X4 FILLER_55_240 ();
 FILLCELL_X2 FILLER_55_244 ();
 FILLCELL_X4 FILLER_55_250 ();
 FILLCELL_X1 FILLER_55_254 ();
 FILLCELL_X8 FILLER_55_261 ();
 FILLCELL_X1 FILLER_55_269 ();
 FILLCELL_X4 FILLER_55_275 ();
 FILLCELL_X1 FILLER_55_279 ();
 FILLCELL_X8 FILLER_55_289 ();
 FILLCELL_X2 FILLER_55_297 ();
 FILLCELL_X1 FILLER_55_299 ();
 FILLCELL_X4 FILLER_55_304 ();
 FILLCELL_X4 FILLER_55_312 ();
 FILLCELL_X4 FILLER_55_320 ();
 FILLCELL_X1 FILLER_55_324 ();
 FILLCELL_X4 FILLER_55_329 ();
 FILLCELL_X4 FILLER_55_339 ();
 FILLCELL_X16 FILLER_55_352 ();
 FILLCELL_X8 FILLER_55_368 ();
 FILLCELL_X4 FILLER_55_376 ();
 FILLCELL_X32 FILLER_55_1518 ();
 FILLCELL_X32 FILLER_55_1550 ();
 FILLCELL_X32 FILLER_55_1582 ();
 FILLCELL_X32 FILLER_55_1614 ();
 FILLCELL_X32 FILLER_55_1646 ();
 FILLCELL_X32 FILLER_55_1678 ();
 FILLCELL_X32 FILLER_55_1710 ();
 FILLCELL_X8 FILLER_55_1742 ();
 FILLCELL_X4 FILLER_55_1750 ();
 FILLCELL_X2 FILLER_55_1754 ();
 FILLCELL_X4 FILLER_56_1 ();
 FILLCELL_X4 FILLER_56_8 ();
 FILLCELL_X1 FILLER_56_12 ();
 FILLCELL_X4 FILLER_56_17 ();
 FILLCELL_X4 FILLER_56_40 ();
 FILLCELL_X8 FILLER_56_53 ();
 FILLCELL_X2 FILLER_56_61 ();
 FILLCELL_X1 FILLER_56_63 ();
 FILLCELL_X4 FILLER_56_68 ();
 FILLCELL_X4 FILLER_56_75 ();
 FILLCELL_X8 FILLER_56_82 ();
 FILLCELL_X1 FILLER_56_90 ();
 FILLCELL_X8 FILLER_56_95 ();
 FILLCELL_X2 FILLER_56_103 ();
 FILLCELL_X4 FILLER_56_108 ();
 FILLCELL_X2 FILLER_56_112 ();
 FILLCELL_X1 FILLER_56_114 ();
 FILLCELL_X4 FILLER_56_118 ();
 FILLCELL_X8 FILLER_56_126 ();
 FILLCELL_X4 FILLER_56_134 ();
 FILLCELL_X1 FILLER_56_138 ();
 FILLCELL_X8 FILLER_56_143 ();
 FILLCELL_X2 FILLER_56_151 ();
 FILLCELL_X1 FILLER_56_153 ();
 FILLCELL_X4 FILLER_56_157 ();
 FILLCELL_X2 FILLER_56_161 ();
 FILLCELL_X4 FILLER_56_168 ();
 FILLCELL_X4 FILLER_56_181 ();
 FILLCELL_X8 FILLER_56_188 ();
 FILLCELL_X4 FILLER_56_196 ();
 FILLCELL_X2 FILLER_56_200 ();
 FILLCELL_X1 FILLER_56_202 ();
 FILLCELL_X8 FILLER_56_207 ();
 FILLCELL_X4 FILLER_56_215 ();
 FILLCELL_X1 FILLER_56_219 ();
 FILLCELL_X4 FILLER_56_224 ();
 FILLCELL_X4 FILLER_56_232 ();
 FILLCELL_X1 FILLER_56_236 ();
 FILLCELL_X4 FILLER_56_240 ();
 FILLCELL_X4 FILLER_56_248 ();
 FILLCELL_X1 FILLER_56_252 ();
 FILLCELL_X4 FILLER_56_256 ();
 FILLCELL_X8 FILLER_56_267 ();
 FILLCELL_X4 FILLER_56_275 ();
 FILLCELL_X2 FILLER_56_279 ();
 FILLCELL_X4 FILLER_56_285 ();
 FILLCELL_X2 FILLER_56_289 ();
 FILLCELL_X32 FILLER_56_295 ();
 FILLCELL_X8 FILLER_56_327 ();
 FILLCELL_X4 FILLER_56_335 ();
 FILLCELL_X2 FILLER_56_339 ();
 FILLCELL_X4 FILLER_56_346 ();
 FILLCELL_X4 FILLER_56_353 ();
 FILLCELL_X1 FILLER_56_357 ();
 FILLCELL_X4 FILLER_56_361 ();
 FILLCELL_X2 FILLER_56_365 ();
 FILLCELL_X8 FILLER_56_371 ();
 FILLCELL_X1 FILLER_56_379 ();
 FILLCELL_X32 FILLER_56_1518 ();
 FILLCELL_X32 FILLER_56_1550 ();
 FILLCELL_X32 FILLER_56_1582 ();
 FILLCELL_X32 FILLER_56_1614 ();
 FILLCELL_X32 FILLER_56_1646 ();
 FILLCELL_X32 FILLER_56_1678 ();
 FILLCELL_X32 FILLER_56_1710 ();
 FILLCELL_X8 FILLER_56_1742 ();
 FILLCELL_X4 FILLER_56_1750 ();
 FILLCELL_X2 FILLER_56_1754 ();
 FILLCELL_X8 FILLER_57_1 ();
 FILLCELL_X8 FILLER_57_13 ();
 FILLCELL_X32 FILLER_57_24 ();
 FILLCELL_X4 FILLER_57_56 ();
 FILLCELL_X1 FILLER_57_60 ();
 FILLCELL_X4 FILLER_57_80 ();
 FILLCELL_X1 FILLER_57_84 ();
 FILLCELL_X4 FILLER_57_90 ();
 FILLCELL_X8 FILLER_57_103 ();
 FILLCELL_X1 FILLER_57_111 ();
 FILLCELL_X4 FILLER_57_116 ();
 FILLCELL_X4 FILLER_57_124 ();
 FILLCELL_X8 FILLER_57_137 ();
 FILLCELL_X2 FILLER_57_145 ();
 FILLCELL_X4 FILLER_57_152 ();
 FILLCELL_X2 FILLER_57_156 ();
 FILLCELL_X8 FILLER_57_162 ();
 FILLCELL_X2 FILLER_57_170 ();
 FILLCELL_X1 FILLER_57_172 ();
 FILLCELL_X4 FILLER_57_182 ();
 FILLCELL_X8 FILLER_57_190 ();
 FILLCELL_X4 FILLER_57_203 ();
 FILLCELL_X16 FILLER_57_210 ();
 FILLCELL_X8 FILLER_57_226 ();
 FILLCELL_X2 FILLER_57_234 ();
 FILLCELL_X1 FILLER_57_236 ();
 FILLCELL_X4 FILLER_57_240 ();
 FILLCELL_X4 FILLER_57_247 ();
 FILLCELL_X4 FILLER_57_255 ();
 FILLCELL_X16 FILLER_57_263 ();
 FILLCELL_X4 FILLER_57_279 ();
 FILLCELL_X4 FILLER_57_287 ();
 FILLCELL_X2 FILLER_57_291 ();
 FILLCELL_X1 FILLER_57_293 ();
 FILLCELL_X4 FILLER_57_298 ();
 FILLCELL_X4 FILLER_57_306 ();
 FILLCELL_X4 FILLER_57_314 ();
 FILLCELL_X2 FILLER_57_318 ();
 FILLCELL_X4 FILLER_57_324 ();
 FILLCELL_X2 FILLER_57_328 ();
 FILLCELL_X4 FILLER_57_333 ();
 FILLCELL_X8 FILLER_57_340 ();
 FILLCELL_X2 FILLER_57_348 ();
 FILLCELL_X1 FILLER_57_350 ();
 FILLCELL_X4 FILLER_57_355 ();
 FILLCELL_X1 FILLER_57_359 ();
 FILLCELL_X4 FILLER_57_365 ();
 FILLCELL_X2 FILLER_57_369 ();
 FILLCELL_X1 FILLER_57_371 ();
 FILLCELL_X4 FILLER_57_376 ();
 FILLCELL_X32 FILLER_57_1518 ();
 FILLCELL_X32 FILLER_57_1550 ();
 FILLCELL_X32 FILLER_57_1582 ();
 FILLCELL_X32 FILLER_57_1614 ();
 FILLCELL_X32 FILLER_57_1646 ();
 FILLCELL_X32 FILLER_57_1678 ();
 FILLCELL_X32 FILLER_57_1710 ();
 FILLCELL_X8 FILLER_57_1742 ();
 FILLCELL_X4 FILLER_57_1750 ();
 FILLCELL_X2 FILLER_57_1754 ();
 FILLCELL_X4 FILLER_58_1 ();
 FILLCELL_X2 FILLER_58_5 ();
 FILLCELL_X1 FILLER_58_7 ();
 FILLCELL_X4 FILLER_58_12 ();
 FILLCELL_X4 FILLER_58_20 ();
 FILLCELL_X2 FILLER_58_24 ();
 FILLCELL_X4 FILLER_58_29 ();
 FILLCELL_X4 FILLER_58_37 ();
 FILLCELL_X4 FILLER_58_50 ();
 FILLCELL_X16 FILLER_58_60 ();
 FILLCELL_X8 FILLER_58_76 ();
 FILLCELL_X1 FILLER_58_84 ();
 FILLCELL_X4 FILLER_58_94 ();
 FILLCELL_X8 FILLER_58_104 ();
 FILLCELL_X1 FILLER_58_112 ();
 FILLCELL_X4 FILLER_58_117 ();
 FILLCELL_X4 FILLER_58_130 ();
 FILLCELL_X4 FILLER_58_143 ();
 FILLCELL_X4 FILLER_58_153 ();
 FILLCELL_X4 FILLER_58_160 ();
 FILLCELL_X4 FILLER_58_168 ();
 FILLCELL_X2 FILLER_58_172 ();
 FILLCELL_X4 FILLER_58_179 ();
 FILLCELL_X4 FILLER_58_187 ();
 FILLCELL_X1 FILLER_58_191 ();
 FILLCELL_X4 FILLER_58_196 ();
 FILLCELL_X4 FILLER_58_206 ();
 FILLCELL_X4 FILLER_58_215 ();
 FILLCELL_X4 FILLER_58_223 ();
 FILLCELL_X4 FILLER_58_231 ();
 FILLCELL_X2 FILLER_58_235 ();
 FILLCELL_X8 FILLER_58_243 ();
 FILLCELL_X2 FILLER_58_251 ();
 FILLCELL_X4 FILLER_58_262 ();
 FILLCELL_X4 FILLER_58_275 ();
 FILLCELL_X4 FILLER_58_288 ();
 FILLCELL_X8 FILLER_58_296 ();
 FILLCELL_X4 FILLER_58_313 ();
 FILLCELL_X4 FILLER_58_322 ();
 FILLCELL_X8 FILLER_58_335 ();
 FILLCELL_X2 FILLER_58_343 ();
 FILLCELL_X4 FILLER_58_349 ();
 FILLCELL_X4 FILLER_58_362 ();
 FILLCELL_X4 FILLER_58_375 ();
 FILLCELL_X1 FILLER_58_379 ();
 FILLCELL_X32 FILLER_58_1518 ();
 FILLCELL_X32 FILLER_58_1550 ();
 FILLCELL_X32 FILLER_58_1582 ();
 FILLCELL_X32 FILLER_58_1614 ();
 FILLCELL_X32 FILLER_58_1646 ();
 FILLCELL_X32 FILLER_58_1678 ();
 FILLCELL_X32 FILLER_58_1710 ();
 FILLCELL_X4 FILLER_58_1742 ();
 FILLCELL_X2 FILLER_58_1746 ();
 FILLCELL_X1 FILLER_58_1748 ();
 FILLCELL_X4 FILLER_58_1752 ();
 FILLCELL_X4 FILLER_59_1 ();
 FILLCELL_X4 FILLER_59_14 ();
 FILLCELL_X4 FILLER_59_23 ();
 FILLCELL_X8 FILLER_59_31 ();
 FILLCELL_X1 FILLER_59_39 ();
 FILLCELL_X4 FILLER_59_49 ();
 FILLCELL_X4 FILLER_59_58 ();
 FILLCELL_X4 FILLER_59_65 ();
 FILLCELL_X4 FILLER_59_75 ();
 FILLCELL_X1 FILLER_59_79 ();
 FILLCELL_X4 FILLER_59_83 ();
 FILLCELL_X2 FILLER_59_87 ();
 FILLCELL_X4 FILLER_59_92 ();
 FILLCELL_X4 FILLER_59_99 ();
 FILLCELL_X32 FILLER_59_107 ();
 FILLCELL_X16 FILLER_59_139 ();
 FILLCELL_X8 FILLER_59_155 ();
 FILLCELL_X16 FILLER_59_167 ();
 FILLCELL_X4 FILLER_59_183 ();
 FILLCELL_X2 FILLER_59_187 ();
 FILLCELL_X4 FILLER_59_198 ();
 FILLCELL_X8 FILLER_59_211 ();
 FILLCELL_X1 FILLER_59_219 ();
 FILLCELL_X4 FILLER_59_229 ();
 FILLCELL_X4 FILLER_59_242 ();
 FILLCELL_X4 FILLER_59_250 ();
 FILLCELL_X8 FILLER_59_257 ();
 FILLCELL_X2 FILLER_59_265 ();
 FILLCELL_X1 FILLER_59_267 ();
 FILLCELL_X4 FILLER_59_273 ();
 FILLCELL_X4 FILLER_59_283 ();
 FILLCELL_X16 FILLER_59_291 ();
 FILLCELL_X8 FILLER_59_307 ();
 FILLCELL_X4 FILLER_59_319 ();
 FILLCELL_X4 FILLER_59_332 ();
 FILLCELL_X8 FILLER_59_342 ();
 FILLCELL_X4 FILLER_59_350 ();
 FILLCELL_X1 FILLER_59_354 ();
 FILLCELL_X4 FILLER_59_358 ();
 FILLCELL_X4 FILLER_59_368 ();
 FILLCELL_X4 FILLER_59_376 ();
 FILLCELL_X32 FILLER_59_1518 ();
 FILLCELL_X32 FILLER_59_1550 ();
 FILLCELL_X32 FILLER_59_1582 ();
 FILLCELL_X32 FILLER_59_1614 ();
 FILLCELL_X32 FILLER_59_1646 ();
 FILLCELL_X32 FILLER_59_1678 ();
 FILLCELL_X32 FILLER_59_1710 ();
 FILLCELL_X8 FILLER_59_1742 ();
 FILLCELL_X4 FILLER_59_1750 ();
 FILLCELL_X2 FILLER_59_1754 ();
 FILLCELL_X8 FILLER_60_1 ();
 FILLCELL_X4 FILLER_60_9 ();
 FILLCELL_X1 FILLER_60_13 ();
 FILLCELL_X4 FILLER_60_23 ();
 FILLCELL_X8 FILLER_60_31 ();
 FILLCELL_X2 FILLER_60_39 ();
 FILLCELL_X4 FILLER_60_46 ();
 FILLCELL_X2 FILLER_60_50 ();
 FILLCELL_X1 FILLER_60_52 ();
 FILLCELL_X4 FILLER_60_56 ();
 FILLCELL_X4 FILLER_60_63 ();
 FILLCELL_X2 FILLER_60_67 ();
 FILLCELL_X4 FILLER_60_78 ();
 FILLCELL_X4 FILLER_60_85 ();
 FILLCELL_X8 FILLER_60_95 ();
 FILLCELL_X1 FILLER_60_103 ();
 FILLCELL_X4 FILLER_60_109 ();
 FILLCELL_X1 FILLER_60_113 ();
 FILLCELL_X8 FILLER_60_118 ();
 FILLCELL_X4 FILLER_60_126 ();
 FILLCELL_X4 FILLER_60_135 ();
 FILLCELL_X8 FILLER_60_148 ();
 FILLCELL_X8 FILLER_60_160 ();
 FILLCELL_X4 FILLER_60_168 ();
 FILLCELL_X2 FILLER_60_172 ();
 FILLCELL_X8 FILLER_60_178 ();
 FILLCELL_X4 FILLER_60_186 ();
 FILLCELL_X4 FILLER_60_194 ();
 FILLCELL_X1 FILLER_60_198 ();
 FILLCELL_X8 FILLER_60_208 ();
 FILLCELL_X4 FILLER_60_216 ();
 FILLCELL_X2 FILLER_60_220 ();
 FILLCELL_X1 FILLER_60_222 ();
 FILLCELL_X4 FILLER_60_227 ();
 FILLCELL_X32 FILLER_60_236 ();
 FILLCELL_X2 FILLER_60_268 ();
 FILLCELL_X1 FILLER_60_270 ();
 FILLCELL_X4 FILLER_60_274 ();
 FILLCELL_X4 FILLER_60_281 ();
 FILLCELL_X1 FILLER_60_285 ();
 FILLCELL_X16 FILLER_60_289 ();
 FILLCELL_X8 FILLER_60_305 ();
 FILLCELL_X4 FILLER_60_313 ();
 FILLCELL_X4 FILLER_60_321 ();
 FILLCELL_X2 FILLER_60_325 ();
 FILLCELL_X4 FILLER_60_331 ();
 FILLCELL_X2 FILLER_60_335 ();
 FILLCELL_X1 FILLER_60_337 ();
 FILLCELL_X8 FILLER_60_343 ();
 FILLCELL_X4 FILLER_60_351 ();
 FILLCELL_X16 FILLER_60_358 ();
 FILLCELL_X4 FILLER_60_374 ();
 FILLCELL_X2 FILLER_60_378 ();
 FILLCELL_X32 FILLER_60_1518 ();
 FILLCELL_X32 FILLER_60_1550 ();
 FILLCELL_X32 FILLER_60_1582 ();
 FILLCELL_X32 FILLER_60_1614 ();
 FILLCELL_X32 FILLER_60_1646 ();
 FILLCELL_X32 FILLER_60_1678 ();
 FILLCELL_X32 FILLER_60_1710 ();
 FILLCELL_X8 FILLER_60_1742 ();
 FILLCELL_X4 FILLER_60_1750 ();
 FILLCELL_X2 FILLER_60_1754 ();
 FILLCELL_X8 FILLER_61_1 ();
 FILLCELL_X4 FILLER_61_9 ();
 FILLCELL_X4 FILLER_61_19 ();
 FILLCELL_X4 FILLER_61_28 ();
 FILLCELL_X1 FILLER_61_32 ();
 FILLCELL_X4 FILLER_61_37 ();
 FILLCELL_X4 FILLER_61_46 ();
 FILLCELL_X2 FILLER_61_50 ();
 FILLCELL_X8 FILLER_61_55 ();
 FILLCELL_X4 FILLER_61_63 ();
 FILLCELL_X1 FILLER_61_67 ();
 FILLCELL_X4 FILLER_61_72 ();
 FILLCELL_X8 FILLER_61_85 ();
 FILLCELL_X2 FILLER_61_93 ();
 FILLCELL_X4 FILLER_61_104 ();
 FILLCELL_X8 FILLER_61_117 ();
 FILLCELL_X4 FILLER_61_125 ();
 FILLCELL_X4 FILLER_61_135 ();
 FILLCELL_X1 FILLER_61_139 ();
 FILLCELL_X4 FILLER_61_149 ();
 FILLCELL_X2 FILLER_61_153 ();
 FILLCELL_X4 FILLER_61_159 ();
 FILLCELL_X1 FILLER_61_163 ();
 FILLCELL_X4 FILLER_61_167 ();
 FILLCELL_X4 FILLER_61_177 ();
 FILLCELL_X4 FILLER_61_185 ();
 FILLCELL_X1 FILLER_61_189 ();
 FILLCELL_X4 FILLER_61_194 ();
 FILLCELL_X4 FILLER_61_202 ();
 FILLCELL_X16 FILLER_61_210 ();
 FILLCELL_X8 FILLER_61_226 ();
 FILLCELL_X4 FILLER_61_234 ();
 FILLCELL_X4 FILLER_61_242 ();
 FILLCELL_X8 FILLER_61_250 ();
 FILLCELL_X2 FILLER_61_258 ();
 FILLCELL_X8 FILLER_61_269 ();
 FILLCELL_X8 FILLER_61_280 ();
 FILLCELL_X4 FILLER_61_288 ();
 FILLCELL_X4 FILLER_61_296 ();
 FILLCELL_X4 FILLER_61_306 ();
 FILLCELL_X16 FILLER_61_315 ();
 FILLCELL_X1 FILLER_61_331 ();
 FILLCELL_X4 FILLER_61_335 ();
 FILLCELL_X4 FILLER_61_342 ();
 FILLCELL_X4 FILLER_61_353 ();
 FILLCELL_X4 FILLER_61_361 ();
 FILLCELL_X8 FILLER_61_368 ();
 FILLCELL_X4 FILLER_61_376 ();
 FILLCELL_X32 FILLER_61_1518 ();
 FILLCELL_X32 FILLER_61_1550 ();
 FILLCELL_X32 FILLER_61_1582 ();
 FILLCELL_X32 FILLER_61_1614 ();
 FILLCELL_X32 FILLER_61_1646 ();
 FILLCELL_X32 FILLER_61_1678 ();
 FILLCELL_X32 FILLER_61_1710 ();
 FILLCELL_X8 FILLER_61_1742 ();
 FILLCELL_X4 FILLER_61_1750 ();
 FILLCELL_X2 FILLER_61_1754 ();
 FILLCELL_X4 FILLER_62_1 ();
 FILLCELL_X4 FILLER_62_12 ();
 FILLCELL_X4 FILLER_62_20 ();
 FILLCELL_X2 FILLER_62_24 ();
 FILLCELL_X1 FILLER_62_26 ();
 FILLCELL_X4 FILLER_62_31 ();
 FILLCELL_X4 FILLER_62_44 ();
 FILLCELL_X4 FILLER_62_57 ();
 FILLCELL_X8 FILLER_62_67 ();
 FILLCELL_X2 FILLER_62_75 ();
 FILLCELL_X1 FILLER_62_77 ();
 FILLCELL_X8 FILLER_62_83 ();
 FILLCELL_X4 FILLER_62_94 ();
 FILLCELL_X4 FILLER_62_102 ();
 FILLCELL_X4 FILLER_62_110 ();
 FILLCELL_X4 FILLER_62_118 ();
 FILLCELL_X4 FILLER_62_127 ();
 FILLCELL_X2 FILLER_62_131 ();
 FILLCELL_X1 FILLER_62_133 ();
 FILLCELL_X4 FILLER_62_138 ();
 FILLCELL_X8 FILLER_62_151 ();
 FILLCELL_X1 FILLER_62_159 ();
 FILLCELL_X4 FILLER_62_169 ();
 FILLCELL_X4 FILLER_62_182 ();
 FILLCELL_X8 FILLER_62_190 ();
 FILLCELL_X1 FILLER_62_198 ();
 FILLCELL_X4 FILLER_62_203 ();
 FILLCELL_X2 FILLER_62_207 ();
 FILLCELL_X1 FILLER_62_209 ();
 FILLCELL_X8 FILLER_62_214 ();
 FILLCELL_X2 FILLER_62_222 ();
 FILLCELL_X8 FILLER_62_233 ();
 FILLCELL_X1 FILLER_62_241 ();
 FILLCELL_X4 FILLER_62_246 ();
 FILLCELL_X8 FILLER_62_259 ();
 FILLCELL_X2 FILLER_62_267 ();
 FILLCELL_X8 FILLER_62_275 ();
 FILLCELL_X1 FILLER_62_283 ();
 FILLCELL_X4 FILLER_62_293 ();
 FILLCELL_X4 FILLER_62_306 ();
 FILLCELL_X8 FILLER_62_313 ();
 FILLCELL_X4 FILLER_62_330 ();
 FILLCELL_X1 FILLER_62_334 ();
 FILLCELL_X4 FILLER_62_341 ();
 FILLCELL_X4 FILLER_62_351 ();
 FILLCELL_X2 FILLER_62_355 ();
 FILLCELL_X4 FILLER_62_376 ();
 FILLCELL_X32 FILLER_62_1518 ();
 FILLCELL_X32 FILLER_62_1550 ();
 FILLCELL_X32 FILLER_62_1582 ();
 FILLCELL_X32 FILLER_62_1614 ();
 FILLCELL_X32 FILLER_62_1646 ();
 FILLCELL_X32 FILLER_62_1678 ();
 FILLCELL_X32 FILLER_62_1710 ();
 FILLCELL_X8 FILLER_62_1742 ();
 FILLCELL_X4 FILLER_62_1750 ();
 FILLCELL_X2 FILLER_62_1754 ();
 FILLCELL_X4 FILLER_63_1 ();
 FILLCELL_X4 FILLER_63_24 ();
 FILLCELL_X1 FILLER_63_28 ();
 FILLCELL_X4 FILLER_63_33 ();
 FILLCELL_X4 FILLER_63_41 ();
 FILLCELL_X2 FILLER_63_45 ();
 FILLCELL_X8 FILLER_63_51 ();
 FILLCELL_X2 FILLER_63_59 ();
 FILLCELL_X4 FILLER_63_64 ();
 FILLCELL_X1 FILLER_63_68 ();
 FILLCELL_X8 FILLER_63_74 ();
 FILLCELL_X4 FILLER_63_82 ();
 FILLCELL_X2 FILLER_63_86 ();
 FILLCELL_X1 FILLER_63_88 ();
 FILLCELL_X4 FILLER_63_93 ();
 FILLCELL_X4 FILLER_63_100 ();
 FILLCELL_X2 FILLER_63_104 ();
 FILLCELL_X16 FILLER_63_110 ();
 FILLCELL_X4 FILLER_63_126 ();
 FILLCELL_X1 FILLER_63_130 ();
 FILLCELL_X16 FILLER_63_134 ();
 FILLCELL_X4 FILLER_63_150 ();
 FILLCELL_X2 FILLER_63_154 ();
 FILLCELL_X1 FILLER_63_156 ();
 FILLCELL_X4 FILLER_63_160 ();
 FILLCELL_X1 FILLER_63_164 ();
 FILLCELL_X4 FILLER_63_170 ();
 FILLCELL_X1 FILLER_63_174 ();
 FILLCELL_X8 FILLER_63_180 ();
 FILLCELL_X2 FILLER_63_188 ();
 FILLCELL_X4 FILLER_63_195 ();
 FILLCELL_X4 FILLER_63_208 ();
 FILLCELL_X2 FILLER_63_212 ();
 FILLCELL_X1 FILLER_63_214 ();
 FILLCELL_X4 FILLER_63_219 ();
 FILLCELL_X4 FILLER_63_227 ();
 FILLCELL_X4 FILLER_63_235 ();
 FILLCELL_X2 FILLER_63_239 ();
 FILLCELL_X1 FILLER_63_241 ();
 FILLCELL_X4 FILLER_63_246 ();
 FILLCELL_X2 FILLER_63_250 ();
 FILLCELL_X1 FILLER_63_252 ();
 FILLCELL_X4 FILLER_63_257 ();
 FILLCELL_X4 FILLER_63_266 ();
 FILLCELL_X16 FILLER_63_273 ();
 FILLCELL_X4 FILLER_63_289 ();
 FILLCELL_X2 FILLER_63_293 ();
 FILLCELL_X4 FILLER_63_300 ();
 FILLCELL_X8 FILLER_63_307 ();
 FILLCELL_X1 FILLER_63_315 ();
 FILLCELL_X4 FILLER_63_320 ();
 FILLCELL_X4 FILLER_63_330 ();
 FILLCELL_X8 FILLER_63_337 ();
 FILLCELL_X4 FILLER_63_345 ();
 FILLCELL_X2 FILLER_63_349 ();
 FILLCELL_X1 FILLER_63_351 ();
 FILLCELL_X4 FILLER_63_357 ();
 FILLCELL_X16 FILLER_63_364 ();
 FILLCELL_X4 FILLER_63_1518 ();
 FILLCELL_X32 FILLER_63_1541 ();
 FILLCELL_X32 FILLER_63_1573 ();
 FILLCELL_X32 FILLER_63_1605 ();
 FILLCELL_X32 FILLER_63_1637 ();
 FILLCELL_X32 FILLER_63_1669 ();
 FILLCELL_X32 FILLER_63_1701 ();
 FILLCELL_X16 FILLER_63_1733 ();
 FILLCELL_X4 FILLER_63_1749 ();
 FILLCELL_X2 FILLER_63_1753 ();
 FILLCELL_X1 FILLER_63_1755 ();
 FILLCELL_X4 FILLER_64_1 ();
 FILLCELL_X4 FILLER_64_11 ();
 FILLCELL_X4 FILLER_64_19 ();
 FILLCELL_X16 FILLER_64_36 ();
 FILLCELL_X8 FILLER_64_52 ();
 FILLCELL_X4 FILLER_64_60 ();
 FILLCELL_X1 FILLER_64_64 ();
 FILLCELL_X4 FILLER_64_71 ();
 FILLCELL_X4 FILLER_64_79 ();
 FILLCELL_X1 FILLER_64_83 ();
 FILLCELL_X4 FILLER_64_88 ();
 FILLCELL_X2 FILLER_64_92 ();
 FILLCELL_X1 FILLER_64_94 ();
 FILLCELL_X8 FILLER_64_104 ();
 FILLCELL_X4 FILLER_64_116 ();
 FILLCELL_X1 FILLER_64_120 ();
 FILLCELL_X4 FILLER_64_125 ();
 FILLCELL_X4 FILLER_64_133 ();
 FILLCELL_X4 FILLER_64_142 ();
 FILLCELL_X4 FILLER_64_151 ();
 FILLCELL_X8 FILLER_64_161 ();
 FILLCELL_X4 FILLER_64_174 ();
 FILLCELL_X8 FILLER_64_182 ();
 FILLCELL_X2 FILLER_64_190 ();
 FILLCELL_X4 FILLER_64_195 ();
 FILLCELL_X32 FILLER_64_208 ();
 FILLCELL_X2 FILLER_64_240 ();
 FILLCELL_X1 FILLER_64_242 ();
 FILLCELL_X8 FILLER_64_247 ();
 FILLCELL_X4 FILLER_64_255 ();
 FILLCELL_X1 FILLER_64_259 ();
 FILLCELL_X4 FILLER_64_263 ();
 FILLCELL_X4 FILLER_64_272 ();
 FILLCELL_X1 FILLER_64_276 ();
 FILLCELL_X4 FILLER_64_286 ();
 FILLCELL_X4 FILLER_64_294 ();
 FILLCELL_X4 FILLER_64_301 ();
 FILLCELL_X4 FILLER_64_308 ();
 FILLCELL_X1 FILLER_64_312 ();
 FILLCELL_X4 FILLER_64_322 ();
 FILLCELL_X4 FILLER_64_331 ();
 FILLCELL_X2 FILLER_64_335 ();
 FILLCELL_X8 FILLER_64_347 ();
 FILLCELL_X4 FILLER_64_355 ();
 FILLCELL_X4 FILLER_64_368 ();
 FILLCELL_X4 FILLER_64_375 ();
 FILLCELL_X1 FILLER_64_379 ();
 FILLCELL_X4 FILLER_64_1518 ();
 FILLCELL_X4 FILLER_64_1526 ();
 FILLCELL_X32 FILLER_64_1534 ();
 FILLCELL_X32 FILLER_64_1566 ();
 FILLCELL_X32 FILLER_64_1598 ();
 FILLCELL_X32 FILLER_64_1630 ();
 FILLCELL_X32 FILLER_64_1662 ();
 FILLCELL_X32 FILLER_64_1694 ();
 FILLCELL_X16 FILLER_64_1726 ();
 FILLCELL_X8 FILLER_64_1742 ();
 FILLCELL_X4 FILLER_64_1750 ();
 FILLCELL_X2 FILLER_64_1754 ();
 FILLCELL_X8 FILLER_65_1 ();
 FILLCELL_X2 FILLER_65_9 ();
 FILLCELL_X1 FILLER_65_11 ();
 FILLCELL_X4 FILLER_65_18 ();
 FILLCELL_X16 FILLER_65_26 ();
 FILLCELL_X8 FILLER_65_42 ();
 FILLCELL_X4 FILLER_65_53 ();
 FILLCELL_X4 FILLER_65_66 ();
 FILLCELL_X8 FILLER_65_79 ();
 FILLCELL_X1 FILLER_65_87 ();
 FILLCELL_X4 FILLER_65_92 ();
 FILLCELL_X8 FILLER_65_105 ();
 FILLCELL_X2 FILLER_65_113 ();
 FILLCELL_X1 FILLER_65_115 ();
 FILLCELL_X4 FILLER_65_125 ();
 FILLCELL_X4 FILLER_65_138 ();
 FILLCELL_X2 FILLER_65_142 ();
 FILLCELL_X8 FILLER_65_153 ();
 FILLCELL_X2 FILLER_65_161 ();
 FILLCELL_X4 FILLER_65_169 ();
 FILLCELL_X4 FILLER_65_182 ();
 FILLCELL_X8 FILLER_65_189 ();
 FILLCELL_X8 FILLER_65_202 ();
 FILLCELL_X4 FILLER_65_214 ();
 FILLCELL_X4 FILLER_65_222 ();
 FILLCELL_X2 FILLER_65_226 ();
 FILLCELL_X4 FILLER_65_234 ();
 FILLCELL_X2 FILLER_65_238 ();
 FILLCELL_X1 FILLER_65_240 ();
 FILLCELL_X4 FILLER_65_244 ();
 FILLCELL_X4 FILLER_65_257 ();
 FILLCELL_X8 FILLER_65_267 ();
 FILLCELL_X2 FILLER_65_275 ();
 FILLCELL_X4 FILLER_65_286 ();
 FILLCELL_X4 FILLER_65_296 ();
 FILLCELL_X2 FILLER_65_300 ();
 FILLCELL_X1 FILLER_65_302 ();
 FILLCELL_X16 FILLER_65_306 ();
 FILLCELL_X8 FILLER_65_322 ();
 FILLCELL_X1 FILLER_65_330 ();
 FILLCELL_X8 FILLER_65_334 ();
 FILLCELL_X4 FILLER_65_345 ();
 FILLCELL_X4 FILLER_65_355 ();
 FILLCELL_X8 FILLER_65_368 ();
 FILLCELL_X4 FILLER_65_376 ();
 FILLCELL_X4 FILLER_65_1518 ();
 FILLCELL_X1 FILLER_65_1522 ();
 FILLCELL_X32 FILLER_65_1542 ();
 FILLCELL_X32 FILLER_65_1574 ();
 FILLCELL_X32 FILLER_65_1606 ();
 FILLCELL_X32 FILLER_65_1638 ();
 FILLCELL_X32 FILLER_65_1670 ();
 FILLCELL_X32 FILLER_65_1702 ();
 FILLCELL_X16 FILLER_65_1734 ();
 FILLCELL_X4 FILLER_65_1750 ();
 FILLCELL_X2 FILLER_65_1754 ();
 FILLCELL_X8 FILLER_66_1 ();
 FILLCELL_X8 FILLER_66_13 ();
 FILLCELL_X4 FILLER_66_21 ();
 FILLCELL_X4 FILLER_66_28 ();
 FILLCELL_X4 FILLER_66_35 ();
 FILLCELL_X4 FILLER_66_48 ();
 FILLCELL_X2 FILLER_66_52 ();
 FILLCELL_X1 FILLER_66_54 ();
 FILLCELL_X4 FILLER_66_58 ();
 FILLCELL_X4 FILLER_66_67 ();
 FILLCELL_X16 FILLER_66_76 ();
 FILLCELL_X1 FILLER_66_92 ();
 FILLCELL_X4 FILLER_66_102 ();
 FILLCELL_X8 FILLER_66_110 ();
 FILLCELL_X4 FILLER_66_118 ();
 FILLCELL_X2 FILLER_66_122 ();
 FILLCELL_X8 FILLER_66_128 ();
 FILLCELL_X4 FILLER_66_136 ();
 FILLCELL_X2 FILLER_66_140 ();
 FILLCELL_X4 FILLER_66_146 ();
 FILLCELL_X8 FILLER_66_153 ();
 FILLCELL_X4 FILLER_66_161 ();
 FILLCELL_X2 FILLER_66_165 ();
 FILLCELL_X1 FILLER_66_167 ();
 FILLCELL_X4 FILLER_66_171 ();
 FILLCELL_X4 FILLER_66_184 ();
 FILLCELL_X1 FILLER_66_188 ();
 FILLCELL_X4 FILLER_66_195 ();
 FILLCELL_X4 FILLER_66_208 ();
 FILLCELL_X2 FILLER_66_212 ();
 FILLCELL_X4 FILLER_66_223 ();
 FILLCELL_X4 FILLER_66_236 ();
 FILLCELL_X8 FILLER_66_244 ();
 FILLCELL_X2 FILLER_66_252 ();
 FILLCELL_X4 FILLER_66_263 ();
 FILLCELL_X4 FILLER_66_271 ();
 FILLCELL_X2 FILLER_66_275 ();
 FILLCELL_X4 FILLER_66_286 ();
 FILLCELL_X2 FILLER_66_290 ();
 FILLCELL_X1 FILLER_66_292 ();
 FILLCELL_X4 FILLER_66_298 ();
 FILLCELL_X4 FILLER_66_308 ();
 FILLCELL_X4 FILLER_66_315 ();
 FILLCELL_X4 FILLER_66_323 ();
 FILLCELL_X16 FILLER_66_333 ();
 FILLCELL_X8 FILLER_66_349 ();
 FILLCELL_X1 FILLER_66_357 ();
 FILLCELL_X16 FILLER_66_362 ();
 FILLCELL_X2 FILLER_66_378 ();
 FILLCELL_X32 FILLER_66_1518 ();
 FILLCELL_X32 FILLER_66_1550 ();
 FILLCELL_X32 FILLER_66_1582 ();
 FILLCELL_X32 FILLER_66_1614 ();
 FILLCELL_X32 FILLER_66_1646 ();
 FILLCELL_X32 FILLER_66_1678 ();
 FILLCELL_X32 FILLER_66_1710 ();
 FILLCELL_X8 FILLER_66_1742 ();
 FILLCELL_X4 FILLER_66_1750 ();
 FILLCELL_X2 FILLER_66_1754 ();
 FILLCELL_X4 FILLER_67_1 ();
 FILLCELL_X4 FILLER_67_24 ();
 FILLCELL_X1 FILLER_67_28 ();
 FILLCELL_X4 FILLER_67_35 ();
 FILLCELL_X4 FILLER_67_48 ();
 FILLCELL_X16 FILLER_67_57 ();
 FILLCELL_X2 FILLER_67_73 ();
 FILLCELL_X4 FILLER_67_78 ();
 FILLCELL_X2 FILLER_67_82 ();
 FILLCELL_X4 FILLER_67_87 ();
 FILLCELL_X4 FILLER_67_97 ();
 FILLCELL_X4 FILLER_67_104 ();
 FILLCELL_X2 FILLER_67_108 ();
 FILLCELL_X4 FILLER_67_114 ();
 FILLCELL_X4 FILLER_67_124 ();
 FILLCELL_X4 FILLER_67_133 ();
 FILLCELL_X2 FILLER_67_137 ();
 FILLCELL_X1 FILLER_67_139 ();
 FILLCELL_X4 FILLER_67_143 ();
 FILLCELL_X1 FILLER_67_147 ();
 FILLCELL_X16 FILLER_67_152 ();
 FILLCELL_X4 FILLER_67_168 ();
 FILLCELL_X16 FILLER_67_181 ();
 FILLCELL_X4 FILLER_67_201 ();
 FILLCELL_X4 FILLER_67_209 ();
 FILLCELL_X2 FILLER_67_213 ();
 FILLCELL_X4 FILLER_67_219 ();
 FILLCELL_X2 FILLER_67_223 ();
 FILLCELL_X1 FILLER_67_225 ();
 FILLCELL_X8 FILLER_67_231 ();
 FILLCELL_X4 FILLER_67_242 ();
 FILLCELL_X1 FILLER_67_246 ();
 FILLCELL_X4 FILLER_67_250 ();
 FILLCELL_X16 FILLER_67_263 ();
 FILLCELL_X8 FILLER_67_279 ();
 FILLCELL_X1 FILLER_67_287 ();
 FILLCELL_X8 FILLER_67_293 ();
 FILLCELL_X2 FILLER_67_301 ();
 FILLCELL_X4 FILLER_67_312 ();
 FILLCELL_X4 FILLER_67_321 ();
 FILLCELL_X2 FILLER_67_325 ();
 FILLCELL_X1 FILLER_67_327 ();
 FILLCELL_X16 FILLER_67_341 ();
 FILLCELL_X2 FILLER_67_357 ();
 FILLCELL_X4 FILLER_67_362 ();
 FILLCELL_X8 FILLER_67_370 ();
 FILLCELL_X2 FILLER_67_378 ();
 FILLCELL_X32 FILLER_67_1518 ();
 FILLCELL_X32 FILLER_67_1550 ();
 FILLCELL_X32 FILLER_67_1582 ();
 FILLCELL_X32 FILLER_67_1614 ();
 FILLCELL_X32 FILLER_67_1646 ();
 FILLCELL_X32 FILLER_67_1678 ();
 FILLCELL_X32 FILLER_67_1710 ();
 FILLCELL_X8 FILLER_67_1742 ();
 FILLCELL_X4 FILLER_67_1750 ();
 FILLCELL_X2 FILLER_67_1754 ();
 FILLCELL_X32 FILLER_68_1 ();
 FILLCELL_X2 FILLER_68_33 ();
 FILLCELL_X1 FILLER_68_35 ();
 FILLCELL_X4 FILLER_68_39 ();
 FILLCELL_X16 FILLER_68_47 ();
 FILLCELL_X1 FILLER_68_63 ();
 FILLCELL_X4 FILLER_68_73 ();
 FILLCELL_X2 FILLER_68_77 ();
 FILLCELL_X1 FILLER_68_79 ();
 FILLCELL_X8 FILLER_68_84 ();
 FILLCELL_X2 FILLER_68_92 ();
 FILLCELL_X4 FILLER_68_99 ();
 FILLCELL_X8 FILLER_68_108 ();
 FILLCELL_X2 FILLER_68_116 ();
 FILLCELL_X4 FILLER_68_127 ();
 FILLCELL_X8 FILLER_68_136 ();
 FILLCELL_X1 FILLER_68_144 ();
 FILLCELL_X8 FILLER_68_154 ();
 FILLCELL_X2 FILLER_68_162 ();
 FILLCELL_X1 FILLER_68_164 ();
 FILLCELL_X4 FILLER_68_170 ();
 FILLCELL_X2 FILLER_68_174 ();
 FILLCELL_X1 FILLER_68_176 ();
 FILLCELL_X4 FILLER_68_180 ();
 FILLCELL_X32 FILLER_68_187 ();
 FILLCELL_X16 FILLER_68_219 ();
 FILLCELL_X1 FILLER_68_235 ();
 FILLCELL_X4 FILLER_68_239 ();
 FILLCELL_X4 FILLER_68_246 ();
 FILLCELL_X2 FILLER_68_250 ();
 FILLCELL_X1 FILLER_68_252 ();
 FILLCELL_X16 FILLER_68_262 ();
 FILLCELL_X4 FILLER_68_282 ();
 FILLCELL_X2 FILLER_68_286 ();
 FILLCELL_X1 FILLER_68_288 ();
 FILLCELL_X4 FILLER_68_296 ();
 FILLCELL_X2 FILLER_68_300 ();
 FILLCELL_X4 FILLER_68_311 ();
 FILLCELL_X4 FILLER_68_319 ();
 FILLCELL_X2 FILLER_68_323 ();
 FILLCELL_X8 FILLER_68_329 ();
 FILLCELL_X1 FILLER_68_337 ();
 FILLCELL_X4 FILLER_68_342 ();
 FILLCELL_X4 FILLER_68_350 ();
 FILLCELL_X4 FILLER_68_357 ();
 FILLCELL_X8 FILLER_68_370 ();
 FILLCELL_X2 FILLER_68_378 ();
 FILLCELL_X4 FILLER_68_1518 ();
 FILLCELL_X2 FILLER_68_1522 ();
 FILLCELL_X1 FILLER_68_1524 ();
 FILLCELL_X32 FILLER_68_1544 ();
 FILLCELL_X32 FILLER_68_1576 ();
 FILLCELL_X32 FILLER_68_1608 ();
 FILLCELL_X32 FILLER_68_1640 ();
 FILLCELL_X32 FILLER_68_1672 ();
 FILLCELL_X32 FILLER_68_1704 ();
 FILLCELL_X8 FILLER_68_1736 ();
 FILLCELL_X4 FILLER_68_1744 ();
 FILLCELL_X1 FILLER_68_1748 ();
 FILLCELL_X4 FILLER_68_1752 ();
 FILLCELL_X4 FILLER_69_1 ();
 FILLCELL_X4 FILLER_69_22 ();
 FILLCELL_X4 FILLER_69_29 ();
 FILLCELL_X1 FILLER_69_33 ();
 FILLCELL_X8 FILLER_69_37 ();
 FILLCELL_X4 FILLER_69_45 ();
 FILLCELL_X2 FILLER_69_49 ();
 FILLCELL_X1 FILLER_69_51 ();
 FILLCELL_X4 FILLER_69_55 ();
 FILLCELL_X4 FILLER_69_65 ();
 FILLCELL_X8 FILLER_69_78 ();
 FILLCELL_X2 FILLER_69_86 ();
 FILLCELL_X1 FILLER_69_88 ();
 FILLCELL_X4 FILLER_69_93 ();
 FILLCELL_X4 FILLER_69_101 ();
 FILLCELL_X4 FILLER_69_114 ();
 FILLCELL_X8 FILLER_69_127 ();
 FILLCELL_X1 FILLER_69_135 ();
 FILLCELL_X4 FILLER_69_142 ();
 FILLCELL_X4 FILLER_69_155 ();
 FILLCELL_X4 FILLER_69_163 ();
 FILLCELL_X4 FILLER_69_173 ();
 FILLCELL_X4 FILLER_69_186 ();
 FILLCELL_X2 FILLER_69_190 ();
 FILLCELL_X1 FILLER_69_192 ();
 FILLCELL_X4 FILLER_69_197 ();
 FILLCELL_X4 FILLER_69_205 ();
 FILLCELL_X8 FILLER_69_213 ();
 FILLCELL_X4 FILLER_69_224 ();
 FILLCELL_X8 FILLER_69_234 ();
 FILLCELL_X1 FILLER_69_242 ();
 FILLCELL_X4 FILLER_69_247 ();
 FILLCELL_X4 FILLER_69_255 ();
 FILLCELL_X4 FILLER_69_263 ();
 FILLCELL_X4 FILLER_69_273 ();
 FILLCELL_X8 FILLER_69_287 ();
 FILLCELL_X4 FILLER_69_295 ();
 FILLCELL_X1 FILLER_69_299 ();
 FILLCELL_X8 FILLER_69_309 ();
 FILLCELL_X8 FILLER_69_321 ();
 FILLCELL_X1 FILLER_69_329 ();
 FILLCELL_X4 FILLER_69_336 ();
 FILLCELL_X4 FILLER_69_347 ();
 FILLCELL_X4 FILLER_69_357 ();
 FILLCELL_X8 FILLER_69_370 ();
 FILLCELL_X2 FILLER_69_378 ();
 FILLCELL_X4 FILLER_69_1518 ();
 FILLCELL_X32 FILLER_69_1526 ();
 FILLCELL_X32 FILLER_69_1558 ();
 FILLCELL_X32 FILLER_69_1590 ();
 FILLCELL_X32 FILLER_69_1622 ();
 FILLCELL_X32 FILLER_69_1654 ();
 FILLCELL_X32 FILLER_69_1686 ();
 FILLCELL_X32 FILLER_69_1718 ();
 FILLCELL_X4 FILLER_69_1750 ();
 FILLCELL_X2 FILLER_69_1754 ();
 FILLCELL_X4 FILLER_70_1 ();
 FILLCELL_X2 FILLER_70_5 ();
 FILLCELL_X4 FILLER_70_11 ();
 FILLCELL_X8 FILLER_70_19 ();
 FILLCELL_X2 FILLER_70_27 ();
 FILLCELL_X4 FILLER_70_36 ();
 FILLCELL_X4 FILLER_70_46 ();
 FILLCELL_X8 FILLER_70_53 ();
 FILLCELL_X4 FILLER_70_61 ();
 FILLCELL_X2 FILLER_70_65 ();
 FILLCELL_X1 FILLER_70_67 ();
 FILLCELL_X4 FILLER_70_73 ();
 FILLCELL_X16 FILLER_70_80 ();
 FILLCELL_X1 FILLER_70_96 ();
 FILLCELL_X4 FILLER_70_101 ();
 FILLCELL_X8 FILLER_70_109 ();
 FILLCELL_X4 FILLER_70_117 ();
 FILLCELL_X2 FILLER_70_121 ();
 FILLCELL_X1 FILLER_70_123 ();
 FILLCELL_X4 FILLER_70_127 ();
 FILLCELL_X8 FILLER_70_134 ();
 FILLCELL_X4 FILLER_70_147 ();
 FILLCELL_X16 FILLER_70_155 ();
 FILLCELL_X4 FILLER_70_180 ();
 FILLCELL_X4 FILLER_70_188 ();
 FILLCELL_X1 FILLER_70_192 ();
 FILLCELL_X4 FILLER_70_197 ();
 FILLCELL_X4 FILLER_70_210 ();
 FILLCELL_X4 FILLER_70_223 ();
 FILLCELL_X4 FILLER_70_236 ();
 FILLCELL_X16 FILLER_70_244 ();
 FILLCELL_X1 FILLER_70_260 ();
 FILLCELL_X4 FILLER_70_266 ();
 FILLCELL_X4 FILLER_70_274 ();
 FILLCELL_X16 FILLER_70_282 ();
 FILLCELL_X4 FILLER_70_302 ();
 FILLCELL_X4 FILLER_70_310 ();
 FILLCELL_X8 FILLER_70_318 ();
 FILLCELL_X2 FILLER_70_326 ();
 FILLCELL_X4 FILLER_70_337 ();
 FILLCELL_X4 FILLER_70_348 ();
 FILLCELL_X4 FILLER_70_358 ();
 FILLCELL_X4 FILLER_70_367 ();
 FILLCELL_X4 FILLER_70_375 ();
 FILLCELL_X1 FILLER_70_379 ();
 FILLCELL_X4 FILLER_70_1518 ();
 FILLCELL_X2 FILLER_70_1522 ();
 FILLCELL_X32 FILLER_70_1543 ();
 FILLCELL_X32 FILLER_70_1575 ();
 FILLCELL_X32 FILLER_70_1607 ();
 FILLCELL_X32 FILLER_70_1639 ();
 FILLCELL_X32 FILLER_70_1671 ();
 FILLCELL_X32 FILLER_70_1703 ();
 FILLCELL_X16 FILLER_70_1735 ();
 FILLCELL_X4 FILLER_70_1751 ();
 FILLCELL_X1 FILLER_70_1755 ();
 FILLCELL_X4 FILLER_71_1 ();
 FILLCELL_X4 FILLER_71_24 ();
 FILLCELL_X4 FILLER_71_34 ();
 FILLCELL_X4 FILLER_71_41 ();
 FILLCELL_X2 FILLER_71_45 ();
 FILLCELL_X1 FILLER_71_47 ();
 FILLCELL_X4 FILLER_71_51 ();
 FILLCELL_X8 FILLER_71_64 ();
 FILLCELL_X1 FILLER_71_72 ();
 FILLCELL_X4 FILLER_71_76 ();
 FILLCELL_X4 FILLER_71_83 ();
 FILLCELL_X4 FILLER_71_96 ();
 FILLCELL_X2 FILLER_71_100 ();
 FILLCELL_X1 FILLER_71_102 ();
 FILLCELL_X4 FILLER_71_107 ();
 FILLCELL_X1 FILLER_71_111 ();
 FILLCELL_X4 FILLER_71_117 ();
 FILLCELL_X4 FILLER_71_126 ();
 FILLCELL_X8 FILLER_71_133 ();
 FILLCELL_X4 FILLER_71_141 ();
 FILLCELL_X8 FILLER_71_154 ();
 FILLCELL_X4 FILLER_71_162 ();
 FILLCELL_X2 FILLER_71_166 ();
 FILLCELL_X8 FILLER_71_177 ();
 FILLCELL_X32 FILLER_71_189 ();
 FILLCELL_X2 FILLER_71_221 ();
 FILLCELL_X1 FILLER_71_223 ();
 FILLCELL_X4 FILLER_71_228 ();
 FILLCELL_X1 FILLER_71_232 ();
 FILLCELL_X8 FILLER_71_238 ();
 FILLCELL_X4 FILLER_71_246 ();
 FILLCELL_X4 FILLER_71_254 ();
 FILLCELL_X8 FILLER_71_264 ();
 FILLCELL_X2 FILLER_71_272 ();
 FILLCELL_X1 FILLER_71_274 ();
 FILLCELL_X8 FILLER_71_279 ();
 FILLCELL_X1 FILLER_71_287 ();
 FILLCELL_X8 FILLER_71_291 ();
 FILLCELL_X2 FILLER_71_299 ();
 FILLCELL_X16 FILLER_71_304 ();
 FILLCELL_X2 FILLER_71_320 ();
 FILLCELL_X1 FILLER_71_322 ();
 FILLCELL_X4 FILLER_71_326 ();
 FILLCELL_X8 FILLER_71_340 ();
 FILLCELL_X2 FILLER_71_348 ();
 FILLCELL_X4 FILLER_71_354 ();
 FILLCELL_X4 FILLER_71_363 ();
 FILLCELL_X8 FILLER_71_371 ();
 FILLCELL_X1 FILLER_71_379 ();
 FILLCELL_X4 FILLER_71_1518 ();
 FILLCELL_X32 FILLER_71_1526 ();
 FILLCELL_X32 FILLER_71_1558 ();
 FILLCELL_X32 FILLER_71_1590 ();
 FILLCELL_X32 FILLER_71_1622 ();
 FILLCELL_X32 FILLER_71_1654 ();
 FILLCELL_X32 FILLER_71_1686 ();
 FILLCELL_X32 FILLER_71_1718 ();
 FILLCELL_X4 FILLER_71_1750 ();
 FILLCELL_X2 FILLER_71_1754 ();
 FILLCELL_X8 FILLER_72_1 ();
 FILLCELL_X4 FILLER_72_9 ();
 FILLCELL_X1 FILLER_72_13 ();
 FILLCELL_X16 FILLER_72_18 ();
 FILLCELL_X1 FILLER_72_34 ();
 FILLCELL_X8 FILLER_72_38 ();
 FILLCELL_X4 FILLER_72_46 ();
 FILLCELL_X1 FILLER_72_50 ();
 FILLCELL_X4 FILLER_72_57 ();
 FILLCELL_X4 FILLER_72_70 ();
 FILLCELL_X2 FILLER_72_74 ();
 FILLCELL_X4 FILLER_72_82 ();
 FILLCELL_X4 FILLER_72_95 ();
 FILLCELL_X2 FILLER_72_99 ();
 FILLCELL_X8 FILLER_72_105 ();
 FILLCELL_X2 FILLER_72_113 ();
 FILLCELL_X1 FILLER_72_115 ();
 FILLCELL_X4 FILLER_72_122 ();
 FILLCELL_X4 FILLER_72_131 ();
 FILLCELL_X8 FILLER_72_139 ();
 FILLCELL_X4 FILLER_72_151 ();
 FILLCELL_X4 FILLER_72_159 ();
 FILLCELL_X1 FILLER_72_163 ();
 FILLCELL_X4 FILLER_72_168 ();
 FILLCELL_X4 FILLER_72_176 ();
 FILLCELL_X4 FILLER_72_184 ();
 FILLCELL_X2 FILLER_72_188 ();
 FILLCELL_X16 FILLER_72_209 ();
 FILLCELL_X4 FILLER_72_225 ();
 FILLCELL_X1 FILLER_72_229 ();
 FILLCELL_X8 FILLER_72_234 ();
 FILLCELL_X1 FILLER_72_242 ();
 FILLCELL_X4 FILLER_72_252 ();
 FILLCELL_X4 FILLER_72_265 ();
 FILLCELL_X4 FILLER_72_278 ();
 FILLCELL_X4 FILLER_72_286 ();
 FILLCELL_X2 FILLER_72_290 ();
 FILLCELL_X1 FILLER_72_292 ();
 FILLCELL_X4 FILLER_72_299 ();
 FILLCELL_X4 FILLER_72_307 ();
 FILLCELL_X4 FILLER_72_314 ();
 FILLCELL_X4 FILLER_72_322 ();
 FILLCELL_X2 FILLER_72_326 ();
 FILLCELL_X1 FILLER_72_328 ();
 FILLCELL_X8 FILLER_72_332 ();
 FILLCELL_X4 FILLER_72_340 ();
 FILLCELL_X2 FILLER_72_344 ();
 FILLCELL_X4 FILLER_72_349 ();
 FILLCELL_X4 FILLER_72_357 ();
 FILLCELL_X8 FILLER_72_365 ();
 FILLCELL_X4 FILLER_72_373 ();
 FILLCELL_X2 FILLER_72_377 ();
 FILLCELL_X1 FILLER_72_379 ();
 FILLCELL_X8 FILLER_72_1518 ();
 FILLCELL_X1 FILLER_72_1526 ();
 FILLCELL_X32 FILLER_72_1546 ();
 FILLCELL_X32 FILLER_72_1578 ();
 FILLCELL_X32 FILLER_72_1610 ();
 FILLCELL_X32 FILLER_72_1642 ();
 FILLCELL_X32 FILLER_72_1674 ();
 FILLCELL_X32 FILLER_72_1706 ();
 FILLCELL_X16 FILLER_72_1738 ();
 FILLCELL_X2 FILLER_72_1754 ();
 FILLCELL_X4 FILLER_73_1 ();
 FILLCELL_X16 FILLER_73_8 ();
 FILLCELL_X2 FILLER_73_24 ();
 FILLCELL_X4 FILLER_73_32 ();
 FILLCELL_X4 FILLER_73_45 ();
 FILLCELL_X2 FILLER_73_49 ();
 FILLCELL_X1 FILLER_73_51 ();
 FILLCELL_X4 FILLER_73_55 ();
 FILLCELL_X4 FILLER_73_64 ();
 FILLCELL_X8 FILLER_73_72 ();
 FILLCELL_X4 FILLER_73_83 ();
 FILLCELL_X8 FILLER_73_92 ();
 FILLCELL_X2 FILLER_73_100 ();
 FILLCELL_X1 FILLER_73_102 ();
 FILLCELL_X4 FILLER_73_112 ();
 FILLCELL_X4 FILLER_73_125 ();
 FILLCELL_X8 FILLER_73_138 ();
 FILLCELL_X2 FILLER_73_146 ();
 FILLCELL_X32 FILLER_73_152 ();
 FILLCELL_X16 FILLER_73_184 ();
 FILLCELL_X4 FILLER_73_203 ();
 FILLCELL_X4 FILLER_73_211 ();
 FILLCELL_X2 FILLER_73_215 ();
 FILLCELL_X8 FILLER_73_226 ();
 FILLCELL_X2 FILLER_73_234 ();
 FILLCELL_X8 FILLER_73_240 ();
 FILLCELL_X2 FILLER_73_248 ();
 FILLCELL_X1 FILLER_73_250 ();
 FILLCELL_X4 FILLER_73_255 ();
 FILLCELL_X2 FILLER_73_259 ();
 FILLCELL_X1 FILLER_73_261 ();
 FILLCELL_X4 FILLER_73_267 ();
 FILLCELL_X8 FILLER_73_274 ();
 FILLCELL_X4 FILLER_73_286 ();
 FILLCELL_X4 FILLER_73_299 ();
 FILLCELL_X4 FILLER_73_312 ();
 FILLCELL_X4 FILLER_73_325 ();
 FILLCELL_X4 FILLER_73_333 ();
 FILLCELL_X4 FILLER_73_340 ();
 FILLCELL_X8 FILLER_73_348 ();
 FILLCELL_X1 FILLER_73_356 ();
 FILLCELL_X4 FILLER_73_376 ();
 FILLCELL_X32 FILLER_73_1518 ();
 FILLCELL_X32 FILLER_73_1550 ();
 FILLCELL_X32 FILLER_73_1582 ();
 FILLCELL_X32 FILLER_73_1614 ();
 FILLCELL_X32 FILLER_73_1646 ();
 FILLCELL_X32 FILLER_73_1678 ();
 FILLCELL_X32 FILLER_73_1710 ();
 FILLCELL_X8 FILLER_73_1742 ();
 FILLCELL_X4 FILLER_73_1750 ();
 FILLCELL_X2 FILLER_73_1754 ();
 FILLCELL_X4 FILLER_74_1 ();
 FILLCELL_X4 FILLER_74_24 ();
 FILLCELL_X1 FILLER_74_28 ();
 FILLCELL_X4 FILLER_74_32 ();
 FILLCELL_X4 FILLER_74_45 ();
 FILLCELL_X4 FILLER_74_54 ();
 FILLCELL_X2 FILLER_74_58 ();
 FILLCELL_X1 FILLER_74_60 ();
 FILLCELL_X16 FILLER_74_64 ();
 FILLCELL_X8 FILLER_74_80 ();
 FILLCELL_X4 FILLER_74_88 ();
 FILLCELL_X2 FILLER_74_92 ();
 FILLCELL_X8 FILLER_74_98 ();
 FILLCELL_X4 FILLER_74_106 ();
 FILLCELL_X2 FILLER_74_110 ();
 FILLCELL_X4 FILLER_74_116 ();
 FILLCELL_X2 FILLER_74_120 ();
 FILLCELL_X1 FILLER_74_122 ();
 FILLCELL_X8 FILLER_74_127 ();
 FILLCELL_X4 FILLER_74_135 ();
 FILLCELL_X1 FILLER_74_139 ();
 FILLCELL_X8 FILLER_74_144 ();
 FILLCELL_X4 FILLER_74_152 ();
 FILLCELL_X2 FILLER_74_156 ();
 FILLCELL_X1 FILLER_74_158 ();
 FILLCELL_X4 FILLER_74_163 ();
 FILLCELL_X4 FILLER_74_171 ();
 FILLCELL_X4 FILLER_74_179 ();
 FILLCELL_X4 FILLER_74_192 ();
 FILLCELL_X4 FILLER_74_202 ();
 FILLCELL_X2 FILLER_74_206 ();
 FILLCELL_X1 FILLER_74_208 ();
 FILLCELL_X4 FILLER_74_213 ();
 FILLCELL_X4 FILLER_74_226 ();
 FILLCELL_X4 FILLER_74_239 ();
 FILLCELL_X4 FILLER_74_249 ();
 FILLCELL_X32 FILLER_74_257 ();
 FILLCELL_X8 FILLER_74_289 ();
 FILLCELL_X2 FILLER_74_297 ();
 FILLCELL_X16 FILLER_74_304 ();
 FILLCELL_X4 FILLER_74_320 ();
 FILLCELL_X1 FILLER_74_324 ();
 FILLCELL_X4 FILLER_74_329 ();
 FILLCELL_X2 FILLER_74_333 ();
 FILLCELL_X1 FILLER_74_335 ();
 FILLCELL_X4 FILLER_74_342 ();
 FILLCELL_X4 FILLER_74_355 ();
 FILLCELL_X16 FILLER_74_362 ();
 FILLCELL_X2 FILLER_74_378 ();
 FILLCELL_X8 FILLER_74_1518 ();
 FILLCELL_X32 FILLER_74_1530 ();
 FILLCELL_X32 FILLER_74_1562 ();
 FILLCELL_X32 FILLER_74_1594 ();
 FILLCELL_X32 FILLER_74_1626 ();
 FILLCELL_X32 FILLER_74_1658 ();
 FILLCELL_X32 FILLER_74_1690 ();
 FILLCELL_X32 FILLER_74_1722 ();
 FILLCELL_X2 FILLER_74_1754 ();
 FILLCELL_X8 FILLER_75_1 ();
 FILLCELL_X1 FILLER_75_9 ();
 FILLCELL_X4 FILLER_75_16 ();
 FILLCELL_X8 FILLER_75_27 ();
 FILLCELL_X4 FILLER_75_35 ();
 FILLCELL_X1 FILLER_75_39 ();
 FILLCELL_X4 FILLER_75_44 ();
 FILLCELL_X4 FILLER_75_53 ();
 FILLCELL_X4 FILLER_75_60 ();
 FILLCELL_X2 FILLER_75_64 ();
 FILLCELL_X4 FILLER_75_72 ();
 FILLCELL_X4 FILLER_75_81 ();
 FILLCELL_X1 FILLER_75_85 ();
 FILLCELL_X4 FILLER_75_89 ();
 FILLCELL_X4 FILLER_75_99 ();
 FILLCELL_X4 FILLER_75_108 ();
 FILLCELL_X16 FILLER_75_116 ();
 FILLCELL_X1 FILLER_75_132 ();
 FILLCELL_X4 FILLER_75_142 ();
 FILLCELL_X4 FILLER_75_155 ();
 FILLCELL_X4 FILLER_75_163 ();
 FILLCELL_X2 FILLER_75_167 ();
 FILLCELL_X4 FILLER_75_173 ();
 FILLCELL_X2 FILLER_75_177 ();
 FILLCELL_X4 FILLER_75_188 ();
 FILLCELL_X2 FILLER_75_192 ();
 FILLCELL_X1 FILLER_75_194 ();
 FILLCELL_X4 FILLER_75_200 ();
 FILLCELL_X4 FILLER_75_209 ();
 FILLCELL_X8 FILLER_75_217 ();
 FILLCELL_X2 FILLER_75_225 ();
 FILLCELL_X8 FILLER_75_232 ();
 FILLCELL_X1 FILLER_75_240 ();
 FILLCELL_X8 FILLER_75_246 ();
 FILLCELL_X1 FILLER_75_254 ();
 FILLCELL_X4 FILLER_75_264 ();
 FILLCELL_X4 FILLER_75_274 ();
 FILLCELL_X4 FILLER_75_283 ();
 FILLCELL_X2 FILLER_75_287 ();
 FILLCELL_X1 FILLER_75_289 ();
 FILLCELL_X4 FILLER_75_294 ();
 FILLCELL_X2 FILLER_75_298 ();
 FILLCELL_X4 FILLER_75_303 ();
 FILLCELL_X4 FILLER_75_310 ();
 FILLCELL_X4 FILLER_75_317 ();
 FILLCELL_X2 FILLER_75_321 ();
 FILLCELL_X8 FILLER_75_326 ();
 FILLCELL_X4 FILLER_75_334 ();
 FILLCELL_X4 FILLER_75_347 ();
 FILLCELL_X8 FILLER_75_356 ();
 FILLCELL_X8 FILLER_75_367 ();
 FILLCELL_X4 FILLER_75_375 ();
 FILLCELL_X1 FILLER_75_379 ();
 FILLCELL_X4 FILLER_75_1518 ();
 FILLCELL_X1 FILLER_75_1522 ();
 FILLCELL_X32 FILLER_75_1542 ();
 FILLCELL_X32 FILLER_75_1574 ();
 FILLCELL_X32 FILLER_75_1606 ();
 FILLCELL_X32 FILLER_75_1638 ();
 FILLCELL_X32 FILLER_75_1670 ();
 FILLCELL_X32 FILLER_75_1702 ();
 FILLCELL_X16 FILLER_75_1734 ();
 FILLCELL_X4 FILLER_75_1750 ();
 FILLCELL_X2 FILLER_75_1754 ();
 FILLCELL_X8 FILLER_76_1 ();
 FILLCELL_X2 FILLER_76_9 ();
 FILLCELL_X1 FILLER_76_11 ();
 FILLCELL_X8 FILLER_76_18 ();
 FILLCELL_X8 FILLER_76_30 ();
 FILLCELL_X2 FILLER_76_38 ();
 FILLCELL_X4 FILLER_76_46 ();
 FILLCELL_X1 FILLER_76_50 ();
 FILLCELL_X4 FILLER_76_54 ();
 FILLCELL_X4 FILLER_76_67 ();
 FILLCELL_X4 FILLER_76_80 ();
 FILLCELL_X2 FILLER_76_84 ();
 FILLCELL_X1 FILLER_76_86 ();
 FILLCELL_X4 FILLER_76_96 ();
 FILLCELL_X4 FILLER_76_109 ();
 FILLCELL_X4 FILLER_76_122 ();
 FILLCELL_X4 FILLER_76_131 ();
 FILLCELL_X4 FILLER_76_141 ();
 FILLCELL_X2 FILLER_76_145 ();
 FILLCELL_X8 FILLER_76_156 ();
 FILLCELL_X4 FILLER_76_164 ();
 FILLCELL_X1 FILLER_76_168 ();
 FILLCELL_X4 FILLER_76_173 ();
 FILLCELL_X2 FILLER_76_177 ();
 FILLCELL_X16 FILLER_76_188 ();
 FILLCELL_X8 FILLER_76_204 ();
 FILLCELL_X4 FILLER_76_212 ();
 FILLCELL_X1 FILLER_76_216 ();
 FILLCELL_X4 FILLER_76_226 ();
 FILLCELL_X1 FILLER_76_230 ();
 FILLCELL_X4 FILLER_76_237 ();
 FILLCELL_X4 FILLER_76_246 ();
 FILLCELL_X4 FILLER_76_253 ();
 FILLCELL_X8 FILLER_76_266 ();
 FILLCELL_X4 FILLER_76_283 ();
 FILLCELL_X4 FILLER_76_296 ();
 FILLCELL_X8 FILLER_76_306 ();
 FILLCELL_X1 FILLER_76_314 ();
 FILLCELL_X4 FILLER_76_321 ();
 FILLCELL_X4 FILLER_76_329 ();
 FILLCELL_X16 FILLER_76_336 ();
 FILLCELL_X1 FILLER_76_352 ();
 FILLCELL_X4 FILLER_76_356 ();
 FILLCELL_X4 FILLER_76_366 ();
 FILLCELL_X4 FILLER_76_375 ();
 FILLCELL_X1 FILLER_76_379 ();
 FILLCELL_X32 FILLER_76_1518 ();
 FILLCELL_X32 FILLER_76_1550 ();
 FILLCELL_X32 FILLER_76_1582 ();
 FILLCELL_X32 FILLER_76_1614 ();
 FILLCELL_X32 FILLER_76_1646 ();
 FILLCELL_X32 FILLER_76_1678 ();
 FILLCELL_X32 FILLER_76_1710 ();
 FILLCELL_X8 FILLER_76_1742 ();
 FILLCELL_X4 FILLER_76_1750 ();
 FILLCELL_X2 FILLER_76_1754 ();
 FILLCELL_X16 FILLER_77_1 ();
 FILLCELL_X2 FILLER_77_17 ();
 FILLCELL_X4 FILLER_77_23 ();
 FILLCELL_X4 FILLER_77_36 ();
 FILLCELL_X4 FILLER_77_49 ();
 FILLCELL_X8 FILLER_77_57 ();
 FILLCELL_X4 FILLER_77_70 ();
 FILLCELL_X16 FILLER_77_78 ();
 FILLCELL_X1 FILLER_77_94 ();
 FILLCELL_X8 FILLER_77_99 ();
 FILLCELL_X2 FILLER_77_107 ();
 FILLCELL_X4 FILLER_77_113 ();
 FILLCELL_X2 FILLER_77_117 ();
 FILLCELL_X4 FILLER_77_124 ();
 FILLCELL_X2 FILLER_77_128 ();
 FILLCELL_X4 FILLER_77_133 ();
 FILLCELL_X8 FILLER_77_142 ();
 FILLCELL_X2 FILLER_77_150 ();
 FILLCELL_X1 FILLER_77_152 ();
 FILLCELL_X4 FILLER_77_157 ();
 FILLCELL_X8 FILLER_77_165 ();
 FILLCELL_X2 FILLER_77_173 ();
 FILLCELL_X1 FILLER_77_175 ();
 FILLCELL_X16 FILLER_77_180 ();
 FILLCELL_X2 FILLER_77_196 ();
 FILLCELL_X4 FILLER_77_202 ();
 FILLCELL_X2 FILLER_77_206 ();
 FILLCELL_X4 FILLER_77_213 ();
 FILLCELL_X4 FILLER_77_226 ();
 FILLCELL_X4 FILLER_77_239 ();
 FILLCELL_X4 FILLER_77_248 ();
 FILLCELL_X2 FILLER_77_252 ();
 FILLCELL_X4 FILLER_77_263 ();
 FILLCELL_X2 FILLER_77_267 ();
 FILLCELL_X4 FILLER_77_274 ();
 FILLCELL_X8 FILLER_77_281 ();
 FILLCELL_X4 FILLER_77_298 ();
 FILLCELL_X2 FILLER_77_302 ();
 FILLCELL_X1 FILLER_77_304 ();
 FILLCELL_X4 FILLER_77_309 ();
 FILLCELL_X4 FILLER_77_322 ();
 FILLCELL_X8 FILLER_77_335 ();
 FILLCELL_X2 FILLER_77_343 ();
 FILLCELL_X1 FILLER_77_345 ();
 FILLCELL_X4 FILLER_77_350 ();
 FILLCELL_X4 FILLER_77_363 ();
 FILLCELL_X4 FILLER_77_376 ();
 FILLCELL_X32 FILLER_77_1518 ();
 FILLCELL_X32 FILLER_77_1550 ();
 FILLCELL_X32 FILLER_77_1582 ();
 FILLCELL_X32 FILLER_77_1614 ();
 FILLCELL_X32 FILLER_77_1646 ();
 FILLCELL_X32 FILLER_77_1678 ();
 FILLCELL_X32 FILLER_77_1710 ();
 FILLCELL_X8 FILLER_77_1742 ();
 FILLCELL_X4 FILLER_77_1750 ();
 FILLCELL_X2 FILLER_77_1754 ();
 FILLCELL_X8 FILLER_78_1 ();
 FILLCELL_X16 FILLER_78_13 ();
 FILLCELL_X8 FILLER_78_29 ();
 FILLCELL_X2 FILLER_78_37 ();
 FILLCELL_X4 FILLER_78_48 ();
 FILLCELL_X2 FILLER_78_52 ();
 FILLCELL_X4 FILLER_78_57 ();
 FILLCELL_X16 FILLER_78_64 ();
 FILLCELL_X8 FILLER_78_80 ();
 FILLCELL_X8 FILLER_78_92 ();
 FILLCELL_X1 FILLER_78_100 ();
 FILLCELL_X8 FILLER_78_104 ();
 FILLCELL_X4 FILLER_78_115 ();
 FILLCELL_X16 FILLER_78_128 ();
 FILLCELL_X2 FILLER_78_144 ();
 FILLCELL_X1 FILLER_78_146 ();
 FILLCELL_X8 FILLER_78_151 ();
 FILLCELL_X4 FILLER_78_159 ();
 FILLCELL_X2 FILLER_78_163 ();
 FILLCELL_X4 FILLER_78_169 ();
 FILLCELL_X4 FILLER_78_182 ();
 FILLCELL_X4 FILLER_78_195 ();
 FILLCELL_X4 FILLER_78_208 ();
 FILLCELL_X8 FILLER_78_218 ();
 FILLCELL_X4 FILLER_78_229 ();
 FILLCELL_X4 FILLER_78_238 ();
 FILLCELL_X8 FILLER_78_246 ();
 FILLCELL_X4 FILLER_78_260 ();
 FILLCELL_X4 FILLER_78_267 ();
 FILLCELL_X2 FILLER_78_271 ();
 FILLCELL_X16 FILLER_78_277 ();
 FILLCELL_X2 FILLER_78_293 ();
 FILLCELL_X8 FILLER_78_300 ();
 FILLCELL_X2 FILLER_78_308 ();
 FILLCELL_X4 FILLER_78_314 ();
 FILLCELL_X32 FILLER_78_323 ();
 FILLCELL_X4 FILLER_78_355 ();
 FILLCELL_X1 FILLER_78_359 ();
 FILLCELL_X8 FILLER_78_369 ();
 FILLCELL_X2 FILLER_78_377 ();
 FILLCELL_X1 FILLER_78_379 ();
 FILLCELL_X32 FILLER_78_1518 ();
 FILLCELL_X32 FILLER_78_1550 ();
 FILLCELL_X32 FILLER_78_1582 ();
 FILLCELL_X32 FILLER_78_1614 ();
 FILLCELL_X32 FILLER_78_1646 ();
 FILLCELL_X32 FILLER_78_1678 ();
 FILLCELL_X32 FILLER_78_1710 ();
 FILLCELL_X4 FILLER_78_1742 ();
 FILLCELL_X2 FILLER_78_1746 ();
 FILLCELL_X1 FILLER_78_1748 ();
 FILLCELL_X4 FILLER_78_1752 ();
 FILLCELL_X4 FILLER_79_1 ();
 FILLCELL_X8 FILLER_79_24 ();
 FILLCELL_X4 FILLER_79_32 ();
 FILLCELL_X2 FILLER_79_36 ();
 FILLCELL_X4 FILLER_79_42 ();
 FILLCELL_X4 FILLER_79_51 ();
 FILLCELL_X2 FILLER_79_55 ();
 FILLCELL_X4 FILLER_79_60 ();
 FILLCELL_X4 FILLER_79_73 ();
 FILLCELL_X4 FILLER_79_81 ();
 FILLCELL_X1 FILLER_79_85 ();
 FILLCELL_X16 FILLER_79_105 ();
 FILLCELL_X1 FILLER_79_121 ();
 FILLCELL_X4 FILLER_79_131 ();
 FILLCELL_X8 FILLER_79_139 ();
 FILLCELL_X1 FILLER_79_147 ();
 FILLCELL_X4 FILLER_79_152 ();
 FILLCELL_X8 FILLER_79_160 ();
 FILLCELL_X1 FILLER_79_168 ();
 FILLCELL_X4 FILLER_79_173 ();
 FILLCELL_X8 FILLER_79_181 ();
 FILLCELL_X4 FILLER_79_189 ();
 FILLCELL_X2 FILLER_79_193 ();
 FILLCELL_X1 FILLER_79_195 ();
 FILLCELL_X4 FILLER_79_200 ();
 FILLCELL_X8 FILLER_79_209 ();
 FILLCELL_X1 FILLER_79_217 ();
 FILLCELL_X16 FILLER_79_221 ();
 FILLCELL_X2 FILLER_79_237 ();
 FILLCELL_X1 FILLER_79_239 ();
 FILLCELL_X4 FILLER_79_245 ();
 FILLCELL_X4 FILLER_79_258 ();
 FILLCELL_X8 FILLER_79_271 ();
 FILLCELL_X4 FILLER_79_283 ();
 FILLCELL_X4 FILLER_79_291 ();
 FILLCELL_X8 FILLER_79_299 ();
 FILLCELL_X4 FILLER_79_307 ();
 FILLCELL_X4 FILLER_79_315 ();
 FILLCELL_X8 FILLER_79_323 ();
 FILLCELL_X2 FILLER_79_331 ();
 FILLCELL_X4 FILLER_79_337 ();
 FILLCELL_X4 FILLER_79_345 ();
 FILLCELL_X4 FILLER_79_353 ();
 FILLCELL_X4 FILLER_79_361 ();
 FILLCELL_X8 FILLER_79_369 ();
 FILLCELL_X2 FILLER_79_377 ();
 FILLCELL_X1 FILLER_79_379 ();
 FILLCELL_X32 FILLER_79_1518 ();
 FILLCELL_X32 FILLER_79_1550 ();
 FILLCELL_X32 FILLER_79_1582 ();
 FILLCELL_X32 FILLER_79_1614 ();
 FILLCELL_X32 FILLER_79_1646 ();
 FILLCELL_X32 FILLER_79_1678 ();
 FILLCELL_X32 FILLER_79_1710 ();
 FILLCELL_X8 FILLER_79_1742 ();
 FILLCELL_X4 FILLER_79_1750 ();
 FILLCELL_X2 FILLER_79_1754 ();
 FILLCELL_X8 FILLER_80_1 ();
 FILLCELL_X4 FILLER_80_9 ();
 FILLCELL_X2 FILLER_80_13 ();
 FILLCELL_X1 FILLER_80_15 ();
 FILLCELL_X8 FILLER_80_20 ();
 FILLCELL_X4 FILLER_80_31 ();
 FILLCELL_X8 FILLER_80_44 ();
 FILLCELL_X2 FILLER_80_52 ();
 FILLCELL_X4 FILLER_80_60 ();
 FILLCELL_X4 FILLER_80_73 ();
 FILLCELL_X4 FILLER_80_82 ();
 FILLCELL_X2 FILLER_80_86 ();
 FILLCELL_X4 FILLER_80_92 ();
 FILLCELL_X4 FILLER_80_100 ();
 FILLCELL_X4 FILLER_80_110 ();
 FILLCELL_X4 FILLER_80_123 ();
 FILLCELL_X2 FILLER_80_127 ();
 FILLCELL_X1 FILLER_80_129 ();
 FILLCELL_X4 FILLER_80_134 ();
 FILLCELL_X4 FILLER_80_142 ();
 FILLCELL_X4 FILLER_80_155 ();
 FILLCELL_X4 FILLER_80_163 ();
 FILLCELL_X2 FILLER_80_167 ();
 FILLCELL_X4 FILLER_80_173 ();
 FILLCELL_X4 FILLER_80_181 ();
 FILLCELL_X8 FILLER_80_189 ();
 FILLCELL_X4 FILLER_80_197 ();
 FILLCELL_X4 FILLER_80_205 ();
 FILLCELL_X16 FILLER_80_213 ();
 FILLCELL_X1 FILLER_80_229 ();
 FILLCELL_X4 FILLER_80_234 ();
 FILLCELL_X4 FILLER_80_242 ();
 FILLCELL_X4 FILLER_80_250 ();
 FILLCELL_X8 FILLER_80_257 ();
 FILLCELL_X2 FILLER_80_265 ();
 FILLCELL_X4 FILLER_80_276 ();
 FILLCELL_X1 FILLER_80_280 ();
 FILLCELL_X8 FILLER_80_286 ();
 FILLCELL_X2 FILLER_80_294 ();
 FILLCELL_X4 FILLER_80_300 ();
 FILLCELL_X8 FILLER_80_308 ();
 FILLCELL_X4 FILLER_80_316 ();
 FILLCELL_X4 FILLER_80_324 ();
 FILLCELL_X4 FILLER_80_333 ();
 FILLCELL_X8 FILLER_80_346 ();
 FILLCELL_X4 FILLER_80_354 ();
 FILLCELL_X1 FILLER_80_358 ();
 FILLCELL_X16 FILLER_80_363 ();
 FILLCELL_X1 FILLER_80_379 ();
 FILLCELL_X32 FILLER_80_1518 ();
 FILLCELL_X32 FILLER_80_1550 ();
 FILLCELL_X32 FILLER_80_1582 ();
 FILLCELL_X32 FILLER_80_1614 ();
 FILLCELL_X32 FILLER_80_1646 ();
 FILLCELL_X32 FILLER_80_1678 ();
 FILLCELL_X32 FILLER_80_1710 ();
 FILLCELL_X8 FILLER_80_1742 ();
 FILLCELL_X4 FILLER_80_1750 ();
 FILLCELL_X2 FILLER_80_1754 ();
 FILLCELL_X4 FILLER_81_1 ();
 FILLCELL_X2 FILLER_81_5 ();
 FILLCELL_X1 FILLER_81_7 ();
 FILLCELL_X4 FILLER_81_12 ();
 FILLCELL_X2 FILLER_81_16 ();
 FILLCELL_X4 FILLER_81_27 ();
 FILLCELL_X4 FILLER_81_40 ();
 FILLCELL_X4 FILLER_81_50 ();
 FILLCELL_X2 FILLER_81_54 ();
 FILLCELL_X1 FILLER_81_56 ();
 FILLCELL_X4 FILLER_81_61 ();
 FILLCELL_X8 FILLER_81_70 ();
 FILLCELL_X4 FILLER_81_82 ();
 FILLCELL_X16 FILLER_81_90 ();
 FILLCELL_X1 FILLER_81_106 ();
 FILLCELL_X8 FILLER_81_112 ();
 FILLCELL_X1 FILLER_81_120 ();
 FILLCELL_X4 FILLER_81_125 ();
 FILLCELL_X4 FILLER_81_133 ();
 FILLCELL_X4 FILLER_81_141 ();
 FILLCELL_X2 FILLER_81_145 ();
 FILLCELL_X16 FILLER_81_156 ();
 FILLCELL_X1 FILLER_81_172 ();
 FILLCELL_X4 FILLER_81_182 ();
 FILLCELL_X1 FILLER_81_186 ();
 FILLCELL_X4 FILLER_81_191 ();
 FILLCELL_X8 FILLER_81_199 ();
 FILLCELL_X8 FILLER_81_211 ();
 FILLCELL_X4 FILLER_81_223 ();
 FILLCELL_X4 FILLER_81_236 ();
 FILLCELL_X1 FILLER_81_240 ();
 FILLCELL_X8 FILLER_81_245 ();
 FILLCELL_X1 FILLER_81_253 ();
 FILLCELL_X16 FILLER_81_258 ();
 FILLCELL_X1 FILLER_81_274 ();
 FILLCELL_X4 FILLER_81_279 ();
 FILLCELL_X8 FILLER_81_292 ();
 FILLCELL_X4 FILLER_81_304 ();
 FILLCELL_X4 FILLER_81_312 ();
 FILLCELL_X4 FILLER_81_325 ();
 FILLCELL_X4 FILLER_81_338 ();
 FILLCELL_X32 FILLER_81_348 ();
 FILLCELL_X32 FILLER_81_1518 ();
 FILLCELL_X32 FILLER_81_1550 ();
 FILLCELL_X32 FILLER_81_1582 ();
 FILLCELL_X32 FILLER_81_1614 ();
 FILLCELL_X32 FILLER_81_1646 ();
 FILLCELL_X32 FILLER_81_1678 ();
 FILLCELL_X32 FILLER_81_1710 ();
 FILLCELL_X8 FILLER_81_1742 ();
 FILLCELL_X4 FILLER_81_1750 ();
 FILLCELL_X2 FILLER_81_1754 ();
 FILLCELL_X4 FILLER_82_1 ();
 FILLCELL_X4 FILLER_82_8 ();
 FILLCELL_X4 FILLER_82_16 ();
 FILLCELL_X4 FILLER_82_24 ();
 FILLCELL_X2 FILLER_82_28 ();
 FILLCELL_X4 FILLER_82_34 ();
 FILLCELL_X2 FILLER_82_38 ();
 FILLCELL_X16 FILLER_82_43 ();
 FILLCELL_X4 FILLER_82_59 ();
 FILLCELL_X4 FILLER_82_68 ();
 FILLCELL_X8 FILLER_82_76 ();
 FILLCELL_X2 FILLER_82_84 ();
 FILLCELL_X4 FILLER_82_90 ();
 FILLCELL_X2 FILLER_82_94 ();
 FILLCELL_X1 FILLER_82_96 ();
 FILLCELL_X4 FILLER_82_101 ();
 FILLCELL_X4 FILLER_82_109 ();
 FILLCELL_X8 FILLER_82_117 ();
 FILLCELL_X2 FILLER_82_125 ();
 FILLCELL_X4 FILLER_82_131 ();
 FILLCELL_X2 FILLER_82_135 ();
 FILLCELL_X1 FILLER_82_137 ();
 FILLCELL_X4 FILLER_82_142 ();
 FILLCELL_X16 FILLER_82_155 ();
 FILLCELL_X2 FILLER_82_171 ();
 FILLCELL_X1 FILLER_82_173 ();
 FILLCELL_X8 FILLER_82_183 ();
 FILLCELL_X2 FILLER_82_191 ();
 FILLCELL_X4 FILLER_82_197 ();
 FILLCELL_X8 FILLER_82_210 ();
 FILLCELL_X4 FILLER_82_218 ();
 FILLCELL_X1 FILLER_82_222 ();
 FILLCELL_X4 FILLER_82_226 ();
 FILLCELL_X8 FILLER_82_239 ();
 FILLCELL_X4 FILLER_82_251 ();
 FILLCELL_X4 FILLER_82_259 ();
 FILLCELL_X16 FILLER_82_267 ();
 FILLCELL_X2 FILLER_82_283 ();
 FILLCELL_X8 FILLER_82_294 ();
 FILLCELL_X2 FILLER_82_302 ();
 FILLCELL_X4 FILLER_82_308 ();
 FILLCELL_X8 FILLER_82_316 ();
 FILLCELL_X4 FILLER_82_324 ();
 FILLCELL_X2 FILLER_82_328 ();
 FILLCELL_X4 FILLER_82_334 ();
 FILLCELL_X4 FILLER_82_342 ();
 FILLCELL_X4 FILLER_82_350 ();
 FILLCELL_X4 FILLER_82_358 ();
 FILLCELL_X8 FILLER_82_366 ();
 FILLCELL_X4 FILLER_82_374 ();
 FILLCELL_X2 FILLER_82_378 ();
 FILLCELL_X32 FILLER_82_1518 ();
 FILLCELL_X32 FILLER_82_1550 ();
 FILLCELL_X32 FILLER_82_1582 ();
 FILLCELL_X32 FILLER_82_1614 ();
 FILLCELL_X32 FILLER_82_1646 ();
 FILLCELL_X32 FILLER_82_1678 ();
 FILLCELL_X32 FILLER_82_1710 ();
 FILLCELL_X8 FILLER_82_1742 ();
 FILLCELL_X4 FILLER_82_1750 ();
 FILLCELL_X2 FILLER_82_1754 ();
 FILLCELL_X4 FILLER_83_1 ();
 FILLCELL_X8 FILLER_83_22 ();
 FILLCELL_X2 FILLER_83_30 ();
 FILLCELL_X4 FILLER_83_36 ();
 FILLCELL_X4 FILLER_83_49 ();
 FILLCELL_X4 FILLER_83_62 ();
 FILLCELL_X8 FILLER_83_75 ();
 FILLCELL_X1 FILLER_83_83 ();
 FILLCELL_X8 FILLER_83_103 ();
 FILLCELL_X2 FILLER_83_111 ();
 FILLCELL_X16 FILLER_83_119 ();
 FILLCELL_X2 FILLER_83_135 ();
 FILLCELL_X4 FILLER_83_140 ();
 FILLCELL_X4 FILLER_83_150 ();
 FILLCELL_X4 FILLER_83_159 ();
 FILLCELL_X1 FILLER_83_163 ();
 FILLCELL_X4 FILLER_83_169 ();
 FILLCELL_X4 FILLER_83_182 ();
 FILLCELL_X8 FILLER_83_192 ();
 FILLCELL_X2 FILLER_83_200 ();
 FILLCELL_X8 FILLER_83_211 ();
 FILLCELL_X1 FILLER_83_219 ();
 FILLCELL_X4 FILLER_83_224 ();
 FILLCELL_X4 FILLER_83_237 ();
 FILLCELL_X2 FILLER_83_241 ();
 FILLCELL_X1 FILLER_83_243 ();
 FILLCELL_X4 FILLER_83_247 ();
 FILLCELL_X2 FILLER_83_251 ();
 FILLCELL_X1 FILLER_83_253 ();
 FILLCELL_X4 FILLER_83_263 ();
 FILLCELL_X2 FILLER_83_267 ();
 FILLCELL_X1 FILLER_83_269 ();
 FILLCELL_X4 FILLER_83_276 ();
 FILLCELL_X4 FILLER_83_289 ();
 FILLCELL_X8 FILLER_83_296 ();
 FILLCELL_X2 FILLER_83_304 ();
 FILLCELL_X8 FILLER_83_315 ();
 FILLCELL_X4 FILLER_83_323 ();
 FILLCELL_X2 FILLER_83_327 ();
 FILLCELL_X4 FILLER_83_334 ();
 FILLCELL_X1 FILLER_83_338 ();
 FILLCELL_X32 FILLER_83_342 ();
 FILLCELL_X4 FILLER_83_374 ();
 FILLCELL_X2 FILLER_83_378 ();
 FILLCELL_X32 FILLER_83_1518 ();
 FILLCELL_X32 FILLER_83_1550 ();
 FILLCELL_X32 FILLER_83_1582 ();
 FILLCELL_X32 FILLER_83_1614 ();
 FILLCELL_X32 FILLER_83_1646 ();
 FILLCELL_X32 FILLER_83_1678 ();
 FILLCELL_X32 FILLER_83_1710 ();
 FILLCELL_X8 FILLER_83_1742 ();
 FILLCELL_X4 FILLER_83_1750 ();
 FILLCELL_X2 FILLER_83_1754 ();
 FILLCELL_X16 FILLER_84_1 ();
 FILLCELL_X8 FILLER_84_17 ();
 FILLCELL_X4 FILLER_84_25 ();
 FILLCELL_X4 FILLER_84_33 ();
 FILLCELL_X4 FILLER_84_46 ();
 FILLCELL_X4 FILLER_84_55 ();
 FILLCELL_X2 FILLER_84_59 ();
 FILLCELL_X1 FILLER_84_61 ();
 FILLCELL_X8 FILLER_84_68 ();
 FILLCELL_X16 FILLER_84_80 ();
 FILLCELL_X4 FILLER_84_96 ();
 FILLCELL_X2 FILLER_84_100 ();
 FILLCELL_X8 FILLER_84_111 ();
 FILLCELL_X4 FILLER_84_128 ();
 FILLCELL_X4 FILLER_84_136 ();
 FILLCELL_X2 FILLER_84_140 ();
 FILLCELL_X16 FILLER_84_147 ();
 FILLCELL_X8 FILLER_84_163 ();
 FILLCELL_X2 FILLER_84_171 ();
 FILLCELL_X1 FILLER_84_173 ();
 FILLCELL_X4 FILLER_84_177 ();
 FILLCELL_X1 FILLER_84_181 ();
 FILLCELL_X8 FILLER_84_187 ();
 FILLCELL_X4 FILLER_84_195 ();
 FILLCELL_X2 FILLER_84_199 ();
 FILLCELL_X8 FILLER_84_210 ();
 FILLCELL_X2 FILLER_84_218 ();
 FILLCELL_X1 FILLER_84_220 ();
 FILLCELL_X4 FILLER_84_226 ();
 FILLCELL_X4 FILLER_84_236 ();
 FILLCELL_X8 FILLER_84_245 ();
 FILLCELL_X2 FILLER_84_253 ();
 FILLCELL_X4 FILLER_84_264 ();
 FILLCELL_X8 FILLER_84_272 ();
 FILLCELL_X4 FILLER_84_280 ();
 FILLCELL_X2 FILLER_84_284 ();
 FILLCELL_X1 FILLER_84_286 ();
 FILLCELL_X4 FILLER_84_292 ();
 FILLCELL_X4 FILLER_84_305 ();
 FILLCELL_X4 FILLER_84_318 ();
 FILLCELL_X8 FILLER_84_326 ();
 FILLCELL_X4 FILLER_84_343 ();
 FILLCELL_X4 FILLER_84_356 ();
 FILLCELL_X16 FILLER_84_364 ();
 FILLCELL_X32 FILLER_84_1518 ();
 FILLCELL_X32 FILLER_84_1550 ();
 FILLCELL_X32 FILLER_84_1582 ();
 FILLCELL_X32 FILLER_84_1614 ();
 FILLCELL_X32 FILLER_84_1646 ();
 FILLCELL_X32 FILLER_84_1678 ();
 FILLCELL_X32 FILLER_84_1710 ();
 FILLCELL_X8 FILLER_84_1742 ();
 FILLCELL_X4 FILLER_84_1750 ();
 FILLCELL_X2 FILLER_84_1754 ();
 FILLCELL_X8 FILLER_85_1 ();
 FILLCELL_X2 FILLER_85_9 ();
 FILLCELL_X1 FILLER_85_11 ();
 FILLCELL_X4 FILLER_85_16 ();
 FILLCELL_X2 FILLER_85_20 ();
 FILLCELL_X4 FILLER_85_25 ();
 FILLCELL_X4 FILLER_85_33 ();
 FILLCELL_X16 FILLER_85_41 ();
 FILLCELL_X8 FILLER_85_60 ();
 FILLCELL_X2 FILLER_85_68 ();
 FILLCELL_X8 FILLER_85_73 ();
 FILLCELL_X2 FILLER_85_81 ();
 FILLCELL_X1 FILLER_85_83 ();
 FILLCELL_X8 FILLER_85_88 ();
 FILLCELL_X4 FILLER_85_99 ();
 FILLCELL_X4 FILLER_85_106 ();
 FILLCELL_X4 FILLER_85_115 ();
 FILLCELL_X2 FILLER_85_119 ();
 FILLCELL_X8 FILLER_85_126 ();
 FILLCELL_X2 FILLER_85_134 ();
 FILLCELL_X4 FILLER_85_140 ();
 FILLCELL_X4 FILLER_85_153 ();
 FILLCELL_X8 FILLER_85_160 ();
 FILLCELL_X2 FILLER_85_168 ();
 FILLCELL_X4 FILLER_85_174 ();
 FILLCELL_X8 FILLER_85_182 ();
 FILLCELL_X2 FILLER_85_190 ();
 FILLCELL_X4 FILLER_85_197 ();
 FILLCELL_X4 FILLER_85_207 ();
 FILLCELL_X8 FILLER_85_216 ();
 FILLCELL_X2 FILLER_85_224 ();
 FILLCELL_X1 FILLER_85_226 ();
 FILLCELL_X4 FILLER_85_231 ();
 FILLCELL_X1 FILLER_85_235 ();
 FILLCELL_X4 FILLER_85_240 ();
 FILLCELL_X2 FILLER_85_244 ();
 FILLCELL_X1 FILLER_85_246 ();
 FILLCELL_X4 FILLER_85_253 ();
 FILLCELL_X8 FILLER_85_266 ();
 FILLCELL_X4 FILLER_85_274 ();
 FILLCELL_X2 FILLER_85_278 ();
 FILLCELL_X1 FILLER_85_280 ();
 FILLCELL_X8 FILLER_85_285 ();
 FILLCELL_X4 FILLER_85_293 ();
 FILLCELL_X2 FILLER_85_297 ();
 FILLCELL_X8 FILLER_85_304 ();
 FILLCELL_X4 FILLER_85_318 ();
 FILLCELL_X4 FILLER_85_327 ();
 FILLCELL_X2 FILLER_85_331 ();
 FILLCELL_X1 FILLER_85_333 ();
 FILLCELL_X4 FILLER_85_337 ();
 FILLCELL_X4 FILLER_85_347 ();
 FILLCELL_X1 FILLER_85_351 ();
 FILLCELL_X16 FILLER_85_361 ();
 FILLCELL_X2 FILLER_85_377 ();
 FILLCELL_X1 FILLER_85_379 ();
 FILLCELL_X32 FILLER_85_1518 ();
 FILLCELL_X32 FILLER_85_1550 ();
 FILLCELL_X32 FILLER_85_1582 ();
 FILLCELL_X32 FILLER_85_1614 ();
 FILLCELL_X32 FILLER_85_1646 ();
 FILLCELL_X32 FILLER_85_1678 ();
 FILLCELL_X32 FILLER_85_1710 ();
 FILLCELL_X8 FILLER_85_1742 ();
 FILLCELL_X4 FILLER_85_1750 ();
 FILLCELL_X2 FILLER_85_1754 ();
 FILLCELL_X8 FILLER_86_1 ();
 FILLCELL_X4 FILLER_86_13 ();
 FILLCELL_X1 FILLER_86_17 ();
 FILLCELL_X4 FILLER_86_27 ();
 FILLCELL_X1 FILLER_86_31 ();
 FILLCELL_X8 FILLER_86_37 ();
 FILLCELL_X2 FILLER_86_45 ();
 FILLCELL_X1 FILLER_86_47 ();
 FILLCELL_X4 FILLER_86_53 ();
 FILLCELL_X4 FILLER_86_61 ();
 FILLCELL_X4 FILLER_86_68 ();
 FILLCELL_X4 FILLER_86_76 ();
 FILLCELL_X4 FILLER_86_86 ();
 FILLCELL_X16 FILLER_86_94 ();
 FILLCELL_X8 FILLER_86_110 ();
 FILLCELL_X2 FILLER_86_118 ();
 FILLCELL_X1 FILLER_86_120 ();
 FILLCELL_X8 FILLER_86_130 ();
 FILLCELL_X4 FILLER_86_138 ();
 FILLCELL_X2 FILLER_86_142 ();
 FILLCELL_X4 FILLER_86_153 ();
 FILLCELL_X4 FILLER_86_166 ();
 FILLCELL_X2 FILLER_86_170 ();
 FILLCELL_X1 FILLER_86_172 ();
 FILLCELL_X4 FILLER_86_178 ();
 FILLCELL_X8 FILLER_86_186 ();
 FILLCELL_X2 FILLER_86_194 ();
 FILLCELL_X1 FILLER_86_196 ();
 FILLCELL_X4 FILLER_86_206 ();
 FILLCELL_X4 FILLER_86_213 ();
 FILLCELL_X4 FILLER_86_221 ();
 FILLCELL_X4 FILLER_86_234 ();
 FILLCELL_X4 FILLER_86_242 ();
 FILLCELL_X2 FILLER_86_246 ();
 FILLCELL_X1 FILLER_86_248 ();
 FILLCELL_X4 FILLER_86_254 ();
 FILLCELL_X2 FILLER_86_258 ();
 FILLCELL_X4 FILLER_86_265 ();
 FILLCELL_X1 FILLER_86_269 ();
 FILLCELL_X4 FILLER_86_274 ();
 FILLCELL_X4 FILLER_86_282 ();
 FILLCELL_X8 FILLER_86_295 ();
 FILLCELL_X2 FILLER_86_303 ();
 FILLCELL_X4 FILLER_86_310 ();
 FILLCELL_X4 FILLER_86_317 ();
 FILLCELL_X8 FILLER_86_325 ();
 FILLCELL_X4 FILLER_86_333 ();
 FILLCELL_X2 FILLER_86_337 ();
 FILLCELL_X4 FILLER_86_344 ();
 FILLCELL_X4 FILLER_86_353 ();
 FILLCELL_X2 FILLER_86_357 ();
 FILLCELL_X4 FILLER_86_363 ();
 FILLCELL_X8 FILLER_86_371 ();
 FILLCELL_X1 FILLER_86_379 ();
 FILLCELL_X32 FILLER_86_1518 ();
 FILLCELL_X32 FILLER_86_1550 ();
 FILLCELL_X32 FILLER_86_1582 ();
 FILLCELL_X32 FILLER_86_1614 ();
 FILLCELL_X32 FILLER_86_1646 ();
 FILLCELL_X32 FILLER_86_1678 ();
 FILLCELL_X32 FILLER_86_1710 ();
 FILLCELL_X8 FILLER_86_1742 ();
 FILLCELL_X4 FILLER_86_1750 ();
 FILLCELL_X2 FILLER_86_1754 ();
 FILLCELL_X8 FILLER_87_1 ();
 FILLCELL_X2 FILLER_87_9 ();
 FILLCELL_X1 FILLER_87_11 ();
 FILLCELL_X4 FILLER_87_21 ();
 FILLCELL_X8 FILLER_87_31 ();
 FILLCELL_X4 FILLER_87_48 ();
 FILLCELL_X4 FILLER_87_61 ();
 FILLCELL_X1 FILLER_87_65 ();
 FILLCELL_X4 FILLER_87_75 ();
 FILLCELL_X4 FILLER_87_88 ();
 FILLCELL_X4 FILLER_87_97 ();
 FILLCELL_X4 FILLER_87_110 ();
 FILLCELL_X4 FILLER_87_123 ();
 FILLCELL_X4 FILLER_87_133 ();
 FILLCELL_X8 FILLER_87_141 ();
 FILLCELL_X4 FILLER_87_149 ();
 FILLCELL_X4 FILLER_87_159 ();
 FILLCELL_X4 FILLER_87_168 ();
 FILLCELL_X8 FILLER_87_176 ();
 FILLCELL_X4 FILLER_87_184 ();
 FILLCELL_X2 FILLER_87_188 ();
 FILLCELL_X1 FILLER_87_190 ();
 FILLCELL_X4 FILLER_87_195 ();
 FILLCELL_X16 FILLER_87_205 ();
 FILLCELL_X4 FILLER_87_221 ();
 FILLCELL_X1 FILLER_87_225 ();
 FILLCELL_X4 FILLER_87_235 ();
 FILLCELL_X2 FILLER_87_239 ();
 FILLCELL_X1 FILLER_87_241 ();
 FILLCELL_X4 FILLER_87_248 ();
 FILLCELL_X4 FILLER_87_257 ();
 FILLCELL_X4 FILLER_87_270 ();
 FILLCELL_X2 FILLER_87_274 ();
 FILLCELL_X1 FILLER_87_276 ();
 FILLCELL_X8 FILLER_87_281 ();
 FILLCELL_X2 FILLER_87_289 ();
 FILLCELL_X16 FILLER_87_295 ();
 FILLCELL_X2 FILLER_87_311 ();
 FILLCELL_X1 FILLER_87_313 ();
 FILLCELL_X4 FILLER_87_323 ();
 FILLCELL_X16 FILLER_87_336 ();
 FILLCELL_X4 FILLER_87_352 ();
 FILLCELL_X4 FILLER_87_365 ();
 FILLCELL_X4 FILLER_87_373 ();
 FILLCELL_X2 FILLER_87_377 ();
 FILLCELL_X1 FILLER_87_379 ();
 FILLCELL_X32 FILLER_87_1518 ();
 FILLCELL_X32 FILLER_87_1550 ();
 FILLCELL_X32 FILLER_87_1582 ();
 FILLCELL_X32 FILLER_87_1614 ();
 FILLCELL_X32 FILLER_87_1646 ();
 FILLCELL_X32 FILLER_87_1678 ();
 FILLCELL_X32 FILLER_87_1710 ();
 FILLCELL_X4 FILLER_87_1742 ();
 FILLCELL_X2 FILLER_87_1746 ();
 FILLCELL_X1 FILLER_87_1748 ();
 FILLCELL_X4 FILLER_87_1752 ();
 FILLCELL_X4 FILLER_88_1 ();
 FILLCELL_X2 FILLER_88_5 ();
 FILLCELL_X1 FILLER_88_7 ();
 FILLCELL_X4 FILLER_88_12 ();
 FILLCELL_X1 FILLER_88_16 ();
 FILLCELL_X4 FILLER_88_22 ();
 FILLCELL_X4 FILLER_88_30 ();
 FILLCELL_X8 FILLER_88_37 ();
 FILLCELL_X4 FILLER_88_48 ();
 FILLCELL_X4 FILLER_88_58 ();
 FILLCELL_X8 FILLER_88_67 ();
 FILLCELL_X1 FILLER_88_75 ();
 FILLCELL_X4 FILLER_88_81 ();
 FILLCELL_X1 FILLER_88_85 ();
 FILLCELL_X4 FILLER_88_90 ();
 FILLCELL_X2 FILLER_88_94 ();
 FILLCELL_X4 FILLER_88_100 ();
 FILLCELL_X4 FILLER_88_107 ();
 FILLCELL_X4 FILLER_88_114 ();
 FILLCELL_X4 FILLER_88_123 ();
 FILLCELL_X2 FILLER_88_127 ();
 FILLCELL_X1 FILLER_88_129 ();
 FILLCELL_X8 FILLER_88_155 ();
 FILLCELL_X2 FILLER_88_163 ();
 FILLCELL_X1 FILLER_88_165 ();
 FILLCELL_X4 FILLER_88_170 ();
 FILLCELL_X4 FILLER_88_183 ();
 FILLCELL_X4 FILLER_88_196 ();
 FILLCELL_X4 FILLER_88_209 ();
 FILLCELL_X8 FILLER_88_216 ();
 FILLCELL_X4 FILLER_88_224 ();
 FILLCELL_X2 FILLER_88_228 ();
 FILLCELL_X1 FILLER_88_230 ();
 FILLCELL_X8 FILLER_88_240 ();
 FILLCELL_X4 FILLER_88_248 ();
 FILLCELL_X1 FILLER_88_252 ();
 FILLCELL_X4 FILLER_88_262 ();
 FILLCELL_X8 FILLER_88_275 ();
 FILLCELL_X2 FILLER_88_283 ();
 FILLCELL_X1 FILLER_88_285 ();
 FILLCELL_X4 FILLER_88_290 ();
 FILLCELL_X4 FILLER_88_303 ();
 FILLCELL_X4 FILLER_88_311 ();
 FILLCELL_X2 FILLER_88_315 ();
 FILLCELL_X4 FILLER_88_323 ();
 FILLCELL_X4 FILLER_88_336 ();
 FILLCELL_X4 FILLER_88_343 ();
 FILLCELL_X2 FILLER_88_347 ();
 FILLCELL_X4 FILLER_88_353 ();
 FILLCELL_X8 FILLER_88_366 ();
 FILLCELL_X4 FILLER_88_374 ();
 FILLCELL_X2 FILLER_88_378 ();
 FILLCELL_X32 FILLER_88_1518 ();
 FILLCELL_X32 FILLER_88_1550 ();
 FILLCELL_X32 FILLER_88_1582 ();
 FILLCELL_X32 FILLER_88_1614 ();
 FILLCELL_X32 FILLER_88_1646 ();
 FILLCELL_X32 FILLER_88_1678 ();
 FILLCELL_X32 FILLER_88_1710 ();
 FILLCELL_X8 FILLER_88_1742 ();
 FILLCELL_X4 FILLER_88_1750 ();
 FILLCELL_X2 FILLER_88_1754 ();
 FILLCELL_X4 FILLER_89_1 ();
 FILLCELL_X2 FILLER_89_5 ();
 FILLCELL_X1 FILLER_89_7 ();
 FILLCELL_X16 FILLER_89_12 ();
 FILLCELL_X8 FILLER_89_28 ();
 FILLCELL_X4 FILLER_89_36 ();
 FILLCELL_X2 FILLER_89_40 ();
 FILLCELL_X1 FILLER_89_42 ();
 FILLCELL_X8 FILLER_89_46 ();
 FILLCELL_X2 FILLER_89_54 ();
 FILLCELL_X4 FILLER_89_60 ();
 FILLCELL_X4 FILLER_89_67 ();
 FILLCELL_X16 FILLER_89_74 ();
 FILLCELL_X4 FILLER_89_90 ();
 FILLCELL_X2 FILLER_89_94 ();
 FILLCELL_X4 FILLER_89_100 ();
 FILLCELL_X2 FILLER_89_104 ();
 FILLCELL_X1 FILLER_89_106 ();
 FILLCELL_X4 FILLER_89_111 ();
 FILLCELL_X8 FILLER_89_119 ();
 FILLCELL_X16 FILLER_89_131 ();
 FILLCELL_X8 FILLER_89_147 ();
 FILLCELL_X2 FILLER_89_155 ();
 FILLCELL_X4 FILLER_89_166 ();
 FILLCELL_X2 FILLER_89_170 ();
 FILLCELL_X1 FILLER_89_172 ();
 FILLCELL_X8 FILLER_89_177 ();
 FILLCELL_X4 FILLER_89_185 ();
 FILLCELL_X2 FILLER_89_189 ();
 FILLCELL_X1 FILLER_89_191 ();
 FILLCELL_X4 FILLER_89_197 ();
 FILLCELL_X8 FILLER_89_204 ();
 FILLCELL_X8 FILLER_89_216 ();
 FILLCELL_X4 FILLER_89_224 ();
 FILLCELL_X1 FILLER_89_228 ();
 FILLCELL_X4 FILLER_89_234 ();
 FILLCELL_X16 FILLER_89_241 ();
 FILLCELL_X1 FILLER_89_257 ();
 FILLCELL_X4 FILLER_89_263 ();
 FILLCELL_X4 FILLER_89_273 ();
 FILLCELL_X4 FILLER_89_280 ();
 FILLCELL_X4 FILLER_89_293 ();
 FILLCELL_X8 FILLER_89_306 ();
 FILLCELL_X2 FILLER_89_314 ();
 FILLCELL_X8 FILLER_89_319 ();
 FILLCELL_X4 FILLER_89_327 ();
 FILLCELL_X2 FILLER_89_331 ();
 FILLCELL_X16 FILLER_89_338 ();
 FILLCELL_X2 FILLER_89_354 ();
 FILLCELL_X8 FILLER_89_365 ();
 FILLCELL_X4 FILLER_89_373 ();
 FILLCELL_X2 FILLER_89_377 ();
 FILLCELL_X1 FILLER_89_379 ();
 FILLCELL_X32 FILLER_89_1518 ();
 FILLCELL_X32 FILLER_89_1550 ();
 FILLCELL_X32 FILLER_89_1582 ();
 FILLCELL_X32 FILLER_89_1614 ();
 FILLCELL_X32 FILLER_89_1646 ();
 FILLCELL_X32 FILLER_89_1678 ();
 FILLCELL_X32 FILLER_89_1710 ();
 FILLCELL_X8 FILLER_89_1742 ();
 FILLCELL_X4 FILLER_89_1750 ();
 FILLCELL_X2 FILLER_89_1754 ();
 FILLCELL_X4 FILLER_90_1 ();
 FILLCELL_X8 FILLER_90_24 ();
 FILLCELL_X8 FILLER_90_41 ();
 FILLCELL_X2 FILLER_90_49 ();
 FILLCELL_X8 FILLER_90_55 ();
 FILLCELL_X2 FILLER_90_63 ();
 FILLCELL_X16 FILLER_90_71 ();
 FILLCELL_X4 FILLER_90_90 ();
 FILLCELL_X4 FILLER_90_103 ();
 FILLCELL_X8 FILLER_90_112 ();
 FILLCELL_X2 FILLER_90_120 ();
 FILLCELL_X1 FILLER_90_122 ();
 FILLCELL_X4 FILLER_90_127 ();
 FILLCELL_X16 FILLER_90_135 ();
 FILLCELL_X4 FILLER_90_155 ();
 FILLCELL_X8 FILLER_90_168 ();
 FILLCELL_X16 FILLER_90_180 ();
 FILLCELL_X4 FILLER_90_196 ();
 FILLCELL_X2 FILLER_90_200 ();
 FILLCELL_X1 FILLER_90_202 ();
 FILLCELL_X4 FILLER_90_212 ();
 FILLCELL_X16 FILLER_90_225 ();
 FILLCELL_X2 FILLER_90_241 ();
 FILLCELL_X16 FILLER_90_247 ();
 FILLCELL_X4 FILLER_90_263 ();
 FILLCELL_X16 FILLER_90_270 ();
 FILLCELL_X4 FILLER_90_286 ();
 FILLCELL_X2 FILLER_90_290 ();
 FILLCELL_X1 FILLER_90_292 ();
 FILLCELL_X16 FILLER_90_296 ();
 FILLCELL_X4 FILLER_90_312 ();
 FILLCELL_X8 FILLER_90_320 ();
 FILLCELL_X2 FILLER_90_328 ();
 FILLCELL_X8 FILLER_90_334 ();
 FILLCELL_X4 FILLER_90_342 ();
 FILLCELL_X4 FILLER_90_351 ();
 FILLCELL_X4 FILLER_90_361 ();
 FILLCELL_X8 FILLER_90_370 ();
 FILLCELL_X2 FILLER_90_378 ();
 FILLCELL_X32 FILLER_90_1518 ();
 FILLCELL_X32 FILLER_90_1550 ();
 FILLCELL_X32 FILLER_90_1582 ();
 FILLCELL_X32 FILLER_90_1614 ();
 FILLCELL_X32 FILLER_90_1646 ();
 FILLCELL_X32 FILLER_90_1678 ();
 FILLCELL_X32 FILLER_90_1710 ();
 FILLCELL_X8 FILLER_90_1742 ();
 FILLCELL_X4 FILLER_90_1750 ();
 FILLCELL_X2 FILLER_90_1754 ();
 FILLCELL_X16 FILLER_91_1 ();
 FILLCELL_X8 FILLER_91_17 ();
 FILLCELL_X4 FILLER_91_28 ();
 FILLCELL_X4 FILLER_91_41 ();
 FILLCELL_X4 FILLER_91_50 ();
 FILLCELL_X2 FILLER_91_54 ();
 FILLCELL_X1 FILLER_91_56 ();
 FILLCELL_X8 FILLER_91_66 ();
 FILLCELL_X4 FILLER_91_83 ();
 FILLCELL_X4 FILLER_91_91 ();
 FILLCELL_X1 FILLER_91_95 ();
 FILLCELL_X4 FILLER_91_100 ();
 FILLCELL_X8 FILLER_91_113 ();
 FILLCELL_X4 FILLER_91_125 ();
 FILLCELL_X4 FILLER_91_134 ();
 FILLCELL_X16 FILLER_91_142 ();
 FILLCELL_X1 FILLER_91_158 ();
 FILLCELL_X8 FILLER_91_168 ();
 FILLCELL_X2 FILLER_91_176 ();
 FILLCELL_X4 FILLER_91_182 ();
 FILLCELL_X4 FILLER_91_190 ();
 FILLCELL_X8 FILLER_91_198 ();
 FILLCELL_X4 FILLER_91_206 ();
 FILLCELL_X2 FILLER_91_210 ();
 FILLCELL_X1 FILLER_91_212 ();
 FILLCELL_X4 FILLER_91_217 ();
 FILLCELL_X4 FILLER_91_230 ();
 FILLCELL_X2 FILLER_91_234 ();
 FILLCELL_X1 FILLER_91_236 ();
 FILLCELL_X4 FILLER_91_241 ();
 FILLCELL_X4 FILLER_91_254 ();
 FILLCELL_X4 FILLER_91_262 ();
 FILLCELL_X4 FILLER_91_270 ();
 FILLCELL_X4 FILLER_91_278 ();
 FILLCELL_X4 FILLER_91_287 ();
 FILLCELL_X4 FILLER_91_297 ();
 FILLCELL_X4 FILLER_91_304 ();
 FILLCELL_X2 FILLER_91_308 ();
 FILLCELL_X1 FILLER_91_310 ();
 FILLCELL_X4 FILLER_91_315 ();
 FILLCELL_X4 FILLER_91_328 ();
 FILLCELL_X2 FILLER_91_332 ();
 FILLCELL_X4 FILLER_91_338 ();
 FILLCELL_X4 FILLER_91_346 ();
 FILLCELL_X2 FILLER_91_350 ();
 FILLCELL_X1 FILLER_91_352 ();
 FILLCELL_X4 FILLER_91_356 ();
 FILLCELL_X16 FILLER_91_364 ();
 FILLCELL_X32 FILLER_91_1518 ();
 FILLCELL_X32 FILLER_91_1550 ();
 FILLCELL_X32 FILLER_91_1582 ();
 FILLCELL_X32 FILLER_91_1614 ();
 FILLCELL_X32 FILLER_91_1646 ();
 FILLCELL_X32 FILLER_91_1678 ();
 FILLCELL_X32 FILLER_91_1710 ();
 FILLCELL_X8 FILLER_91_1742 ();
 FILLCELL_X4 FILLER_91_1750 ();
 FILLCELL_X2 FILLER_91_1754 ();
 FILLCELL_X4 FILLER_92_1 ();
 FILLCELL_X16 FILLER_92_8 ();
 FILLCELL_X4 FILLER_92_24 ();
 FILLCELL_X1 FILLER_92_28 ();
 FILLCELL_X4 FILLER_92_35 ();
 FILLCELL_X4 FILLER_92_43 ();
 FILLCELL_X2 FILLER_92_47 ();
 FILLCELL_X1 FILLER_92_49 ();
 FILLCELL_X4 FILLER_92_53 ();
 FILLCELL_X4 FILLER_92_60 ();
 FILLCELL_X4 FILLER_92_69 ();
 FILLCELL_X8 FILLER_92_77 ();
 FILLCELL_X2 FILLER_92_85 ();
 FILLCELL_X1 FILLER_92_87 ();
 FILLCELL_X4 FILLER_92_91 ();
 FILLCELL_X4 FILLER_92_101 ();
 FILLCELL_X8 FILLER_92_110 ();
 FILLCELL_X2 FILLER_92_118 ();
 FILLCELL_X1 FILLER_92_120 ();
 FILLCELL_X4 FILLER_92_130 ();
 FILLCELL_X4 FILLER_92_143 ();
 FILLCELL_X4 FILLER_92_152 ();
 FILLCELL_X4 FILLER_92_162 ();
 FILLCELL_X8 FILLER_92_171 ();
 FILLCELL_X4 FILLER_92_179 ();
 FILLCELL_X8 FILLER_92_192 ();
 FILLCELL_X2 FILLER_92_200 ();
 FILLCELL_X4 FILLER_92_207 ();
 FILLCELL_X4 FILLER_92_217 ();
 FILLCELL_X4 FILLER_92_224 ();
 FILLCELL_X2 FILLER_92_228 ();
 FILLCELL_X1 FILLER_92_230 ();
 FILLCELL_X4 FILLER_92_235 ();
 FILLCELL_X2 FILLER_92_239 ();
 FILLCELL_X1 FILLER_92_241 ();
 FILLCELL_X4 FILLER_92_245 ();
 FILLCELL_X4 FILLER_92_255 ();
 FILLCELL_X32 FILLER_92_268 ();
 FILLCELL_X4 FILLER_92_300 ();
 FILLCELL_X4 FILLER_92_313 ();
 FILLCELL_X4 FILLER_92_320 ();
 FILLCELL_X4 FILLER_92_329 ();
 FILLCELL_X16 FILLER_92_342 ();
 FILLCELL_X2 FILLER_92_358 ();
 FILLCELL_X16 FILLER_92_364 ();
 FILLCELL_X32 FILLER_92_1518 ();
 FILLCELL_X32 FILLER_92_1550 ();
 FILLCELL_X32 FILLER_92_1582 ();
 FILLCELL_X32 FILLER_92_1614 ();
 FILLCELL_X32 FILLER_92_1646 ();
 FILLCELL_X32 FILLER_92_1678 ();
 FILLCELL_X32 FILLER_92_1710 ();
 FILLCELL_X8 FILLER_92_1742 ();
 FILLCELL_X4 FILLER_92_1750 ();
 FILLCELL_X2 FILLER_92_1754 ();
 FILLCELL_X32 FILLER_93_1 ();
 FILLCELL_X4 FILLER_93_33 ();
 FILLCELL_X16 FILLER_93_40 ();
 FILLCELL_X8 FILLER_93_56 ();
 FILLCELL_X4 FILLER_93_64 ();
 FILLCELL_X2 FILLER_93_68 ();
 FILLCELL_X1 FILLER_93_70 ();
 FILLCELL_X8 FILLER_93_74 ();
 FILLCELL_X4 FILLER_93_82 ();
 FILLCELL_X1 FILLER_93_86 ();
 FILLCELL_X4 FILLER_93_91 ();
 FILLCELL_X16 FILLER_93_99 ();
 FILLCELL_X8 FILLER_93_115 ();
 FILLCELL_X4 FILLER_93_123 ();
 FILLCELL_X1 FILLER_93_127 ();
 FILLCELL_X4 FILLER_93_131 ();
 FILLCELL_X4 FILLER_93_138 ();
 FILLCELL_X4 FILLER_93_145 ();
 FILLCELL_X4 FILLER_93_153 ();
 FILLCELL_X1 FILLER_93_157 ();
 FILLCELL_X4 FILLER_93_161 ();
 FILLCELL_X1 FILLER_93_165 ();
 FILLCELL_X8 FILLER_93_170 ();
 FILLCELL_X4 FILLER_93_178 ();
 FILLCELL_X4 FILLER_93_187 ();
 FILLCELL_X4 FILLER_93_200 ();
 FILLCELL_X4 FILLER_93_210 ();
 FILLCELL_X8 FILLER_93_217 ();
 FILLCELL_X4 FILLER_93_225 ();
 FILLCELL_X16 FILLER_93_233 ();
 FILLCELL_X2 FILLER_93_249 ();
 FILLCELL_X1 FILLER_93_251 ();
 FILLCELL_X8 FILLER_93_257 ();
 FILLCELL_X16 FILLER_93_268 ();
 FILLCELL_X8 FILLER_93_284 ();
 FILLCELL_X4 FILLER_93_292 ();
 FILLCELL_X2 FILLER_93_296 ();
 FILLCELL_X1 FILLER_93_298 ();
 FILLCELL_X4 FILLER_93_305 ();
 FILLCELL_X4 FILLER_93_314 ();
 FILLCELL_X4 FILLER_93_322 ();
 FILLCELL_X1 FILLER_93_326 ();
 FILLCELL_X4 FILLER_93_333 ();
 FILLCELL_X8 FILLER_93_340 ();
 FILLCELL_X2 FILLER_93_348 ();
 FILLCELL_X4 FILLER_93_354 ();
 FILLCELL_X8 FILLER_93_367 ();
 FILLCELL_X4 FILLER_93_375 ();
 FILLCELL_X1 FILLER_93_379 ();
 FILLCELL_X32 FILLER_93_1518 ();
 FILLCELL_X32 FILLER_93_1550 ();
 FILLCELL_X32 FILLER_93_1582 ();
 FILLCELL_X32 FILLER_93_1614 ();
 FILLCELL_X32 FILLER_93_1646 ();
 FILLCELL_X32 FILLER_93_1678 ();
 FILLCELL_X32 FILLER_93_1710 ();
 FILLCELL_X8 FILLER_93_1742 ();
 FILLCELL_X4 FILLER_93_1750 ();
 FILLCELL_X2 FILLER_93_1754 ();
 FILLCELL_X16 FILLER_94_1 ();
 FILLCELL_X8 FILLER_94_17 ();
 FILLCELL_X2 FILLER_94_25 ();
 FILLCELL_X1 FILLER_94_27 ();
 FILLCELL_X4 FILLER_94_31 ();
 FILLCELL_X1 FILLER_94_35 ();
 FILLCELL_X4 FILLER_94_45 ();
 FILLCELL_X8 FILLER_94_54 ();
 FILLCELL_X1 FILLER_94_62 ();
 FILLCELL_X4 FILLER_94_72 ();
 FILLCELL_X4 FILLER_94_81 ();
 FILLCELL_X1 FILLER_94_85 ();
 FILLCELL_X4 FILLER_94_90 ();
 FILLCELL_X4 FILLER_94_98 ();
 FILLCELL_X8 FILLER_94_107 ();
 FILLCELL_X2 FILLER_94_115 ();
 FILLCELL_X1 FILLER_94_117 ();
 FILLCELL_X4 FILLER_94_127 ();
 FILLCELL_X4 FILLER_94_134 ();
 FILLCELL_X1 FILLER_94_138 ();
 FILLCELL_X8 FILLER_94_145 ();
 FILLCELL_X2 FILLER_94_153 ();
 FILLCELL_X4 FILLER_94_159 ();
 FILLCELL_X2 FILLER_94_163 ();
 FILLCELL_X8 FILLER_94_169 ();
 FILLCELL_X1 FILLER_94_177 ();
 FILLCELL_X4 FILLER_94_181 ();
 FILLCELL_X4 FILLER_94_188 ();
 FILLCELL_X4 FILLER_94_196 ();
 FILLCELL_X16 FILLER_94_203 ();
 FILLCELL_X2 FILLER_94_219 ();
 FILLCELL_X1 FILLER_94_221 ();
 FILLCELL_X4 FILLER_94_226 ();
 FILLCELL_X4 FILLER_94_239 ();
 FILLCELL_X8 FILLER_94_247 ();
 FILLCELL_X4 FILLER_94_255 ();
 FILLCELL_X8 FILLER_94_262 ();
 FILLCELL_X4 FILLER_94_275 ();
 FILLCELL_X4 FILLER_94_288 ();
 FILLCELL_X8 FILLER_94_296 ();
 FILLCELL_X2 FILLER_94_304 ();
 FILLCELL_X4 FILLER_94_315 ();
 FILLCELL_X4 FILLER_94_324 ();
 FILLCELL_X1 FILLER_94_328 ();
 FILLCELL_X8 FILLER_94_332 ();
 FILLCELL_X4 FILLER_94_340 ();
 FILLCELL_X2 FILLER_94_344 ();
 FILLCELL_X1 FILLER_94_346 ();
 FILLCELL_X4 FILLER_94_352 ();
 FILLCELL_X8 FILLER_94_361 ();
 FILLCELL_X4 FILLER_94_373 ();
 FILLCELL_X2 FILLER_94_377 ();
 FILLCELL_X1 FILLER_94_379 ();
 FILLCELL_X32 FILLER_94_1518 ();
 FILLCELL_X32 FILLER_94_1550 ();
 FILLCELL_X32 FILLER_94_1582 ();
 FILLCELL_X32 FILLER_94_1614 ();
 FILLCELL_X32 FILLER_94_1646 ();
 FILLCELL_X32 FILLER_94_1678 ();
 FILLCELL_X32 FILLER_94_1710 ();
 FILLCELL_X8 FILLER_94_1742 ();
 FILLCELL_X4 FILLER_94_1750 ();
 FILLCELL_X2 FILLER_94_1754 ();
 FILLCELL_X16 FILLER_95_1 ();
 FILLCELL_X8 FILLER_95_17 ();
 FILLCELL_X1 FILLER_95_25 ();
 FILLCELL_X4 FILLER_95_32 ();
 FILLCELL_X4 FILLER_95_45 ();
 FILLCELL_X4 FILLER_95_53 ();
 FILLCELL_X2 FILLER_95_57 ();
 FILLCELL_X1 FILLER_95_59 ();
 FILLCELL_X4 FILLER_95_63 ();
 FILLCELL_X4 FILLER_95_76 ();
 FILLCELL_X4 FILLER_95_84 ();
 FILLCELL_X2 FILLER_95_88 ();
 FILLCELL_X1 FILLER_95_90 ();
 FILLCELL_X4 FILLER_95_100 ();
 FILLCELL_X1 FILLER_95_104 ();
 FILLCELL_X4 FILLER_95_108 ();
 FILLCELL_X4 FILLER_95_117 ();
 FILLCELL_X4 FILLER_95_130 ();
 FILLCELL_X16 FILLER_95_138 ();
 FILLCELL_X8 FILLER_95_154 ();
 FILLCELL_X4 FILLER_95_162 ();
 FILLCELL_X1 FILLER_95_166 ();
 FILLCELL_X4 FILLER_95_172 ();
 FILLCELL_X4 FILLER_95_179 ();
 FILLCELL_X8 FILLER_95_186 ();
 FILLCELL_X4 FILLER_95_194 ();
 FILLCELL_X8 FILLER_95_207 ();
 FILLCELL_X4 FILLER_95_219 ();
 FILLCELL_X4 FILLER_95_228 ();
 FILLCELL_X4 FILLER_95_238 ();
 FILLCELL_X4 FILLER_95_245 ();
 FILLCELL_X4 FILLER_95_254 ();
 FILLCELL_X8 FILLER_95_267 ();
 FILLCELL_X1 FILLER_95_275 ();
 FILLCELL_X4 FILLER_95_285 ();
 FILLCELL_X8 FILLER_95_295 ();
 FILLCELL_X4 FILLER_95_306 ();
 FILLCELL_X8 FILLER_95_313 ();
 FILLCELL_X2 FILLER_95_321 ();
 FILLCELL_X4 FILLER_95_329 ();
 FILLCELL_X8 FILLER_95_338 ();
 FILLCELL_X4 FILLER_95_352 ();
 FILLCELL_X4 FILLER_95_365 ();
 FILLCELL_X4 FILLER_95_373 ();
 FILLCELL_X2 FILLER_95_377 ();
 FILLCELL_X1 FILLER_95_379 ();
 FILLCELL_X32 FILLER_95_1518 ();
 FILLCELL_X32 FILLER_95_1550 ();
 FILLCELL_X32 FILLER_95_1582 ();
 FILLCELL_X32 FILLER_95_1614 ();
 FILLCELL_X32 FILLER_95_1646 ();
 FILLCELL_X32 FILLER_95_1678 ();
 FILLCELL_X32 FILLER_95_1710 ();
 FILLCELL_X8 FILLER_95_1742 ();
 FILLCELL_X4 FILLER_95_1750 ();
 FILLCELL_X2 FILLER_95_1754 ();
 FILLCELL_X32 FILLER_96_1 ();
 FILLCELL_X8 FILLER_96_36 ();
 FILLCELL_X1 FILLER_96_44 ();
 FILLCELL_X8 FILLER_96_48 ();
 FILLCELL_X1 FILLER_96_56 ();
 FILLCELL_X8 FILLER_96_60 ();
 FILLCELL_X16 FILLER_96_74 ();
 FILLCELL_X2 FILLER_96_90 ();
 FILLCELL_X4 FILLER_96_101 ();
 FILLCELL_X4 FILLER_96_109 ();
 FILLCELL_X4 FILLER_96_116 ();
 FILLCELL_X1 FILLER_96_120 ();
 FILLCELL_X8 FILLER_96_127 ();
 FILLCELL_X1 FILLER_96_135 ();
 FILLCELL_X4 FILLER_96_139 ();
 FILLCELL_X8 FILLER_96_146 ();
 FILLCELL_X4 FILLER_96_154 ();
 FILLCELL_X1 FILLER_96_158 ();
 FILLCELL_X4 FILLER_96_168 ();
 FILLCELL_X4 FILLER_96_181 ();
 FILLCELL_X8 FILLER_96_191 ();
 FILLCELL_X2 FILLER_96_199 ();
 FILLCELL_X4 FILLER_96_210 ();
 FILLCELL_X8 FILLER_96_218 ();
 FILLCELL_X8 FILLER_96_235 ();
 FILLCELL_X4 FILLER_96_246 ();
 FILLCELL_X2 FILLER_96_250 ();
 FILLCELL_X4 FILLER_96_261 ();
 FILLCELL_X4 FILLER_96_269 ();
 FILLCELL_X4 FILLER_96_276 ();
 FILLCELL_X8 FILLER_96_283 ();
 FILLCELL_X2 FILLER_96_291 ();
 FILLCELL_X4 FILLER_96_298 ();
 FILLCELL_X4 FILLER_96_305 ();
 FILLCELL_X2 FILLER_96_309 ();
 FILLCELL_X1 FILLER_96_311 ();
 FILLCELL_X4 FILLER_96_315 ();
 FILLCELL_X4 FILLER_96_328 ();
 FILLCELL_X8 FILLER_96_341 ();
 FILLCELL_X4 FILLER_96_352 ();
 FILLCELL_X16 FILLER_96_359 ();
 FILLCELL_X4 FILLER_96_375 ();
 FILLCELL_X1 FILLER_96_379 ();
 FILLCELL_X8 FILLER_96_1518 ();
 FILLCELL_X4 FILLER_96_1526 ();
 FILLCELL_X2 FILLER_96_1530 ();
 FILLCELL_X32 FILLER_96_1551 ();
 FILLCELL_X32 FILLER_96_1583 ();
 FILLCELL_X32 FILLER_96_1615 ();
 FILLCELL_X32 FILLER_96_1647 ();
 FILLCELL_X32 FILLER_96_1679 ();
 FILLCELL_X32 FILLER_96_1711 ();
 FILLCELL_X8 FILLER_96_1743 ();
 FILLCELL_X4 FILLER_96_1751 ();
 FILLCELL_X1 FILLER_96_1755 ();
 FILLCELL_X32 FILLER_97_1 ();
 FILLCELL_X8 FILLER_97_33 ();
 FILLCELL_X8 FILLER_97_60 ();
 FILLCELL_X4 FILLER_97_71 ();
 FILLCELL_X4 FILLER_97_80 ();
 FILLCELL_X2 FILLER_97_84 ();
 FILLCELL_X1 FILLER_97_86 ();
 FILLCELL_X4 FILLER_97_90 ();
 FILLCELL_X4 FILLER_97_100 ();
 FILLCELL_X16 FILLER_97_109 ();
 FILLCELL_X8 FILLER_97_125 ();
 FILLCELL_X2 FILLER_97_133 ();
 FILLCELL_X4 FILLER_97_140 ();
 FILLCELL_X4 FILLER_97_153 ();
 FILLCELL_X8 FILLER_97_161 ();
 FILLCELL_X2 FILLER_97_169 ();
 FILLCELL_X1 FILLER_97_171 ();
 FILLCELL_X4 FILLER_97_176 ();
 FILLCELL_X8 FILLER_97_183 ();
 FILLCELL_X2 FILLER_97_191 ();
 FILLCELL_X1 FILLER_97_193 ();
 FILLCELL_X4 FILLER_97_199 ();
 FILLCELL_X2 FILLER_97_203 ();
 FILLCELL_X1 FILLER_97_205 ();
 FILLCELL_X4 FILLER_97_212 ();
 FILLCELL_X16 FILLER_97_221 ();
 FILLCELL_X1 FILLER_97_237 ();
 FILLCELL_X4 FILLER_97_241 ();
 FILLCELL_X2 FILLER_97_245 ();
 FILLCELL_X4 FILLER_97_250 ();
 FILLCELL_X16 FILLER_97_260 ();
 FILLCELL_X8 FILLER_97_276 ();
 FILLCELL_X4 FILLER_97_293 ();
 FILLCELL_X4 FILLER_97_306 ();
 FILLCELL_X8 FILLER_97_314 ();
 FILLCELL_X2 FILLER_97_322 ();
 FILLCELL_X4 FILLER_97_327 ();
 FILLCELL_X1 FILLER_97_331 ();
 FILLCELL_X32 FILLER_97_336 ();
 FILLCELL_X8 FILLER_97_368 ();
 FILLCELL_X4 FILLER_97_376 ();
 FILLCELL_X8 FILLER_97_1518 ();
 FILLCELL_X2 FILLER_97_1526 ();
 FILLCELL_X1 FILLER_97_1528 ();
 FILLCELL_X32 FILLER_97_1533 ();
 FILLCELL_X32 FILLER_97_1565 ();
 FILLCELL_X32 FILLER_97_1597 ();
 FILLCELL_X32 FILLER_97_1629 ();
 FILLCELL_X32 FILLER_97_1661 ();
 FILLCELL_X32 FILLER_97_1693 ();
 FILLCELL_X16 FILLER_97_1725 ();
 FILLCELL_X8 FILLER_97_1741 ();
 FILLCELL_X4 FILLER_97_1752 ();
 FILLCELL_X32 FILLER_98_1 ();
 FILLCELL_X4 FILLER_98_33 ();
 FILLCELL_X2 FILLER_98_37 ();
 FILLCELL_X8 FILLER_98_43 ();
 FILLCELL_X1 FILLER_98_51 ();
 FILLCELL_X4 FILLER_98_55 ();
 FILLCELL_X8 FILLER_98_66 ();
 FILLCELL_X2 FILLER_98_74 ();
 FILLCELL_X32 FILLER_98_80 ();
 FILLCELL_X2 FILLER_98_112 ();
 FILLCELL_X4 FILLER_98_117 ();
 FILLCELL_X2 FILLER_98_121 ();
 FILLCELL_X1 FILLER_98_123 ();
 FILLCELL_X8 FILLER_98_130 ();
 FILLCELL_X1 FILLER_98_138 ();
 FILLCELL_X4 FILLER_98_142 ();
 FILLCELL_X4 FILLER_98_155 ();
 FILLCELL_X32 FILLER_98_165 ();
 FILLCELL_X1 FILLER_98_197 ();
 FILLCELL_X4 FILLER_98_201 ();
 FILLCELL_X4 FILLER_98_208 ();
 FILLCELL_X2 FILLER_98_212 ();
 FILLCELL_X8 FILLER_98_217 ();
 FILLCELL_X4 FILLER_98_225 ();
 FILLCELL_X8 FILLER_98_235 ();
 FILLCELL_X2 FILLER_98_243 ();
 FILLCELL_X1 FILLER_98_245 ();
 FILLCELL_X8 FILLER_98_249 ();
 FILLCELL_X4 FILLER_98_260 ();
 FILLCELL_X4 FILLER_98_269 ();
 FILLCELL_X8 FILLER_98_277 ();
 FILLCELL_X4 FILLER_98_285 ();
 FILLCELL_X4 FILLER_98_292 ();
 FILLCELL_X4 FILLER_98_302 ();
 FILLCELL_X4 FILLER_98_309 ();
 FILLCELL_X1 FILLER_98_313 ();
 FILLCELL_X8 FILLER_98_317 ();
 FILLCELL_X2 FILLER_98_325 ();
 FILLCELL_X32 FILLER_98_330 ();
 FILLCELL_X16 FILLER_98_362 ();
 FILLCELL_X2 FILLER_98_378 ();
 FILLCELL_X4 FILLER_98_1518 ();
 FILLCELL_X1 FILLER_98_1522 ();
 FILLCELL_X4 FILLER_98_1527 ();
 FILLCELL_X32 FILLER_98_1550 ();
 FILLCELL_X32 FILLER_98_1582 ();
 FILLCELL_X32 FILLER_98_1614 ();
 FILLCELL_X32 FILLER_98_1646 ();
 FILLCELL_X32 FILLER_98_1678 ();
 FILLCELL_X32 FILLER_98_1710 ();
 FILLCELL_X8 FILLER_98_1742 ();
 FILLCELL_X4 FILLER_98_1750 ();
 FILLCELL_X2 FILLER_98_1754 ();
 FILLCELL_X32 FILLER_99_1 ();
 FILLCELL_X16 FILLER_99_33 ();
 FILLCELL_X8 FILLER_99_49 ();
 FILLCELL_X1 FILLER_99_57 ();
 FILLCELL_X4 FILLER_99_64 ();
 FILLCELL_X4 FILLER_99_74 ();
 FILLCELL_X8 FILLER_99_95 ();
 FILLCELL_X4 FILLER_99_103 ();
 FILLCELL_X4 FILLER_99_110 ();
 FILLCELL_X4 FILLER_99_123 ();
 FILLCELL_X4 FILLER_99_136 ();
 FILLCELL_X8 FILLER_99_143 ();
 FILLCELL_X4 FILLER_99_151 ();
 FILLCELL_X1 FILLER_99_155 ();
 FILLCELL_X4 FILLER_99_161 ();
 FILLCELL_X2 FILLER_99_165 ();
 FILLCELL_X1 FILLER_99_167 ();
 FILLCELL_X4 FILLER_99_171 ();
 FILLCELL_X4 FILLER_99_184 ();
 FILLCELL_X4 FILLER_99_193 ();
 FILLCELL_X4 FILLER_99_201 ();
 FILLCELL_X1 FILLER_99_205 ();
 FILLCELL_X4 FILLER_99_212 ();
 FILLCELL_X1 FILLER_99_216 ();
 FILLCELL_X4 FILLER_99_221 ();
 FILLCELL_X4 FILLER_99_232 ();
 FILLCELL_X8 FILLER_99_246 ();
 FILLCELL_X1 FILLER_99_254 ();
 FILLCELL_X4 FILLER_99_264 ();
 FILLCELL_X8 FILLER_99_277 ();
 FILLCELL_X4 FILLER_99_285 ();
 FILLCELL_X2 FILLER_99_289 ();
 FILLCELL_X1 FILLER_99_291 ();
 FILLCELL_X4 FILLER_99_295 ();
 FILLCELL_X2 FILLER_99_299 ();
 FILLCELL_X4 FILLER_99_304 ();
 FILLCELL_X4 FILLER_99_317 ();
 FILLCELL_X32 FILLER_99_331 ();
 FILLCELL_X16 FILLER_99_363 ();
 FILLCELL_X1 FILLER_99_379 ();
 FILLCELL_X32 FILLER_99_1518 ();
 FILLCELL_X32 FILLER_99_1550 ();
 FILLCELL_X32 FILLER_99_1582 ();
 FILLCELL_X32 FILLER_99_1614 ();
 FILLCELL_X32 FILLER_99_1646 ();
 FILLCELL_X32 FILLER_99_1678 ();
 FILLCELL_X32 FILLER_99_1710 ();
 FILLCELL_X8 FILLER_99_1742 ();
 FILLCELL_X4 FILLER_99_1750 ();
 FILLCELL_X2 FILLER_99_1754 ();
 FILLCELL_X32 FILLER_100_1 ();
 FILLCELL_X32 FILLER_100_33 ();
 FILLCELL_X32 FILLER_100_65 ();
 FILLCELL_X16 FILLER_100_97 ();
 FILLCELL_X8 FILLER_100_113 ();
 FILLCELL_X4 FILLER_100_126 ();
 FILLCELL_X8 FILLER_100_134 ();
 FILLCELL_X4 FILLER_100_142 ();
 FILLCELL_X2 FILLER_100_146 ();
 FILLCELL_X1 FILLER_100_148 ();
 FILLCELL_X8 FILLER_100_153 ();
 FILLCELL_X2 FILLER_100_161 ();
 FILLCELL_X4 FILLER_100_166 ();
 FILLCELL_X4 FILLER_100_176 ();
 FILLCELL_X4 FILLER_100_189 ();
 FILLCELL_X4 FILLER_100_202 ();
 FILLCELL_X4 FILLER_100_215 ();
 FILLCELL_X4 FILLER_100_223 ();
 FILLCELL_X1 FILLER_100_227 ();
 FILLCELL_X16 FILLER_100_232 ();
 FILLCELL_X8 FILLER_100_248 ();
 FILLCELL_X2 FILLER_100_256 ();
 FILLCELL_X4 FILLER_100_261 ();
 FILLCELL_X4 FILLER_100_271 ();
 FILLCELL_X8 FILLER_100_278 ();
 FILLCELL_X1 FILLER_100_286 ();
 FILLCELL_X16 FILLER_100_291 ();
 FILLCELL_X4 FILLER_100_307 ();
 FILLCELL_X2 FILLER_100_311 ();
 FILLCELL_X1 FILLER_100_313 ();
 FILLCELL_X32 FILLER_100_321 ();
 FILLCELL_X16 FILLER_100_353 ();
 FILLCELL_X8 FILLER_100_369 ();
 FILLCELL_X2 FILLER_100_377 ();
 FILLCELL_X1 FILLER_100_379 ();
 FILLCELL_X32 FILLER_100_1518 ();
 FILLCELL_X32 FILLER_100_1550 ();
 FILLCELL_X32 FILLER_100_1582 ();
 FILLCELL_X32 FILLER_100_1614 ();
 FILLCELL_X32 FILLER_100_1646 ();
 FILLCELL_X32 FILLER_100_1678 ();
 FILLCELL_X32 FILLER_100_1710 ();
 FILLCELL_X8 FILLER_100_1742 ();
 FILLCELL_X4 FILLER_100_1750 ();
 FILLCELL_X2 FILLER_100_1754 ();
 FILLCELL_X32 FILLER_101_1 ();
 FILLCELL_X32 FILLER_101_33 ();
 FILLCELL_X32 FILLER_101_65 ();
 FILLCELL_X32 FILLER_101_97 ();
 FILLCELL_X16 FILLER_101_129 ();
 FILLCELL_X4 FILLER_101_145 ();
 FILLCELL_X2 FILLER_101_149 ();
 FILLCELL_X16 FILLER_101_170 ();
 FILLCELL_X2 FILLER_101_186 ();
 FILLCELL_X8 FILLER_101_191 ();
 FILLCELL_X4 FILLER_101_199 ();
 FILLCELL_X2 FILLER_101_203 ();
 FILLCELL_X1 FILLER_101_205 ();
 FILLCELL_X4 FILLER_101_211 ();
 FILLCELL_X4 FILLER_101_218 ();
 FILLCELL_X1 FILLER_101_222 ();
 FILLCELL_X4 FILLER_101_226 ();
 FILLCELL_X4 FILLER_101_233 ();
 FILLCELL_X4 FILLER_101_244 ();
 FILLCELL_X4 FILLER_101_251 ();
 FILLCELL_X2 FILLER_101_255 ();
 FILLCELL_X16 FILLER_101_260 ();
 FILLCELL_X2 FILLER_101_276 ();
 FILLCELL_X4 FILLER_101_284 ();
 FILLCELL_X4 FILLER_101_295 ();
 FILLCELL_X32 FILLER_101_303 ();
 FILLCELL_X32 FILLER_101_335 ();
 FILLCELL_X8 FILLER_101_367 ();
 FILLCELL_X4 FILLER_101_375 ();
 FILLCELL_X1 FILLER_101_379 ();
 FILLCELL_X32 FILLER_101_1518 ();
 FILLCELL_X32 FILLER_101_1550 ();
 FILLCELL_X32 FILLER_101_1582 ();
 FILLCELL_X32 FILLER_101_1614 ();
 FILLCELL_X32 FILLER_101_1646 ();
 FILLCELL_X32 FILLER_101_1678 ();
 FILLCELL_X32 FILLER_101_1710 ();
 FILLCELL_X8 FILLER_101_1742 ();
 FILLCELL_X4 FILLER_101_1750 ();
 FILLCELL_X2 FILLER_101_1754 ();
 FILLCELL_X4 FILLER_102_1 ();
 FILLCELL_X32 FILLER_102_8 ();
 FILLCELL_X32 FILLER_102_40 ();
 FILLCELL_X32 FILLER_102_72 ();
 FILLCELL_X32 FILLER_102_104 ();
 FILLCELL_X32 FILLER_102_136 ();
 FILLCELL_X32 FILLER_102_168 ();
 FILLCELL_X16 FILLER_102_200 ();
 FILLCELL_X8 FILLER_102_216 ();
 FILLCELL_X4 FILLER_102_224 ();
 FILLCELL_X4 FILLER_102_234 ();
 FILLCELL_X32 FILLER_102_244 ();
 FILLCELL_X8 FILLER_102_276 ();
 FILLCELL_X4 FILLER_102_284 ();
 FILLCELL_X32 FILLER_102_294 ();
 FILLCELL_X32 FILLER_102_326 ();
 FILLCELL_X16 FILLER_102_358 ();
 FILLCELL_X4 FILLER_102_374 ();
 FILLCELL_X2 FILLER_102_378 ();
 FILLCELL_X32 FILLER_102_1518 ();
 FILLCELL_X32 FILLER_102_1550 ();
 FILLCELL_X32 FILLER_102_1582 ();
 FILLCELL_X32 FILLER_102_1614 ();
 FILLCELL_X32 FILLER_102_1646 ();
 FILLCELL_X32 FILLER_102_1678 ();
 FILLCELL_X32 FILLER_102_1710 ();
 FILLCELL_X8 FILLER_102_1742 ();
 FILLCELL_X4 FILLER_102_1750 ();
 FILLCELL_X2 FILLER_102_1754 ();
 FILLCELL_X32 FILLER_103_1 ();
 FILLCELL_X32 FILLER_103_33 ();
 FILLCELL_X32 FILLER_103_65 ();
 FILLCELL_X32 FILLER_103_97 ();
 FILLCELL_X32 FILLER_103_129 ();
 FILLCELL_X32 FILLER_103_161 ();
 FILLCELL_X32 FILLER_103_193 ();
 FILLCELL_X8 FILLER_103_225 ();
 FILLCELL_X4 FILLER_103_233 ();
 FILLCELL_X2 FILLER_103_237 ();
 FILLCELL_X1 FILLER_103_239 ();
 FILLCELL_X32 FILLER_103_244 ();
 FILLCELL_X8 FILLER_103_276 ();
 FILLCELL_X2 FILLER_103_284 ();
 FILLCELL_X1 FILLER_103_286 ();
 FILLCELL_X32 FILLER_103_291 ();
 FILLCELL_X32 FILLER_103_323 ();
 FILLCELL_X16 FILLER_103_355 ();
 FILLCELL_X8 FILLER_103_371 ();
 FILLCELL_X1 FILLER_103_379 ();
 FILLCELL_X32 FILLER_103_1518 ();
 FILLCELL_X32 FILLER_103_1550 ();
 FILLCELL_X32 FILLER_103_1582 ();
 FILLCELL_X32 FILLER_103_1614 ();
 FILLCELL_X32 FILLER_103_1646 ();
 FILLCELL_X32 FILLER_103_1678 ();
 FILLCELL_X32 FILLER_103_1710 ();
 FILLCELL_X8 FILLER_103_1742 ();
 FILLCELL_X4 FILLER_103_1750 ();
 FILLCELL_X2 FILLER_103_1754 ();
 FILLCELL_X32 FILLER_104_1 ();
 FILLCELL_X32 FILLER_104_33 ();
 FILLCELL_X32 FILLER_104_65 ();
 FILLCELL_X32 FILLER_104_97 ();
 FILLCELL_X32 FILLER_104_129 ();
 FILLCELL_X32 FILLER_104_161 ();
 FILLCELL_X32 FILLER_104_193 ();
 FILLCELL_X32 FILLER_104_225 ();
 FILLCELL_X16 FILLER_104_257 ();
 FILLCELL_X8 FILLER_104_273 ();
 FILLCELL_X1 FILLER_104_281 ();
 FILLCELL_X32 FILLER_104_301 ();
 FILLCELL_X32 FILLER_104_333 ();
 FILLCELL_X8 FILLER_104_365 ();
 FILLCELL_X4 FILLER_104_373 ();
 FILLCELL_X2 FILLER_104_377 ();
 FILLCELL_X1 FILLER_104_379 ();
 FILLCELL_X32 FILLER_104_1518 ();
 FILLCELL_X32 FILLER_104_1550 ();
 FILLCELL_X32 FILLER_104_1582 ();
 FILLCELL_X32 FILLER_104_1614 ();
 FILLCELL_X32 FILLER_104_1646 ();
 FILLCELL_X32 FILLER_104_1678 ();
 FILLCELL_X32 FILLER_104_1710 ();
 FILLCELL_X8 FILLER_104_1742 ();
 FILLCELL_X4 FILLER_104_1750 ();
 FILLCELL_X2 FILLER_104_1754 ();
 FILLCELL_X32 FILLER_105_1 ();
 FILLCELL_X32 FILLER_105_33 ();
 FILLCELL_X32 FILLER_105_65 ();
 FILLCELL_X32 FILLER_105_97 ();
 FILLCELL_X32 FILLER_105_129 ();
 FILLCELL_X32 FILLER_105_161 ();
 FILLCELL_X32 FILLER_105_193 ();
 FILLCELL_X8 FILLER_105_225 ();
 FILLCELL_X4 FILLER_105_233 ();
 FILLCELL_X2 FILLER_105_237 ();
 FILLCELL_X8 FILLER_105_256 ();
 FILLCELL_X2 FILLER_105_264 ();
 FILLCELL_X1 FILLER_105_266 ();
 FILLCELL_X4 FILLER_105_270 ();
 FILLCELL_X1 FILLER_105_274 ();
 FILLCELL_X8 FILLER_105_278 ();
 FILLCELL_X4 FILLER_105_286 ();
 FILLCELL_X2 FILLER_105_290 ();
 FILLCELL_X4 FILLER_105_294 ();
 FILLCELL_X2 FILLER_105_298 ();
 FILLCELL_X1 FILLER_105_300 ();
 FILLCELL_X4 FILLER_105_306 ();
 FILLCELL_X4 FILLER_105_313 ();
 FILLCELL_X32 FILLER_105_322 ();
 FILLCELL_X16 FILLER_105_354 ();
 FILLCELL_X8 FILLER_105_370 ();
 FILLCELL_X2 FILLER_105_378 ();
 FILLCELL_X32 FILLER_105_1518 ();
 FILLCELL_X32 FILLER_105_1550 ();
 FILLCELL_X32 FILLER_105_1582 ();
 FILLCELL_X32 FILLER_105_1614 ();
 FILLCELL_X32 FILLER_105_1646 ();
 FILLCELL_X32 FILLER_105_1678 ();
 FILLCELL_X32 FILLER_105_1710 ();
 FILLCELL_X8 FILLER_105_1742 ();
 FILLCELL_X4 FILLER_105_1750 ();
 FILLCELL_X2 FILLER_105_1754 ();
 FILLCELL_X32 FILLER_106_1 ();
 FILLCELL_X32 FILLER_106_33 ();
 FILLCELL_X32 FILLER_106_65 ();
 FILLCELL_X32 FILLER_106_97 ();
 FILLCELL_X32 FILLER_106_129 ();
 FILLCELL_X32 FILLER_106_161 ();
 FILLCELL_X32 FILLER_106_193 ();
 FILLCELL_X32 FILLER_106_225 ();
 FILLCELL_X2 FILLER_106_257 ();
 FILLCELL_X1 FILLER_106_259 ();
 FILLCELL_X4 FILLER_106_277 ();
 FILLCELL_X2 FILLER_106_281 ();
 FILLCELL_X1 FILLER_106_283 ();
 FILLCELL_X4 FILLER_106_303 ();
 FILLCELL_X1 FILLER_106_307 ();
 FILLCELL_X4 FILLER_106_325 ();
 FILLCELL_X32 FILLER_106_332 ();
 FILLCELL_X16 FILLER_106_364 ();
 FILLCELL_X32 FILLER_106_1518 ();
 FILLCELL_X32 FILLER_106_1550 ();
 FILLCELL_X32 FILLER_106_1582 ();
 FILLCELL_X32 FILLER_106_1614 ();
 FILLCELL_X32 FILLER_106_1646 ();
 FILLCELL_X32 FILLER_106_1678 ();
 FILLCELL_X32 FILLER_106_1710 ();
 FILLCELL_X4 FILLER_106_1742 ();
 FILLCELL_X2 FILLER_106_1746 ();
 FILLCELL_X1 FILLER_106_1748 ();
 FILLCELL_X4 FILLER_106_1752 ();
 FILLCELL_X32 FILLER_107_1 ();
 FILLCELL_X32 FILLER_107_33 ();
 FILLCELL_X32 FILLER_107_65 ();
 FILLCELL_X32 FILLER_107_97 ();
 FILLCELL_X32 FILLER_107_129 ();
 FILLCELL_X32 FILLER_107_161 ();
 FILLCELL_X32 FILLER_107_193 ();
 FILLCELL_X16 FILLER_107_225 ();
 FILLCELL_X8 FILLER_107_241 ();
 FILLCELL_X4 FILLER_107_249 ();
 FILLCELL_X2 FILLER_107_253 ();
 FILLCELL_X1 FILLER_107_255 ();
 FILLCELL_X4 FILLER_107_259 ();
 FILLCELL_X4 FILLER_107_266 ();
 FILLCELL_X4 FILLER_107_273 ();
 FILLCELL_X4 FILLER_107_280 ();
 FILLCELL_X8 FILLER_107_288 ();
 FILLCELL_X1 FILLER_107_296 ();
 FILLCELL_X4 FILLER_107_300 ();
 FILLCELL_X8 FILLER_107_308 ();
 FILLCELL_X4 FILLER_107_320 ();
 FILLCELL_X4 FILLER_107_327 ();
 FILLCELL_X2 FILLER_107_331 ();
 FILLCELL_X4 FILLER_107_336 ();
 FILLCELL_X2 FILLER_107_340 ();
 FILLCELL_X1 FILLER_107_342 ();
 FILLCELL_X32 FILLER_107_346 ();
 FILLCELL_X2 FILLER_107_378 ();
 FILLCELL_X32 FILLER_107_1518 ();
 FILLCELL_X32 FILLER_107_1550 ();
 FILLCELL_X32 FILLER_107_1582 ();
 FILLCELL_X32 FILLER_107_1614 ();
 FILLCELL_X32 FILLER_107_1646 ();
 FILLCELL_X32 FILLER_107_1678 ();
 FILLCELL_X32 FILLER_107_1710 ();
 FILLCELL_X8 FILLER_107_1742 ();
 FILLCELL_X4 FILLER_107_1750 ();
 FILLCELL_X2 FILLER_107_1754 ();
 FILLCELL_X32 FILLER_108_1 ();
 FILLCELL_X32 FILLER_108_33 ();
 FILLCELL_X32 FILLER_108_65 ();
 FILLCELL_X32 FILLER_108_97 ();
 FILLCELL_X32 FILLER_108_129 ();
 FILLCELL_X32 FILLER_108_161 ();
 FILLCELL_X32 FILLER_108_193 ();
 FILLCELL_X8 FILLER_108_225 ();
 FILLCELL_X4 FILLER_108_233 ();
 FILLCELL_X2 FILLER_108_237 ();
 FILLCELL_X4 FILLER_108_241 ();
 FILLCELL_X8 FILLER_108_250 ();
 FILLCELL_X4 FILLER_108_263 ();
 FILLCELL_X8 FILLER_108_272 ();
 FILLCELL_X2 FILLER_108_280 ();
 FILLCELL_X4 FILLER_108_287 ();
 FILLCELL_X4 FILLER_108_295 ();
 FILLCELL_X8 FILLER_108_302 ();
 FILLCELL_X1 FILLER_108_310 ();
 FILLCELL_X4 FILLER_108_314 ();
 FILLCELL_X1 FILLER_108_318 ();
 FILLCELL_X4 FILLER_108_322 ();
 FILLCELL_X4 FILLER_108_335 ();
 FILLCELL_X2 FILLER_108_339 ();
 FILLCELL_X4 FILLER_108_346 ();
 FILLCELL_X4 FILLER_108_353 ();
 FILLCELL_X16 FILLER_108_360 ();
 FILLCELL_X4 FILLER_108_376 ();
 FILLCELL_X32 FILLER_108_1518 ();
 FILLCELL_X32 FILLER_108_1550 ();
 FILLCELL_X32 FILLER_108_1582 ();
 FILLCELL_X32 FILLER_108_1614 ();
 FILLCELL_X32 FILLER_108_1646 ();
 FILLCELL_X32 FILLER_108_1678 ();
 FILLCELL_X32 FILLER_108_1710 ();
 FILLCELL_X8 FILLER_108_1742 ();
 FILLCELL_X4 FILLER_108_1750 ();
 FILLCELL_X2 FILLER_108_1754 ();
 FILLCELL_X32 FILLER_109_1 ();
 FILLCELL_X32 FILLER_109_33 ();
 FILLCELL_X32 FILLER_109_65 ();
 FILLCELL_X32 FILLER_109_97 ();
 FILLCELL_X32 FILLER_109_129 ();
 FILLCELL_X32 FILLER_109_161 ();
 FILLCELL_X32 FILLER_109_193 ();
 FILLCELL_X8 FILLER_109_225 ();
 FILLCELL_X4 FILLER_109_233 ();
 FILLCELL_X2 FILLER_109_237 ();
 FILLCELL_X1 FILLER_109_239 ();
 FILLCELL_X4 FILLER_109_243 ();
 FILLCELL_X4 FILLER_109_264 ();
 FILLCELL_X4 FILLER_109_273 ();
 FILLCELL_X4 FILLER_109_281 ();
 FILLCELL_X2 FILLER_109_285 ();
 FILLCELL_X4 FILLER_109_291 ();
 FILLCELL_X4 FILLER_109_297 ();
 FILLCELL_X4 FILLER_109_306 ();
 FILLCELL_X8 FILLER_109_329 ();
 FILLCELL_X1 FILLER_109_337 ();
 FILLCELL_X8 FILLER_109_355 ();
 FILLCELL_X1 FILLER_109_363 ();
 FILLCELL_X8 FILLER_109_367 ();
 FILLCELL_X4 FILLER_109_375 ();
 FILLCELL_X1 FILLER_109_379 ();
 FILLCELL_X32 FILLER_109_1518 ();
 FILLCELL_X32 FILLER_109_1550 ();
 FILLCELL_X32 FILLER_109_1582 ();
 FILLCELL_X32 FILLER_109_1614 ();
 FILLCELL_X32 FILLER_109_1646 ();
 FILLCELL_X32 FILLER_109_1678 ();
 FILLCELL_X32 FILLER_109_1710 ();
 FILLCELL_X8 FILLER_109_1742 ();
 FILLCELL_X4 FILLER_109_1750 ();
 FILLCELL_X2 FILLER_109_1754 ();
 FILLCELL_X32 FILLER_110_1 ();
 FILLCELL_X32 FILLER_110_33 ();
 FILLCELL_X32 FILLER_110_65 ();
 FILLCELL_X32 FILLER_110_97 ();
 FILLCELL_X32 FILLER_110_129 ();
 FILLCELL_X32 FILLER_110_161 ();
 FILLCELL_X32 FILLER_110_193 ();
 FILLCELL_X16 FILLER_110_225 ();
 FILLCELL_X8 FILLER_110_241 ();
 FILLCELL_X4 FILLER_110_249 ();
 FILLCELL_X4 FILLER_110_256 ();
 FILLCELL_X4 FILLER_110_263 ();
 FILLCELL_X8 FILLER_110_270 ();
 FILLCELL_X2 FILLER_110_278 ();
 FILLCELL_X1 FILLER_110_280 ();
 FILLCELL_X4 FILLER_110_283 ();
 FILLCELL_X1 FILLER_110_287 ();
 FILLCELL_X4 FILLER_110_293 ();
 FILLCELL_X4 FILLER_110_310 ();
 FILLCELL_X2 FILLER_110_314 ();
 FILLCELL_X4 FILLER_110_320 ();
 FILLCELL_X4 FILLER_110_329 ();
 FILLCELL_X2 FILLER_110_333 ();
 FILLCELL_X4 FILLER_110_338 ();
 FILLCELL_X4 FILLER_110_346 ();
 FILLCELL_X1 FILLER_110_350 ();
 FILLCELL_X4 FILLER_110_354 ();
 FILLCELL_X4 FILLER_110_361 ();
 FILLCELL_X1 FILLER_110_365 ();
 FILLCELL_X4 FILLER_110_369 ();
 FILLCELL_X4 FILLER_110_376 ();
 FILLCELL_X32 FILLER_110_1518 ();
 FILLCELL_X32 FILLER_110_1550 ();
 FILLCELL_X32 FILLER_110_1582 ();
 FILLCELL_X32 FILLER_110_1614 ();
 FILLCELL_X32 FILLER_110_1646 ();
 FILLCELL_X32 FILLER_110_1678 ();
 FILLCELL_X32 FILLER_110_1710 ();
 FILLCELL_X8 FILLER_110_1742 ();
 FILLCELL_X4 FILLER_110_1750 ();
 FILLCELL_X2 FILLER_110_1754 ();
 FILLCELL_X4 FILLER_111_1 ();
 FILLCELL_X32 FILLER_111_8 ();
 FILLCELL_X32 FILLER_111_40 ();
 FILLCELL_X32 FILLER_111_72 ();
 FILLCELL_X32 FILLER_111_104 ();
 FILLCELL_X32 FILLER_111_136 ();
 FILLCELL_X32 FILLER_111_168 ();
 FILLCELL_X32 FILLER_111_200 ();
 FILLCELL_X8 FILLER_111_232 ();
 FILLCELL_X2 FILLER_111_240 ();
 FILLCELL_X4 FILLER_111_245 ();
 FILLCELL_X4 FILLER_111_252 ();
 FILLCELL_X4 FILLER_111_259 ();
 FILLCELL_X8 FILLER_111_269 ();
 FILLCELL_X4 FILLER_111_277 ();
 FILLCELL_X1 FILLER_111_281 ();
 FILLCELL_X4 FILLER_111_286 ();
 FILLCELL_X1 FILLER_111_290 ();
 FILLCELL_X8 FILLER_111_293 ();
 FILLCELL_X4 FILLER_111_301 ();
 FILLCELL_X4 FILLER_111_308 ();
 FILLCELL_X4 FILLER_111_315 ();
 FILLCELL_X4 FILLER_111_323 ();
 FILLCELL_X2 FILLER_111_327 ();
 FILLCELL_X4 FILLER_111_332 ();
 FILLCELL_X4 FILLER_111_341 ();
 FILLCELL_X1 FILLER_111_345 ();
 FILLCELL_X4 FILLER_111_350 ();
 FILLCELL_X4 FILLER_111_356 ();
 FILLCELL_X4 FILLER_111_363 ();
 FILLCELL_X8 FILLER_111_370 ();
 FILLCELL_X2 FILLER_111_378 ();
 FILLCELL_X32 FILLER_111_1518 ();
 FILLCELL_X32 FILLER_111_1550 ();
 FILLCELL_X32 FILLER_111_1582 ();
 FILLCELL_X32 FILLER_111_1614 ();
 FILLCELL_X32 FILLER_111_1646 ();
 FILLCELL_X32 FILLER_111_1678 ();
 FILLCELL_X32 FILLER_111_1710 ();
 FILLCELL_X8 FILLER_111_1742 ();
 FILLCELL_X4 FILLER_111_1750 ();
 FILLCELL_X2 FILLER_111_1754 ();
 FILLCELL_X32 FILLER_112_1 ();
 FILLCELL_X32 FILLER_112_33 ();
 FILLCELL_X32 FILLER_112_65 ();
 FILLCELL_X32 FILLER_112_97 ();
 FILLCELL_X32 FILLER_112_129 ();
 FILLCELL_X32 FILLER_112_161 ();
 FILLCELL_X32 FILLER_112_193 ();
 FILLCELL_X16 FILLER_112_225 ();
 FILLCELL_X2 FILLER_112_241 ();
 FILLCELL_X1 FILLER_112_243 ();
 FILLCELL_X4 FILLER_112_261 ();
 FILLCELL_X2 FILLER_112_265 ();
 FILLCELL_X1 FILLER_112_267 ();
 FILLCELL_X4 FILLER_112_279 ();
 FILLCELL_X4 FILLER_112_290 ();
 FILLCELL_X2 FILLER_112_294 ();
 FILLCELL_X1 FILLER_112_296 ();
 FILLCELL_X4 FILLER_112_300 ();
 FILLCELL_X4 FILLER_112_307 ();
 FILLCELL_X4 FILLER_112_316 ();
 FILLCELL_X4 FILLER_112_325 ();
 FILLCELL_X4 FILLER_112_334 ();
 FILLCELL_X1 FILLER_112_338 ();
 FILLCELL_X4 FILLER_112_342 ();
 FILLCELL_X4 FILLER_112_363 ();
 FILLCELL_X4 FILLER_112_373 ();
 FILLCELL_X2 FILLER_112_377 ();
 FILLCELL_X1 FILLER_112_379 ();
 FILLCELL_X32 FILLER_112_1518 ();
 FILLCELL_X32 FILLER_112_1550 ();
 FILLCELL_X32 FILLER_112_1582 ();
 FILLCELL_X32 FILLER_112_1614 ();
 FILLCELL_X32 FILLER_112_1646 ();
 FILLCELL_X32 FILLER_112_1678 ();
 FILLCELL_X32 FILLER_112_1710 ();
 FILLCELL_X8 FILLER_112_1742 ();
 FILLCELL_X4 FILLER_112_1750 ();
 FILLCELL_X2 FILLER_112_1754 ();
 FILLCELL_X32 FILLER_113_1 ();
 FILLCELL_X32 FILLER_113_33 ();
 FILLCELL_X32 FILLER_113_65 ();
 FILLCELL_X32 FILLER_113_97 ();
 FILLCELL_X32 FILLER_113_129 ();
 FILLCELL_X32 FILLER_113_161 ();
 FILLCELL_X32 FILLER_113_193 ();
 FILLCELL_X16 FILLER_113_225 ();
 FILLCELL_X8 FILLER_113_241 ();
 FILLCELL_X1 FILLER_113_249 ();
 FILLCELL_X4 FILLER_113_253 ();
 FILLCELL_X4 FILLER_113_262 ();
 FILLCELL_X4 FILLER_113_269 ();
 FILLCELL_X1 FILLER_113_273 ();
 FILLCELL_X4 FILLER_113_279 ();
 FILLCELL_X4 FILLER_113_287 ();
 FILLCELL_X8 FILLER_113_295 ();
 FILLCELL_X1 FILLER_113_303 ();
 FILLCELL_X4 FILLER_113_321 ();
 FILLCELL_X2 FILLER_113_325 ();
 FILLCELL_X4 FILLER_113_332 ();
 FILLCELL_X4 FILLER_113_340 ();
 FILLCELL_X4 FILLER_113_348 ();
 FILLCELL_X8 FILLER_113_356 ();
 FILLCELL_X2 FILLER_113_364 ();
 FILLCELL_X4 FILLER_113_369 ();
 FILLCELL_X4 FILLER_113_376 ();
 FILLCELL_X32 FILLER_113_1518 ();
 FILLCELL_X32 FILLER_113_1550 ();
 FILLCELL_X32 FILLER_113_1582 ();
 FILLCELL_X32 FILLER_113_1614 ();
 FILLCELL_X32 FILLER_113_1646 ();
 FILLCELL_X32 FILLER_113_1678 ();
 FILLCELL_X32 FILLER_113_1710 ();
 FILLCELL_X8 FILLER_113_1742 ();
 FILLCELL_X4 FILLER_113_1750 ();
 FILLCELL_X2 FILLER_113_1754 ();
 FILLCELL_X32 FILLER_114_1 ();
 FILLCELL_X32 FILLER_114_33 ();
 FILLCELL_X32 FILLER_114_65 ();
 FILLCELL_X32 FILLER_114_97 ();
 FILLCELL_X32 FILLER_114_129 ();
 FILLCELL_X32 FILLER_114_161 ();
 FILLCELL_X32 FILLER_114_193 ();
 FILLCELL_X16 FILLER_114_225 ();
 FILLCELL_X8 FILLER_114_241 ();
 FILLCELL_X2 FILLER_114_249 ();
 FILLCELL_X1 FILLER_114_251 ();
 FILLCELL_X4 FILLER_114_269 ();
 FILLCELL_X8 FILLER_114_278 ();
 FILLCELL_X4 FILLER_114_291 ();
 FILLCELL_X4 FILLER_114_300 ();
 FILLCELL_X1 FILLER_114_304 ();
 FILLCELL_X4 FILLER_114_308 ();
 FILLCELL_X4 FILLER_114_317 ();
 FILLCELL_X8 FILLER_114_324 ();
 FILLCELL_X4 FILLER_114_339 ();
 FILLCELL_X2 FILLER_114_343 ();
 FILLCELL_X4 FILLER_114_350 ();
 FILLCELL_X4 FILLER_114_357 ();
 FILLCELL_X4 FILLER_114_367 ();
 FILLCELL_X2 FILLER_114_371 ();
 FILLCELL_X4 FILLER_114_376 ();
 FILLCELL_X32 FILLER_114_1518 ();
 FILLCELL_X32 FILLER_114_1550 ();
 FILLCELL_X32 FILLER_114_1582 ();
 FILLCELL_X32 FILLER_114_1614 ();
 FILLCELL_X32 FILLER_114_1646 ();
 FILLCELL_X32 FILLER_114_1678 ();
 FILLCELL_X32 FILLER_114_1710 ();
 FILLCELL_X8 FILLER_114_1742 ();
 FILLCELL_X4 FILLER_114_1750 ();
 FILLCELL_X2 FILLER_114_1754 ();
 FILLCELL_X32 FILLER_115_1 ();
 FILLCELL_X32 FILLER_115_33 ();
 FILLCELL_X32 FILLER_115_65 ();
 FILLCELL_X32 FILLER_115_97 ();
 FILLCELL_X32 FILLER_115_129 ();
 FILLCELL_X32 FILLER_115_161 ();
 FILLCELL_X32 FILLER_115_193 ();
 FILLCELL_X32 FILLER_115_225 ();
 FILLCELL_X8 FILLER_115_257 ();
 FILLCELL_X4 FILLER_115_268 ();
 FILLCELL_X4 FILLER_115_275 ();
 FILLCELL_X2 FILLER_115_279 ();
 FILLCELL_X1 FILLER_115_281 ();
 FILLCELL_X4 FILLER_115_299 ();
 FILLCELL_X4 FILLER_115_306 ();
 FILLCELL_X2 FILLER_115_310 ();
 FILLCELL_X4 FILLER_115_315 ();
 FILLCELL_X4 FILLER_115_322 ();
 FILLCELL_X4 FILLER_115_329 ();
 FILLCELL_X1 FILLER_115_333 ();
 FILLCELL_X4 FILLER_115_337 ();
 FILLCELL_X2 FILLER_115_341 ();
 FILLCELL_X1 FILLER_115_343 ();
 FILLCELL_X4 FILLER_115_348 ();
 FILLCELL_X1 FILLER_115_352 ();
 FILLCELL_X8 FILLER_115_370 ();
 FILLCELL_X2 FILLER_115_378 ();
 FILLCELL_X32 FILLER_115_1518 ();
 FILLCELL_X32 FILLER_115_1550 ();
 FILLCELL_X32 FILLER_115_1582 ();
 FILLCELL_X32 FILLER_115_1614 ();
 FILLCELL_X32 FILLER_115_1646 ();
 FILLCELL_X32 FILLER_115_1678 ();
 FILLCELL_X32 FILLER_115_1710 ();
 FILLCELL_X8 FILLER_115_1742 ();
 FILLCELL_X4 FILLER_115_1750 ();
 FILLCELL_X2 FILLER_115_1754 ();
 FILLCELL_X32 FILLER_116_1 ();
 FILLCELL_X32 FILLER_116_33 ();
 FILLCELL_X32 FILLER_116_65 ();
 FILLCELL_X32 FILLER_116_97 ();
 FILLCELL_X32 FILLER_116_129 ();
 FILLCELL_X32 FILLER_116_161 ();
 FILLCELL_X32 FILLER_116_193 ();
 FILLCELL_X32 FILLER_116_225 ();
 FILLCELL_X8 FILLER_116_257 ();
 FILLCELL_X1 FILLER_116_265 ();
 FILLCELL_X4 FILLER_116_269 ();
 FILLCELL_X2 FILLER_116_273 ();
 FILLCELL_X1 FILLER_116_275 ();
 FILLCELL_X8 FILLER_116_278 ();
 FILLCELL_X4 FILLER_116_286 ();
 FILLCELL_X2 FILLER_116_290 ();
 FILLCELL_X4 FILLER_116_295 ();
 FILLCELL_X4 FILLER_116_302 ();
 FILLCELL_X4 FILLER_116_311 ();
 FILLCELL_X4 FILLER_116_321 ();
 FILLCELL_X4 FILLER_116_330 ();
 FILLCELL_X4 FILLER_116_337 ();
 FILLCELL_X1 FILLER_116_341 ();
 FILLCELL_X4 FILLER_116_348 ();
 FILLCELL_X4 FILLER_116_355 ();
 FILLCELL_X4 FILLER_116_362 ();
 FILLCELL_X4 FILLER_116_369 ();
 FILLCELL_X4 FILLER_116_376 ();
 FILLCELL_X32 FILLER_116_1518 ();
 FILLCELL_X32 FILLER_116_1550 ();
 FILLCELL_X32 FILLER_116_1582 ();
 FILLCELL_X32 FILLER_116_1614 ();
 FILLCELL_X32 FILLER_116_1646 ();
 FILLCELL_X32 FILLER_116_1678 ();
 FILLCELL_X32 FILLER_116_1710 ();
 FILLCELL_X4 FILLER_116_1742 ();
 FILLCELL_X2 FILLER_116_1746 ();
 FILLCELL_X1 FILLER_116_1748 ();
 FILLCELL_X4 FILLER_116_1752 ();
 FILLCELL_X32 FILLER_117_1 ();
 FILLCELL_X32 FILLER_117_33 ();
 FILLCELL_X32 FILLER_117_65 ();
 FILLCELL_X32 FILLER_117_97 ();
 FILLCELL_X32 FILLER_117_129 ();
 FILLCELL_X32 FILLER_117_161 ();
 FILLCELL_X32 FILLER_117_193 ();
 FILLCELL_X32 FILLER_117_225 ();
 FILLCELL_X32 FILLER_117_257 ();
 FILLCELL_X16 FILLER_117_289 ();
 FILLCELL_X4 FILLER_117_322 ();
 FILLCELL_X1 FILLER_117_326 ();
 FILLCELL_X4 FILLER_117_333 ();
 FILLCELL_X2 FILLER_117_337 ();
 FILLCELL_X1 FILLER_117_339 ();
 FILLCELL_X4 FILLER_117_344 ();
 FILLCELL_X4 FILLER_117_351 ();
 FILLCELL_X8 FILLER_117_357 ();
 FILLCELL_X1 FILLER_117_365 ();
 FILLCELL_X4 FILLER_117_369 ();
 FILLCELL_X4 FILLER_117_376 ();
 FILLCELL_X32 FILLER_117_1518 ();
 FILLCELL_X32 FILLER_117_1550 ();
 FILLCELL_X32 FILLER_117_1582 ();
 FILLCELL_X32 FILLER_117_1614 ();
 FILLCELL_X32 FILLER_117_1646 ();
 FILLCELL_X32 FILLER_117_1678 ();
 FILLCELL_X32 FILLER_117_1710 ();
 FILLCELL_X8 FILLER_117_1742 ();
 FILLCELL_X4 FILLER_117_1750 ();
 FILLCELL_X2 FILLER_117_1754 ();
 FILLCELL_X32 FILLER_118_1 ();
 FILLCELL_X32 FILLER_118_33 ();
 FILLCELL_X32 FILLER_118_65 ();
 FILLCELL_X32 FILLER_118_97 ();
 FILLCELL_X32 FILLER_118_129 ();
 FILLCELL_X32 FILLER_118_161 ();
 FILLCELL_X32 FILLER_118_193 ();
 FILLCELL_X32 FILLER_118_225 ();
 FILLCELL_X32 FILLER_118_257 ();
 FILLCELL_X16 FILLER_118_289 ();
 FILLCELL_X4 FILLER_118_305 ();
 FILLCELL_X4 FILLER_118_312 ();
 FILLCELL_X1 FILLER_118_316 ();
 FILLCELL_X4 FILLER_118_321 ();
 FILLCELL_X4 FILLER_118_342 ();
 FILLCELL_X1 FILLER_118_346 ();
 FILLCELL_X4 FILLER_118_364 ();
 FILLCELL_X8 FILLER_118_371 ();
 FILLCELL_X1 FILLER_118_379 ();
 FILLCELL_X32 FILLER_118_1518 ();
 FILLCELL_X32 FILLER_118_1550 ();
 FILLCELL_X32 FILLER_118_1582 ();
 FILLCELL_X32 FILLER_118_1614 ();
 FILLCELL_X32 FILLER_118_1646 ();
 FILLCELL_X32 FILLER_118_1678 ();
 FILLCELL_X32 FILLER_118_1710 ();
 FILLCELL_X8 FILLER_118_1742 ();
 FILLCELL_X4 FILLER_118_1750 ();
 FILLCELL_X2 FILLER_118_1754 ();
 FILLCELL_X32 FILLER_119_1 ();
 FILLCELL_X32 FILLER_119_33 ();
 FILLCELL_X32 FILLER_119_65 ();
 FILLCELL_X32 FILLER_119_97 ();
 FILLCELL_X32 FILLER_119_129 ();
 FILLCELL_X32 FILLER_119_161 ();
 FILLCELL_X32 FILLER_119_193 ();
 FILLCELL_X32 FILLER_119_225 ();
 FILLCELL_X32 FILLER_119_257 ();
 FILLCELL_X32 FILLER_119_289 ();
 FILLCELL_X8 FILLER_119_321 ();
 FILLCELL_X4 FILLER_119_329 ();
 FILLCELL_X2 FILLER_119_333 ();
 FILLCELL_X16 FILLER_119_338 ();
 FILLCELL_X8 FILLER_119_354 ();
 FILLCELL_X4 FILLER_119_362 ();
 FILLCELL_X2 FILLER_119_366 ();
 FILLCELL_X1 FILLER_119_368 ();
 FILLCELL_X8 FILLER_119_372 ();
 FILLCELL_X32 FILLER_119_1518 ();
 FILLCELL_X32 FILLER_119_1550 ();
 FILLCELL_X32 FILLER_119_1582 ();
 FILLCELL_X32 FILLER_119_1614 ();
 FILLCELL_X32 FILLER_119_1646 ();
 FILLCELL_X32 FILLER_119_1678 ();
 FILLCELL_X32 FILLER_119_1710 ();
 FILLCELL_X8 FILLER_119_1742 ();
 FILLCELL_X4 FILLER_119_1750 ();
 FILLCELL_X2 FILLER_119_1754 ();
 FILLCELL_X32 FILLER_120_1 ();
 FILLCELL_X32 FILLER_120_33 ();
 FILLCELL_X32 FILLER_120_65 ();
 FILLCELL_X32 FILLER_120_97 ();
 FILLCELL_X32 FILLER_120_129 ();
 FILLCELL_X32 FILLER_120_161 ();
 FILLCELL_X32 FILLER_120_193 ();
 FILLCELL_X32 FILLER_120_225 ();
 FILLCELL_X32 FILLER_120_257 ();
 FILLCELL_X32 FILLER_120_289 ();
 FILLCELL_X16 FILLER_120_321 ();
 FILLCELL_X2 FILLER_120_337 ();
 FILLCELL_X1 FILLER_120_339 ();
 FILLCELL_X16 FILLER_120_343 ();
 FILLCELL_X8 FILLER_120_359 ();
 FILLCELL_X4 FILLER_120_367 ();
 FILLCELL_X2 FILLER_120_371 ();
 FILLCELL_X4 FILLER_120_376 ();
 FILLCELL_X32 FILLER_120_1518 ();
 FILLCELL_X32 FILLER_120_1550 ();
 FILLCELL_X32 FILLER_120_1582 ();
 FILLCELL_X32 FILLER_120_1614 ();
 FILLCELL_X32 FILLER_120_1646 ();
 FILLCELL_X32 FILLER_120_1678 ();
 FILLCELL_X32 FILLER_120_1710 ();
 FILLCELL_X8 FILLER_120_1742 ();
 FILLCELL_X4 FILLER_120_1750 ();
 FILLCELL_X2 FILLER_120_1754 ();
 FILLCELL_X4 FILLER_121_1 ();
 FILLCELL_X32 FILLER_121_8 ();
 FILLCELL_X32 FILLER_121_40 ();
 FILLCELL_X32 FILLER_121_72 ();
 FILLCELL_X32 FILLER_121_104 ();
 FILLCELL_X32 FILLER_121_136 ();
 FILLCELL_X32 FILLER_121_168 ();
 FILLCELL_X32 FILLER_121_200 ();
 FILLCELL_X32 FILLER_121_232 ();
 FILLCELL_X32 FILLER_121_264 ();
 FILLCELL_X32 FILLER_121_296 ();
 FILLCELL_X16 FILLER_121_328 ();
 FILLCELL_X8 FILLER_121_344 ();
 FILLCELL_X4 FILLER_121_352 ();
 FILLCELL_X1 FILLER_121_356 ();
 FILLCELL_X4 FILLER_121_360 ();
 FILLCELL_X4 FILLER_121_367 ();
 FILLCELL_X2 FILLER_121_371 ();
 FILLCELL_X4 FILLER_121_376 ();
 FILLCELL_X32 FILLER_121_1518 ();
 FILLCELL_X32 FILLER_121_1550 ();
 FILLCELL_X32 FILLER_121_1582 ();
 FILLCELL_X32 FILLER_121_1614 ();
 FILLCELL_X32 FILLER_121_1646 ();
 FILLCELL_X32 FILLER_121_1678 ();
 FILLCELL_X32 FILLER_121_1710 ();
 FILLCELL_X8 FILLER_121_1742 ();
 FILLCELL_X4 FILLER_121_1750 ();
 FILLCELL_X2 FILLER_121_1754 ();
 FILLCELL_X32 FILLER_122_1 ();
 FILLCELL_X32 FILLER_122_33 ();
 FILLCELL_X32 FILLER_122_65 ();
 FILLCELL_X32 FILLER_122_97 ();
 FILLCELL_X32 FILLER_122_129 ();
 FILLCELL_X32 FILLER_122_161 ();
 FILLCELL_X32 FILLER_122_193 ();
 FILLCELL_X32 FILLER_122_225 ();
 FILLCELL_X32 FILLER_122_257 ();
 FILLCELL_X32 FILLER_122_289 ();
 FILLCELL_X32 FILLER_122_321 ();
 FILLCELL_X16 FILLER_122_353 ();
 FILLCELL_X8 FILLER_122_369 ();
 FILLCELL_X2 FILLER_122_377 ();
 FILLCELL_X1 FILLER_122_379 ();
 FILLCELL_X32 FILLER_122_1518 ();
 FILLCELL_X32 FILLER_122_1550 ();
 FILLCELL_X32 FILLER_122_1582 ();
 FILLCELL_X32 FILLER_122_1614 ();
 FILLCELL_X32 FILLER_122_1646 ();
 FILLCELL_X32 FILLER_122_1678 ();
 FILLCELL_X32 FILLER_122_1710 ();
 FILLCELL_X8 FILLER_122_1742 ();
 FILLCELL_X4 FILLER_122_1750 ();
 FILLCELL_X2 FILLER_122_1754 ();
 FILLCELL_X32 FILLER_123_1 ();
 FILLCELL_X32 FILLER_123_33 ();
 FILLCELL_X32 FILLER_123_65 ();
 FILLCELL_X32 FILLER_123_97 ();
 FILLCELL_X32 FILLER_123_129 ();
 FILLCELL_X32 FILLER_123_161 ();
 FILLCELL_X32 FILLER_123_193 ();
 FILLCELL_X32 FILLER_123_225 ();
 FILLCELL_X32 FILLER_123_257 ();
 FILLCELL_X32 FILLER_123_289 ();
 FILLCELL_X32 FILLER_123_321 ();
 FILLCELL_X8 FILLER_123_353 ();
 FILLCELL_X4 FILLER_123_361 ();
 FILLCELL_X1 FILLER_123_365 ();
 FILLCELL_X4 FILLER_123_369 ();
 FILLCELL_X4 FILLER_123_376 ();
 FILLCELL_X32 FILLER_123_1518 ();
 FILLCELL_X32 FILLER_123_1550 ();
 FILLCELL_X32 FILLER_123_1582 ();
 FILLCELL_X32 FILLER_123_1614 ();
 FILLCELL_X32 FILLER_123_1646 ();
 FILLCELL_X32 FILLER_123_1678 ();
 FILLCELL_X32 FILLER_123_1710 ();
 FILLCELL_X8 FILLER_123_1742 ();
 FILLCELL_X4 FILLER_123_1750 ();
 FILLCELL_X2 FILLER_123_1754 ();
 FILLCELL_X32 FILLER_124_1 ();
 FILLCELL_X32 FILLER_124_33 ();
 FILLCELL_X32 FILLER_124_65 ();
 FILLCELL_X32 FILLER_124_97 ();
 FILLCELL_X32 FILLER_124_129 ();
 FILLCELL_X32 FILLER_124_161 ();
 FILLCELL_X32 FILLER_124_193 ();
 FILLCELL_X32 FILLER_124_225 ();
 FILLCELL_X32 FILLER_124_257 ();
 FILLCELL_X32 FILLER_124_289 ();
 FILLCELL_X32 FILLER_124_321 ();
 FILLCELL_X16 FILLER_124_353 ();
 FILLCELL_X8 FILLER_124_369 ();
 FILLCELL_X2 FILLER_124_377 ();
 FILLCELL_X1 FILLER_124_379 ();
 FILLCELL_X32 FILLER_124_1518 ();
 FILLCELL_X32 FILLER_124_1550 ();
 FILLCELL_X32 FILLER_124_1582 ();
 FILLCELL_X32 FILLER_124_1614 ();
 FILLCELL_X32 FILLER_124_1646 ();
 FILLCELL_X32 FILLER_124_1678 ();
 FILLCELL_X32 FILLER_124_1710 ();
 FILLCELL_X8 FILLER_124_1742 ();
 FILLCELL_X4 FILLER_124_1750 ();
 FILLCELL_X2 FILLER_124_1754 ();
 FILLCELL_X32 FILLER_125_1 ();
 FILLCELL_X32 FILLER_125_33 ();
 FILLCELL_X32 FILLER_125_65 ();
 FILLCELL_X32 FILLER_125_97 ();
 FILLCELL_X32 FILLER_125_129 ();
 FILLCELL_X32 FILLER_125_161 ();
 FILLCELL_X32 FILLER_125_193 ();
 FILLCELL_X32 FILLER_125_225 ();
 FILLCELL_X32 FILLER_125_257 ();
 FILLCELL_X32 FILLER_125_289 ();
 FILLCELL_X32 FILLER_125_321 ();
 FILLCELL_X16 FILLER_125_353 ();
 FILLCELL_X8 FILLER_125_369 ();
 FILLCELL_X2 FILLER_125_377 ();
 FILLCELL_X1 FILLER_125_379 ();
 FILLCELL_X32 FILLER_125_1518 ();
 FILLCELL_X32 FILLER_125_1550 ();
 FILLCELL_X32 FILLER_125_1582 ();
 FILLCELL_X32 FILLER_125_1614 ();
 FILLCELL_X32 FILLER_125_1646 ();
 FILLCELL_X32 FILLER_125_1678 ();
 FILLCELL_X32 FILLER_125_1710 ();
 FILLCELL_X8 FILLER_125_1742 ();
 FILLCELL_X4 FILLER_125_1750 ();
 FILLCELL_X2 FILLER_125_1754 ();
 FILLCELL_X32 FILLER_126_1 ();
 FILLCELL_X32 FILLER_126_33 ();
 FILLCELL_X32 FILLER_126_65 ();
 FILLCELL_X32 FILLER_126_97 ();
 FILLCELL_X32 FILLER_126_129 ();
 FILLCELL_X32 FILLER_126_161 ();
 FILLCELL_X32 FILLER_126_193 ();
 FILLCELL_X32 FILLER_126_225 ();
 FILLCELL_X32 FILLER_126_257 ();
 FILLCELL_X32 FILLER_126_289 ();
 FILLCELL_X32 FILLER_126_321 ();
 FILLCELL_X16 FILLER_126_353 ();
 FILLCELL_X4 FILLER_126_369 ();
 FILLCELL_X4 FILLER_126_376 ();
 FILLCELL_X32 FILLER_126_1518 ();
 FILLCELL_X32 FILLER_126_1550 ();
 FILLCELL_X32 FILLER_126_1582 ();
 FILLCELL_X32 FILLER_126_1614 ();
 FILLCELL_X32 FILLER_126_1646 ();
 FILLCELL_X32 FILLER_126_1678 ();
 FILLCELL_X32 FILLER_126_1710 ();
 FILLCELL_X4 FILLER_126_1742 ();
 FILLCELL_X2 FILLER_126_1746 ();
 FILLCELL_X4 FILLER_126_1752 ();
 FILLCELL_X32 FILLER_127_1 ();
 FILLCELL_X32 FILLER_127_33 ();
 FILLCELL_X32 FILLER_127_65 ();
 FILLCELL_X32 FILLER_127_97 ();
 FILLCELL_X32 FILLER_127_129 ();
 FILLCELL_X32 FILLER_127_161 ();
 FILLCELL_X32 FILLER_127_193 ();
 FILLCELL_X32 FILLER_127_225 ();
 FILLCELL_X32 FILLER_127_257 ();
 FILLCELL_X32 FILLER_127_289 ();
 FILLCELL_X32 FILLER_127_321 ();
 FILLCELL_X16 FILLER_127_353 ();
 FILLCELL_X8 FILLER_127_369 ();
 FILLCELL_X2 FILLER_127_377 ();
 FILLCELL_X1 FILLER_127_379 ();
 FILLCELL_X32 FILLER_127_1518 ();
 FILLCELL_X32 FILLER_127_1550 ();
 FILLCELL_X32 FILLER_127_1582 ();
 FILLCELL_X32 FILLER_127_1614 ();
 FILLCELL_X32 FILLER_127_1646 ();
 FILLCELL_X32 FILLER_127_1678 ();
 FILLCELL_X32 FILLER_127_1710 ();
 FILLCELL_X8 FILLER_127_1742 ();
 FILLCELL_X4 FILLER_127_1750 ();
 FILLCELL_X2 FILLER_127_1754 ();
 FILLCELL_X32 FILLER_128_1 ();
 FILLCELL_X32 FILLER_128_33 ();
 FILLCELL_X32 FILLER_128_65 ();
 FILLCELL_X32 FILLER_128_97 ();
 FILLCELL_X32 FILLER_128_129 ();
 FILLCELL_X32 FILLER_128_161 ();
 FILLCELL_X32 FILLER_128_193 ();
 FILLCELL_X32 FILLER_128_225 ();
 FILLCELL_X32 FILLER_128_257 ();
 FILLCELL_X32 FILLER_128_289 ();
 FILLCELL_X32 FILLER_128_321 ();
 FILLCELL_X16 FILLER_128_353 ();
 FILLCELL_X8 FILLER_128_369 ();
 FILLCELL_X2 FILLER_128_377 ();
 FILLCELL_X1 FILLER_128_379 ();
 FILLCELL_X32 FILLER_128_1518 ();
 FILLCELL_X32 FILLER_128_1550 ();
 FILLCELL_X32 FILLER_128_1582 ();
 FILLCELL_X32 FILLER_128_1614 ();
 FILLCELL_X32 FILLER_128_1646 ();
 FILLCELL_X32 FILLER_128_1678 ();
 FILLCELL_X32 FILLER_128_1710 ();
 FILLCELL_X8 FILLER_128_1742 ();
 FILLCELL_X4 FILLER_128_1750 ();
 FILLCELL_X2 FILLER_128_1754 ();
 FILLCELL_X32 FILLER_129_1 ();
 FILLCELL_X32 FILLER_129_33 ();
 FILLCELL_X32 FILLER_129_65 ();
 FILLCELL_X32 FILLER_129_97 ();
 FILLCELL_X32 FILLER_129_129 ();
 FILLCELL_X32 FILLER_129_161 ();
 FILLCELL_X32 FILLER_129_193 ();
 FILLCELL_X32 FILLER_129_225 ();
 FILLCELL_X32 FILLER_129_257 ();
 FILLCELL_X32 FILLER_129_289 ();
 FILLCELL_X32 FILLER_129_321 ();
 FILLCELL_X16 FILLER_129_353 ();
 FILLCELL_X8 FILLER_129_369 ();
 FILLCELL_X2 FILLER_129_377 ();
 FILLCELL_X1 FILLER_129_379 ();
 FILLCELL_X32 FILLER_129_1518 ();
 FILLCELL_X32 FILLER_129_1550 ();
 FILLCELL_X32 FILLER_129_1582 ();
 FILLCELL_X32 FILLER_129_1614 ();
 FILLCELL_X32 FILLER_129_1646 ();
 FILLCELL_X32 FILLER_129_1678 ();
 FILLCELL_X32 FILLER_129_1710 ();
 FILLCELL_X8 FILLER_129_1742 ();
 FILLCELL_X4 FILLER_129_1750 ();
 FILLCELL_X2 FILLER_129_1754 ();
 FILLCELL_X4 FILLER_130_1 ();
 FILLCELL_X32 FILLER_130_8 ();
 FILLCELL_X32 FILLER_130_40 ();
 FILLCELL_X32 FILLER_130_72 ();
 FILLCELL_X32 FILLER_130_104 ();
 FILLCELL_X32 FILLER_130_136 ();
 FILLCELL_X32 FILLER_130_168 ();
 FILLCELL_X32 FILLER_130_200 ();
 FILLCELL_X32 FILLER_130_232 ();
 FILLCELL_X32 FILLER_130_264 ();
 FILLCELL_X32 FILLER_130_296 ();
 FILLCELL_X32 FILLER_130_328 ();
 FILLCELL_X16 FILLER_130_360 ();
 FILLCELL_X4 FILLER_130_376 ();
 FILLCELL_X32 FILLER_130_1518 ();
 FILLCELL_X32 FILLER_130_1550 ();
 FILLCELL_X32 FILLER_130_1582 ();
 FILLCELL_X32 FILLER_130_1614 ();
 FILLCELL_X32 FILLER_130_1646 ();
 FILLCELL_X32 FILLER_130_1678 ();
 FILLCELL_X32 FILLER_130_1710 ();
 FILLCELL_X8 FILLER_130_1742 ();
 FILLCELL_X4 FILLER_130_1750 ();
 FILLCELL_X2 FILLER_130_1754 ();
 FILLCELL_X32 FILLER_131_1 ();
 FILLCELL_X32 FILLER_131_33 ();
 FILLCELL_X32 FILLER_131_65 ();
 FILLCELL_X32 FILLER_131_97 ();
 FILLCELL_X32 FILLER_131_129 ();
 FILLCELL_X32 FILLER_131_161 ();
 FILLCELL_X32 FILLER_131_193 ();
 FILLCELL_X32 FILLER_131_225 ();
 FILLCELL_X32 FILLER_131_257 ();
 FILLCELL_X32 FILLER_131_289 ();
 FILLCELL_X32 FILLER_131_321 ();
 FILLCELL_X16 FILLER_131_353 ();
 FILLCELL_X8 FILLER_131_369 ();
 FILLCELL_X2 FILLER_131_377 ();
 FILLCELL_X1 FILLER_131_379 ();
 FILLCELL_X32 FILLER_131_1518 ();
 FILLCELL_X32 FILLER_131_1550 ();
 FILLCELL_X32 FILLER_131_1582 ();
 FILLCELL_X32 FILLER_131_1614 ();
 FILLCELL_X32 FILLER_131_1646 ();
 FILLCELL_X32 FILLER_131_1678 ();
 FILLCELL_X32 FILLER_131_1710 ();
 FILLCELL_X8 FILLER_131_1742 ();
 FILLCELL_X4 FILLER_131_1750 ();
 FILLCELL_X2 FILLER_131_1754 ();
 FILLCELL_X32 FILLER_132_1 ();
 FILLCELL_X32 FILLER_132_33 ();
 FILLCELL_X32 FILLER_132_65 ();
 FILLCELL_X32 FILLER_132_97 ();
 FILLCELL_X32 FILLER_132_129 ();
 FILLCELL_X32 FILLER_132_161 ();
 FILLCELL_X32 FILLER_132_193 ();
 FILLCELL_X32 FILLER_132_225 ();
 FILLCELL_X32 FILLER_132_257 ();
 FILLCELL_X32 FILLER_132_289 ();
 FILLCELL_X32 FILLER_132_321 ();
 FILLCELL_X16 FILLER_132_353 ();
 FILLCELL_X8 FILLER_132_369 ();
 FILLCELL_X2 FILLER_132_377 ();
 FILLCELL_X1 FILLER_132_379 ();
 FILLCELL_X32 FILLER_132_1518 ();
 FILLCELL_X32 FILLER_132_1550 ();
 FILLCELL_X32 FILLER_132_1582 ();
 FILLCELL_X32 FILLER_132_1614 ();
 FILLCELL_X32 FILLER_132_1646 ();
 FILLCELL_X32 FILLER_132_1678 ();
 FILLCELL_X32 FILLER_132_1710 ();
 FILLCELL_X8 FILLER_132_1742 ();
 FILLCELL_X4 FILLER_132_1750 ();
 FILLCELL_X2 FILLER_132_1754 ();
 FILLCELL_X32 FILLER_133_1 ();
 FILLCELL_X32 FILLER_133_33 ();
 FILLCELL_X32 FILLER_133_65 ();
 FILLCELL_X32 FILLER_133_97 ();
 FILLCELL_X32 FILLER_133_129 ();
 FILLCELL_X32 FILLER_133_161 ();
 FILLCELL_X32 FILLER_133_193 ();
 FILLCELL_X32 FILLER_133_225 ();
 FILLCELL_X32 FILLER_133_257 ();
 FILLCELL_X32 FILLER_133_289 ();
 FILLCELL_X32 FILLER_133_321 ();
 FILLCELL_X16 FILLER_133_353 ();
 FILLCELL_X8 FILLER_133_369 ();
 FILLCELL_X2 FILLER_133_377 ();
 FILLCELL_X1 FILLER_133_379 ();
 FILLCELL_X32 FILLER_133_1518 ();
 FILLCELL_X32 FILLER_133_1550 ();
 FILLCELL_X32 FILLER_133_1582 ();
 FILLCELL_X32 FILLER_133_1614 ();
 FILLCELL_X32 FILLER_133_1646 ();
 FILLCELL_X32 FILLER_133_1678 ();
 FILLCELL_X32 FILLER_133_1710 ();
 FILLCELL_X8 FILLER_133_1742 ();
 FILLCELL_X4 FILLER_133_1750 ();
 FILLCELL_X2 FILLER_133_1754 ();
 FILLCELL_X32 FILLER_134_1 ();
 FILLCELL_X32 FILLER_134_33 ();
 FILLCELL_X32 FILLER_134_65 ();
 FILLCELL_X32 FILLER_134_97 ();
 FILLCELL_X32 FILLER_134_129 ();
 FILLCELL_X32 FILLER_134_161 ();
 FILLCELL_X32 FILLER_134_193 ();
 FILLCELL_X32 FILLER_134_225 ();
 FILLCELL_X32 FILLER_134_257 ();
 FILLCELL_X32 FILLER_134_289 ();
 FILLCELL_X32 FILLER_134_321 ();
 FILLCELL_X16 FILLER_134_353 ();
 FILLCELL_X8 FILLER_134_369 ();
 FILLCELL_X2 FILLER_134_377 ();
 FILLCELL_X1 FILLER_134_379 ();
 FILLCELL_X32 FILLER_134_1518 ();
 FILLCELL_X32 FILLER_134_1550 ();
 FILLCELL_X32 FILLER_134_1582 ();
 FILLCELL_X32 FILLER_134_1614 ();
 FILLCELL_X32 FILLER_134_1646 ();
 FILLCELL_X32 FILLER_134_1678 ();
 FILLCELL_X32 FILLER_134_1710 ();
 FILLCELL_X8 FILLER_134_1742 ();
 FILLCELL_X4 FILLER_134_1750 ();
 FILLCELL_X2 FILLER_134_1754 ();
 FILLCELL_X32 FILLER_135_1 ();
 FILLCELL_X32 FILLER_135_33 ();
 FILLCELL_X32 FILLER_135_65 ();
 FILLCELL_X32 FILLER_135_97 ();
 FILLCELL_X32 FILLER_135_129 ();
 FILLCELL_X32 FILLER_135_161 ();
 FILLCELL_X32 FILLER_135_193 ();
 FILLCELL_X32 FILLER_135_225 ();
 FILLCELL_X32 FILLER_135_257 ();
 FILLCELL_X32 FILLER_135_289 ();
 FILLCELL_X32 FILLER_135_321 ();
 FILLCELL_X16 FILLER_135_353 ();
 FILLCELL_X8 FILLER_135_369 ();
 FILLCELL_X2 FILLER_135_377 ();
 FILLCELL_X1 FILLER_135_379 ();
 FILLCELL_X32 FILLER_135_1518 ();
 FILLCELL_X32 FILLER_135_1550 ();
 FILLCELL_X32 FILLER_135_1582 ();
 FILLCELL_X32 FILLER_135_1614 ();
 FILLCELL_X32 FILLER_135_1646 ();
 FILLCELL_X32 FILLER_135_1678 ();
 FILLCELL_X32 FILLER_135_1710 ();
 FILLCELL_X4 FILLER_135_1742 ();
 FILLCELL_X2 FILLER_135_1746 ();
 FILLCELL_X1 FILLER_135_1748 ();
 FILLCELL_X4 FILLER_135_1752 ();
 FILLCELL_X32 FILLER_136_1 ();
 FILLCELL_X32 FILLER_136_33 ();
 FILLCELL_X32 FILLER_136_65 ();
 FILLCELL_X32 FILLER_136_97 ();
 FILLCELL_X32 FILLER_136_129 ();
 FILLCELL_X32 FILLER_136_161 ();
 FILLCELL_X32 FILLER_136_193 ();
 FILLCELL_X32 FILLER_136_225 ();
 FILLCELL_X32 FILLER_136_257 ();
 FILLCELL_X32 FILLER_136_289 ();
 FILLCELL_X32 FILLER_136_321 ();
 FILLCELL_X16 FILLER_136_353 ();
 FILLCELL_X8 FILLER_136_369 ();
 FILLCELL_X2 FILLER_136_377 ();
 FILLCELL_X1 FILLER_136_379 ();
 FILLCELL_X32 FILLER_136_1518 ();
 FILLCELL_X32 FILLER_136_1550 ();
 FILLCELL_X32 FILLER_136_1582 ();
 FILLCELL_X32 FILLER_136_1614 ();
 FILLCELL_X32 FILLER_136_1646 ();
 FILLCELL_X32 FILLER_136_1678 ();
 FILLCELL_X32 FILLER_136_1710 ();
 FILLCELL_X8 FILLER_136_1742 ();
 FILLCELL_X4 FILLER_136_1750 ();
 FILLCELL_X2 FILLER_136_1754 ();
 FILLCELL_X32 FILLER_137_1 ();
 FILLCELL_X32 FILLER_137_33 ();
 FILLCELL_X32 FILLER_137_65 ();
 FILLCELL_X32 FILLER_137_97 ();
 FILLCELL_X32 FILLER_137_129 ();
 FILLCELL_X32 FILLER_137_161 ();
 FILLCELL_X32 FILLER_137_193 ();
 FILLCELL_X32 FILLER_137_225 ();
 FILLCELL_X32 FILLER_137_257 ();
 FILLCELL_X32 FILLER_137_289 ();
 FILLCELL_X32 FILLER_137_321 ();
 FILLCELL_X16 FILLER_137_353 ();
 FILLCELL_X8 FILLER_137_369 ();
 FILLCELL_X2 FILLER_137_377 ();
 FILLCELL_X1 FILLER_137_379 ();
 FILLCELL_X32 FILLER_137_1518 ();
 FILLCELL_X32 FILLER_137_1550 ();
 FILLCELL_X32 FILLER_137_1582 ();
 FILLCELL_X32 FILLER_137_1614 ();
 FILLCELL_X32 FILLER_137_1646 ();
 FILLCELL_X32 FILLER_137_1678 ();
 FILLCELL_X32 FILLER_137_1710 ();
 FILLCELL_X8 FILLER_137_1742 ();
 FILLCELL_X4 FILLER_137_1750 ();
 FILLCELL_X2 FILLER_137_1754 ();
 FILLCELL_X32 FILLER_138_1 ();
 FILLCELL_X32 FILLER_138_33 ();
 FILLCELL_X32 FILLER_138_65 ();
 FILLCELL_X32 FILLER_138_97 ();
 FILLCELL_X32 FILLER_138_129 ();
 FILLCELL_X32 FILLER_138_161 ();
 FILLCELL_X32 FILLER_138_193 ();
 FILLCELL_X32 FILLER_138_225 ();
 FILLCELL_X32 FILLER_138_257 ();
 FILLCELL_X32 FILLER_138_289 ();
 FILLCELL_X32 FILLER_138_321 ();
 FILLCELL_X16 FILLER_138_353 ();
 FILLCELL_X8 FILLER_138_369 ();
 FILLCELL_X2 FILLER_138_377 ();
 FILLCELL_X1 FILLER_138_379 ();
 FILLCELL_X32 FILLER_138_1518 ();
 FILLCELL_X32 FILLER_138_1550 ();
 FILLCELL_X32 FILLER_138_1582 ();
 FILLCELL_X32 FILLER_138_1614 ();
 FILLCELL_X32 FILLER_138_1646 ();
 FILLCELL_X32 FILLER_138_1678 ();
 FILLCELL_X32 FILLER_138_1710 ();
 FILLCELL_X8 FILLER_138_1742 ();
 FILLCELL_X4 FILLER_138_1750 ();
 FILLCELL_X2 FILLER_138_1754 ();
 FILLCELL_X32 FILLER_139_1 ();
 FILLCELL_X32 FILLER_139_33 ();
 FILLCELL_X32 FILLER_139_65 ();
 FILLCELL_X32 FILLER_139_97 ();
 FILLCELL_X32 FILLER_139_129 ();
 FILLCELL_X32 FILLER_139_161 ();
 FILLCELL_X32 FILLER_139_193 ();
 FILLCELL_X32 FILLER_139_225 ();
 FILLCELL_X32 FILLER_139_257 ();
 FILLCELL_X32 FILLER_139_289 ();
 FILLCELL_X32 FILLER_139_321 ();
 FILLCELL_X16 FILLER_139_353 ();
 FILLCELL_X8 FILLER_139_369 ();
 FILLCELL_X2 FILLER_139_377 ();
 FILLCELL_X1 FILLER_139_379 ();
 FILLCELL_X32 FILLER_139_1518 ();
 FILLCELL_X32 FILLER_139_1550 ();
 FILLCELL_X32 FILLER_139_1582 ();
 FILLCELL_X32 FILLER_139_1614 ();
 FILLCELL_X32 FILLER_139_1646 ();
 FILLCELL_X32 FILLER_139_1678 ();
 FILLCELL_X32 FILLER_139_1710 ();
 FILLCELL_X8 FILLER_139_1742 ();
 FILLCELL_X4 FILLER_139_1750 ();
 FILLCELL_X2 FILLER_139_1754 ();
 FILLCELL_X4 FILLER_140_1 ();
 FILLCELL_X32 FILLER_140_8 ();
 FILLCELL_X32 FILLER_140_40 ();
 FILLCELL_X32 FILLER_140_72 ();
 FILLCELL_X32 FILLER_140_104 ();
 FILLCELL_X32 FILLER_140_136 ();
 FILLCELL_X32 FILLER_140_168 ();
 FILLCELL_X32 FILLER_140_200 ();
 FILLCELL_X32 FILLER_140_232 ();
 FILLCELL_X32 FILLER_140_264 ();
 FILLCELL_X32 FILLER_140_296 ();
 FILLCELL_X32 FILLER_140_328 ();
 FILLCELL_X16 FILLER_140_360 ();
 FILLCELL_X4 FILLER_140_376 ();
 FILLCELL_X32 FILLER_140_1518 ();
 FILLCELL_X32 FILLER_140_1550 ();
 FILLCELL_X32 FILLER_140_1582 ();
 FILLCELL_X32 FILLER_140_1614 ();
 FILLCELL_X32 FILLER_140_1646 ();
 FILLCELL_X32 FILLER_140_1678 ();
 FILLCELL_X32 FILLER_140_1710 ();
 FILLCELL_X8 FILLER_140_1742 ();
 FILLCELL_X4 FILLER_140_1750 ();
 FILLCELL_X2 FILLER_140_1754 ();
 FILLCELL_X32 FILLER_141_1 ();
 FILLCELL_X32 FILLER_141_33 ();
 FILLCELL_X32 FILLER_141_65 ();
 FILLCELL_X32 FILLER_141_97 ();
 FILLCELL_X32 FILLER_141_129 ();
 FILLCELL_X32 FILLER_141_161 ();
 FILLCELL_X32 FILLER_141_193 ();
 FILLCELL_X32 FILLER_141_225 ();
 FILLCELL_X32 FILLER_141_257 ();
 FILLCELL_X32 FILLER_141_289 ();
 FILLCELL_X32 FILLER_141_321 ();
 FILLCELL_X16 FILLER_141_353 ();
 FILLCELL_X8 FILLER_141_369 ();
 FILLCELL_X2 FILLER_141_377 ();
 FILLCELL_X1 FILLER_141_379 ();
 FILLCELL_X32 FILLER_141_1518 ();
 FILLCELL_X32 FILLER_141_1550 ();
 FILLCELL_X32 FILLER_141_1582 ();
 FILLCELL_X32 FILLER_141_1614 ();
 FILLCELL_X32 FILLER_141_1646 ();
 FILLCELL_X32 FILLER_141_1678 ();
 FILLCELL_X32 FILLER_141_1710 ();
 FILLCELL_X8 FILLER_141_1742 ();
 FILLCELL_X4 FILLER_141_1750 ();
 FILLCELL_X2 FILLER_141_1754 ();
 FILLCELL_X32 FILLER_142_1 ();
 FILLCELL_X32 FILLER_142_33 ();
 FILLCELL_X32 FILLER_142_65 ();
 FILLCELL_X32 FILLER_142_97 ();
 FILLCELL_X32 FILLER_142_129 ();
 FILLCELL_X32 FILLER_142_161 ();
 FILLCELL_X32 FILLER_142_193 ();
 FILLCELL_X32 FILLER_142_225 ();
 FILLCELL_X32 FILLER_142_257 ();
 FILLCELL_X32 FILLER_142_289 ();
 FILLCELL_X32 FILLER_142_321 ();
 FILLCELL_X16 FILLER_142_353 ();
 FILLCELL_X8 FILLER_142_369 ();
 FILLCELL_X2 FILLER_142_377 ();
 FILLCELL_X1 FILLER_142_379 ();
 FILLCELL_X32 FILLER_142_1518 ();
 FILLCELL_X32 FILLER_142_1550 ();
 FILLCELL_X32 FILLER_142_1582 ();
 FILLCELL_X32 FILLER_142_1614 ();
 FILLCELL_X32 FILLER_142_1646 ();
 FILLCELL_X32 FILLER_142_1678 ();
 FILLCELL_X32 FILLER_142_1710 ();
 FILLCELL_X8 FILLER_142_1742 ();
 FILLCELL_X4 FILLER_142_1750 ();
 FILLCELL_X2 FILLER_142_1754 ();
 FILLCELL_X32 FILLER_143_1 ();
 FILLCELL_X32 FILLER_143_33 ();
 FILLCELL_X32 FILLER_143_65 ();
 FILLCELL_X32 FILLER_143_97 ();
 FILLCELL_X32 FILLER_143_129 ();
 FILLCELL_X32 FILLER_143_161 ();
 FILLCELL_X32 FILLER_143_193 ();
 FILLCELL_X32 FILLER_143_225 ();
 FILLCELL_X32 FILLER_143_257 ();
 FILLCELL_X32 FILLER_143_289 ();
 FILLCELL_X32 FILLER_143_321 ();
 FILLCELL_X16 FILLER_143_353 ();
 FILLCELL_X8 FILLER_143_369 ();
 FILLCELL_X2 FILLER_143_377 ();
 FILLCELL_X1 FILLER_143_379 ();
 FILLCELL_X32 FILLER_143_1518 ();
 FILLCELL_X32 FILLER_143_1550 ();
 FILLCELL_X32 FILLER_143_1582 ();
 FILLCELL_X32 FILLER_143_1614 ();
 FILLCELL_X32 FILLER_143_1646 ();
 FILLCELL_X32 FILLER_143_1678 ();
 FILLCELL_X32 FILLER_143_1710 ();
 FILLCELL_X8 FILLER_143_1742 ();
 FILLCELL_X4 FILLER_143_1750 ();
 FILLCELL_X2 FILLER_143_1754 ();
 FILLCELL_X32 FILLER_144_1 ();
 FILLCELL_X32 FILLER_144_33 ();
 FILLCELL_X32 FILLER_144_65 ();
 FILLCELL_X32 FILLER_144_97 ();
 FILLCELL_X32 FILLER_144_129 ();
 FILLCELL_X32 FILLER_144_161 ();
 FILLCELL_X32 FILLER_144_193 ();
 FILLCELL_X32 FILLER_144_225 ();
 FILLCELL_X32 FILLER_144_257 ();
 FILLCELL_X32 FILLER_144_289 ();
 FILLCELL_X32 FILLER_144_321 ();
 FILLCELL_X16 FILLER_144_353 ();
 FILLCELL_X8 FILLER_144_369 ();
 FILLCELL_X2 FILLER_144_377 ();
 FILLCELL_X1 FILLER_144_379 ();
 FILLCELL_X32 FILLER_144_1518 ();
 FILLCELL_X32 FILLER_144_1550 ();
 FILLCELL_X32 FILLER_144_1582 ();
 FILLCELL_X32 FILLER_144_1614 ();
 FILLCELL_X32 FILLER_144_1646 ();
 FILLCELL_X32 FILLER_144_1678 ();
 FILLCELL_X32 FILLER_144_1710 ();
 FILLCELL_X8 FILLER_144_1742 ();
 FILLCELL_X4 FILLER_144_1750 ();
 FILLCELL_X2 FILLER_144_1754 ();
 FILLCELL_X32 FILLER_145_1 ();
 FILLCELL_X32 FILLER_145_33 ();
 FILLCELL_X32 FILLER_145_65 ();
 FILLCELL_X32 FILLER_145_97 ();
 FILLCELL_X32 FILLER_145_129 ();
 FILLCELL_X32 FILLER_145_161 ();
 FILLCELL_X32 FILLER_145_193 ();
 FILLCELL_X32 FILLER_145_225 ();
 FILLCELL_X32 FILLER_145_257 ();
 FILLCELL_X32 FILLER_145_289 ();
 FILLCELL_X32 FILLER_145_321 ();
 FILLCELL_X16 FILLER_145_353 ();
 FILLCELL_X8 FILLER_145_369 ();
 FILLCELL_X2 FILLER_145_377 ();
 FILLCELL_X1 FILLER_145_379 ();
 FILLCELL_X32 FILLER_145_1518 ();
 FILLCELL_X32 FILLER_145_1550 ();
 FILLCELL_X32 FILLER_145_1582 ();
 FILLCELL_X32 FILLER_145_1614 ();
 FILLCELL_X32 FILLER_145_1646 ();
 FILLCELL_X32 FILLER_145_1678 ();
 FILLCELL_X32 FILLER_145_1710 ();
 FILLCELL_X4 FILLER_145_1742 ();
 FILLCELL_X2 FILLER_145_1746 ();
 FILLCELL_X1 FILLER_145_1748 ();
 FILLCELL_X4 FILLER_145_1752 ();
 FILLCELL_X32 FILLER_146_1 ();
 FILLCELL_X32 FILLER_146_33 ();
 FILLCELL_X32 FILLER_146_65 ();
 FILLCELL_X32 FILLER_146_97 ();
 FILLCELL_X32 FILLER_146_129 ();
 FILLCELL_X32 FILLER_146_161 ();
 FILLCELL_X32 FILLER_146_193 ();
 FILLCELL_X32 FILLER_146_225 ();
 FILLCELL_X32 FILLER_146_257 ();
 FILLCELL_X32 FILLER_146_289 ();
 FILLCELL_X32 FILLER_146_321 ();
 FILLCELL_X16 FILLER_146_353 ();
 FILLCELL_X8 FILLER_146_369 ();
 FILLCELL_X2 FILLER_146_377 ();
 FILLCELL_X1 FILLER_146_379 ();
 FILLCELL_X32 FILLER_146_1518 ();
 FILLCELL_X32 FILLER_146_1550 ();
 FILLCELL_X32 FILLER_146_1582 ();
 FILLCELL_X32 FILLER_146_1614 ();
 FILLCELL_X32 FILLER_146_1646 ();
 FILLCELL_X32 FILLER_146_1678 ();
 FILLCELL_X32 FILLER_146_1710 ();
 FILLCELL_X8 FILLER_146_1742 ();
 FILLCELL_X4 FILLER_146_1750 ();
 FILLCELL_X2 FILLER_146_1754 ();
 FILLCELL_X32 FILLER_147_1 ();
 FILLCELL_X32 FILLER_147_33 ();
 FILLCELL_X32 FILLER_147_65 ();
 FILLCELL_X32 FILLER_147_97 ();
 FILLCELL_X32 FILLER_147_129 ();
 FILLCELL_X32 FILLER_147_161 ();
 FILLCELL_X32 FILLER_147_193 ();
 FILLCELL_X32 FILLER_147_225 ();
 FILLCELL_X32 FILLER_147_257 ();
 FILLCELL_X32 FILLER_147_289 ();
 FILLCELL_X32 FILLER_147_321 ();
 FILLCELL_X16 FILLER_147_353 ();
 FILLCELL_X8 FILLER_147_369 ();
 FILLCELL_X2 FILLER_147_377 ();
 FILLCELL_X1 FILLER_147_379 ();
 FILLCELL_X32 FILLER_147_1518 ();
 FILLCELL_X32 FILLER_147_1550 ();
 FILLCELL_X32 FILLER_147_1582 ();
 FILLCELL_X32 FILLER_147_1614 ();
 FILLCELL_X32 FILLER_147_1646 ();
 FILLCELL_X32 FILLER_147_1678 ();
 FILLCELL_X32 FILLER_147_1710 ();
 FILLCELL_X8 FILLER_147_1742 ();
 FILLCELL_X4 FILLER_147_1750 ();
 FILLCELL_X2 FILLER_147_1754 ();
 FILLCELL_X32 FILLER_148_1 ();
 FILLCELL_X32 FILLER_148_33 ();
 FILLCELL_X32 FILLER_148_65 ();
 FILLCELL_X32 FILLER_148_97 ();
 FILLCELL_X32 FILLER_148_129 ();
 FILLCELL_X32 FILLER_148_161 ();
 FILLCELL_X32 FILLER_148_193 ();
 FILLCELL_X32 FILLER_148_225 ();
 FILLCELL_X32 FILLER_148_257 ();
 FILLCELL_X32 FILLER_148_289 ();
 FILLCELL_X32 FILLER_148_321 ();
 FILLCELL_X16 FILLER_148_353 ();
 FILLCELL_X8 FILLER_148_369 ();
 FILLCELL_X2 FILLER_148_377 ();
 FILLCELL_X1 FILLER_148_379 ();
 FILLCELL_X32 FILLER_148_1518 ();
 FILLCELL_X32 FILLER_148_1550 ();
 FILLCELL_X32 FILLER_148_1582 ();
 FILLCELL_X32 FILLER_148_1614 ();
 FILLCELL_X32 FILLER_148_1646 ();
 FILLCELL_X32 FILLER_148_1678 ();
 FILLCELL_X32 FILLER_148_1710 ();
 FILLCELL_X8 FILLER_148_1742 ();
 FILLCELL_X4 FILLER_148_1750 ();
 FILLCELL_X2 FILLER_148_1754 ();
 FILLCELL_X32 FILLER_149_1 ();
 FILLCELL_X32 FILLER_149_33 ();
 FILLCELL_X32 FILLER_149_65 ();
 FILLCELL_X32 FILLER_149_97 ();
 FILLCELL_X32 FILLER_149_129 ();
 FILLCELL_X32 FILLER_149_161 ();
 FILLCELL_X32 FILLER_149_193 ();
 FILLCELL_X32 FILLER_149_225 ();
 FILLCELL_X32 FILLER_149_257 ();
 FILLCELL_X32 FILLER_149_289 ();
 FILLCELL_X32 FILLER_149_321 ();
 FILLCELL_X16 FILLER_149_353 ();
 FILLCELL_X8 FILLER_149_369 ();
 FILLCELL_X2 FILLER_149_377 ();
 FILLCELL_X1 FILLER_149_379 ();
 FILLCELL_X32 FILLER_149_1518 ();
 FILLCELL_X32 FILLER_149_1550 ();
 FILLCELL_X32 FILLER_149_1582 ();
 FILLCELL_X32 FILLER_149_1614 ();
 FILLCELL_X32 FILLER_149_1646 ();
 FILLCELL_X32 FILLER_149_1678 ();
 FILLCELL_X32 FILLER_149_1710 ();
 FILLCELL_X8 FILLER_149_1742 ();
 FILLCELL_X4 FILLER_149_1750 ();
 FILLCELL_X2 FILLER_149_1754 ();
 FILLCELL_X4 FILLER_150_1 ();
 FILLCELL_X32 FILLER_150_9 ();
 FILLCELL_X32 FILLER_150_41 ();
 FILLCELL_X32 FILLER_150_73 ();
 FILLCELL_X32 FILLER_150_105 ();
 FILLCELL_X32 FILLER_150_137 ();
 FILLCELL_X32 FILLER_150_169 ();
 FILLCELL_X32 FILLER_150_201 ();
 FILLCELL_X32 FILLER_150_233 ();
 FILLCELL_X32 FILLER_150_265 ();
 FILLCELL_X32 FILLER_150_297 ();
 FILLCELL_X32 FILLER_150_329 ();
 FILLCELL_X16 FILLER_150_361 ();
 FILLCELL_X2 FILLER_150_377 ();
 FILLCELL_X1 FILLER_150_379 ();
 FILLCELL_X32 FILLER_150_1518 ();
 FILLCELL_X32 FILLER_150_1550 ();
 FILLCELL_X32 FILLER_150_1582 ();
 FILLCELL_X32 FILLER_150_1614 ();
 FILLCELL_X32 FILLER_150_1646 ();
 FILLCELL_X32 FILLER_150_1678 ();
 FILLCELL_X32 FILLER_150_1710 ();
 FILLCELL_X8 FILLER_150_1742 ();
 FILLCELL_X4 FILLER_150_1750 ();
 FILLCELL_X2 FILLER_150_1754 ();
 FILLCELL_X32 FILLER_151_1 ();
 FILLCELL_X32 FILLER_151_33 ();
 FILLCELL_X32 FILLER_151_65 ();
 FILLCELL_X32 FILLER_151_97 ();
 FILLCELL_X32 FILLER_151_129 ();
 FILLCELL_X32 FILLER_151_161 ();
 FILLCELL_X32 FILLER_151_193 ();
 FILLCELL_X32 FILLER_151_225 ();
 FILLCELL_X32 FILLER_151_257 ();
 FILLCELL_X32 FILLER_151_289 ();
 FILLCELL_X32 FILLER_151_321 ();
 FILLCELL_X16 FILLER_151_353 ();
 FILLCELL_X8 FILLER_151_369 ();
 FILLCELL_X2 FILLER_151_377 ();
 FILLCELL_X1 FILLER_151_379 ();
 FILLCELL_X32 FILLER_151_1518 ();
 FILLCELL_X32 FILLER_151_1550 ();
 FILLCELL_X32 FILLER_151_1582 ();
 FILLCELL_X32 FILLER_151_1614 ();
 FILLCELL_X32 FILLER_151_1646 ();
 FILLCELL_X32 FILLER_151_1678 ();
 FILLCELL_X32 FILLER_151_1710 ();
 FILLCELL_X8 FILLER_151_1742 ();
 FILLCELL_X4 FILLER_151_1750 ();
 FILLCELL_X2 FILLER_151_1754 ();
 FILLCELL_X32 FILLER_152_1 ();
 FILLCELL_X32 FILLER_152_33 ();
 FILLCELL_X32 FILLER_152_65 ();
 FILLCELL_X32 FILLER_152_97 ();
 FILLCELL_X32 FILLER_152_129 ();
 FILLCELL_X32 FILLER_152_161 ();
 FILLCELL_X32 FILLER_152_193 ();
 FILLCELL_X32 FILLER_152_225 ();
 FILLCELL_X32 FILLER_152_257 ();
 FILLCELL_X32 FILLER_152_289 ();
 FILLCELL_X32 FILLER_152_321 ();
 FILLCELL_X16 FILLER_152_353 ();
 FILLCELL_X8 FILLER_152_369 ();
 FILLCELL_X2 FILLER_152_377 ();
 FILLCELL_X1 FILLER_152_379 ();
 FILLCELL_X32 FILLER_152_1518 ();
 FILLCELL_X32 FILLER_152_1550 ();
 FILLCELL_X32 FILLER_152_1582 ();
 FILLCELL_X32 FILLER_152_1614 ();
 FILLCELL_X32 FILLER_152_1646 ();
 FILLCELL_X32 FILLER_152_1678 ();
 FILLCELL_X32 FILLER_152_1710 ();
 FILLCELL_X8 FILLER_152_1742 ();
 FILLCELL_X4 FILLER_152_1750 ();
 FILLCELL_X2 FILLER_152_1754 ();
 FILLCELL_X32 FILLER_153_1 ();
 FILLCELL_X32 FILLER_153_33 ();
 FILLCELL_X32 FILLER_153_65 ();
 FILLCELL_X32 FILLER_153_97 ();
 FILLCELL_X32 FILLER_153_129 ();
 FILLCELL_X32 FILLER_153_161 ();
 FILLCELL_X32 FILLER_153_193 ();
 FILLCELL_X32 FILLER_153_225 ();
 FILLCELL_X32 FILLER_153_257 ();
 FILLCELL_X32 FILLER_153_289 ();
 FILLCELL_X32 FILLER_153_321 ();
 FILLCELL_X16 FILLER_153_353 ();
 FILLCELL_X8 FILLER_153_369 ();
 FILLCELL_X2 FILLER_153_377 ();
 FILLCELL_X1 FILLER_153_379 ();
 FILLCELL_X32 FILLER_153_1518 ();
 FILLCELL_X32 FILLER_153_1550 ();
 FILLCELL_X32 FILLER_153_1582 ();
 FILLCELL_X32 FILLER_153_1614 ();
 FILLCELL_X32 FILLER_153_1646 ();
 FILLCELL_X32 FILLER_153_1678 ();
 FILLCELL_X32 FILLER_153_1710 ();
 FILLCELL_X8 FILLER_153_1742 ();
 FILLCELL_X4 FILLER_153_1750 ();
 FILLCELL_X2 FILLER_153_1754 ();
 FILLCELL_X32 FILLER_154_1 ();
 FILLCELL_X32 FILLER_154_33 ();
 FILLCELL_X32 FILLER_154_65 ();
 FILLCELL_X32 FILLER_154_97 ();
 FILLCELL_X32 FILLER_154_129 ();
 FILLCELL_X32 FILLER_154_161 ();
 FILLCELL_X32 FILLER_154_193 ();
 FILLCELL_X32 FILLER_154_225 ();
 FILLCELL_X32 FILLER_154_257 ();
 FILLCELL_X32 FILLER_154_289 ();
 FILLCELL_X32 FILLER_154_321 ();
 FILLCELL_X16 FILLER_154_353 ();
 FILLCELL_X8 FILLER_154_369 ();
 FILLCELL_X2 FILLER_154_377 ();
 FILLCELL_X1 FILLER_154_379 ();
 FILLCELL_X32 FILLER_154_1518 ();
 FILLCELL_X32 FILLER_154_1550 ();
 FILLCELL_X32 FILLER_154_1582 ();
 FILLCELL_X32 FILLER_154_1614 ();
 FILLCELL_X32 FILLER_154_1646 ();
 FILLCELL_X32 FILLER_154_1678 ();
 FILLCELL_X32 FILLER_154_1710 ();
 FILLCELL_X4 FILLER_154_1742 ();
 FILLCELL_X2 FILLER_154_1746 ();
 FILLCELL_X1 FILLER_154_1748 ();
 FILLCELL_X4 FILLER_154_1752 ();
 FILLCELL_X32 FILLER_155_1 ();
 FILLCELL_X32 FILLER_155_33 ();
 FILLCELL_X32 FILLER_155_65 ();
 FILLCELL_X32 FILLER_155_97 ();
 FILLCELL_X32 FILLER_155_129 ();
 FILLCELL_X32 FILLER_155_161 ();
 FILLCELL_X32 FILLER_155_193 ();
 FILLCELL_X32 FILLER_155_225 ();
 FILLCELL_X32 FILLER_155_257 ();
 FILLCELL_X32 FILLER_155_289 ();
 FILLCELL_X32 FILLER_155_321 ();
 FILLCELL_X16 FILLER_155_353 ();
 FILLCELL_X8 FILLER_155_369 ();
 FILLCELL_X2 FILLER_155_377 ();
 FILLCELL_X1 FILLER_155_379 ();
 FILLCELL_X32 FILLER_155_1518 ();
 FILLCELL_X32 FILLER_155_1550 ();
 FILLCELL_X32 FILLER_155_1582 ();
 FILLCELL_X32 FILLER_155_1614 ();
 FILLCELL_X32 FILLER_155_1646 ();
 FILLCELL_X32 FILLER_155_1678 ();
 FILLCELL_X32 FILLER_155_1710 ();
 FILLCELL_X8 FILLER_155_1742 ();
 FILLCELL_X4 FILLER_155_1750 ();
 FILLCELL_X2 FILLER_155_1754 ();
 FILLCELL_X32 FILLER_156_1 ();
 FILLCELL_X32 FILLER_156_33 ();
 FILLCELL_X32 FILLER_156_65 ();
 FILLCELL_X32 FILLER_156_97 ();
 FILLCELL_X32 FILLER_156_129 ();
 FILLCELL_X32 FILLER_156_161 ();
 FILLCELL_X32 FILLER_156_193 ();
 FILLCELL_X32 FILLER_156_225 ();
 FILLCELL_X32 FILLER_156_257 ();
 FILLCELL_X32 FILLER_156_289 ();
 FILLCELL_X32 FILLER_156_321 ();
 FILLCELL_X16 FILLER_156_353 ();
 FILLCELL_X8 FILLER_156_369 ();
 FILLCELL_X2 FILLER_156_377 ();
 FILLCELL_X1 FILLER_156_379 ();
 FILLCELL_X32 FILLER_156_1518 ();
 FILLCELL_X32 FILLER_156_1550 ();
 FILLCELL_X32 FILLER_156_1582 ();
 FILLCELL_X32 FILLER_156_1614 ();
 FILLCELL_X32 FILLER_156_1646 ();
 FILLCELL_X32 FILLER_156_1678 ();
 FILLCELL_X32 FILLER_156_1710 ();
 FILLCELL_X8 FILLER_156_1742 ();
 FILLCELL_X4 FILLER_156_1750 ();
 FILLCELL_X2 FILLER_156_1754 ();
 FILLCELL_X32 FILLER_157_1 ();
 FILLCELL_X32 FILLER_157_33 ();
 FILLCELL_X32 FILLER_157_65 ();
 FILLCELL_X32 FILLER_157_97 ();
 FILLCELL_X32 FILLER_157_129 ();
 FILLCELL_X32 FILLER_157_161 ();
 FILLCELL_X32 FILLER_157_193 ();
 FILLCELL_X32 FILLER_157_225 ();
 FILLCELL_X32 FILLER_157_257 ();
 FILLCELL_X32 FILLER_157_289 ();
 FILLCELL_X32 FILLER_157_321 ();
 FILLCELL_X16 FILLER_157_353 ();
 FILLCELL_X8 FILLER_157_369 ();
 FILLCELL_X2 FILLER_157_377 ();
 FILLCELL_X1 FILLER_157_379 ();
 FILLCELL_X32 FILLER_157_1518 ();
 FILLCELL_X32 FILLER_157_1550 ();
 FILLCELL_X32 FILLER_157_1582 ();
 FILLCELL_X32 FILLER_157_1614 ();
 FILLCELL_X32 FILLER_157_1646 ();
 FILLCELL_X32 FILLER_157_1678 ();
 FILLCELL_X32 FILLER_157_1710 ();
 FILLCELL_X8 FILLER_157_1742 ();
 FILLCELL_X4 FILLER_157_1750 ();
 FILLCELL_X2 FILLER_157_1754 ();
 FILLCELL_X32 FILLER_158_1 ();
 FILLCELL_X32 FILLER_158_33 ();
 FILLCELL_X32 FILLER_158_65 ();
 FILLCELL_X32 FILLER_158_97 ();
 FILLCELL_X32 FILLER_158_129 ();
 FILLCELL_X32 FILLER_158_161 ();
 FILLCELL_X32 FILLER_158_193 ();
 FILLCELL_X32 FILLER_158_225 ();
 FILLCELL_X32 FILLER_158_257 ();
 FILLCELL_X32 FILLER_158_289 ();
 FILLCELL_X32 FILLER_158_321 ();
 FILLCELL_X16 FILLER_158_353 ();
 FILLCELL_X8 FILLER_158_369 ();
 FILLCELL_X2 FILLER_158_377 ();
 FILLCELL_X1 FILLER_158_379 ();
 FILLCELL_X32 FILLER_158_1518 ();
 FILLCELL_X32 FILLER_158_1550 ();
 FILLCELL_X32 FILLER_158_1582 ();
 FILLCELL_X32 FILLER_158_1614 ();
 FILLCELL_X32 FILLER_158_1646 ();
 FILLCELL_X32 FILLER_158_1678 ();
 FILLCELL_X32 FILLER_158_1710 ();
 FILLCELL_X8 FILLER_158_1742 ();
 FILLCELL_X4 FILLER_158_1750 ();
 FILLCELL_X2 FILLER_158_1754 ();
 FILLCELL_X4 FILLER_159_1 ();
 FILLCELL_X32 FILLER_159_9 ();
 FILLCELL_X32 FILLER_159_41 ();
 FILLCELL_X32 FILLER_159_73 ();
 FILLCELL_X32 FILLER_159_105 ();
 FILLCELL_X32 FILLER_159_137 ();
 FILLCELL_X32 FILLER_159_169 ();
 FILLCELL_X32 FILLER_159_201 ();
 FILLCELL_X32 FILLER_159_233 ();
 FILLCELL_X32 FILLER_159_265 ();
 FILLCELL_X32 FILLER_159_297 ();
 FILLCELL_X32 FILLER_159_329 ();
 FILLCELL_X16 FILLER_159_361 ();
 FILLCELL_X2 FILLER_159_377 ();
 FILLCELL_X1 FILLER_159_379 ();
 FILLCELL_X32 FILLER_159_1518 ();
 FILLCELL_X32 FILLER_159_1550 ();
 FILLCELL_X32 FILLER_159_1582 ();
 FILLCELL_X32 FILLER_159_1614 ();
 FILLCELL_X32 FILLER_159_1646 ();
 FILLCELL_X32 FILLER_159_1678 ();
 FILLCELL_X32 FILLER_159_1710 ();
 FILLCELL_X8 FILLER_159_1742 ();
 FILLCELL_X4 FILLER_159_1750 ();
 FILLCELL_X2 FILLER_159_1754 ();
 FILLCELL_X32 FILLER_160_1 ();
 FILLCELL_X32 FILLER_160_33 ();
 FILLCELL_X32 FILLER_160_65 ();
 FILLCELL_X32 FILLER_160_97 ();
 FILLCELL_X32 FILLER_160_129 ();
 FILLCELL_X32 FILLER_160_161 ();
 FILLCELL_X32 FILLER_160_193 ();
 FILLCELL_X32 FILLER_160_225 ();
 FILLCELL_X32 FILLER_160_257 ();
 FILLCELL_X32 FILLER_160_289 ();
 FILLCELL_X32 FILLER_160_321 ();
 FILLCELL_X16 FILLER_160_353 ();
 FILLCELL_X8 FILLER_160_369 ();
 FILLCELL_X2 FILLER_160_377 ();
 FILLCELL_X1 FILLER_160_379 ();
 FILLCELL_X32 FILLER_160_1518 ();
 FILLCELL_X32 FILLER_160_1550 ();
 FILLCELL_X32 FILLER_160_1582 ();
 FILLCELL_X32 FILLER_160_1614 ();
 FILLCELL_X32 FILLER_160_1646 ();
 FILLCELL_X32 FILLER_160_1678 ();
 FILLCELL_X32 FILLER_160_1710 ();
 FILLCELL_X8 FILLER_160_1742 ();
 FILLCELL_X4 FILLER_160_1750 ();
 FILLCELL_X2 FILLER_160_1754 ();
 FILLCELL_X32 FILLER_161_1 ();
 FILLCELL_X32 FILLER_161_33 ();
 FILLCELL_X32 FILLER_161_65 ();
 FILLCELL_X32 FILLER_161_97 ();
 FILLCELL_X32 FILLER_161_129 ();
 FILLCELL_X32 FILLER_161_161 ();
 FILLCELL_X32 FILLER_161_193 ();
 FILLCELL_X32 FILLER_161_225 ();
 FILLCELL_X32 FILLER_161_257 ();
 FILLCELL_X32 FILLER_161_289 ();
 FILLCELL_X32 FILLER_161_321 ();
 FILLCELL_X16 FILLER_161_353 ();
 FILLCELL_X8 FILLER_161_369 ();
 FILLCELL_X2 FILLER_161_377 ();
 FILLCELL_X1 FILLER_161_379 ();
 FILLCELL_X32 FILLER_161_1518 ();
 FILLCELL_X32 FILLER_161_1550 ();
 FILLCELL_X32 FILLER_161_1582 ();
 FILLCELL_X32 FILLER_161_1614 ();
 FILLCELL_X32 FILLER_161_1646 ();
 FILLCELL_X32 FILLER_161_1678 ();
 FILLCELL_X32 FILLER_161_1710 ();
 FILLCELL_X8 FILLER_161_1742 ();
 FILLCELL_X4 FILLER_161_1750 ();
 FILLCELL_X2 FILLER_161_1754 ();
 FILLCELL_X32 FILLER_162_1 ();
 FILLCELL_X32 FILLER_162_33 ();
 FILLCELL_X32 FILLER_162_65 ();
 FILLCELL_X32 FILLER_162_97 ();
 FILLCELL_X32 FILLER_162_129 ();
 FILLCELL_X32 FILLER_162_161 ();
 FILLCELL_X32 FILLER_162_193 ();
 FILLCELL_X32 FILLER_162_225 ();
 FILLCELL_X32 FILLER_162_257 ();
 FILLCELL_X32 FILLER_162_289 ();
 FILLCELL_X32 FILLER_162_321 ();
 FILLCELL_X16 FILLER_162_353 ();
 FILLCELL_X8 FILLER_162_369 ();
 FILLCELL_X2 FILLER_162_377 ();
 FILLCELL_X1 FILLER_162_379 ();
 FILLCELL_X32 FILLER_162_1518 ();
 FILLCELL_X32 FILLER_162_1550 ();
 FILLCELL_X32 FILLER_162_1582 ();
 FILLCELL_X32 FILLER_162_1614 ();
 FILLCELL_X32 FILLER_162_1646 ();
 FILLCELL_X32 FILLER_162_1678 ();
 FILLCELL_X32 FILLER_162_1710 ();
 FILLCELL_X8 FILLER_162_1742 ();
 FILLCELL_X4 FILLER_162_1750 ();
 FILLCELL_X2 FILLER_162_1754 ();
 FILLCELL_X32 FILLER_163_1 ();
 FILLCELL_X32 FILLER_163_33 ();
 FILLCELL_X32 FILLER_163_65 ();
 FILLCELL_X32 FILLER_163_97 ();
 FILLCELL_X32 FILLER_163_129 ();
 FILLCELL_X32 FILLER_163_161 ();
 FILLCELL_X32 FILLER_163_193 ();
 FILLCELL_X32 FILLER_163_225 ();
 FILLCELL_X32 FILLER_163_257 ();
 FILLCELL_X32 FILLER_163_289 ();
 FILLCELL_X32 FILLER_163_321 ();
 FILLCELL_X16 FILLER_163_353 ();
 FILLCELL_X8 FILLER_163_369 ();
 FILLCELL_X2 FILLER_163_377 ();
 FILLCELL_X1 FILLER_163_379 ();
 FILLCELL_X32 FILLER_163_1518 ();
 FILLCELL_X32 FILLER_163_1550 ();
 FILLCELL_X32 FILLER_163_1582 ();
 FILLCELL_X32 FILLER_163_1614 ();
 FILLCELL_X32 FILLER_163_1646 ();
 FILLCELL_X32 FILLER_163_1678 ();
 FILLCELL_X32 FILLER_163_1710 ();
 FILLCELL_X8 FILLER_163_1742 ();
 FILLCELL_X4 FILLER_163_1750 ();
 FILLCELL_X2 FILLER_163_1754 ();
 FILLCELL_X32 FILLER_164_1 ();
 FILLCELL_X32 FILLER_164_33 ();
 FILLCELL_X32 FILLER_164_65 ();
 FILLCELL_X32 FILLER_164_97 ();
 FILLCELL_X32 FILLER_164_129 ();
 FILLCELL_X32 FILLER_164_161 ();
 FILLCELL_X32 FILLER_164_193 ();
 FILLCELL_X32 FILLER_164_225 ();
 FILLCELL_X32 FILLER_164_257 ();
 FILLCELL_X32 FILLER_164_289 ();
 FILLCELL_X32 FILLER_164_321 ();
 FILLCELL_X16 FILLER_164_353 ();
 FILLCELL_X8 FILLER_164_369 ();
 FILLCELL_X2 FILLER_164_377 ();
 FILLCELL_X1 FILLER_164_379 ();
 FILLCELL_X32 FILLER_164_1518 ();
 FILLCELL_X32 FILLER_164_1550 ();
 FILLCELL_X32 FILLER_164_1582 ();
 FILLCELL_X32 FILLER_164_1614 ();
 FILLCELL_X32 FILLER_164_1646 ();
 FILLCELL_X32 FILLER_164_1678 ();
 FILLCELL_X32 FILLER_164_1710 ();
 FILLCELL_X4 FILLER_164_1742 ();
 FILLCELL_X2 FILLER_164_1746 ();
 FILLCELL_X1 FILLER_164_1748 ();
 FILLCELL_X4 FILLER_164_1752 ();
 FILLCELL_X32 FILLER_165_1 ();
 FILLCELL_X32 FILLER_165_33 ();
 FILLCELL_X32 FILLER_165_65 ();
 FILLCELL_X32 FILLER_165_97 ();
 FILLCELL_X32 FILLER_165_129 ();
 FILLCELL_X32 FILLER_165_161 ();
 FILLCELL_X32 FILLER_165_193 ();
 FILLCELL_X32 FILLER_165_225 ();
 FILLCELL_X32 FILLER_165_257 ();
 FILLCELL_X32 FILLER_165_289 ();
 FILLCELL_X32 FILLER_165_321 ();
 FILLCELL_X16 FILLER_165_353 ();
 FILLCELL_X8 FILLER_165_369 ();
 FILLCELL_X2 FILLER_165_377 ();
 FILLCELL_X1 FILLER_165_379 ();
 FILLCELL_X32 FILLER_165_1518 ();
 FILLCELL_X32 FILLER_165_1550 ();
 FILLCELL_X32 FILLER_165_1582 ();
 FILLCELL_X32 FILLER_165_1614 ();
 FILLCELL_X32 FILLER_165_1646 ();
 FILLCELL_X32 FILLER_165_1678 ();
 FILLCELL_X32 FILLER_165_1710 ();
 FILLCELL_X8 FILLER_165_1742 ();
 FILLCELL_X4 FILLER_165_1750 ();
 FILLCELL_X2 FILLER_165_1754 ();
 FILLCELL_X32 FILLER_166_1 ();
 FILLCELL_X32 FILLER_166_33 ();
 FILLCELL_X32 FILLER_166_65 ();
 FILLCELL_X32 FILLER_166_97 ();
 FILLCELL_X32 FILLER_166_129 ();
 FILLCELL_X32 FILLER_166_161 ();
 FILLCELL_X32 FILLER_166_193 ();
 FILLCELL_X32 FILLER_166_225 ();
 FILLCELL_X32 FILLER_166_257 ();
 FILLCELL_X32 FILLER_166_289 ();
 FILLCELL_X32 FILLER_166_321 ();
 FILLCELL_X16 FILLER_166_353 ();
 FILLCELL_X8 FILLER_166_369 ();
 FILLCELL_X2 FILLER_166_377 ();
 FILLCELL_X1 FILLER_166_379 ();
 FILLCELL_X32 FILLER_166_1518 ();
 FILLCELL_X32 FILLER_166_1550 ();
 FILLCELL_X32 FILLER_166_1582 ();
 FILLCELL_X32 FILLER_166_1614 ();
 FILLCELL_X32 FILLER_166_1646 ();
 FILLCELL_X32 FILLER_166_1678 ();
 FILLCELL_X32 FILLER_166_1710 ();
 FILLCELL_X8 FILLER_166_1742 ();
 FILLCELL_X4 FILLER_166_1750 ();
 FILLCELL_X2 FILLER_166_1754 ();
 FILLCELL_X32 FILLER_167_1 ();
 FILLCELL_X32 FILLER_167_33 ();
 FILLCELL_X32 FILLER_167_65 ();
 FILLCELL_X32 FILLER_167_97 ();
 FILLCELL_X32 FILLER_167_129 ();
 FILLCELL_X32 FILLER_167_161 ();
 FILLCELL_X32 FILLER_167_193 ();
 FILLCELL_X32 FILLER_167_225 ();
 FILLCELL_X32 FILLER_167_257 ();
 FILLCELL_X32 FILLER_167_289 ();
 FILLCELL_X32 FILLER_167_321 ();
 FILLCELL_X16 FILLER_167_353 ();
 FILLCELL_X8 FILLER_167_369 ();
 FILLCELL_X2 FILLER_167_377 ();
 FILLCELL_X1 FILLER_167_379 ();
 FILLCELL_X32 FILLER_167_1518 ();
 FILLCELL_X32 FILLER_167_1550 ();
 FILLCELL_X32 FILLER_167_1582 ();
 FILLCELL_X32 FILLER_167_1614 ();
 FILLCELL_X32 FILLER_167_1646 ();
 FILLCELL_X32 FILLER_167_1678 ();
 FILLCELL_X32 FILLER_167_1710 ();
 FILLCELL_X8 FILLER_167_1742 ();
 FILLCELL_X4 FILLER_167_1750 ();
 FILLCELL_X2 FILLER_167_1754 ();
 FILLCELL_X32 FILLER_168_1 ();
 FILLCELL_X32 FILLER_168_33 ();
 FILLCELL_X32 FILLER_168_65 ();
 FILLCELL_X32 FILLER_168_97 ();
 FILLCELL_X32 FILLER_168_129 ();
 FILLCELL_X32 FILLER_168_161 ();
 FILLCELL_X32 FILLER_168_193 ();
 FILLCELL_X32 FILLER_168_225 ();
 FILLCELL_X32 FILLER_168_257 ();
 FILLCELL_X32 FILLER_168_289 ();
 FILLCELL_X32 FILLER_168_321 ();
 FILLCELL_X16 FILLER_168_353 ();
 FILLCELL_X8 FILLER_168_369 ();
 FILLCELL_X2 FILLER_168_377 ();
 FILLCELL_X1 FILLER_168_379 ();
 FILLCELL_X32 FILLER_168_1518 ();
 FILLCELL_X32 FILLER_168_1550 ();
 FILLCELL_X32 FILLER_168_1582 ();
 FILLCELL_X32 FILLER_168_1614 ();
 FILLCELL_X32 FILLER_168_1646 ();
 FILLCELL_X32 FILLER_168_1678 ();
 FILLCELL_X32 FILLER_168_1710 ();
 FILLCELL_X8 FILLER_168_1742 ();
 FILLCELL_X4 FILLER_168_1750 ();
 FILLCELL_X2 FILLER_168_1754 ();
 FILLCELL_X4 FILLER_169_1 ();
 FILLCELL_X32 FILLER_169_8 ();
 FILLCELL_X32 FILLER_169_40 ();
 FILLCELL_X32 FILLER_169_72 ();
 FILLCELL_X32 FILLER_169_104 ();
 FILLCELL_X32 FILLER_169_136 ();
 FILLCELL_X32 FILLER_169_168 ();
 FILLCELL_X32 FILLER_169_200 ();
 FILLCELL_X32 FILLER_169_232 ();
 FILLCELL_X32 FILLER_169_264 ();
 FILLCELL_X32 FILLER_169_296 ();
 FILLCELL_X32 FILLER_169_328 ();
 FILLCELL_X16 FILLER_169_360 ();
 FILLCELL_X4 FILLER_169_376 ();
 FILLCELL_X32 FILLER_169_1518 ();
 FILLCELL_X32 FILLER_169_1550 ();
 FILLCELL_X32 FILLER_169_1582 ();
 FILLCELL_X32 FILLER_169_1614 ();
 FILLCELL_X32 FILLER_169_1646 ();
 FILLCELL_X32 FILLER_169_1678 ();
 FILLCELL_X32 FILLER_169_1710 ();
 FILLCELL_X8 FILLER_169_1742 ();
 FILLCELL_X4 FILLER_169_1750 ();
 FILLCELL_X2 FILLER_169_1754 ();
 FILLCELL_X32 FILLER_170_1 ();
 FILLCELL_X32 FILLER_170_33 ();
 FILLCELL_X32 FILLER_170_65 ();
 FILLCELL_X32 FILLER_170_97 ();
 FILLCELL_X32 FILLER_170_129 ();
 FILLCELL_X32 FILLER_170_161 ();
 FILLCELL_X32 FILLER_170_193 ();
 FILLCELL_X32 FILLER_170_225 ();
 FILLCELL_X32 FILLER_170_257 ();
 FILLCELL_X32 FILLER_170_289 ();
 FILLCELL_X32 FILLER_170_321 ();
 FILLCELL_X16 FILLER_170_353 ();
 FILLCELL_X8 FILLER_170_369 ();
 FILLCELL_X2 FILLER_170_377 ();
 FILLCELL_X1 FILLER_170_379 ();
 FILLCELL_X32 FILLER_170_1518 ();
 FILLCELL_X32 FILLER_170_1550 ();
 FILLCELL_X32 FILLER_170_1582 ();
 FILLCELL_X32 FILLER_170_1614 ();
 FILLCELL_X32 FILLER_170_1646 ();
 FILLCELL_X32 FILLER_170_1678 ();
 FILLCELL_X32 FILLER_170_1710 ();
 FILLCELL_X8 FILLER_170_1742 ();
 FILLCELL_X4 FILLER_170_1750 ();
 FILLCELL_X2 FILLER_170_1754 ();
 FILLCELL_X32 FILLER_171_1 ();
 FILLCELL_X32 FILLER_171_33 ();
 FILLCELL_X32 FILLER_171_65 ();
 FILLCELL_X32 FILLER_171_97 ();
 FILLCELL_X32 FILLER_171_129 ();
 FILLCELL_X32 FILLER_171_161 ();
 FILLCELL_X32 FILLER_171_193 ();
 FILLCELL_X32 FILLER_171_225 ();
 FILLCELL_X32 FILLER_171_257 ();
 FILLCELL_X32 FILLER_171_289 ();
 FILLCELL_X32 FILLER_171_321 ();
 FILLCELL_X16 FILLER_171_353 ();
 FILLCELL_X8 FILLER_171_369 ();
 FILLCELL_X2 FILLER_171_377 ();
 FILLCELL_X1 FILLER_171_379 ();
 FILLCELL_X32 FILLER_171_1518 ();
 FILLCELL_X32 FILLER_171_1550 ();
 FILLCELL_X32 FILLER_171_1582 ();
 FILLCELL_X32 FILLER_171_1614 ();
 FILLCELL_X32 FILLER_171_1646 ();
 FILLCELL_X32 FILLER_171_1678 ();
 FILLCELL_X32 FILLER_171_1710 ();
 FILLCELL_X8 FILLER_171_1742 ();
 FILLCELL_X4 FILLER_171_1750 ();
 FILLCELL_X2 FILLER_171_1754 ();
 FILLCELL_X32 FILLER_172_1 ();
 FILLCELL_X32 FILLER_172_33 ();
 FILLCELL_X32 FILLER_172_65 ();
 FILLCELL_X32 FILLER_172_97 ();
 FILLCELL_X32 FILLER_172_129 ();
 FILLCELL_X32 FILLER_172_161 ();
 FILLCELL_X32 FILLER_172_193 ();
 FILLCELL_X32 FILLER_172_225 ();
 FILLCELL_X32 FILLER_172_257 ();
 FILLCELL_X32 FILLER_172_289 ();
 FILLCELL_X32 FILLER_172_321 ();
 FILLCELL_X16 FILLER_172_353 ();
 FILLCELL_X8 FILLER_172_369 ();
 FILLCELL_X2 FILLER_172_377 ();
 FILLCELL_X1 FILLER_172_379 ();
 FILLCELL_X32 FILLER_172_1518 ();
 FILLCELL_X32 FILLER_172_1550 ();
 FILLCELL_X32 FILLER_172_1582 ();
 FILLCELL_X32 FILLER_172_1614 ();
 FILLCELL_X32 FILLER_172_1646 ();
 FILLCELL_X32 FILLER_172_1678 ();
 FILLCELL_X32 FILLER_172_1710 ();
 FILLCELL_X8 FILLER_172_1742 ();
 FILLCELL_X4 FILLER_172_1750 ();
 FILLCELL_X2 FILLER_172_1754 ();
 FILLCELL_X32 FILLER_173_1 ();
 FILLCELL_X32 FILLER_173_33 ();
 FILLCELL_X32 FILLER_173_65 ();
 FILLCELL_X32 FILLER_173_97 ();
 FILLCELL_X32 FILLER_173_129 ();
 FILLCELL_X32 FILLER_173_161 ();
 FILLCELL_X32 FILLER_173_193 ();
 FILLCELL_X32 FILLER_173_225 ();
 FILLCELL_X32 FILLER_173_257 ();
 FILLCELL_X32 FILLER_173_289 ();
 FILLCELL_X32 FILLER_173_321 ();
 FILLCELL_X16 FILLER_173_353 ();
 FILLCELL_X8 FILLER_173_369 ();
 FILLCELL_X2 FILLER_173_377 ();
 FILLCELL_X1 FILLER_173_379 ();
 FILLCELL_X32 FILLER_173_1518 ();
 FILLCELL_X32 FILLER_173_1550 ();
 FILLCELL_X32 FILLER_173_1582 ();
 FILLCELL_X32 FILLER_173_1614 ();
 FILLCELL_X32 FILLER_173_1646 ();
 FILLCELL_X32 FILLER_173_1678 ();
 FILLCELL_X32 FILLER_173_1710 ();
 FILLCELL_X8 FILLER_173_1742 ();
 FILLCELL_X4 FILLER_173_1750 ();
 FILLCELL_X2 FILLER_173_1754 ();
 FILLCELL_X32 FILLER_174_1 ();
 FILLCELL_X32 FILLER_174_33 ();
 FILLCELL_X32 FILLER_174_65 ();
 FILLCELL_X32 FILLER_174_97 ();
 FILLCELL_X32 FILLER_174_129 ();
 FILLCELL_X32 FILLER_174_161 ();
 FILLCELL_X32 FILLER_174_193 ();
 FILLCELL_X32 FILLER_174_225 ();
 FILLCELL_X32 FILLER_174_257 ();
 FILLCELL_X32 FILLER_174_289 ();
 FILLCELL_X32 FILLER_174_321 ();
 FILLCELL_X16 FILLER_174_353 ();
 FILLCELL_X8 FILLER_174_369 ();
 FILLCELL_X2 FILLER_174_377 ();
 FILLCELL_X1 FILLER_174_379 ();
 FILLCELL_X32 FILLER_174_1518 ();
 FILLCELL_X32 FILLER_174_1550 ();
 FILLCELL_X32 FILLER_174_1582 ();
 FILLCELL_X32 FILLER_174_1614 ();
 FILLCELL_X32 FILLER_174_1646 ();
 FILLCELL_X32 FILLER_174_1678 ();
 FILLCELL_X32 FILLER_174_1710 ();
 FILLCELL_X2 FILLER_174_1742 ();
 FILLCELL_X1 FILLER_174_1744 ();
 FILLCELL_X4 FILLER_174_1752 ();
 FILLCELL_X32 FILLER_175_1 ();
 FILLCELL_X32 FILLER_175_33 ();
 FILLCELL_X32 FILLER_175_65 ();
 FILLCELL_X32 FILLER_175_97 ();
 FILLCELL_X32 FILLER_175_129 ();
 FILLCELL_X32 FILLER_175_161 ();
 FILLCELL_X32 FILLER_175_193 ();
 FILLCELL_X32 FILLER_175_225 ();
 FILLCELL_X32 FILLER_175_257 ();
 FILLCELL_X32 FILLER_175_289 ();
 FILLCELL_X32 FILLER_175_321 ();
 FILLCELL_X16 FILLER_175_353 ();
 FILLCELL_X8 FILLER_175_369 ();
 FILLCELL_X2 FILLER_175_377 ();
 FILLCELL_X1 FILLER_175_379 ();
 FILLCELL_X32 FILLER_175_1518 ();
 FILLCELL_X32 FILLER_175_1550 ();
 FILLCELL_X32 FILLER_175_1582 ();
 FILLCELL_X32 FILLER_175_1614 ();
 FILLCELL_X32 FILLER_175_1646 ();
 FILLCELL_X32 FILLER_175_1678 ();
 FILLCELL_X32 FILLER_175_1710 ();
 FILLCELL_X8 FILLER_175_1742 ();
 FILLCELL_X4 FILLER_175_1750 ();
 FILLCELL_X2 FILLER_175_1754 ();
 FILLCELL_X32 FILLER_176_1 ();
 FILLCELL_X32 FILLER_176_33 ();
 FILLCELL_X32 FILLER_176_65 ();
 FILLCELL_X32 FILLER_176_97 ();
 FILLCELL_X32 FILLER_176_129 ();
 FILLCELL_X32 FILLER_176_161 ();
 FILLCELL_X32 FILLER_176_193 ();
 FILLCELL_X32 FILLER_176_225 ();
 FILLCELL_X32 FILLER_176_257 ();
 FILLCELL_X32 FILLER_176_289 ();
 FILLCELL_X32 FILLER_176_321 ();
 FILLCELL_X16 FILLER_176_353 ();
 FILLCELL_X8 FILLER_176_369 ();
 FILLCELL_X2 FILLER_176_377 ();
 FILLCELL_X1 FILLER_176_379 ();
 FILLCELL_X32 FILLER_176_1518 ();
 FILLCELL_X32 FILLER_176_1550 ();
 FILLCELL_X32 FILLER_176_1582 ();
 FILLCELL_X32 FILLER_176_1614 ();
 FILLCELL_X32 FILLER_176_1646 ();
 FILLCELL_X32 FILLER_176_1678 ();
 FILLCELL_X32 FILLER_176_1710 ();
 FILLCELL_X8 FILLER_176_1742 ();
 FILLCELL_X4 FILLER_176_1750 ();
 FILLCELL_X2 FILLER_176_1754 ();
 FILLCELL_X32 FILLER_177_1 ();
 FILLCELL_X32 FILLER_177_33 ();
 FILLCELL_X32 FILLER_177_65 ();
 FILLCELL_X32 FILLER_177_97 ();
 FILLCELL_X32 FILLER_177_129 ();
 FILLCELL_X32 FILLER_177_161 ();
 FILLCELL_X32 FILLER_177_193 ();
 FILLCELL_X32 FILLER_177_225 ();
 FILLCELL_X32 FILLER_177_257 ();
 FILLCELL_X32 FILLER_177_289 ();
 FILLCELL_X32 FILLER_177_321 ();
 FILLCELL_X16 FILLER_177_353 ();
 FILLCELL_X8 FILLER_177_369 ();
 FILLCELL_X2 FILLER_177_377 ();
 FILLCELL_X1 FILLER_177_379 ();
 FILLCELL_X32 FILLER_177_1518 ();
 FILLCELL_X32 FILLER_177_1550 ();
 FILLCELL_X32 FILLER_177_1582 ();
 FILLCELL_X32 FILLER_177_1614 ();
 FILLCELL_X32 FILLER_177_1646 ();
 FILLCELL_X32 FILLER_177_1678 ();
 FILLCELL_X32 FILLER_177_1710 ();
 FILLCELL_X8 FILLER_177_1742 ();
 FILLCELL_X4 FILLER_177_1750 ();
 FILLCELL_X2 FILLER_177_1754 ();
 FILLCELL_X4 FILLER_178_1 ();
 FILLCELL_X32 FILLER_178_9 ();
 FILLCELL_X32 FILLER_178_41 ();
 FILLCELL_X32 FILLER_178_73 ();
 FILLCELL_X32 FILLER_178_105 ();
 FILLCELL_X32 FILLER_178_137 ();
 FILLCELL_X32 FILLER_178_169 ();
 FILLCELL_X32 FILLER_178_201 ();
 FILLCELL_X32 FILLER_178_233 ();
 FILLCELL_X32 FILLER_178_265 ();
 FILLCELL_X32 FILLER_178_297 ();
 FILLCELL_X32 FILLER_178_329 ();
 FILLCELL_X16 FILLER_178_361 ();
 FILLCELL_X2 FILLER_178_377 ();
 FILLCELL_X1 FILLER_178_379 ();
 FILLCELL_X32 FILLER_178_1518 ();
 FILLCELL_X32 FILLER_178_1550 ();
 FILLCELL_X32 FILLER_178_1582 ();
 FILLCELL_X32 FILLER_178_1614 ();
 FILLCELL_X32 FILLER_178_1646 ();
 FILLCELL_X32 FILLER_178_1678 ();
 FILLCELL_X32 FILLER_178_1710 ();
 FILLCELL_X8 FILLER_178_1742 ();
 FILLCELL_X4 FILLER_178_1750 ();
 FILLCELL_X2 FILLER_178_1754 ();
 FILLCELL_X32 FILLER_179_1 ();
 FILLCELL_X32 FILLER_179_33 ();
 FILLCELL_X32 FILLER_179_65 ();
 FILLCELL_X32 FILLER_179_97 ();
 FILLCELL_X32 FILLER_179_129 ();
 FILLCELL_X32 FILLER_179_161 ();
 FILLCELL_X32 FILLER_179_193 ();
 FILLCELL_X32 FILLER_179_225 ();
 FILLCELL_X32 FILLER_179_257 ();
 FILLCELL_X32 FILLER_179_289 ();
 FILLCELL_X32 FILLER_179_321 ();
 FILLCELL_X16 FILLER_179_353 ();
 FILLCELL_X8 FILLER_179_369 ();
 FILLCELL_X2 FILLER_179_377 ();
 FILLCELL_X1 FILLER_179_379 ();
 FILLCELL_X32 FILLER_179_1518 ();
 FILLCELL_X32 FILLER_179_1550 ();
 FILLCELL_X32 FILLER_179_1582 ();
 FILLCELL_X32 FILLER_179_1614 ();
 FILLCELL_X32 FILLER_179_1646 ();
 FILLCELL_X32 FILLER_179_1678 ();
 FILLCELL_X32 FILLER_179_1710 ();
 FILLCELL_X8 FILLER_179_1742 ();
 FILLCELL_X4 FILLER_179_1750 ();
 FILLCELL_X2 FILLER_179_1754 ();
 FILLCELL_X32 FILLER_180_1 ();
 FILLCELL_X32 FILLER_180_33 ();
 FILLCELL_X32 FILLER_180_65 ();
 FILLCELL_X32 FILLER_180_97 ();
 FILLCELL_X32 FILLER_180_129 ();
 FILLCELL_X32 FILLER_180_161 ();
 FILLCELL_X32 FILLER_180_193 ();
 FILLCELL_X32 FILLER_180_225 ();
 FILLCELL_X32 FILLER_180_257 ();
 FILLCELL_X32 FILLER_180_289 ();
 FILLCELL_X32 FILLER_180_321 ();
 FILLCELL_X16 FILLER_180_353 ();
 FILLCELL_X8 FILLER_180_369 ();
 FILLCELL_X2 FILLER_180_377 ();
 FILLCELL_X1 FILLER_180_379 ();
 FILLCELL_X32 FILLER_180_1518 ();
 FILLCELL_X32 FILLER_180_1550 ();
 FILLCELL_X32 FILLER_180_1582 ();
 FILLCELL_X32 FILLER_180_1614 ();
 FILLCELL_X32 FILLER_180_1646 ();
 FILLCELL_X32 FILLER_180_1678 ();
 FILLCELL_X32 FILLER_180_1710 ();
 FILLCELL_X8 FILLER_180_1742 ();
 FILLCELL_X4 FILLER_180_1750 ();
 FILLCELL_X2 FILLER_180_1754 ();
 FILLCELL_X32 FILLER_181_1 ();
 FILLCELL_X32 FILLER_181_33 ();
 FILLCELL_X32 FILLER_181_65 ();
 FILLCELL_X32 FILLER_181_97 ();
 FILLCELL_X32 FILLER_181_129 ();
 FILLCELL_X32 FILLER_181_161 ();
 FILLCELL_X32 FILLER_181_193 ();
 FILLCELL_X32 FILLER_181_225 ();
 FILLCELL_X32 FILLER_181_257 ();
 FILLCELL_X32 FILLER_181_289 ();
 FILLCELL_X32 FILLER_181_321 ();
 FILLCELL_X16 FILLER_181_353 ();
 FILLCELL_X8 FILLER_181_369 ();
 FILLCELL_X2 FILLER_181_377 ();
 FILLCELL_X1 FILLER_181_379 ();
 FILLCELL_X32 FILLER_181_1518 ();
 FILLCELL_X32 FILLER_181_1550 ();
 FILLCELL_X32 FILLER_181_1582 ();
 FILLCELL_X32 FILLER_181_1614 ();
 FILLCELL_X32 FILLER_181_1646 ();
 FILLCELL_X32 FILLER_181_1678 ();
 FILLCELL_X32 FILLER_181_1710 ();
 FILLCELL_X8 FILLER_181_1742 ();
 FILLCELL_X4 FILLER_181_1750 ();
 FILLCELL_X2 FILLER_181_1754 ();
 FILLCELL_X32 FILLER_182_1 ();
 FILLCELL_X32 FILLER_182_33 ();
 FILLCELL_X32 FILLER_182_65 ();
 FILLCELL_X32 FILLER_182_97 ();
 FILLCELL_X32 FILLER_182_129 ();
 FILLCELL_X32 FILLER_182_161 ();
 FILLCELL_X32 FILLER_182_193 ();
 FILLCELL_X32 FILLER_182_225 ();
 FILLCELL_X32 FILLER_182_257 ();
 FILLCELL_X32 FILLER_182_289 ();
 FILLCELL_X32 FILLER_182_321 ();
 FILLCELL_X16 FILLER_182_353 ();
 FILLCELL_X8 FILLER_182_369 ();
 FILLCELL_X2 FILLER_182_377 ();
 FILLCELL_X1 FILLER_182_379 ();
 FILLCELL_X32 FILLER_182_1518 ();
 FILLCELL_X32 FILLER_182_1550 ();
 FILLCELL_X32 FILLER_182_1582 ();
 FILLCELL_X32 FILLER_182_1614 ();
 FILLCELL_X32 FILLER_182_1646 ();
 FILLCELL_X32 FILLER_182_1678 ();
 FILLCELL_X32 FILLER_182_1710 ();
 FILLCELL_X8 FILLER_182_1742 ();
 FILLCELL_X4 FILLER_182_1750 ();
 FILLCELL_X2 FILLER_182_1754 ();
 FILLCELL_X32 FILLER_183_1 ();
 FILLCELL_X32 FILLER_183_33 ();
 FILLCELL_X32 FILLER_183_65 ();
 FILLCELL_X32 FILLER_183_97 ();
 FILLCELL_X32 FILLER_183_129 ();
 FILLCELL_X32 FILLER_183_161 ();
 FILLCELL_X32 FILLER_183_193 ();
 FILLCELL_X32 FILLER_183_225 ();
 FILLCELL_X32 FILLER_183_257 ();
 FILLCELL_X32 FILLER_183_289 ();
 FILLCELL_X32 FILLER_183_321 ();
 FILLCELL_X16 FILLER_183_353 ();
 FILLCELL_X8 FILLER_183_369 ();
 FILLCELL_X2 FILLER_183_377 ();
 FILLCELL_X1 FILLER_183_379 ();
 FILLCELL_X32 FILLER_183_1518 ();
 FILLCELL_X32 FILLER_183_1550 ();
 FILLCELL_X32 FILLER_183_1582 ();
 FILLCELL_X32 FILLER_183_1614 ();
 FILLCELL_X32 FILLER_183_1646 ();
 FILLCELL_X32 FILLER_183_1678 ();
 FILLCELL_X32 FILLER_183_1710 ();
 FILLCELL_X4 FILLER_183_1742 ();
 FILLCELL_X2 FILLER_183_1746 ();
 FILLCELL_X1 FILLER_183_1748 ();
 FILLCELL_X4 FILLER_183_1752 ();
 FILLCELL_X32 FILLER_184_1 ();
 FILLCELL_X32 FILLER_184_33 ();
 FILLCELL_X32 FILLER_184_65 ();
 FILLCELL_X32 FILLER_184_97 ();
 FILLCELL_X32 FILLER_184_129 ();
 FILLCELL_X32 FILLER_184_161 ();
 FILLCELL_X32 FILLER_184_193 ();
 FILLCELL_X32 FILLER_184_225 ();
 FILLCELL_X32 FILLER_184_257 ();
 FILLCELL_X32 FILLER_184_289 ();
 FILLCELL_X32 FILLER_184_321 ();
 FILLCELL_X16 FILLER_184_353 ();
 FILLCELL_X8 FILLER_184_369 ();
 FILLCELL_X2 FILLER_184_377 ();
 FILLCELL_X1 FILLER_184_379 ();
 FILLCELL_X32 FILLER_184_1518 ();
 FILLCELL_X32 FILLER_184_1550 ();
 FILLCELL_X32 FILLER_184_1582 ();
 FILLCELL_X32 FILLER_184_1614 ();
 FILLCELL_X32 FILLER_184_1646 ();
 FILLCELL_X32 FILLER_184_1678 ();
 FILLCELL_X32 FILLER_184_1710 ();
 FILLCELL_X8 FILLER_184_1742 ();
 FILLCELL_X4 FILLER_184_1750 ();
 FILLCELL_X2 FILLER_184_1754 ();
 FILLCELL_X32 FILLER_185_1 ();
 FILLCELL_X32 FILLER_185_33 ();
 FILLCELL_X32 FILLER_185_65 ();
 FILLCELL_X32 FILLER_185_97 ();
 FILLCELL_X32 FILLER_185_129 ();
 FILLCELL_X32 FILLER_185_161 ();
 FILLCELL_X32 FILLER_185_193 ();
 FILLCELL_X32 FILLER_185_225 ();
 FILLCELL_X32 FILLER_185_257 ();
 FILLCELL_X32 FILLER_185_289 ();
 FILLCELL_X32 FILLER_185_321 ();
 FILLCELL_X16 FILLER_185_353 ();
 FILLCELL_X8 FILLER_185_369 ();
 FILLCELL_X2 FILLER_185_377 ();
 FILLCELL_X1 FILLER_185_379 ();
 FILLCELL_X32 FILLER_185_1518 ();
 FILLCELL_X32 FILLER_185_1550 ();
 FILLCELL_X32 FILLER_185_1582 ();
 FILLCELL_X32 FILLER_185_1614 ();
 FILLCELL_X32 FILLER_185_1646 ();
 FILLCELL_X32 FILLER_185_1678 ();
 FILLCELL_X32 FILLER_185_1710 ();
 FILLCELL_X8 FILLER_185_1742 ();
 FILLCELL_X4 FILLER_185_1750 ();
 FILLCELL_X2 FILLER_185_1754 ();
 FILLCELL_X32 FILLER_186_1 ();
 FILLCELL_X32 FILLER_186_33 ();
 FILLCELL_X32 FILLER_186_65 ();
 FILLCELL_X32 FILLER_186_97 ();
 FILLCELL_X32 FILLER_186_129 ();
 FILLCELL_X32 FILLER_186_161 ();
 FILLCELL_X32 FILLER_186_193 ();
 FILLCELL_X32 FILLER_186_225 ();
 FILLCELL_X32 FILLER_186_257 ();
 FILLCELL_X32 FILLER_186_289 ();
 FILLCELL_X32 FILLER_186_321 ();
 FILLCELL_X16 FILLER_186_353 ();
 FILLCELL_X8 FILLER_186_369 ();
 FILLCELL_X2 FILLER_186_377 ();
 FILLCELL_X1 FILLER_186_379 ();
 FILLCELL_X32 FILLER_186_1518 ();
 FILLCELL_X32 FILLER_186_1550 ();
 FILLCELL_X32 FILLER_186_1582 ();
 FILLCELL_X32 FILLER_186_1614 ();
 FILLCELL_X32 FILLER_186_1646 ();
 FILLCELL_X32 FILLER_186_1678 ();
 FILLCELL_X32 FILLER_186_1710 ();
 FILLCELL_X8 FILLER_186_1742 ();
 FILLCELL_X4 FILLER_186_1750 ();
 FILLCELL_X2 FILLER_186_1754 ();
 FILLCELL_X32 FILLER_187_1 ();
 FILLCELL_X32 FILLER_187_33 ();
 FILLCELL_X32 FILLER_187_65 ();
 FILLCELL_X32 FILLER_187_97 ();
 FILLCELL_X32 FILLER_187_129 ();
 FILLCELL_X32 FILLER_187_161 ();
 FILLCELL_X32 FILLER_187_193 ();
 FILLCELL_X32 FILLER_187_225 ();
 FILLCELL_X32 FILLER_187_257 ();
 FILLCELL_X32 FILLER_187_289 ();
 FILLCELL_X32 FILLER_187_321 ();
 FILLCELL_X16 FILLER_187_353 ();
 FILLCELL_X8 FILLER_187_369 ();
 FILLCELL_X2 FILLER_187_377 ();
 FILLCELL_X1 FILLER_187_379 ();
 FILLCELL_X32 FILLER_187_1518 ();
 FILLCELL_X32 FILLER_187_1550 ();
 FILLCELL_X32 FILLER_187_1582 ();
 FILLCELL_X32 FILLER_187_1614 ();
 FILLCELL_X32 FILLER_187_1646 ();
 FILLCELL_X32 FILLER_187_1678 ();
 FILLCELL_X32 FILLER_187_1710 ();
 FILLCELL_X8 FILLER_187_1742 ();
 FILLCELL_X4 FILLER_187_1750 ();
 FILLCELL_X2 FILLER_187_1754 ();
 FILLCELL_X4 FILLER_188_1 ();
 FILLCELL_X32 FILLER_188_10 ();
 FILLCELL_X32 FILLER_188_42 ();
 FILLCELL_X32 FILLER_188_74 ();
 FILLCELL_X32 FILLER_188_106 ();
 FILLCELL_X32 FILLER_188_138 ();
 FILLCELL_X32 FILLER_188_170 ();
 FILLCELL_X32 FILLER_188_202 ();
 FILLCELL_X32 FILLER_188_234 ();
 FILLCELL_X32 FILLER_188_266 ();
 FILLCELL_X32 FILLER_188_298 ();
 FILLCELL_X32 FILLER_188_330 ();
 FILLCELL_X16 FILLER_188_362 ();
 FILLCELL_X2 FILLER_188_378 ();
 FILLCELL_X32 FILLER_188_1518 ();
 FILLCELL_X32 FILLER_188_1550 ();
 FILLCELL_X32 FILLER_188_1582 ();
 FILLCELL_X32 FILLER_188_1614 ();
 FILLCELL_X32 FILLER_188_1646 ();
 FILLCELL_X32 FILLER_188_1678 ();
 FILLCELL_X32 FILLER_188_1710 ();
 FILLCELL_X8 FILLER_188_1742 ();
 FILLCELL_X4 FILLER_188_1750 ();
 FILLCELL_X2 FILLER_188_1754 ();
 FILLCELL_X32 FILLER_189_1 ();
 FILLCELL_X32 FILLER_189_33 ();
 FILLCELL_X32 FILLER_189_65 ();
 FILLCELL_X32 FILLER_189_97 ();
 FILLCELL_X32 FILLER_189_129 ();
 FILLCELL_X32 FILLER_189_161 ();
 FILLCELL_X32 FILLER_189_193 ();
 FILLCELL_X32 FILLER_189_225 ();
 FILLCELL_X32 FILLER_189_257 ();
 FILLCELL_X32 FILLER_189_289 ();
 FILLCELL_X32 FILLER_189_321 ();
 FILLCELL_X16 FILLER_189_353 ();
 FILLCELL_X8 FILLER_189_369 ();
 FILLCELL_X2 FILLER_189_377 ();
 FILLCELL_X1 FILLER_189_379 ();
 FILLCELL_X32 FILLER_189_1518 ();
 FILLCELL_X32 FILLER_189_1550 ();
 FILLCELL_X32 FILLER_189_1582 ();
 FILLCELL_X32 FILLER_189_1614 ();
 FILLCELL_X32 FILLER_189_1646 ();
 FILLCELL_X32 FILLER_189_1678 ();
 FILLCELL_X32 FILLER_189_1710 ();
 FILLCELL_X8 FILLER_189_1742 ();
 FILLCELL_X4 FILLER_189_1750 ();
 FILLCELL_X2 FILLER_189_1754 ();
 FILLCELL_X32 FILLER_190_1 ();
 FILLCELL_X32 FILLER_190_33 ();
 FILLCELL_X32 FILLER_190_65 ();
 FILLCELL_X32 FILLER_190_97 ();
 FILLCELL_X32 FILLER_190_129 ();
 FILLCELL_X32 FILLER_190_161 ();
 FILLCELL_X32 FILLER_190_193 ();
 FILLCELL_X32 FILLER_190_225 ();
 FILLCELL_X32 FILLER_190_257 ();
 FILLCELL_X32 FILLER_190_289 ();
 FILLCELL_X32 FILLER_190_321 ();
 FILLCELL_X16 FILLER_190_353 ();
 FILLCELL_X8 FILLER_190_369 ();
 FILLCELL_X2 FILLER_190_377 ();
 FILLCELL_X1 FILLER_190_379 ();
 FILLCELL_X32 FILLER_190_1518 ();
 FILLCELL_X32 FILLER_190_1550 ();
 FILLCELL_X32 FILLER_190_1582 ();
 FILLCELL_X32 FILLER_190_1614 ();
 FILLCELL_X32 FILLER_190_1646 ();
 FILLCELL_X32 FILLER_190_1678 ();
 FILLCELL_X32 FILLER_190_1710 ();
 FILLCELL_X8 FILLER_190_1742 ();
 FILLCELL_X4 FILLER_190_1750 ();
 FILLCELL_X2 FILLER_190_1754 ();
 FILLCELL_X32 FILLER_191_1 ();
 FILLCELL_X32 FILLER_191_33 ();
 FILLCELL_X32 FILLER_191_65 ();
 FILLCELL_X32 FILLER_191_97 ();
 FILLCELL_X32 FILLER_191_129 ();
 FILLCELL_X32 FILLER_191_161 ();
 FILLCELL_X32 FILLER_191_193 ();
 FILLCELL_X32 FILLER_191_225 ();
 FILLCELL_X32 FILLER_191_257 ();
 FILLCELL_X32 FILLER_191_289 ();
 FILLCELL_X32 FILLER_191_321 ();
 FILLCELL_X16 FILLER_191_353 ();
 FILLCELL_X8 FILLER_191_369 ();
 FILLCELL_X2 FILLER_191_377 ();
 FILLCELL_X1 FILLER_191_379 ();
 FILLCELL_X32 FILLER_191_1518 ();
 FILLCELL_X32 FILLER_191_1550 ();
 FILLCELL_X32 FILLER_191_1582 ();
 FILLCELL_X32 FILLER_191_1614 ();
 FILLCELL_X32 FILLER_191_1646 ();
 FILLCELL_X32 FILLER_191_1678 ();
 FILLCELL_X32 FILLER_191_1710 ();
 FILLCELL_X8 FILLER_191_1742 ();
 FILLCELL_X4 FILLER_191_1750 ();
 FILLCELL_X2 FILLER_191_1754 ();
 FILLCELL_X32 FILLER_192_1 ();
 FILLCELL_X32 FILLER_192_33 ();
 FILLCELL_X32 FILLER_192_65 ();
 FILLCELL_X32 FILLER_192_97 ();
 FILLCELL_X32 FILLER_192_129 ();
 FILLCELL_X32 FILLER_192_161 ();
 FILLCELL_X32 FILLER_192_193 ();
 FILLCELL_X32 FILLER_192_225 ();
 FILLCELL_X32 FILLER_192_257 ();
 FILLCELL_X32 FILLER_192_289 ();
 FILLCELL_X32 FILLER_192_321 ();
 FILLCELL_X16 FILLER_192_353 ();
 FILLCELL_X8 FILLER_192_369 ();
 FILLCELL_X2 FILLER_192_377 ();
 FILLCELL_X1 FILLER_192_379 ();
 FILLCELL_X32 FILLER_192_1518 ();
 FILLCELL_X32 FILLER_192_1550 ();
 FILLCELL_X32 FILLER_192_1582 ();
 FILLCELL_X32 FILLER_192_1614 ();
 FILLCELL_X32 FILLER_192_1646 ();
 FILLCELL_X32 FILLER_192_1678 ();
 FILLCELL_X32 FILLER_192_1710 ();
 FILLCELL_X8 FILLER_192_1742 ();
 FILLCELL_X4 FILLER_192_1750 ();
 FILLCELL_X2 FILLER_192_1754 ();
 FILLCELL_X32 FILLER_193_1 ();
 FILLCELL_X32 FILLER_193_33 ();
 FILLCELL_X32 FILLER_193_65 ();
 FILLCELL_X32 FILLER_193_97 ();
 FILLCELL_X32 FILLER_193_129 ();
 FILLCELL_X32 FILLER_193_161 ();
 FILLCELL_X32 FILLER_193_193 ();
 FILLCELL_X32 FILLER_193_225 ();
 FILLCELL_X32 FILLER_193_257 ();
 FILLCELL_X32 FILLER_193_289 ();
 FILLCELL_X32 FILLER_193_321 ();
 FILLCELL_X16 FILLER_193_353 ();
 FILLCELL_X8 FILLER_193_369 ();
 FILLCELL_X2 FILLER_193_377 ();
 FILLCELL_X1 FILLER_193_379 ();
 FILLCELL_X32 FILLER_193_1518 ();
 FILLCELL_X32 FILLER_193_1550 ();
 FILLCELL_X32 FILLER_193_1582 ();
 FILLCELL_X32 FILLER_193_1614 ();
 FILLCELL_X32 FILLER_193_1646 ();
 FILLCELL_X32 FILLER_193_1678 ();
 FILLCELL_X32 FILLER_193_1710 ();
 FILLCELL_X4 FILLER_193_1742 ();
 FILLCELL_X2 FILLER_193_1746 ();
 FILLCELL_X1 FILLER_193_1748 ();
 FILLCELL_X4 FILLER_193_1752 ();
 FILLCELL_X32 FILLER_194_1 ();
 FILLCELL_X32 FILLER_194_33 ();
 FILLCELL_X32 FILLER_194_65 ();
 FILLCELL_X32 FILLER_194_97 ();
 FILLCELL_X32 FILLER_194_129 ();
 FILLCELL_X32 FILLER_194_161 ();
 FILLCELL_X32 FILLER_194_193 ();
 FILLCELL_X32 FILLER_194_225 ();
 FILLCELL_X32 FILLER_194_257 ();
 FILLCELL_X32 FILLER_194_289 ();
 FILLCELL_X32 FILLER_194_321 ();
 FILLCELL_X16 FILLER_194_353 ();
 FILLCELL_X8 FILLER_194_369 ();
 FILLCELL_X2 FILLER_194_377 ();
 FILLCELL_X1 FILLER_194_379 ();
 FILLCELL_X32 FILLER_194_1518 ();
 FILLCELL_X32 FILLER_194_1550 ();
 FILLCELL_X32 FILLER_194_1582 ();
 FILLCELL_X32 FILLER_194_1614 ();
 FILLCELL_X32 FILLER_194_1646 ();
 FILLCELL_X32 FILLER_194_1678 ();
 FILLCELL_X32 FILLER_194_1710 ();
 FILLCELL_X8 FILLER_194_1742 ();
 FILLCELL_X4 FILLER_194_1750 ();
 FILLCELL_X2 FILLER_194_1754 ();
 FILLCELL_X32 FILLER_195_1 ();
 FILLCELL_X32 FILLER_195_33 ();
 FILLCELL_X32 FILLER_195_65 ();
 FILLCELL_X32 FILLER_195_97 ();
 FILLCELL_X32 FILLER_195_129 ();
 FILLCELL_X32 FILLER_195_161 ();
 FILLCELL_X32 FILLER_195_193 ();
 FILLCELL_X32 FILLER_195_225 ();
 FILLCELL_X32 FILLER_195_257 ();
 FILLCELL_X32 FILLER_195_289 ();
 FILLCELL_X32 FILLER_195_321 ();
 FILLCELL_X16 FILLER_195_353 ();
 FILLCELL_X8 FILLER_195_369 ();
 FILLCELL_X2 FILLER_195_377 ();
 FILLCELL_X1 FILLER_195_379 ();
 FILLCELL_X32 FILLER_195_1518 ();
 FILLCELL_X32 FILLER_195_1550 ();
 FILLCELL_X32 FILLER_195_1582 ();
 FILLCELL_X32 FILLER_195_1614 ();
 FILLCELL_X32 FILLER_195_1646 ();
 FILLCELL_X32 FILLER_195_1678 ();
 FILLCELL_X32 FILLER_195_1710 ();
 FILLCELL_X8 FILLER_195_1742 ();
 FILLCELL_X4 FILLER_195_1750 ();
 FILLCELL_X2 FILLER_195_1754 ();
 FILLCELL_X32 FILLER_196_1 ();
 FILLCELL_X32 FILLER_196_33 ();
 FILLCELL_X32 FILLER_196_65 ();
 FILLCELL_X32 FILLER_196_97 ();
 FILLCELL_X32 FILLER_196_129 ();
 FILLCELL_X32 FILLER_196_161 ();
 FILLCELL_X32 FILLER_196_193 ();
 FILLCELL_X32 FILLER_196_225 ();
 FILLCELL_X32 FILLER_196_257 ();
 FILLCELL_X32 FILLER_196_289 ();
 FILLCELL_X32 FILLER_196_321 ();
 FILLCELL_X16 FILLER_196_353 ();
 FILLCELL_X8 FILLER_196_369 ();
 FILLCELL_X2 FILLER_196_377 ();
 FILLCELL_X1 FILLER_196_379 ();
 FILLCELL_X32 FILLER_196_1518 ();
 FILLCELL_X32 FILLER_196_1550 ();
 FILLCELL_X32 FILLER_196_1582 ();
 FILLCELL_X32 FILLER_196_1614 ();
 FILLCELL_X32 FILLER_196_1646 ();
 FILLCELL_X32 FILLER_196_1678 ();
 FILLCELL_X32 FILLER_196_1710 ();
 FILLCELL_X8 FILLER_196_1742 ();
 FILLCELL_X4 FILLER_196_1750 ();
 FILLCELL_X2 FILLER_196_1754 ();
 FILLCELL_X32 FILLER_197_1 ();
 FILLCELL_X32 FILLER_197_33 ();
 FILLCELL_X32 FILLER_197_65 ();
 FILLCELL_X32 FILLER_197_97 ();
 FILLCELL_X32 FILLER_197_129 ();
 FILLCELL_X32 FILLER_197_161 ();
 FILLCELL_X32 FILLER_197_193 ();
 FILLCELL_X32 FILLER_197_225 ();
 FILLCELL_X32 FILLER_197_257 ();
 FILLCELL_X32 FILLER_197_289 ();
 FILLCELL_X32 FILLER_197_321 ();
 FILLCELL_X16 FILLER_197_353 ();
 FILLCELL_X8 FILLER_197_369 ();
 FILLCELL_X2 FILLER_197_377 ();
 FILLCELL_X1 FILLER_197_379 ();
 FILLCELL_X32 FILLER_197_1518 ();
 FILLCELL_X32 FILLER_197_1550 ();
 FILLCELL_X32 FILLER_197_1582 ();
 FILLCELL_X32 FILLER_197_1614 ();
 FILLCELL_X32 FILLER_197_1646 ();
 FILLCELL_X32 FILLER_197_1678 ();
 FILLCELL_X32 FILLER_197_1710 ();
 FILLCELL_X8 FILLER_197_1742 ();
 FILLCELL_X4 FILLER_197_1750 ();
 FILLCELL_X2 FILLER_197_1754 ();
 FILLCELL_X4 FILLER_198_1 ();
 FILLCELL_X32 FILLER_198_8 ();
 FILLCELL_X32 FILLER_198_40 ();
 FILLCELL_X32 FILLER_198_72 ();
 FILLCELL_X32 FILLER_198_104 ();
 FILLCELL_X32 FILLER_198_136 ();
 FILLCELL_X32 FILLER_198_168 ();
 FILLCELL_X32 FILLER_198_200 ();
 FILLCELL_X32 FILLER_198_232 ();
 FILLCELL_X32 FILLER_198_264 ();
 FILLCELL_X32 FILLER_198_296 ();
 FILLCELL_X32 FILLER_198_328 ();
 FILLCELL_X16 FILLER_198_360 ();
 FILLCELL_X4 FILLER_198_376 ();
 FILLCELL_X32 FILLER_198_1518 ();
 FILLCELL_X32 FILLER_198_1550 ();
 FILLCELL_X32 FILLER_198_1582 ();
 FILLCELL_X32 FILLER_198_1614 ();
 FILLCELL_X32 FILLER_198_1646 ();
 FILLCELL_X32 FILLER_198_1678 ();
 FILLCELL_X32 FILLER_198_1710 ();
 FILLCELL_X8 FILLER_198_1742 ();
 FILLCELL_X4 FILLER_198_1750 ();
 FILLCELL_X2 FILLER_198_1754 ();
 FILLCELL_X32 FILLER_199_1 ();
 FILLCELL_X32 FILLER_199_33 ();
 FILLCELL_X32 FILLER_199_65 ();
 FILLCELL_X32 FILLER_199_97 ();
 FILLCELL_X32 FILLER_199_129 ();
 FILLCELL_X32 FILLER_199_161 ();
 FILLCELL_X32 FILLER_199_193 ();
 FILLCELL_X32 FILLER_199_225 ();
 FILLCELL_X32 FILLER_199_257 ();
 FILLCELL_X32 FILLER_199_289 ();
 FILLCELL_X32 FILLER_199_321 ();
 FILLCELL_X16 FILLER_199_353 ();
 FILLCELL_X8 FILLER_199_369 ();
 FILLCELL_X2 FILLER_199_377 ();
 FILLCELL_X1 FILLER_199_379 ();
 FILLCELL_X32 FILLER_199_1518 ();
 FILLCELL_X32 FILLER_199_1550 ();
 FILLCELL_X32 FILLER_199_1582 ();
 FILLCELL_X32 FILLER_199_1614 ();
 FILLCELL_X32 FILLER_199_1646 ();
 FILLCELL_X32 FILLER_199_1678 ();
 FILLCELL_X32 FILLER_199_1710 ();
 FILLCELL_X8 FILLER_199_1742 ();
 FILLCELL_X4 FILLER_199_1750 ();
 FILLCELL_X2 FILLER_199_1754 ();
 FILLCELL_X32 FILLER_200_1 ();
 FILLCELL_X32 FILLER_200_33 ();
 FILLCELL_X32 FILLER_200_65 ();
 FILLCELL_X32 FILLER_200_97 ();
 FILLCELL_X32 FILLER_200_129 ();
 FILLCELL_X32 FILLER_200_161 ();
 FILLCELL_X32 FILLER_200_193 ();
 FILLCELL_X32 FILLER_200_225 ();
 FILLCELL_X32 FILLER_200_257 ();
 FILLCELL_X32 FILLER_200_289 ();
 FILLCELL_X32 FILLER_200_321 ();
 FILLCELL_X16 FILLER_200_353 ();
 FILLCELL_X8 FILLER_200_369 ();
 FILLCELL_X2 FILLER_200_377 ();
 FILLCELL_X1 FILLER_200_379 ();
 FILLCELL_X32 FILLER_200_1518 ();
 FILLCELL_X32 FILLER_200_1550 ();
 FILLCELL_X32 FILLER_200_1582 ();
 FILLCELL_X32 FILLER_200_1614 ();
 FILLCELL_X32 FILLER_200_1646 ();
 FILLCELL_X32 FILLER_200_1678 ();
 FILLCELL_X32 FILLER_200_1710 ();
 FILLCELL_X8 FILLER_200_1742 ();
 FILLCELL_X4 FILLER_200_1750 ();
 FILLCELL_X2 FILLER_200_1754 ();
 FILLCELL_X32 FILLER_201_1 ();
 FILLCELL_X32 FILLER_201_33 ();
 FILLCELL_X32 FILLER_201_65 ();
 FILLCELL_X32 FILLER_201_97 ();
 FILLCELL_X32 FILLER_201_129 ();
 FILLCELL_X32 FILLER_201_161 ();
 FILLCELL_X32 FILLER_201_193 ();
 FILLCELL_X32 FILLER_201_225 ();
 FILLCELL_X32 FILLER_201_257 ();
 FILLCELL_X32 FILLER_201_289 ();
 FILLCELL_X32 FILLER_201_321 ();
 FILLCELL_X16 FILLER_201_353 ();
 FILLCELL_X8 FILLER_201_369 ();
 FILLCELL_X2 FILLER_201_377 ();
 FILLCELL_X1 FILLER_201_379 ();
 FILLCELL_X32 FILLER_201_1518 ();
 FILLCELL_X32 FILLER_201_1550 ();
 FILLCELL_X32 FILLER_201_1582 ();
 FILLCELL_X32 FILLER_201_1614 ();
 FILLCELL_X32 FILLER_201_1646 ();
 FILLCELL_X32 FILLER_201_1678 ();
 FILLCELL_X32 FILLER_201_1710 ();
 FILLCELL_X8 FILLER_201_1742 ();
 FILLCELL_X4 FILLER_201_1750 ();
 FILLCELL_X2 FILLER_201_1754 ();
 FILLCELL_X32 FILLER_202_1 ();
 FILLCELL_X32 FILLER_202_33 ();
 FILLCELL_X32 FILLER_202_65 ();
 FILLCELL_X32 FILLER_202_97 ();
 FILLCELL_X32 FILLER_202_129 ();
 FILLCELL_X32 FILLER_202_161 ();
 FILLCELL_X32 FILLER_202_193 ();
 FILLCELL_X32 FILLER_202_225 ();
 FILLCELL_X32 FILLER_202_257 ();
 FILLCELL_X32 FILLER_202_289 ();
 FILLCELL_X32 FILLER_202_321 ();
 FILLCELL_X16 FILLER_202_353 ();
 FILLCELL_X8 FILLER_202_369 ();
 FILLCELL_X2 FILLER_202_377 ();
 FILLCELL_X1 FILLER_202_379 ();
 FILLCELL_X32 FILLER_202_1518 ();
 FILLCELL_X32 FILLER_202_1550 ();
 FILLCELL_X32 FILLER_202_1582 ();
 FILLCELL_X32 FILLER_202_1614 ();
 FILLCELL_X32 FILLER_202_1646 ();
 FILLCELL_X32 FILLER_202_1678 ();
 FILLCELL_X32 FILLER_202_1710 ();
 FILLCELL_X4 FILLER_202_1742 ();
 FILLCELL_X2 FILLER_202_1746 ();
 FILLCELL_X1 FILLER_202_1748 ();
 FILLCELL_X4 FILLER_202_1752 ();
 FILLCELL_X32 FILLER_203_1 ();
 FILLCELL_X32 FILLER_203_33 ();
 FILLCELL_X32 FILLER_203_65 ();
 FILLCELL_X32 FILLER_203_97 ();
 FILLCELL_X32 FILLER_203_129 ();
 FILLCELL_X32 FILLER_203_161 ();
 FILLCELL_X32 FILLER_203_193 ();
 FILLCELL_X32 FILLER_203_225 ();
 FILLCELL_X32 FILLER_203_257 ();
 FILLCELL_X32 FILLER_203_289 ();
 FILLCELL_X32 FILLER_203_321 ();
 FILLCELL_X16 FILLER_203_353 ();
 FILLCELL_X8 FILLER_203_369 ();
 FILLCELL_X2 FILLER_203_377 ();
 FILLCELL_X1 FILLER_203_379 ();
 FILLCELL_X32 FILLER_203_1518 ();
 FILLCELL_X32 FILLER_203_1550 ();
 FILLCELL_X32 FILLER_203_1582 ();
 FILLCELL_X32 FILLER_203_1614 ();
 FILLCELL_X32 FILLER_203_1646 ();
 FILLCELL_X32 FILLER_203_1678 ();
 FILLCELL_X32 FILLER_203_1710 ();
 FILLCELL_X8 FILLER_203_1742 ();
 FILLCELL_X4 FILLER_203_1750 ();
 FILLCELL_X2 FILLER_203_1754 ();
 FILLCELL_X32 FILLER_204_1 ();
 FILLCELL_X32 FILLER_204_33 ();
 FILLCELL_X32 FILLER_204_65 ();
 FILLCELL_X32 FILLER_204_97 ();
 FILLCELL_X32 FILLER_204_129 ();
 FILLCELL_X32 FILLER_204_161 ();
 FILLCELL_X32 FILLER_204_193 ();
 FILLCELL_X32 FILLER_204_225 ();
 FILLCELL_X32 FILLER_204_257 ();
 FILLCELL_X32 FILLER_204_289 ();
 FILLCELL_X32 FILLER_204_321 ();
 FILLCELL_X16 FILLER_204_353 ();
 FILLCELL_X8 FILLER_204_369 ();
 FILLCELL_X2 FILLER_204_377 ();
 FILLCELL_X1 FILLER_204_379 ();
 FILLCELL_X32 FILLER_204_1518 ();
 FILLCELL_X32 FILLER_204_1550 ();
 FILLCELL_X32 FILLER_204_1582 ();
 FILLCELL_X32 FILLER_204_1614 ();
 FILLCELL_X32 FILLER_204_1646 ();
 FILLCELL_X32 FILLER_204_1678 ();
 FILLCELL_X32 FILLER_204_1710 ();
 FILLCELL_X8 FILLER_204_1742 ();
 FILLCELL_X4 FILLER_204_1750 ();
 FILLCELL_X2 FILLER_204_1754 ();
 FILLCELL_X32 FILLER_205_1 ();
 FILLCELL_X32 FILLER_205_33 ();
 FILLCELL_X32 FILLER_205_65 ();
 FILLCELL_X32 FILLER_205_97 ();
 FILLCELL_X32 FILLER_205_129 ();
 FILLCELL_X32 FILLER_205_161 ();
 FILLCELL_X32 FILLER_205_193 ();
 FILLCELL_X32 FILLER_205_225 ();
 FILLCELL_X32 FILLER_205_257 ();
 FILLCELL_X32 FILLER_205_289 ();
 FILLCELL_X32 FILLER_205_321 ();
 FILLCELL_X16 FILLER_205_353 ();
 FILLCELL_X8 FILLER_205_369 ();
 FILLCELL_X2 FILLER_205_377 ();
 FILLCELL_X1 FILLER_205_379 ();
 FILLCELL_X32 FILLER_205_1518 ();
 FILLCELL_X32 FILLER_205_1550 ();
 FILLCELL_X32 FILLER_205_1582 ();
 FILLCELL_X32 FILLER_205_1614 ();
 FILLCELL_X32 FILLER_205_1646 ();
 FILLCELL_X32 FILLER_205_1678 ();
 FILLCELL_X32 FILLER_205_1710 ();
 FILLCELL_X8 FILLER_205_1742 ();
 FILLCELL_X4 FILLER_205_1750 ();
 FILLCELL_X2 FILLER_205_1754 ();
 FILLCELL_X32 FILLER_206_1 ();
 FILLCELL_X32 FILLER_206_33 ();
 FILLCELL_X32 FILLER_206_65 ();
 FILLCELL_X32 FILLER_206_97 ();
 FILLCELL_X32 FILLER_206_129 ();
 FILLCELL_X32 FILLER_206_161 ();
 FILLCELL_X32 FILLER_206_193 ();
 FILLCELL_X32 FILLER_206_225 ();
 FILLCELL_X32 FILLER_206_257 ();
 FILLCELL_X32 FILLER_206_289 ();
 FILLCELL_X32 FILLER_206_321 ();
 FILLCELL_X16 FILLER_206_353 ();
 FILLCELL_X8 FILLER_206_369 ();
 FILLCELL_X2 FILLER_206_377 ();
 FILLCELL_X1 FILLER_206_379 ();
 FILLCELL_X32 FILLER_206_1518 ();
 FILLCELL_X32 FILLER_206_1550 ();
 FILLCELL_X32 FILLER_206_1582 ();
 FILLCELL_X32 FILLER_206_1614 ();
 FILLCELL_X32 FILLER_206_1646 ();
 FILLCELL_X32 FILLER_206_1678 ();
 FILLCELL_X32 FILLER_206_1710 ();
 FILLCELL_X8 FILLER_206_1742 ();
 FILLCELL_X4 FILLER_206_1750 ();
 FILLCELL_X2 FILLER_206_1754 ();
 FILLCELL_X4 FILLER_207_1 ();
 FILLCELL_X32 FILLER_207_18 ();
 FILLCELL_X32 FILLER_207_50 ();
 FILLCELL_X32 FILLER_207_82 ();
 FILLCELL_X32 FILLER_207_114 ();
 FILLCELL_X32 FILLER_207_146 ();
 FILLCELL_X32 FILLER_207_178 ();
 FILLCELL_X32 FILLER_207_210 ();
 FILLCELL_X32 FILLER_207_242 ();
 FILLCELL_X32 FILLER_207_274 ();
 FILLCELL_X32 FILLER_207_306 ();
 FILLCELL_X32 FILLER_207_338 ();
 FILLCELL_X8 FILLER_207_370 ();
 FILLCELL_X2 FILLER_207_378 ();
 FILLCELL_X32 FILLER_207_1518 ();
 FILLCELL_X32 FILLER_207_1550 ();
 FILLCELL_X32 FILLER_207_1582 ();
 FILLCELL_X32 FILLER_207_1614 ();
 FILLCELL_X32 FILLER_207_1646 ();
 FILLCELL_X32 FILLER_207_1678 ();
 FILLCELL_X32 FILLER_207_1710 ();
 FILLCELL_X8 FILLER_207_1742 ();
 FILLCELL_X4 FILLER_207_1750 ();
 FILLCELL_X2 FILLER_207_1754 ();
 FILLCELL_X32 FILLER_208_1 ();
 FILLCELL_X32 FILLER_208_33 ();
 FILLCELL_X32 FILLER_208_65 ();
 FILLCELL_X32 FILLER_208_97 ();
 FILLCELL_X32 FILLER_208_129 ();
 FILLCELL_X32 FILLER_208_161 ();
 FILLCELL_X32 FILLER_208_193 ();
 FILLCELL_X32 FILLER_208_225 ();
 FILLCELL_X32 FILLER_208_257 ();
 FILLCELL_X32 FILLER_208_289 ();
 FILLCELL_X32 FILLER_208_321 ();
 FILLCELL_X32 FILLER_208_353 ();
 FILLCELL_X32 FILLER_208_385 ();
 FILLCELL_X32 FILLER_208_417 ();
 FILLCELL_X32 FILLER_208_449 ();
 FILLCELL_X32 FILLER_208_481 ();
 FILLCELL_X32 FILLER_208_513 ();
 FILLCELL_X32 FILLER_208_545 ();
 FILLCELL_X32 FILLER_208_577 ();
 FILLCELL_X16 FILLER_208_609 ();
 FILLCELL_X4 FILLER_208_625 ();
 FILLCELL_X2 FILLER_208_629 ();
 FILLCELL_X32 FILLER_208_632 ();
 FILLCELL_X32 FILLER_208_664 ();
 FILLCELL_X32 FILLER_208_696 ();
 FILLCELL_X32 FILLER_208_728 ();
 FILLCELL_X32 FILLER_208_760 ();
 FILLCELL_X32 FILLER_208_792 ();
 FILLCELL_X32 FILLER_208_824 ();
 FILLCELL_X32 FILLER_208_856 ();
 FILLCELL_X32 FILLER_208_888 ();
 FILLCELL_X32 FILLER_208_920 ();
 FILLCELL_X32 FILLER_208_952 ();
 FILLCELL_X32 FILLER_208_984 ();
 FILLCELL_X32 FILLER_208_1016 ();
 FILLCELL_X32 FILLER_208_1048 ();
 FILLCELL_X32 FILLER_208_1080 ();
 FILLCELL_X32 FILLER_208_1112 ();
 FILLCELL_X32 FILLER_208_1144 ();
 FILLCELL_X32 FILLER_208_1176 ();
 FILLCELL_X32 FILLER_208_1208 ();
 FILLCELL_X16 FILLER_208_1240 ();
 FILLCELL_X4 FILLER_208_1256 ();
 FILLCELL_X2 FILLER_208_1260 ();
 FILLCELL_X32 FILLER_208_1263 ();
 FILLCELL_X32 FILLER_208_1295 ();
 FILLCELL_X32 FILLER_208_1327 ();
 FILLCELL_X32 FILLER_208_1359 ();
 FILLCELL_X32 FILLER_208_1391 ();
 FILLCELL_X32 FILLER_208_1423 ();
 FILLCELL_X32 FILLER_208_1455 ();
 FILLCELL_X32 FILLER_208_1487 ();
 FILLCELL_X32 FILLER_208_1519 ();
 FILLCELL_X32 FILLER_208_1551 ();
 FILLCELL_X32 FILLER_208_1583 ();
 FILLCELL_X32 FILLER_208_1615 ();
 FILLCELL_X32 FILLER_208_1647 ();
 FILLCELL_X32 FILLER_208_1679 ();
 FILLCELL_X32 FILLER_208_1711 ();
 FILLCELL_X8 FILLER_208_1743 ();
 FILLCELL_X4 FILLER_208_1751 ();
 FILLCELL_X1 FILLER_208_1755 ();
 FILLCELL_X32 FILLER_209_1 ();
 FILLCELL_X32 FILLER_209_33 ();
 FILLCELL_X32 FILLER_209_65 ();
 FILLCELL_X32 FILLER_209_97 ();
 FILLCELL_X32 FILLER_209_129 ();
 FILLCELL_X32 FILLER_209_161 ();
 FILLCELL_X32 FILLER_209_193 ();
 FILLCELL_X32 FILLER_209_225 ();
 FILLCELL_X32 FILLER_209_257 ();
 FILLCELL_X32 FILLER_209_289 ();
 FILLCELL_X32 FILLER_209_321 ();
 FILLCELL_X32 FILLER_209_353 ();
 FILLCELL_X32 FILLER_209_385 ();
 FILLCELL_X32 FILLER_209_417 ();
 FILLCELL_X32 FILLER_209_449 ();
 FILLCELL_X32 FILLER_209_481 ();
 FILLCELL_X32 FILLER_209_513 ();
 FILLCELL_X32 FILLER_209_545 ();
 FILLCELL_X32 FILLER_209_577 ();
 FILLCELL_X32 FILLER_209_609 ();
 FILLCELL_X32 FILLER_209_641 ();
 FILLCELL_X32 FILLER_209_673 ();
 FILLCELL_X32 FILLER_209_705 ();
 FILLCELL_X32 FILLER_209_737 ();
 FILLCELL_X32 FILLER_209_769 ();
 FILLCELL_X32 FILLER_209_801 ();
 FILLCELL_X32 FILLER_209_833 ();
 FILLCELL_X32 FILLER_209_865 ();
 FILLCELL_X32 FILLER_209_897 ();
 FILLCELL_X32 FILLER_209_929 ();
 FILLCELL_X32 FILLER_209_961 ();
 FILLCELL_X32 FILLER_209_993 ();
 FILLCELL_X32 FILLER_209_1025 ();
 FILLCELL_X32 FILLER_209_1057 ();
 FILLCELL_X32 FILLER_209_1089 ();
 FILLCELL_X32 FILLER_209_1121 ();
 FILLCELL_X32 FILLER_209_1153 ();
 FILLCELL_X32 FILLER_209_1185 ();
 FILLCELL_X32 FILLER_209_1217 ();
 FILLCELL_X8 FILLER_209_1249 ();
 FILLCELL_X4 FILLER_209_1257 ();
 FILLCELL_X2 FILLER_209_1261 ();
 FILLCELL_X32 FILLER_209_1264 ();
 FILLCELL_X32 FILLER_209_1296 ();
 FILLCELL_X32 FILLER_209_1328 ();
 FILLCELL_X32 FILLER_209_1360 ();
 FILLCELL_X32 FILLER_209_1392 ();
 FILLCELL_X32 FILLER_209_1424 ();
 FILLCELL_X32 FILLER_209_1456 ();
 FILLCELL_X32 FILLER_209_1488 ();
 FILLCELL_X32 FILLER_209_1520 ();
 FILLCELL_X32 FILLER_209_1552 ();
 FILLCELL_X32 FILLER_209_1584 ();
 FILLCELL_X32 FILLER_209_1616 ();
 FILLCELL_X32 FILLER_209_1648 ();
 FILLCELL_X32 FILLER_209_1680 ();
 FILLCELL_X32 FILLER_209_1712 ();
 FILLCELL_X8 FILLER_209_1744 ();
 FILLCELL_X4 FILLER_209_1752 ();
 FILLCELL_X32 FILLER_210_1 ();
 FILLCELL_X32 FILLER_210_33 ();
 FILLCELL_X32 FILLER_210_65 ();
 FILLCELL_X32 FILLER_210_97 ();
 FILLCELL_X32 FILLER_210_129 ();
 FILLCELL_X32 FILLER_210_161 ();
 FILLCELL_X32 FILLER_210_193 ();
 FILLCELL_X32 FILLER_210_225 ();
 FILLCELL_X32 FILLER_210_257 ();
 FILLCELL_X32 FILLER_210_289 ();
 FILLCELL_X32 FILLER_210_321 ();
 FILLCELL_X32 FILLER_210_353 ();
 FILLCELL_X32 FILLER_210_385 ();
 FILLCELL_X32 FILLER_210_417 ();
 FILLCELL_X32 FILLER_210_449 ();
 FILLCELL_X32 FILLER_210_481 ();
 FILLCELL_X32 FILLER_210_513 ();
 FILLCELL_X32 FILLER_210_545 ();
 FILLCELL_X32 FILLER_210_577 ();
 FILLCELL_X16 FILLER_210_609 ();
 FILLCELL_X4 FILLER_210_625 ();
 FILLCELL_X2 FILLER_210_629 ();
 FILLCELL_X32 FILLER_210_632 ();
 FILLCELL_X32 FILLER_210_664 ();
 FILLCELL_X32 FILLER_210_696 ();
 FILLCELL_X32 FILLER_210_728 ();
 FILLCELL_X32 FILLER_210_760 ();
 FILLCELL_X32 FILLER_210_792 ();
 FILLCELL_X32 FILLER_210_824 ();
 FILLCELL_X32 FILLER_210_856 ();
 FILLCELL_X32 FILLER_210_888 ();
 FILLCELL_X32 FILLER_210_920 ();
 FILLCELL_X32 FILLER_210_952 ();
 FILLCELL_X32 FILLER_210_984 ();
 FILLCELL_X32 FILLER_210_1016 ();
 FILLCELL_X32 FILLER_210_1048 ();
 FILLCELL_X32 FILLER_210_1080 ();
 FILLCELL_X32 FILLER_210_1112 ();
 FILLCELL_X32 FILLER_210_1144 ();
 FILLCELL_X32 FILLER_210_1176 ();
 FILLCELL_X32 FILLER_210_1208 ();
 FILLCELL_X32 FILLER_210_1240 ();
 FILLCELL_X32 FILLER_210_1272 ();
 FILLCELL_X32 FILLER_210_1304 ();
 FILLCELL_X32 FILLER_210_1336 ();
 FILLCELL_X32 FILLER_210_1368 ();
 FILLCELL_X32 FILLER_210_1400 ();
 FILLCELL_X32 FILLER_210_1432 ();
 FILLCELL_X32 FILLER_210_1464 ();
 FILLCELL_X32 FILLER_210_1496 ();
 FILLCELL_X32 FILLER_210_1528 ();
 FILLCELL_X32 FILLER_210_1560 ();
 FILLCELL_X32 FILLER_210_1592 ();
 FILLCELL_X32 FILLER_210_1624 ();
 FILLCELL_X32 FILLER_210_1656 ();
 FILLCELL_X32 FILLER_210_1688 ();
 FILLCELL_X32 FILLER_210_1720 ();
 FILLCELL_X4 FILLER_210_1752 ();
 FILLCELL_X32 FILLER_211_1 ();
 FILLCELL_X32 FILLER_211_33 ();
 FILLCELL_X32 FILLER_211_65 ();
 FILLCELL_X32 FILLER_211_97 ();
 FILLCELL_X32 FILLER_211_129 ();
 FILLCELL_X32 FILLER_211_161 ();
 FILLCELL_X32 FILLER_211_193 ();
 FILLCELL_X32 FILLER_211_225 ();
 FILLCELL_X32 FILLER_211_257 ();
 FILLCELL_X32 FILLER_211_289 ();
 FILLCELL_X32 FILLER_211_321 ();
 FILLCELL_X32 FILLER_211_353 ();
 FILLCELL_X32 FILLER_211_385 ();
 FILLCELL_X32 FILLER_211_417 ();
 FILLCELL_X32 FILLER_211_449 ();
 FILLCELL_X32 FILLER_211_481 ();
 FILLCELL_X32 FILLER_211_513 ();
 FILLCELL_X32 FILLER_211_545 ();
 FILLCELL_X32 FILLER_211_577 ();
 FILLCELL_X32 FILLER_211_609 ();
 FILLCELL_X32 FILLER_211_641 ();
 FILLCELL_X32 FILLER_211_673 ();
 FILLCELL_X32 FILLER_211_705 ();
 FILLCELL_X32 FILLER_211_737 ();
 FILLCELL_X32 FILLER_211_769 ();
 FILLCELL_X32 FILLER_211_801 ();
 FILLCELL_X32 FILLER_211_833 ();
 FILLCELL_X32 FILLER_211_865 ();
 FILLCELL_X32 FILLER_211_897 ();
 FILLCELL_X32 FILLER_211_929 ();
 FILLCELL_X32 FILLER_211_961 ();
 FILLCELL_X32 FILLER_211_993 ();
 FILLCELL_X32 FILLER_211_1025 ();
 FILLCELL_X32 FILLER_211_1057 ();
 FILLCELL_X32 FILLER_211_1089 ();
 FILLCELL_X32 FILLER_211_1121 ();
 FILLCELL_X32 FILLER_211_1153 ();
 FILLCELL_X32 FILLER_211_1185 ();
 FILLCELL_X32 FILLER_211_1217 ();
 FILLCELL_X8 FILLER_211_1249 ();
 FILLCELL_X4 FILLER_211_1257 ();
 FILLCELL_X2 FILLER_211_1261 ();
 FILLCELL_X32 FILLER_211_1264 ();
 FILLCELL_X32 FILLER_211_1296 ();
 FILLCELL_X32 FILLER_211_1328 ();
 FILLCELL_X32 FILLER_211_1360 ();
 FILLCELL_X32 FILLER_211_1392 ();
 FILLCELL_X32 FILLER_211_1424 ();
 FILLCELL_X32 FILLER_211_1456 ();
 FILLCELL_X32 FILLER_211_1488 ();
 FILLCELL_X32 FILLER_211_1520 ();
 FILLCELL_X32 FILLER_211_1552 ();
 FILLCELL_X32 FILLER_211_1584 ();
 FILLCELL_X32 FILLER_211_1616 ();
 FILLCELL_X32 FILLER_211_1648 ();
 FILLCELL_X32 FILLER_211_1680 ();
 FILLCELL_X32 FILLER_211_1712 ();
 FILLCELL_X8 FILLER_211_1744 ();
 FILLCELL_X4 FILLER_211_1752 ();
 FILLCELL_X32 FILLER_212_1 ();
 FILLCELL_X32 FILLER_212_33 ();
 FILLCELL_X32 FILLER_212_65 ();
 FILLCELL_X32 FILLER_212_97 ();
 FILLCELL_X32 FILLER_212_129 ();
 FILLCELL_X32 FILLER_212_161 ();
 FILLCELL_X32 FILLER_212_193 ();
 FILLCELL_X32 FILLER_212_225 ();
 FILLCELL_X32 FILLER_212_257 ();
 FILLCELL_X32 FILLER_212_289 ();
 FILLCELL_X32 FILLER_212_321 ();
 FILLCELL_X32 FILLER_212_353 ();
 FILLCELL_X32 FILLER_212_385 ();
 FILLCELL_X32 FILLER_212_417 ();
 FILLCELL_X32 FILLER_212_449 ();
 FILLCELL_X32 FILLER_212_481 ();
 FILLCELL_X32 FILLER_212_513 ();
 FILLCELL_X32 FILLER_212_545 ();
 FILLCELL_X32 FILLER_212_577 ();
 FILLCELL_X16 FILLER_212_609 ();
 FILLCELL_X4 FILLER_212_625 ();
 FILLCELL_X2 FILLER_212_629 ();
 FILLCELL_X32 FILLER_212_632 ();
 FILLCELL_X32 FILLER_212_664 ();
 FILLCELL_X32 FILLER_212_696 ();
 FILLCELL_X32 FILLER_212_728 ();
 FILLCELL_X32 FILLER_212_760 ();
 FILLCELL_X32 FILLER_212_792 ();
 FILLCELL_X32 FILLER_212_824 ();
 FILLCELL_X32 FILLER_212_856 ();
 FILLCELL_X32 FILLER_212_888 ();
 FILLCELL_X32 FILLER_212_920 ();
 FILLCELL_X32 FILLER_212_952 ();
 FILLCELL_X32 FILLER_212_984 ();
 FILLCELL_X32 FILLER_212_1016 ();
 FILLCELL_X32 FILLER_212_1048 ();
 FILLCELL_X32 FILLER_212_1080 ();
 FILLCELL_X32 FILLER_212_1112 ();
 FILLCELL_X32 FILLER_212_1144 ();
 FILLCELL_X32 FILLER_212_1176 ();
 FILLCELL_X32 FILLER_212_1208 ();
 FILLCELL_X32 FILLER_212_1240 ();
 FILLCELL_X32 FILLER_212_1272 ();
 FILLCELL_X32 FILLER_212_1304 ();
 FILLCELL_X32 FILLER_212_1336 ();
 FILLCELL_X32 FILLER_212_1368 ();
 FILLCELL_X32 FILLER_212_1400 ();
 FILLCELL_X32 FILLER_212_1432 ();
 FILLCELL_X32 FILLER_212_1464 ();
 FILLCELL_X32 FILLER_212_1496 ();
 FILLCELL_X32 FILLER_212_1528 ();
 FILLCELL_X32 FILLER_212_1560 ();
 FILLCELL_X32 FILLER_212_1592 ();
 FILLCELL_X32 FILLER_212_1624 ();
 FILLCELL_X32 FILLER_212_1656 ();
 FILLCELL_X32 FILLER_212_1688 ();
 FILLCELL_X16 FILLER_212_1720 ();
 FILLCELL_X8 FILLER_212_1736 ();
 FILLCELL_X1 FILLER_212_1744 ();
 FILLCELL_X4 FILLER_212_1752 ();
 FILLCELL_X32 FILLER_213_1 ();
 FILLCELL_X32 FILLER_213_33 ();
 FILLCELL_X32 FILLER_213_65 ();
 FILLCELL_X32 FILLER_213_97 ();
 FILLCELL_X32 FILLER_213_129 ();
 FILLCELL_X32 FILLER_213_161 ();
 FILLCELL_X32 FILLER_213_193 ();
 FILLCELL_X32 FILLER_213_225 ();
 FILLCELL_X32 FILLER_213_257 ();
 FILLCELL_X32 FILLER_213_289 ();
 FILLCELL_X32 FILLER_213_321 ();
 FILLCELL_X32 FILLER_213_353 ();
 FILLCELL_X32 FILLER_213_385 ();
 FILLCELL_X32 FILLER_213_417 ();
 FILLCELL_X32 FILLER_213_449 ();
 FILLCELL_X32 FILLER_213_481 ();
 FILLCELL_X32 FILLER_213_513 ();
 FILLCELL_X32 FILLER_213_545 ();
 FILLCELL_X32 FILLER_213_577 ();
 FILLCELL_X32 FILLER_213_609 ();
 FILLCELL_X32 FILLER_213_641 ();
 FILLCELL_X32 FILLER_213_673 ();
 FILLCELL_X32 FILLER_213_705 ();
 FILLCELL_X32 FILLER_213_737 ();
 FILLCELL_X32 FILLER_213_769 ();
 FILLCELL_X32 FILLER_213_801 ();
 FILLCELL_X32 FILLER_213_833 ();
 FILLCELL_X32 FILLER_213_865 ();
 FILLCELL_X32 FILLER_213_897 ();
 FILLCELL_X32 FILLER_213_929 ();
 FILLCELL_X32 FILLER_213_961 ();
 FILLCELL_X32 FILLER_213_993 ();
 FILLCELL_X32 FILLER_213_1025 ();
 FILLCELL_X32 FILLER_213_1057 ();
 FILLCELL_X32 FILLER_213_1089 ();
 FILLCELL_X32 FILLER_213_1121 ();
 FILLCELL_X32 FILLER_213_1153 ();
 FILLCELL_X32 FILLER_213_1185 ();
 FILLCELL_X32 FILLER_213_1217 ();
 FILLCELL_X8 FILLER_213_1249 ();
 FILLCELL_X4 FILLER_213_1257 ();
 FILLCELL_X2 FILLER_213_1261 ();
 FILLCELL_X32 FILLER_213_1264 ();
 FILLCELL_X32 FILLER_213_1296 ();
 FILLCELL_X32 FILLER_213_1328 ();
 FILLCELL_X32 FILLER_213_1360 ();
 FILLCELL_X32 FILLER_213_1392 ();
 FILLCELL_X32 FILLER_213_1424 ();
 FILLCELL_X32 FILLER_213_1456 ();
 FILLCELL_X32 FILLER_213_1488 ();
 FILLCELL_X32 FILLER_213_1520 ();
 FILLCELL_X32 FILLER_213_1552 ();
 FILLCELL_X32 FILLER_213_1584 ();
 FILLCELL_X32 FILLER_213_1616 ();
 FILLCELL_X32 FILLER_213_1648 ();
 FILLCELL_X32 FILLER_213_1680 ();
 FILLCELL_X32 FILLER_213_1712 ();
 FILLCELL_X8 FILLER_213_1744 ();
 FILLCELL_X4 FILLER_213_1752 ();
 FILLCELL_X32 FILLER_214_1 ();
 FILLCELL_X32 FILLER_214_33 ();
 FILLCELL_X32 FILLER_214_65 ();
 FILLCELL_X32 FILLER_214_97 ();
 FILLCELL_X32 FILLER_214_129 ();
 FILLCELL_X32 FILLER_214_161 ();
 FILLCELL_X32 FILLER_214_193 ();
 FILLCELL_X32 FILLER_214_225 ();
 FILLCELL_X32 FILLER_214_257 ();
 FILLCELL_X32 FILLER_214_289 ();
 FILLCELL_X32 FILLER_214_321 ();
 FILLCELL_X32 FILLER_214_353 ();
 FILLCELL_X32 FILLER_214_385 ();
 FILLCELL_X32 FILLER_214_417 ();
 FILLCELL_X32 FILLER_214_449 ();
 FILLCELL_X32 FILLER_214_481 ();
 FILLCELL_X32 FILLER_214_513 ();
 FILLCELL_X32 FILLER_214_545 ();
 FILLCELL_X32 FILLER_214_577 ();
 FILLCELL_X16 FILLER_214_609 ();
 FILLCELL_X4 FILLER_214_625 ();
 FILLCELL_X2 FILLER_214_629 ();
 FILLCELL_X32 FILLER_214_632 ();
 FILLCELL_X32 FILLER_214_664 ();
 FILLCELL_X32 FILLER_214_696 ();
 FILLCELL_X32 FILLER_214_728 ();
 FILLCELL_X32 FILLER_214_760 ();
 FILLCELL_X32 FILLER_214_792 ();
 FILLCELL_X32 FILLER_214_824 ();
 FILLCELL_X32 FILLER_214_856 ();
 FILLCELL_X32 FILLER_214_888 ();
 FILLCELL_X32 FILLER_214_920 ();
 FILLCELL_X32 FILLER_214_952 ();
 FILLCELL_X32 FILLER_214_984 ();
 FILLCELL_X32 FILLER_214_1016 ();
 FILLCELL_X32 FILLER_214_1048 ();
 FILLCELL_X32 FILLER_214_1080 ();
 FILLCELL_X32 FILLER_214_1112 ();
 FILLCELL_X32 FILLER_214_1144 ();
 FILLCELL_X32 FILLER_214_1176 ();
 FILLCELL_X32 FILLER_214_1208 ();
 FILLCELL_X32 FILLER_214_1240 ();
 FILLCELL_X32 FILLER_214_1272 ();
 FILLCELL_X32 FILLER_214_1304 ();
 FILLCELL_X32 FILLER_214_1336 ();
 FILLCELL_X32 FILLER_214_1368 ();
 FILLCELL_X32 FILLER_214_1400 ();
 FILLCELL_X32 FILLER_214_1432 ();
 FILLCELL_X32 FILLER_214_1464 ();
 FILLCELL_X32 FILLER_214_1496 ();
 FILLCELL_X32 FILLER_214_1528 ();
 FILLCELL_X32 FILLER_214_1560 ();
 FILLCELL_X32 FILLER_214_1592 ();
 FILLCELL_X32 FILLER_214_1624 ();
 FILLCELL_X32 FILLER_214_1656 ();
 FILLCELL_X32 FILLER_214_1688 ();
 FILLCELL_X32 FILLER_214_1720 ();
 FILLCELL_X4 FILLER_214_1752 ();
 FILLCELL_X32 FILLER_215_1 ();
 FILLCELL_X32 FILLER_215_33 ();
 FILLCELL_X32 FILLER_215_65 ();
 FILLCELL_X32 FILLER_215_97 ();
 FILLCELL_X32 FILLER_215_129 ();
 FILLCELL_X32 FILLER_215_161 ();
 FILLCELL_X32 FILLER_215_193 ();
 FILLCELL_X32 FILLER_215_225 ();
 FILLCELL_X32 FILLER_215_257 ();
 FILLCELL_X32 FILLER_215_289 ();
 FILLCELL_X32 FILLER_215_321 ();
 FILLCELL_X32 FILLER_215_353 ();
 FILLCELL_X32 FILLER_215_385 ();
 FILLCELL_X32 FILLER_215_417 ();
 FILLCELL_X32 FILLER_215_449 ();
 FILLCELL_X32 FILLER_215_481 ();
 FILLCELL_X32 FILLER_215_513 ();
 FILLCELL_X32 FILLER_215_545 ();
 FILLCELL_X32 FILLER_215_577 ();
 FILLCELL_X32 FILLER_215_609 ();
 FILLCELL_X32 FILLER_215_641 ();
 FILLCELL_X32 FILLER_215_673 ();
 FILLCELL_X32 FILLER_215_705 ();
 FILLCELL_X32 FILLER_215_737 ();
 FILLCELL_X32 FILLER_215_769 ();
 FILLCELL_X32 FILLER_215_801 ();
 FILLCELL_X32 FILLER_215_833 ();
 FILLCELL_X32 FILLER_215_865 ();
 FILLCELL_X32 FILLER_215_897 ();
 FILLCELL_X32 FILLER_215_929 ();
 FILLCELL_X32 FILLER_215_961 ();
 FILLCELL_X32 FILLER_215_993 ();
 FILLCELL_X32 FILLER_215_1025 ();
 FILLCELL_X32 FILLER_215_1057 ();
 FILLCELL_X32 FILLER_215_1089 ();
 FILLCELL_X32 FILLER_215_1121 ();
 FILLCELL_X32 FILLER_215_1153 ();
 FILLCELL_X32 FILLER_215_1185 ();
 FILLCELL_X32 FILLER_215_1217 ();
 FILLCELL_X8 FILLER_215_1249 ();
 FILLCELL_X4 FILLER_215_1257 ();
 FILLCELL_X2 FILLER_215_1261 ();
 FILLCELL_X32 FILLER_215_1264 ();
 FILLCELL_X32 FILLER_215_1296 ();
 FILLCELL_X32 FILLER_215_1328 ();
 FILLCELL_X32 FILLER_215_1360 ();
 FILLCELL_X32 FILLER_215_1392 ();
 FILLCELL_X32 FILLER_215_1424 ();
 FILLCELL_X32 FILLER_215_1456 ();
 FILLCELL_X32 FILLER_215_1488 ();
 FILLCELL_X32 FILLER_215_1520 ();
 FILLCELL_X32 FILLER_215_1552 ();
 FILLCELL_X32 FILLER_215_1584 ();
 FILLCELL_X32 FILLER_215_1616 ();
 FILLCELL_X32 FILLER_215_1648 ();
 FILLCELL_X32 FILLER_215_1680 ();
 FILLCELL_X32 FILLER_215_1712 ();
 FILLCELL_X8 FILLER_215_1744 ();
 FILLCELL_X4 FILLER_215_1752 ();
 FILLCELL_X32 FILLER_216_1 ();
 FILLCELL_X32 FILLER_216_33 ();
 FILLCELL_X32 FILLER_216_65 ();
 FILLCELL_X32 FILLER_216_97 ();
 FILLCELL_X32 FILLER_216_129 ();
 FILLCELL_X32 FILLER_216_161 ();
 FILLCELL_X32 FILLER_216_193 ();
 FILLCELL_X32 FILLER_216_225 ();
 FILLCELL_X32 FILLER_216_257 ();
 FILLCELL_X32 FILLER_216_289 ();
 FILLCELL_X32 FILLER_216_321 ();
 FILLCELL_X32 FILLER_216_353 ();
 FILLCELL_X32 FILLER_216_385 ();
 FILLCELL_X32 FILLER_216_417 ();
 FILLCELL_X32 FILLER_216_449 ();
 FILLCELL_X32 FILLER_216_481 ();
 FILLCELL_X32 FILLER_216_513 ();
 FILLCELL_X32 FILLER_216_545 ();
 FILLCELL_X32 FILLER_216_577 ();
 FILLCELL_X16 FILLER_216_609 ();
 FILLCELL_X4 FILLER_216_625 ();
 FILLCELL_X2 FILLER_216_629 ();
 FILLCELL_X32 FILLER_216_632 ();
 FILLCELL_X32 FILLER_216_664 ();
 FILLCELL_X32 FILLER_216_696 ();
 FILLCELL_X32 FILLER_216_728 ();
 FILLCELL_X32 FILLER_216_760 ();
 FILLCELL_X32 FILLER_216_792 ();
 FILLCELL_X32 FILLER_216_824 ();
 FILLCELL_X32 FILLER_216_856 ();
 FILLCELL_X32 FILLER_216_888 ();
 FILLCELL_X32 FILLER_216_920 ();
 FILLCELL_X32 FILLER_216_952 ();
 FILLCELL_X32 FILLER_216_984 ();
 FILLCELL_X32 FILLER_216_1016 ();
 FILLCELL_X32 FILLER_216_1048 ();
 FILLCELL_X32 FILLER_216_1080 ();
 FILLCELL_X32 FILLER_216_1112 ();
 FILLCELL_X32 FILLER_216_1144 ();
 FILLCELL_X32 FILLER_216_1176 ();
 FILLCELL_X32 FILLER_216_1208 ();
 FILLCELL_X32 FILLER_216_1240 ();
 FILLCELL_X32 FILLER_216_1272 ();
 FILLCELL_X32 FILLER_216_1304 ();
 FILLCELL_X32 FILLER_216_1336 ();
 FILLCELL_X32 FILLER_216_1368 ();
 FILLCELL_X32 FILLER_216_1400 ();
 FILLCELL_X32 FILLER_216_1432 ();
 FILLCELL_X32 FILLER_216_1464 ();
 FILLCELL_X32 FILLER_216_1496 ();
 FILLCELL_X32 FILLER_216_1528 ();
 FILLCELL_X32 FILLER_216_1560 ();
 FILLCELL_X32 FILLER_216_1592 ();
 FILLCELL_X32 FILLER_216_1624 ();
 FILLCELL_X32 FILLER_216_1656 ();
 FILLCELL_X32 FILLER_216_1688 ();
 FILLCELL_X32 FILLER_216_1720 ();
 FILLCELL_X4 FILLER_216_1752 ();
 FILLCELL_X4 FILLER_217_1 ();
 FILLCELL_X32 FILLER_217_10 ();
 FILLCELL_X32 FILLER_217_42 ();
 FILLCELL_X32 FILLER_217_74 ();
 FILLCELL_X32 FILLER_217_106 ();
 FILLCELL_X32 FILLER_217_138 ();
 FILLCELL_X32 FILLER_217_170 ();
 FILLCELL_X32 FILLER_217_202 ();
 FILLCELL_X32 FILLER_217_234 ();
 FILLCELL_X32 FILLER_217_266 ();
 FILLCELL_X32 FILLER_217_298 ();
 FILLCELL_X32 FILLER_217_330 ();
 FILLCELL_X32 FILLER_217_362 ();
 FILLCELL_X32 FILLER_217_394 ();
 FILLCELL_X32 FILLER_217_426 ();
 FILLCELL_X32 FILLER_217_458 ();
 FILLCELL_X32 FILLER_217_490 ();
 FILLCELL_X32 FILLER_217_522 ();
 FILLCELL_X32 FILLER_217_554 ();
 FILLCELL_X32 FILLER_217_586 ();
 FILLCELL_X32 FILLER_217_618 ();
 FILLCELL_X32 FILLER_217_650 ();
 FILLCELL_X32 FILLER_217_682 ();
 FILLCELL_X32 FILLER_217_714 ();
 FILLCELL_X32 FILLER_217_746 ();
 FILLCELL_X32 FILLER_217_778 ();
 FILLCELL_X32 FILLER_217_810 ();
 FILLCELL_X32 FILLER_217_842 ();
 FILLCELL_X32 FILLER_217_874 ();
 FILLCELL_X32 FILLER_217_906 ();
 FILLCELL_X32 FILLER_217_938 ();
 FILLCELL_X32 FILLER_217_970 ();
 FILLCELL_X32 FILLER_217_1002 ();
 FILLCELL_X32 FILLER_217_1034 ();
 FILLCELL_X32 FILLER_217_1066 ();
 FILLCELL_X32 FILLER_217_1098 ();
 FILLCELL_X32 FILLER_217_1130 ();
 FILLCELL_X32 FILLER_217_1162 ();
 FILLCELL_X32 FILLER_217_1194 ();
 FILLCELL_X32 FILLER_217_1226 ();
 FILLCELL_X4 FILLER_217_1258 ();
 FILLCELL_X1 FILLER_217_1262 ();
 FILLCELL_X32 FILLER_217_1264 ();
 FILLCELL_X32 FILLER_217_1296 ();
 FILLCELL_X32 FILLER_217_1328 ();
 FILLCELL_X32 FILLER_217_1360 ();
 FILLCELL_X32 FILLER_217_1392 ();
 FILLCELL_X32 FILLER_217_1424 ();
 FILLCELL_X32 FILLER_217_1456 ();
 FILLCELL_X32 FILLER_217_1488 ();
 FILLCELL_X32 FILLER_217_1520 ();
 FILLCELL_X32 FILLER_217_1552 ();
 FILLCELL_X32 FILLER_217_1584 ();
 FILLCELL_X32 FILLER_217_1616 ();
 FILLCELL_X32 FILLER_217_1648 ();
 FILLCELL_X32 FILLER_217_1680 ();
 FILLCELL_X32 FILLER_217_1712 ();
 FILLCELL_X8 FILLER_217_1744 ();
 FILLCELL_X4 FILLER_217_1752 ();
 FILLCELL_X32 FILLER_218_1 ();
 FILLCELL_X32 FILLER_218_33 ();
 FILLCELL_X32 FILLER_218_65 ();
 FILLCELL_X32 FILLER_218_97 ();
 FILLCELL_X32 FILLER_218_129 ();
 FILLCELL_X32 FILLER_218_161 ();
 FILLCELL_X32 FILLER_218_193 ();
 FILLCELL_X32 FILLER_218_225 ();
 FILLCELL_X32 FILLER_218_257 ();
 FILLCELL_X32 FILLER_218_289 ();
 FILLCELL_X32 FILLER_218_321 ();
 FILLCELL_X32 FILLER_218_353 ();
 FILLCELL_X32 FILLER_218_385 ();
 FILLCELL_X32 FILLER_218_417 ();
 FILLCELL_X32 FILLER_218_449 ();
 FILLCELL_X32 FILLER_218_481 ();
 FILLCELL_X32 FILLER_218_513 ();
 FILLCELL_X32 FILLER_218_545 ();
 FILLCELL_X32 FILLER_218_577 ();
 FILLCELL_X16 FILLER_218_609 ();
 FILLCELL_X4 FILLER_218_625 ();
 FILLCELL_X2 FILLER_218_629 ();
 FILLCELL_X32 FILLER_218_632 ();
 FILLCELL_X32 FILLER_218_664 ();
 FILLCELL_X32 FILLER_218_696 ();
 FILLCELL_X32 FILLER_218_728 ();
 FILLCELL_X32 FILLER_218_760 ();
 FILLCELL_X32 FILLER_218_792 ();
 FILLCELL_X32 FILLER_218_824 ();
 FILLCELL_X32 FILLER_218_856 ();
 FILLCELL_X32 FILLER_218_888 ();
 FILLCELL_X32 FILLER_218_920 ();
 FILLCELL_X32 FILLER_218_952 ();
 FILLCELL_X32 FILLER_218_984 ();
 FILLCELL_X32 FILLER_218_1016 ();
 FILLCELL_X32 FILLER_218_1048 ();
 FILLCELL_X32 FILLER_218_1080 ();
 FILLCELL_X32 FILLER_218_1112 ();
 FILLCELL_X32 FILLER_218_1144 ();
 FILLCELL_X32 FILLER_218_1176 ();
 FILLCELL_X32 FILLER_218_1208 ();
 FILLCELL_X32 FILLER_218_1240 ();
 FILLCELL_X32 FILLER_218_1272 ();
 FILLCELL_X32 FILLER_218_1304 ();
 FILLCELL_X32 FILLER_218_1336 ();
 FILLCELL_X32 FILLER_218_1368 ();
 FILLCELL_X32 FILLER_218_1400 ();
 FILLCELL_X32 FILLER_218_1432 ();
 FILLCELL_X32 FILLER_218_1464 ();
 FILLCELL_X32 FILLER_218_1496 ();
 FILLCELL_X32 FILLER_218_1528 ();
 FILLCELL_X32 FILLER_218_1560 ();
 FILLCELL_X32 FILLER_218_1592 ();
 FILLCELL_X32 FILLER_218_1624 ();
 FILLCELL_X32 FILLER_218_1656 ();
 FILLCELL_X32 FILLER_218_1688 ();
 FILLCELL_X32 FILLER_218_1720 ();
 FILLCELL_X4 FILLER_218_1752 ();
 FILLCELL_X32 FILLER_219_1 ();
 FILLCELL_X32 FILLER_219_33 ();
 FILLCELL_X32 FILLER_219_65 ();
 FILLCELL_X32 FILLER_219_97 ();
 FILLCELL_X32 FILLER_219_129 ();
 FILLCELL_X32 FILLER_219_161 ();
 FILLCELL_X32 FILLER_219_193 ();
 FILLCELL_X32 FILLER_219_225 ();
 FILLCELL_X32 FILLER_219_257 ();
 FILLCELL_X32 FILLER_219_289 ();
 FILLCELL_X32 FILLER_219_321 ();
 FILLCELL_X32 FILLER_219_353 ();
 FILLCELL_X32 FILLER_219_385 ();
 FILLCELL_X32 FILLER_219_417 ();
 FILLCELL_X32 FILLER_219_449 ();
 FILLCELL_X32 FILLER_219_481 ();
 FILLCELL_X32 FILLER_219_513 ();
 FILLCELL_X32 FILLER_219_545 ();
 FILLCELL_X32 FILLER_219_577 ();
 FILLCELL_X32 FILLER_219_609 ();
 FILLCELL_X32 FILLER_219_641 ();
 FILLCELL_X32 FILLER_219_673 ();
 FILLCELL_X32 FILLER_219_705 ();
 FILLCELL_X32 FILLER_219_737 ();
 FILLCELL_X32 FILLER_219_769 ();
 FILLCELL_X32 FILLER_219_801 ();
 FILLCELL_X32 FILLER_219_833 ();
 FILLCELL_X32 FILLER_219_865 ();
 FILLCELL_X32 FILLER_219_897 ();
 FILLCELL_X32 FILLER_219_929 ();
 FILLCELL_X32 FILLER_219_961 ();
 FILLCELL_X32 FILLER_219_993 ();
 FILLCELL_X32 FILLER_219_1025 ();
 FILLCELL_X32 FILLER_219_1057 ();
 FILLCELL_X32 FILLER_219_1089 ();
 FILLCELL_X32 FILLER_219_1121 ();
 FILLCELL_X32 FILLER_219_1153 ();
 FILLCELL_X32 FILLER_219_1185 ();
 FILLCELL_X32 FILLER_219_1217 ();
 FILLCELL_X8 FILLER_219_1249 ();
 FILLCELL_X4 FILLER_219_1257 ();
 FILLCELL_X2 FILLER_219_1261 ();
 FILLCELL_X32 FILLER_219_1264 ();
 FILLCELL_X32 FILLER_219_1296 ();
 FILLCELL_X32 FILLER_219_1328 ();
 FILLCELL_X32 FILLER_219_1360 ();
 FILLCELL_X32 FILLER_219_1392 ();
 FILLCELL_X32 FILLER_219_1424 ();
 FILLCELL_X32 FILLER_219_1456 ();
 FILLCELL_X32 FILLER_219_1488 ();
 FILLCELL_X32 FILLER_219_1520 ();
 FILLCELL_X32 FILLER_219_1552 ();
 FILLCELL_X32 FILLER_219_1584 ();
 FILLCELL_X32 FILLER_219_1616 ();
 FILLCELL_X32 FILLER_219_1648 ();
 FILLCELL_X32 FILLER_219_1680 ();
 FILLCELL_X32 FILLER_219_1712 ();
 FILLCELL_X8 FILLER_219_1744 ();
 FILLCELL_X4 FILLER_219_1752 ();
 FILLCELL_X32 FILLER_220_1 ();
 FILLCELL_X32 FILLER_220_33 ();
 FILLCELL_X32 FILLER_220_65 ();
 FILLCELL_X32 FILLER_220_97 ();
 FILLCELL_X32 FILLER_220_129 ();
 FILLCELL_X32 FILLER_220_161 ();
 FILLCELL_X32 FILLER_220_193 ();
 FILLCELL_X32 FILLER_220_225 ();
 FILLCELL_X32 FILLER_220_257 ();
 FILLCELL_X32 FILLER_220_289 ();
 FILLCELL_X32 FILLER_220_321 ();
 FILLCELL_X32 FILLER_220_353 ();
 FILLCELL_X32 FILLER_220_385 ();
 FILLCELL_X32 FILLER_220_417 ();
 FILLCELL_X32 FILLER_220_449 ();
 FILLCELL_X32 FILLER_220_481 ();
 FILLCELL_X32 FILLER_220_513 ();
 FILLCELL_X32 FILLER_220_545 ();
 FILLCELL_X32 FILLER_220_577 ();
 FILLCELL_X16 FILLER_220_609 ();
 FILLCELL_X4 FILLER_220_625 ();
 FILLCELL_X2 FILLER_220_629 ();
 FILLCELL_X32 FILLER_220_632 ();
 FILLCELL_X32 FILLER_220_664 ();
 FILLCELL_X32 FILLER_220_696 ();
 FILLCELL_X32 FILLER_220_728 ();
 FILLCELL_X32 FILLER_220_760 ();
 FILLCELL_X32 FILLER_220_792 ();
 FILLCELL_X32 FILLER_220_824 ();
 FILLCELL_X32 FILLER_220_856 ();
 FILLCELL_X32 FILLER_220_888 ();
 FILLCELL_X32 FILLER_220_920 ();
 FILLCELL_X32 FILLER_220_952 ();
 FILLCELL_X32 FILLER_220_984 ();
 FILLCELL_X32 FILLER_220_1016 ();
 FILLCELL_X32 FILLER_220_1048 ();
 FILLCELL_X32 FILLER_220_1080 ();
 FILLCELL_X32 FILLER_220_1112 ();
 FILLCELL_X32 FILLER_220_1144 ();
 FILLCELL_X32 FILLER_220_1176 ();
 FILLCELL_X32 FILLER_220_1208 ();
 FILLCELL_X32 FILLER_220_1240 ();
 FILLCELL_X32 FILLER_220_1272 ();
 FILLCELL_X32 FILLER_220_1304 ();
 FILLCELL_X32 FILLER_220_1336 ();
 FILLCELL_X32 FILLER_220_1368 ();
 FILLCELL_X32 FILLER_220_1400 ();
 FILLCELL_X32 FILLER_220_1432 ();
 FILLCELL_X32 FILLER_220_1464 ();
 FILLCELL_X32 FILLER_220_1496 ();
 FILLCELL_X32 FILLER_220_1528 ();
 FILLCELL_X32 FILLER_220_1560 ();
 FILLCELL_X32 FILLER_220_1592 ();
 FILLCELL_X32 FILLER_220_1624 ();
 FILLCELL_X32 FILLER_220_1656 ();
 FILLCELL_X32 FILLER_220_1688 ();
 FILLCELL_X32 FILLER_220_1720 ();
 FILLCELL_X4 FILLER_220_1752 ();
 FILLCELL_X32 FILLER_221_1 ();
 FILLCELL_X32 FILLER_221_33 ();
 FILLCELL_X32 FILLER_221_65 ();
 FILLCELL_X32 FILLER_221_97 ();
 FILLCELL_X32 FILLER_221_129 ();
 FILLCELL_X32 FILLER_221_161 ();
 FILLCELL_X32 FILLER_221_193 ();
 FILLCELL_X32 FILLER_221_225 ();
 FILLCELL_X32 FILLER_221_257 ();
 FILLCELL_X32 FILLER_221_289 ();
 FILLCELL_X32 FILLER_221_321 ();
 FILLCELL_X32 FILLER_221_353 ();
 FILLCELL_X32 FILLER_221_385 ();
 FILLCELL_X32 FILLER_221_417 ();
 FILLCELL_X32 FILLER_221_449 ();
 FILLCELL_X32 FILLER_221_481 ();
 FILLCELL_X32 FILLER_221_513 ();
 FILLCELL_X32 FILLER_221_545 ();
 FILLCELL_X32 FILLER_221_577 ();
 FILLCELL_X32 FILLER_221_609 ();
 FILLCELL_X32 FILLER_221_641 ();
 FILLCELL_X32 FILLER_221_673 ();
 FILLCELL_X32 FILLER_221_705 ();
 FILLCELL_X32 FILLER_221_737 ();
 FILLCELL_X32 FILLER_221_769 ();
 FILLCELL_X32 FILLER_221_801 ();
 FILLCELL_X32 FILLER_221_833 ();
 FILLCELL_X32 FILLER_221_865 ();
 FILLCELL_X32 FILLER_221_897 ();
 FILLCELL_X32 FILLER_221_929 ();
 FILLCELL_X32 FILLER_221_961 ();
 FILLCELL_X32 FILLER_221_993 ();
 FILLCELL_X32 FILLER_221_1025 ();
 FILLCELL_X32 FILLER_221_1057 ();
 FILLCELL_X32 FILLER_221_1089 ();
 FILLCELL_X32 FILLER_221_1121 ();
 FILLCELL_X32 FILLER_221_1153 ();
 FILLCELL_X32 FILLER_221_1185 ();
 FILLCELL_X32 FILLER_221_1217 ();
 FILLCELL_X8 FILLER_221_1249 ();
 FILLCELL_X4 FILLER_221_1257 ();
 FILLCELL_X2 FILLER_221_1261 ();
 FILLCELL_X32 FILLER_221_1264 ();
 FILLCELL_X32 FILLER_221_1296 ();
 FILLCELL_X32 FILLER_221_1328 ();
 FILLCELL_X32 FILLER_221_1360 ();
 FILLCELL_X32 FILLER_221_1392 ();
 FILLCELL_X32 FILLER_221_1424 ();
 FILLCELL_X32 FILLER_221_1456 ();
 FILLCELL_X32 FILLER_221_1488 ();
 FILLCELL_X32 FILLER_221_1520 ();
 FILLCELL_X32 FILLER_221_1552 ();
 FILLCELL_X32 FILLER_221_1584 ();
 FILLCELL_X32 FILLER_221_1616 ();
 FILLCELL_X32 FILLER_221_1648 ();
 FILLCELL_X32 FILLER_221_1680 ();
 FILLCELL_X32 FILLER_221_1712 ();
 FILLCELL_X8 FILLER_221_1744 ();
 FILLCELL_X4 FILLER_221_1752 ();
 FILLCELL_X32 FILLER_222_1 ();
 FILLCELL_X32 FILLER_222_33 ();
 FILLCELL_X32 FILLER_222_65 ();
 FILLCELL_X32 FILLER_222_97 ();
 FILLCELL_X32 FILLER_222_129 ();
 FILLCELL_X32 FILLER_222_161 ();
 FILLCELL_X32 FILLER_222_193 ();
 FILLCELL_X32 FILLER_222_225 ();
 FILLCELL_X32 FILLER_222_257 ();
 FILLCELL_X32 FILLER_222_289 ();
 FILLCELL_X32 FILLER_222_321 ();
 FILLCELL_X32 FILLER_222_353 ();
 FILLCELL_X32 FILLER_222_385 ();
 FILLCELL_X32 FILLER_222_417 ();
 FILLCELL_X32 FILLER_222_449 ();
 FILLCELL_X32 FILLER_222_481 ();
 FILLCELL_X32 FILLER_222_513 ();
 FILLCELL_X32 FILLER_222_545 ();
 FILLCELL_X32 FILLER_222_577 ();
 FILLCELL_X16 FILLER_222_609 ();
 FILLCELL_X4 FILLER_222_625 ();
 FILLCELL_X2 FILLER_222_629 ();
 FILLCELL_X32 FILLER_222_632 ();
 FILLCELL_X32 FILLER_222_664 ();
 FILLCELL_X32 FILLER_222_696 ();
 FILLCELL_X32 FILLER_222_728 ();
 FILLCELL_X32 FILLER_222_760 ();
 FILLCELL_X32 FILLER_222_792 ();
 FILLCELL_X32 FILLER_222_824 ();
 FILLCELL_X32 FILLER_222_856 ();
 FILLCELL_X32 FILLER_222_888 ();
 FILLCELL_X32 FILLER_222_920 ();
 FILLCELL_X32 FILLER_222_952 ();
 FILLCELL_X32 FILLER_222_984 ();
 FILLCELL_X32 FILLER_222_1016 ();
 FILLCELL_X32 FILLER_222_1048 ();
 FILLCELL_X32 FILLER_222_1080 ();
 FILLCELL_X32 FILLER_222_1112 ();
 FILLCELL_X32 FILLER_222_1144 ();
 FILLCELL_X32 FILLER_222_1176 ();
 FILLCELL_X32 FILLER_222_1208 ();
 FILLCELL_X32 FILLER_222_1240 ();
 FILLCELL_X32 FILLER_222_1272 ();
 FILLCELL_X32 FILLER_222_1304 ();
 FILLCELL_X32 FILLER_222_1336 ();
 FILLCELL_X32 FILLER_222_1368 ();
 FILLCELL_X32 FILLER_222_1400 ();
 FILLCELL_X32 FILLER_222_1432 ();
 FILLCELL_X32 FILLER_222_1464 ();
 FILLCELL_X32 FILLER_222_1496 ();
 FILLCELL_X32 FILLER_222_1528 ();
 FILLCELL_X32 FILLER_222_1560 ();
 FILLCELL_X32 FILLER_222_1592 ();
 FILLCELL_X32 FILLER_222_1624 ();
 FILLCELL_X32 FILLER_222_1656 ();
 FILLCELL_X32 FILLER_222_1688 ();
 FILLCELL_X16 FILLER_222_1720 ();
 FILLCELL_X8 FILLER_222_1736 ();
 FILLCELL_X2 FILLER_222_1744 ();
 FILLCELL_X1 FILLER_222_1746 ();
 FILLCELL_X4 FILLER_222_1752 ();
 FILLCELL_X32 FILLER_223_1 ();
 FILLCELL_X32 FILLER_223_33 ();
 FILLCELL_X32 FILLER_223_65 ();
 FILLCELL_X32 FILLER_223_97 ();
 FILLCELL_X32 FILLER_223_129 ();
 FILLCELL_X32 FILLER_223_161 ();
 FILLCELL_X32 FILLER_223_193 ();
 FILLCELL_X32 FILLER_223_225 ();
 FILLCELL_X32 FILLER_223_257 ();
 FILLCELL_X32 FILLER_223_289 ();
 FILLCELL_X32 FILLER_223_321 ();
 FILLCELL_X32 FILLER_223_353 ();
 FILLCELL_X32 FILLER_223_385 ();
 FILLCELL_X32 FILLER_223_417 ();
 FILLCELL_X32 FILLER_223_449 ();
 FILLCELL_X32 FILLER_223_481 ();
 FILLCELL_X32 FILLER_223_513 ();
 FILLCELL_X32 FILLER_223_545 ();
 FILLCELL_X32 FILLER_223_577 ();
 FILLCELL_X32 FILLER_223_609 ();
 FILLCELL_X32 FILLER_223_641 ();
 FILLCELL_X32 FILLER_223_673 ();
 FILLCELL_X32 FILLER_223_705 ();
 FILLCELL_X32 FILLER_223_737 ();
 FILLCELL_X32 FILLER_223_769 ();
 FILLCELL_X32 FILLER_223_801 ();
 FILLCELL_X32 FILLER_223_833 ();
 FILLCELL_X32 FILLER_223_865 ();
 FILLCELL_X32 FILLER_223_897 ();
 FILLCELL_X32 FILLER_223_929 ();
 FILLCELL_X32 FILLER_223_961 ();
 FILLCELL_X32 FILLER_223_993 ();
 FILLCELL_X32 FILLER_223_1025 ();
 FILLCELL_X32 FILLER_223_1057 ();
 FILLCELL_X32 FILLER_223_1089 ();
 FILLCELL_X32 FILLER_223_1121 ();
 FILLCELL_X32 FILLER_223_1153 ();
 FILLCELL_X32 FILLER_223_1185 ();
 FILLCELL_X32 FILLER_223_1217 ();
 FILLCELL_X8 FILLER_223_1249 ();
 FILLCELL_X4 FILLER_223_1257 ();
 FILLCELL_X2 FILLER_223_1261 ();
 FILLCELL_X32 FILLER_223_1264 ();
 FILLCELL_X32 FILLER_223_1296 ();
 FILLCELL_X32 FILLER_223_1328 ();
 FILLCELL_X32 FILLER_223_1360 ();
 FILLCELL_X32 FILLER_223_1392 ();
 FILLCELL_X32 FILLER_223_1424 ();
 FILLCELL_X32 FILLER_223_1456 ();
 FILLCELL_X32 FILLER_223_1488 ();
 FILLCELL_X32 FILLER_223_1520 ();
 FILLCELL_X32 FILLER_223_1552 ();
 FILLCELL_X32 FILLER_223_1584 ();
 FILLCELL_X32 FILLER_223_1616 ();
 FILLCELL_X32 FILLER_223_1648 ();
 FILLCELL_X32 FILLER_223_1680 ();
 FILLCELL_X32 FILLER_223_1712 ();
 FILLCELL_X8 FILLER_223_1744 ();
 FILLCELL_X4 FILLER_223_1752 ();
 FILLCELL_X32 FILLER_224_1 ();
 FILLCELL_X32 FILLER_224_33 ();
 FILLCELL_X32 FILLER_224_65 ();
 FILLCELL_X32 FILLER_224_97 ();
 FILLCELL_X32 FILLER_224_129 ();
 FILLCELL_X32 FILLER_224_161 ();
 FILLCELL_X32 FILLER_224_193 ();
 FILLCELL_X32 FILLER_224_225 ();
 FILLCELL_X32 FILLER_224_257 ();
 FILLCELL_X32 FILLER_224_289 ();
 FILLCELL_X32 FILLER_224_321 ();
 FILLCELL_X32 FILLER_224_353 ();
 FILLCELL_X32 FILLER_224_385 ();
 FILLCELL_X32 FILLER_224_417 ();
 FILLCELL_X32 FILLER_224_449 ();
 FILLCELL_X32 FILLER_224_481 ();
 FILLCELL_X32 FILLER_224_513 ();
 FILLCELL_X32 FILLER_224_545 ();
 FILLCELL_X32 FILLER_224_577 ();
 FILLCELL_X16 FILLER_224_609 ();
 FILLCELL_X4 FILLER_224_625 ();
 FILLCELL_X2 FILLER_224_629 ();
 FILLCELL_X32 FILLER_224_632 ();
 FILLCELL_X32 FILLER_224_664 ();
 FILLCELL_X32 FILLER_224_696 ();
 FILLCELL_X32 FILLER_224_728 ();
 FILLCELL_X32 FILLER_224_760 ();
 FILLCELL_X32 FILLER_224_792 ();
 FILLCELL_X32 FILLER_224_824 ();
 FILLCELL_X32 FILLER_224_856 ();
 FILLCELL_X32 FILLER_224_888 ();
 FILLCELL_X32 FILLER_224_920 ();
 FILLCELL_X32 FILLER_224_952 ();
 FILLCELL_X32 FILLER_224_984 ();
 FILLCELL_X32 FILLER_224_1016 ();
 FILLCELL_X32 FILLER_224_1048 ();
 FILLCELL_X32 FILLER_224_1080 ();
 FILLCELL_X32 FILLER_224_1112 ();
 FILLCELL_X32 FILLER_224_1144 ();
 FILLCELL_X32 FILLER_224_1176 ();
 FILLCELL_X32 FILLER_224_1208 ();
 FILLCELL_X32 FILLER_224_1240 ();
 FILLCELL_X32 FILLER_224_1272 ();
 FILLCELL_X32 FILLER_224_1304 ();
 FILLCELL_X32 FILLER_224_1336 ();
 FILLCELL_X32 FILLER_224_1368 ();
 FILLCELL_X32 FILLER_224_1400 ();
 FILLCELL_X32 FILLER_224_1432 ();
 FILLCELL_X32 FILLER_224_1464 ();
 FILLCELL_X32 FILLER_224_1496 ();
 FILLCELL_X32 FILLER_224_1528 ();
 FILLCELL_X32 FILLER_224_1560 ();
 FILLCELL_X32 FILLER_224_1592 ();
 FILLCELL_X32 FILLER_224_1624 ();
 FILLCELL_X32 FILLER_224_1656 ();
 FILLCELL_X32 FILLER_224_1688 ();
 FILLCELL_X32 FILLER_224_1720 ();
 FILLCELL_X4 FILLER_224_1752 ();
 FILLCELL_X32 FILLER_225_1 ();
 FILLCELL_X32 FILLER_225_33 ();
 FILLCELL_X32 FILLER_225_65 ();
 FILLCELL_X32 FILLER_225_97 ();
 FILLCELL_X32 FILLER_225_129 ();
 FILLCELL_X32 FILLER_225_161 ();
 FILLCELL_X32 FILLER_225_193 ();
 FILLCELL_X32 FILLER_225_225 ();
 FILLCELL_X32 FILLER_225_257 ();
 FILLCELL_X32 FILLER_225_289 ();
 FILLCELL_X32 FILLER_225_321 ();
 FILLCELL_X32 FILLER_225_353 ();
 FILLCELL_X32 FILLER_225_385 ();
 FILLCELL_X32 FILLER_225_417 ();
 FILLCELL_X32 FILLER_225_449 ();
 FILLCELL_X32 FILLER_225_481 ();
 FILLCELL_X32 FILLER_225_513 ();
 FILLCELL_X32 FILLER_225_545 ();
 FILLCELL_X32 FILLER_225_577 ();
 FILLCELL_X32 FILLER_225_609 ();
 FILLCELL_X32 FILLER_225_641 ();
 FILLCELL_X32 FILLER_225_673 ();
 FILLCELL_X32 FILLER_225_705 ();
 FILLCELL_X32 FILLER_225_737 ();
 FILLCELL_X32 FILLER_225_769 ();
 FILLCELL_X32 FILLER_225_801 ();
 FILLCELL_X32 FILLER_225_833 ();
 FILLCELL_X32 FILLER_225_865 ();
 FILLCELL_X32 FILLER_225_897 ();
 FILLCELL_X32 FILLER_225_929 ();
 FILLCELL_X32 FILLER_225_961 ();
 FILLCELL_X32 FILLER_225_993 ();
 FILLCELL_X32 FILLER_225_1025 ();
 FILLCELL_X32 FILLER_225_1057 ();
 FILLCELL_X32 FILLER_225_1089 ();
 FILLCELL_X32 FILLER_225_1121 ();
 FILLCELL_X32 FILLER_225_1153 ();
 FILLCELL_X32 FILLER_225_1185 ();
 FILLCELL_X32 FILLER_225_1217 ();
 FILLCELL_X8 FILLER_225_1249 ();
 FILLCELL_X4 FILLER_225_1257 ();
 FILLCELL_X2 FILLER_225_1261 ();
 FILLCELL_X32 FILLER_225_1264 ();
 FILLCELL_X32 FILLER_225_1296 ();
 FILLCELL_X32 FILLER_225_1328 ();
 FILLCELL_X32 FILLER_225_1360 ();
 FILLCELL_X32 FILLER_225_1392 ();
 FILLCELL_X32 FILLER_225_1424 ();
 FILLCELL_X32 FILLER_225_1456 ();
 FILLCELL_X32 FILLER_225_1488 ();
 FILLCELL_X32 FILLER_225_1520 ();
 FILLCELL_X32 FILLER_225_1552 ();
 FILLCELL_X32 FILLER_225_1584 ();
 FILLCELL_X32 FILLER_225_1616 ();
 FILLCELL_X32 FILLER_225_1648 ();
 FILLCELL_X32 FILLER_225_1680 ();
 FILLCELL_X32 FILLER_225_1712 ();
 FILLCELL_X8 FILLER_225_1744 ();
 FILLCELL_X4 FILLER_225_1752 ();
 FILLCELL_X4 FILLER_226_1 ();
 FILLCELL_X32 FILLER_226_12 ();
 FILLCELL_X32 FILLER_226_44 ();
 FILLCELL_X32 FILLER_226_76 ();
 FILLCELL_X32 FILLER_226_108 ();
 FILLCELL_X32 FILLER_226_140 ();
 FILLCELL_X32 FILLER_226_172 ();
 FILLCELL_X32 FILLER_226_204 ();
 FILLCELL_X32 FILLER_226_236 ();
 FILLCELL_X32 FILLER_226_268 ();
 FILLCELL_X32 FILLER_226_300 ();
 FILLCELL_X32 FILLER_226_332 ();
 FILLCELL_X32 FILLER_226_364 ();
 FILLCELL_X32 FILLER_226_396 ();
 FILLCELL_X32 FILLER_226_428 ();
 FILLCELL_X32 FILLER_226_460 ();
 FILLCELL_X32 FILLER_226_492 ();
 FILLCELL_X32 FILLER_226_524 ();
 FILLCELL_X32 FILLER_226_556 ();
 FILLCELL_X32 FILLER_226_588 ();
 FILLCELL_X8 FILLER_226_620 ();
 FILLCELL_X2 FILLER_226_628 ();
 FILLCELL_X1 FILLER_226_630 ();
 FILLCELL_X32 FILLER_226_632 ();
 FILLCELL_X32 FILLER_226_664 ();
 FILLCELL_X32 FILLER_226_696 ();
 FILLCELL_X32 FILLER_226_728 ();
 FILLCELL_X32 FILLER_226_760 ();
 FILLCELL_X32 FILLER_226_792 ();
 FILLCELL_X32 FILLER_226_824 ();
 FILLCELL_X32 FILLER_226_856 ();
 FILLCELL_X32 FILLER_226_888 ();
 FILLCELL_X32 FILLER_226_920 ();
 FILLCELL_X32 FILLER_226_952 ();
 FILLCELL_X32 FILLER_226_984 ();
 FILLCELL_X32 FILLER_226_1016 ();
 FILLCELL_X32 FILLER_226_1048 ();
 FILLCELL_X32 FILLER_226_1080 ();
 FILLCELL_X32 FILLER_226_1112 ();
 FILLCELL_X32 FILLER_226_1144 ();
 FILLCELL_X32 FILLER_226_1176 ();
 FILLCELL_X32 FILLER_226_1208 ();
 FILLCELL_X32 FILLER_226_1240 ();
 FILLCELL_X32 FILLER_226_1272 ();
 FILLCELL_X32 FILLER_226_1304 ();
 FILLCELL_X32 FILLER_226_1336 ();
 FILLCELL_X32 FILLER_226_1368 ();
 FILLCELL_X32 FILLER_226_1400 ();
 FILLCELL_X32 FILLER_226_1432 ();
 FILLCELL_X32 FILLER_226_1464 ();
 FILLCELL_X32 FILLER_226_1496 ();
 FILLCELL_X32 FILLER_226_1528 ();
 FILLCELL_X32 FILLER_226_1560 ();
 FILLCELL_X32 FILLER_226_1592 ();
 FILLCELL_X32 FILLER_226_1624 ();
 FILLCELL_X32 FILLER_226_1656 ();
 FILLCELL_X32 FILLER_226_1688 ();
 FILLCELL_X32 FILLER_226_1720 ();
 FILLCELL_X4 FILLER_226_1752 ();
 FILLCELL_X32 FILLER_227_1 ();
 FILLCELL_X32 FILLER_227_33 ();
 FILLCELL_X32 FILLER_227_65 ();
 FILLCELL_X32 FILLER_227_97 ();
 FILLCELL_X32 FILLER_227_129 ();
 FILLCELL_X32 FILLER_227_161 ();
 FILLCELL_X32 FILLER_227_193 ();
 FILLCELL_X32 FILLER_227_225 ();
 FILLCELL_X32 FILLER_227_257 ();
 FILLCELL_X32 FILLER_227_289 ();
 FILLCELL_X32 FILLER_227_321 ();
 FILLCELL_X32 FILLER_227_353 ();
 FILLCELL_X32 FILLER_227_385 ();
 FILLCELL_X32 FILLER_227_417 ();
 FILLCELL_X32 FILLER_227_449 ();
 FILLCELL_X32 FILLER_227_481 ();
 FILLCELL_X32 FILLER_227_513 ();
 FILLCELL_X32 FILLER_227_545 ();
 FILLCELL_X32 FILLER_227_577 ();
 FILLCELL_X32 FILLER_227_609 ();
 FILLCELL_X32 FILLER_227_641 ();
 FILLCELL_X32 FILLER_227_673 ();
 FILLCELL_X32 FILLER_227_705 ();
 FILLCELL_X32 FILLER_227_737 ();
 FILLCELL_X32 FILLER_227_769 ();
 FILLCELL_X32 FILLER_227_801 ();
 FILLCELL_X32 FILLER_227_833 ();
 FILLCELL_X32 FILLER_227_865 ();
 FILLCELL_X32 FILLER_227_897 ();
 FILLCELL_X32 FILLER_227_929 ();
 FILLCELL_X32 FILLER_227_961 ();
 FILLCELL_X32 FILLER_227_993 ();
 FILLCELL_X32 FILLER_227_1025 ();
 FILLCELL_X32 FILLER_227_1057 ();
 FILLCELL_X32 FILLER_227_1089 ();
 FILLCELL_X32 FILLER_227_1121 ();
 FILLCELL_X32 FILLER_227_1153 ();
 FILLCELL_X32 FILLER_227_1185 ();
 FILLCELL_X32 FILLER_227_1217 ();
 FILLCELL_X8 FILLER_227_1249 ();
 FILLCELL_X4 FILLER_227_1257 ();
 FILLCELL_X2 FILLER_227_1261 ();
 FILLCELL_X32 FILLER_227_1264 ();
 FILLCELL_X32 FILLER_227_1296 ();
 FILLCELL_X32 FILLER_227_1328 ();
 FILLCELL_X32 FILLER_227_1360 ();
 FILLCELL_X32 FILLER_227_1392 ();
 FILLCELL_X32 FILLER_227_1424 ();
 FILLCELL_X32 FILLER_227_1456 ();
 FILLCELL_X32 FILLER_227_1488 ();
 FILLCELL_X32 FILLER_227_1520 ();
 FILLCELL_X32 FILLER_227_1552 ();
 FILLCELL_X32 FILLER_227_1584 ();
 FILLCELL_X32 FILLER_227_1616 ();
 FILLCELL_X32 FILLER_227_1648 ();
 FILLCELL_X32 FILLER_227_1680 ();
 FILLCELL_X32 FILLER_227_1712 ();
 FILLCELL_X8 FILLER_227_1744 ();
 FILLCELL_X4 FILLER_227_1752 ();
 FILLCELL_X32 FILLER_228_1 ();
 FILLCELL_X32 FILLER_228_33 ();
 FILLCELL_X32 FILLER_228_65 ();
 FILLCELL_X32 FILLER_228_97 ();
 FILLCELL_X32 FILLER_228_129 ();
 FILLCELL_X32 FILLER_228_161 ();
 FILLCELL_X32 FILLER_228_193 ();
 FILLCELL_X32 FILLER_228_225 ();
 FILLCELL_X32 FILLER_228_257 ();
 FILLCELL_X32 FILLER_228_289 ();
 FILLCELL_X32 FILLER_228_321 ();
 FILLCELL_X32 FILLER_228_353 ();
 FILLCELL_X32 FILLER_228_385 ();
 FILLCELL_X32 FILLER_228_417 ();
 FILLCELL_X32 FILLER_228_449 ();
 FILLCELL_X32 FILLER_228_481 ();
 FILLCELL_X32 FILLER_228_513 ();
 FILLCELL_X32 FILLER_228_545 ();
 FILLCELL_X32 FILLER_228_577 ();
 FILLCELL_X16 FILLER_228_609 ();
 FILLCELL_X4 FILLER_228_625 ();
 FILLCELL_X2 FILLER_228_629 ();
 FILLCELL_X32 FILLER_228_632 ();
 FILLCELL_X32 FILLER_228_664 ();
 FILLCELL_X32 FILLER_228_696 ();
 FILLCELL_X32 FILLER_228_728 ();
 FILLCELL_X32 FILLER_228_760 ();
 FILLCELL_X32 FILLER_228_792 ();
 FILLCELL_X32 FILLER_228_824 ();
 FILLCELL_X32 FILLER_228_856 ();
 FILLCELL_X32 FILLER_228_888 ();
 FILLCELL_X32 FILLER_228_920 ();
 FILLCELL_X32 FILLER_228_952 ();
 FILLCELL_X32 FILLER_228_984 ();
 FILLCELL_X32 FILLER_228_1016 ();
 FILLCELL_X32 FILLER_228_1048 ();
 FILLCELL_X32 FILLER_228_1080 ();
 FILLCELL_X32 FILLER_228_1112 ();
 FILLCELL_X32 FILLER_228_1144 ();
 FILLCELL_X32 FILLER_228_1176 ();
 FILLCELL_X32 FILLER_228_1208 ();
 FILLCELL_X32 FILLER_228_1240 ();
 FILLCELL_X32 FILLER_228_1272 ();
 FILLCELL_X32 FILLER_228_1304 ();
 FILLCELL_X32 FILLER_228_1336 ();
 FILLCELL_X32 FILLER_228_1368 ();
 FILLCELL_X32 FILLER_228_1400 ();
 FILLCELL_X32 FILLER_228_1432 ();
 FILLCELL_X32 FILLER_228_1464 ();
 FILLCELL_X32 FILLER_228_1496 ();
 FILLCELL_X32 FILLER_228_1528 ();
 FILLCELL_X32 FILLER_228_1560 ();
 FILLCELL_X32 FILLER_228_1592 ();
 FILLCELL_X32 FILLER_228_1624 ();
 FILLCELL_X32 FILLER_228_1656 ();
 FILLCELL_X32 FILLER_228_1688 ();
 FILLCELL_X32 FILLER_228_1720 ();
 FILLCELL_X4 FILLER_228_1752 ();
 FILLCELL_X32 FILLER_229_1 ();
 FILLCELL_X32 FILLER_229_33 ();
 FILLCELL_X32 FILLER_229_65 ();
 FILLCELL_X32 FILLER_229_97 ();
 FILLCELL_X32 FILLER_229_129 ();
 FILLCELL_X32 FILLER_229_161 ();
 FILLCELL_X32 FILLER_229_193 ();
 FILLCELL_X32 FILLER_229_225 ();
 FILLCELL_X32 FILLER_229_257 ();
 FILLCELL_X32 FILLER_229_289 ();
 FILLCELL_X32 FILLER_229_321 ();
 FILLCELL_X32 FILLER_229_353 ();
 FILLCELL_X32 FILLER_229_385 ();
 FILLCELL_X32 FILLER_229_417 ();
 FILLCELL_X32 FILLER_229_449 ();
 FILLCELL_X32 FILLER_229_481 ();
 FILLCELL_X32 FILLER_229_513 ();
 FILLCELL_X32 FILLER_229_545 ();
 FILLCELL_X32 FILLER_229_577 ();
 FILLCELL_X32 FILLER_229_609 ();
 FILLCELL_X32 FILLER_229_641 ();
 FILLCELL_X32 FILLER_229_673 ();
 FILLCELL_X32 FILLER_229_705 ();
 FILLCELL_X32 FILLER_229_737 ();
 FILLCELL_X32 FILLER_229_769 ();
 FILLCELL_X32 FILLER_229_801 ();
 FILLCELL_X32 FILLER_229_833 ();
 FILLCELL_X32 FILLER_229_865 ();
 FILLCELL_X32 FILLER_229_897 ();
 FILLCELL_X32 FILLER_229_929 ();
 FILLCELL_X32 FILLER_229_961 ();
 FILLCELL_X32 FILLER_229_993 ();
 FILLCELL_X32 FILLER_229_1025 ();
 FILLCELL_X32 FILLER_229_1057 ();
 FILLCELL_X32 FILLER_229_1089 ();
 FILLCELL_X32 FILLER_229_1121 ();
 FILLCELL_X32 FILLER_229_1153 ();
 FILLCELL_X32 FILLER_229_1185 ();
 FILLCELL_X32 FILLER_229_1217 ();
 FILLCELL_X8 FILLER_229_1249 ();
 FILLCELL_X4 FILLER_229_1257 ();
 FILLCELL_X2 FILLER_229_1261 ();
 FILLCELL_X32 FILLER_229_1264 ();
 FILLCELL_X32 FILLER_229_1296 ();
 FILLCELL_X32 FILLER_229_1328 ();
 FILLCELL_X32 FILLER_229_1360 ();
 FILLCELL_X32 FILLER_229_1392 ();
 FILLCELL_X32 FILLER_229_1424 ();
 FILLCELL_X32 FILLER_229_1456 ();
 FILLCELL_X32 FILLER_229_1488 ();
 FILLCELL_X32 FILLER_229_1520 ();
 FILLCELL_X32 FILLER_229_1552 ();
 FILLCELL_X32 FILLER_229_1584 ();
 FILLCELL_X32 FILLER_229_1616 ();
 FILLCELL_X32 FILLER_229_1648 ();
 FILLCELL_X32 FILLER_229_1680 ();
 FILLCELL_X32 FILLER_229_1712 ();
 FILLCELL_X8 FILLER_229_1744 ();
 FILLCELL_X4 FILLER_229_1752 ();
 FILLCELL_X32 FILLER_230_1 ();
 FILLCELL_X32 FILLER_230_33 ();
 FILLCELL_X32 FILLER_230_65 ();
 FILLCELL_X32 FILLER_230_97 ();
 FILLCELL_X32 FILLER_230_129 ();
 FILLCELL_X32 FILLER_230_161 ();
 FILLCELL_X32 FILLER_230_193 ();
 FILLCELL_X32 FILLER_230_225 ();
 FILLCELL_X32 FILLER_230_257 ();
 FILLCELL_X32 FILLER_230_289 ();
 FILLCELL_X32 FILLER_230_321 ();
 FILLCELL_X32 FILLER_230_353 ();
 FILLCELL_X32 FILLER_230_385 ();
 FILLCELL_X32 FILLER_230_417 ();
 FILLCELL_X32 FILLER_230_449 ();
 FILLCELL_X32 FILLER_230_481 ();
 FILLCELL_X32 FILLER_230_513 ();
 FILLCELL_X32 FILLER_230_545 ();
 FILLCELL_X32 FILLER_230_577 ();
 FILLCELL_X16 FILLER_230_609 ();
 FILLCELL_X4 FILLER_230_625 ();
 FILLCELL_X2 FILLER_230_629 ();
 FILLCELL_X32 FILLER_230_632 ();
 FILLCELL_X32 FILLER_230_664 ();
 FILLCELL_X32 FILLER_230_696 ();
 FILLCELL_X32 FILLER_230_728 ();
 FILLCELL_X32 FILLER_230_760 ();
 FILLCELL_X32 FILLER_230_792 ();
 FILLCELL_X32 FILLER_230_824 ();
 FILLCELL_X32 FILLER_230_856 ();
 FILLCELL_X32 FILLER_230_888 ();
 FILLCELL_X32 FILLER_230_920 ();
 FILLCELL_X32 FILLER_230_952 ();
 FILLCELL_X32 FILLER_230_984 ();
 FILLCELL_X32 FILLER_230_1016 ();
 FILLCELL_X32 FILLER_230_1048 ();
 FILLCELL_X32 FILLER_230_1080 ();
 FILLCELL_X32 FILLER_230_1112 ();
 FILLCELL_X32 FILLER_230_1144 ();
 FILLCELL_X32 FILLER_230_1176 ();
 FILLCELL_X32 FILLER_230_1208 ();
 FILLCELL_X32 FILLER_230_1240 ();
 FILLCELL_X32 FILLER_230_1272 ();
 FILLCELL_X32 FILLER_230_1304 ();
 FILLCELL_X32 FILLER_230_1336 ();
 FILLCELL_X32 FILLER_230_1368 ();
 FILLCELL_X32 FILLER_230_1400 ();
 FILLCELL_X32 FILLER_230_1432 ();
 FILLCELL_X32 FILLER_230_1464 ();
 FILLCELL_X32 FILLER_230_1496 ();
 FILLCELL_X32 FILLER_230_1528 ();
 FILLCELL_X32 FILLER_230_1560 ();
 FILLCELL_X32 FILLER_230_1592 ();
 FILLCELL_X32 FILLER_230_1624 ();
 FILLCELL_X32 FILLER_230_1656 ();
 FILLCELL_X32 FILLER_230_1688 ();
 FILLCELL_X32 FILLER_230_1720 ();
 FILLCELL_X4 FILLER_230_1752 ();
 FILLCELL_X32 FILLER_231_1 ();
 FILLCELL_X32 FILLER_231_33 ();
 FILLCELL_X32 FILLER_231_65 ();
 FILLCELL_X32 FILLER_231_97 ();
 FILLCELL_X32 FILLER_231_129 ();
 FILLCELL_X32 FILLER_231_161 ();
 FILLCELL_X32 FILLER_231_193 ();
 FILLCELL_X32 FILLER_231_225 ();
 FILLCELL_X32 FILLER_231_257 ();
 FILLCELL_X32 FILLER_231_289 ();
 FILLCELL_X32 FILLER_231_321 ();
 FILLCELL_X32 FILLER_231_353 ();
 FILLCELL_X32 FILLER_231_385 ();
 FILLCELL_X32 FILLER_231_417 ();
 FILLCELL_X32 FILLER_231_449 ();
 FILLCELL_X32 FILLER_231_481 ();
 FILLCELL_X32 FILLER_231_513 ();
 FILLCELL_X32 FILLER_231_545 ();
 FILLCELL_X32 FILLER_231_577 ();
 FILLCELL_X32 FILLER_231_609 ();
 FILLCELL_X32 FILLER_231_641 ();
 FILLCELL_X32 FILLER_231_673 ();
 FILLCELL_X32 FILLER_231_705 ();
 FILLCELL_X32 FILLER_231_737 ();
 FILLCELL_X32 FILLER_231_769 ();
 FILLCELL_X32 FILLER_231_801 ();
 FILLCELL_X32 FILLER_231_833 ();
 FILLCELL_X32 FILLER_231_865 ();
 FILLCELL_X32 FILLER_231_897 ();
 FILLCELL_X32 FILLER_231_929 ();
 FILLCELL_X32 FILLER_231_961 ();
 FILLCELL_X32 FILLER_231_993 ();
 FILLCELL_X32 FILLER_231_1025 ();
 FILLCELL_X32 FILLER_231_1057 ();
 FILLCELL_X32 FILLER_231_1089 ();
 FILLCELL_X32 FILLER_231_1121 ();
 FILLCELL_X32 FILLER_231_1153 ();
 FILLCELL_X32 FILLER_231_1185 ();
 FILLCELL_X32 FILLER_231_1217 ();
 FILLCELL_X8 FILLER_231_1249 ();
 FILLCELL_X4 FILLER_231_1257 ();
 FILLCELL_X2 FILLER_231_1261 ();
 FILLCELL_X32 FILLER_231_1264 ();
 FILLCELL_X32 FILLER_231_1296 ();
 FILLCELL_X32 FILLER_231_1328 ();
 FILLCELL_X32 FILLER_231_1360 ();
 FILLCELL_X32 FILLER_231_1392 ();
 FILLCELL_X32 FILLER_231_1424 ();
 FILLCELL_X32 FILLER_231_1456 ();
 FILLCELL_X32 FILLER_231_1488 ();
 FILLCELL_X32 FILLER_231_1520 ();
 FILLCELL_X32 FILLER_231_1552 ();
 FILLCELL_X32 FILLER_231_1584 ();
 FILLCELL_X32 FILLER_231_1616 ();
 FILLCELL_X32 FILLER_231_1648 ();
 FILLCELL_X32 FILLER_231_1680 ();
 FILLCELL_X32 FILLER_231_1712 ();
 FILLCELL_X1 FILLER_231_1744 ();
 FILLCELL_X4 FILLER_231_1752 ();
 FILLCELL_X32 FILLER_232_1 ();
 FILLCELL_X32 FILLER_232_33 ();
 FILLCELL_X32 FILLER_232_65 ();
 FILLCELL_X32 FILLER_232_97 ();
 FILLCELL_X32 FILLER_232_129 ();
 FILLCELL_X32 FILLER_232_161 ();
 FILLCELL_X32 FILLER_232_193 ();
 FILLCELL_X32 FILLER_232_225 ();
 FILLCELL_X32 FILLER_232_257 ();
 FILLCELL_X32 FILLER_232_289 ();
 FILLCELL_X32 FILLER_232_321 ();
 FILLCELL_X32 FILLER_232_353 ();
 FILLCELL_X32 FILLER_232_385 ();
 FILLCELL_X32 FILLER_232_417 ();
 FILLCELL_X32 FILLER_232_449 ();
 FILLCELL_X32 FILLER_232_481 ();
 FILLCELL_X32 FILLER_232_513 ();
 FILLCELL_X32 FILLER_232_545 ();
 FILLCELL_X32 FILLER_232_577 ();
 FILLCELL_X16 FILLER_232_609 ();
 FILLCELL_X4 FILLER_232_625 ();
 FILLCELL_X2 FILLER_232_629 ();
 FILLCELL_X32 FILLER_232_632 ();
 FILLCELL_X32 FILLER_232_664 ();
 FILLCELL_X32 FILLER_232_696 ();
 FILLCELL_X32 FILLER_232_728 ();
 FILLCELL_X32 FILLER_232_760 ();
 FILLCELL_X32 FILLER_232_792 ();
 FILLCELL_X32 FILLER_232_824 ();
 FILLCELL_X32 FILLER_232_856 ();
 FILLCELL_X32 FILLER_232_888 ();
 FILLCELL_X32 FILLER_232_920 ();
 FILLCELL_X32 FILLER_232_952 ();
 FILLCELL_X32 FILLER_232_984 ();
 FILLCELL_X32 FILLER_232_1016 ();
 FILLCELL_X32 FILLER_232_1048 ();
 FILLCELL_X32 FILLER_232_1080 ();
 FILLCELL_X32 FILLER_232_1112 ();
 FILLCELL_X32 FILLER_232_1144 ();
 FILLCELL_X32 FILLER_232_1176 ();
 FILLCELL_X32 FILLER_232_1208 ();
 FILLCELL_X32 FILLER_232_1240 ();
 FILLCELL_X32 FILLER_232_1272 ();
 FILLCELL_X32 FILLER_232_1304 ();
 FILLCELL_X32 FILLER_232_1336 ();
 FILLCELL_X32 FILLER_232_1368 ();
 FILLCELL_X32 FILLER_232_1400 ();
 FILLCELL_X32 FILLER_232_1432 ();
 FILLCELL_X32 FILLER_232_1464 ();
 FILLCELL_X32 FILLER_232_1496 ();
 FILLCELL_X32 FILLER_232_1528 ();
 FILLCELL_X32 FILLER_232_1560 ();
 FILLCELL_X32 FILLER_232_1592 ();
 FILLCELL_X32 FILLER_232_1624 ();
 FILLCELL_X32 FILLER_232_1656 ();
 FILLCELL_X32 FILLER_232_1688 ();
 FILLCELL_X32 FILLER_232_1720 ();
 FILLCELL_X4 FILLER_232_1752 ();
 FILLCELL_X32 FILLER_233_1 ();
 FILLCELL_X32 FILLER_233_33 ();
 FILLCELL_X32 FILLER_233_65 ();
 FILLCELL_X32 FILLER_233_97 ();
 FILLCELL_X32 FILLER_233_129 ();
 FILLCELL_X32 FILLER_233_161 ();
 FILLCELL_X32 FILLER_233_193 ();
 FILLCELL_X32 FILLER_233_225 ();
 FILLCELL_X32 FILLER_233_257 ();
 FILLCELL_X32 FILLER_233_289 ();
 FILLCELL_X32 FILLER_233_321 ();
 FILLCELL_X32 FILLER_233_353 ();
 FILLCELL_X32 FILLER_233_385 ();
 FILLCELL_X32 FILLER_233_417 ();
 FILLCELL_X32 FILLER_233_449 ();
 FILLCELL_X32 FILLER_233_481 ();
 FILLCELL_X32 FILLER_233_513 ();
 FILLCELL_X32 FILLER_233_545 ();
 FILLCELL_X32 FILLER_233_577 ();
 FILLCELL_X32 FILLER_233_609 ();
 FILLCELL_X32 FILLER_233_641 ();
 FILLCELL_X32 FILLER_233_673 ();
 FILLCELL_X32 FILLER_233_705 ();
 FILLCELL_X32 FILLER_233_737 ();
 FILLCELL_X32 FILLER_233_769 ();
 FILLCELL_X32 FILLER_233_801 ();
 FILLCELL_X32 FILLER_233_833 ();
 FILLCELL_X32 FILLER_233_865 ();
 FILLCELL_X32 FILLER_233_897 ();
 FILLCELL_X32 FILLER_233_929 ();
 FILLCELL_X32 FILLER_233_961 ();
 FILLCELL_X32 FILLER_233_993 ();
 FILLCELL_X32 FILLER_233_1025 ();
 FILLCELL_X32 FILLER_233_1057 ();
 FILLCELL_X32 FILLER_233_1089 ();
 FILLCELL_X32 FILLER_233_1121 ();
 FILLCELL_X32 FILLER_233_1153 ();
 FILLCELL_X32 FILLER_233_1185 ();
 FILLCELL_X32 FILLER_233_1217 ();
 FILLCELL_X8 FILLER_233_1249 ();
 FILLCELL_X4 FILLER_233_1257 ();
 FILLCELL_X2 FILLER_233_1261 ();
 FILLCELL_X32 FILLER_233_1264 ();
 FILLCELL_X32 FILLER_233_1296 ();
 FILLCELL_X32 FILLER_233_1328 ();
 FILLCELL_X32 FILLER_233_1360 ();
 FILLCELL_X32 FILLER_233_1392 ();
 FILLCELL_X32 FILLER_233_1424 ();
 FILLCELL_X32 FILLER_233_1456 ();
 FILLCELL_X32 FILLER_233_1488 ();
 FILLCELL_X32 FILLER_233_1520 ();
 FILLCELL_X32 FILLER_233_1552 ();
 FILLCELL_X32 FILLER_233_1584 ();
 FILLCELL_X32 FILLER_233_1616 ();
 FILLCELL_X32 FILLER_233_1648 ();
 FILLCELL_X32 FILLER_233_1680 ();
 FILLCELL_X32 FILLER_233_1712 ();
 FILLCELL_X8 FILLER_233_1744 ();
 FILLCELL_X4 FILLER_233_1752 ();
 FILLCELL_X32 FILLER_234_1 ();
 FILLCELL_X32 FILLER_234_33 ();
 FILLCELL_X32 FILLER_234_65 ();
 FILLCELL_X32 FILLER_234_97 ();
 FILLCELL_X32 FILLER_234_129 ();
 FILLCELL_X32 FILLER_234_161 ();
 FILLCELL_X32 FILLER_234_193 ();
 FILLCELL_X32 FILLER_234_225 ();
 FILLCELL_X32 FILLER_234_257 ();
 FILLCELL_X32 FILLER_234_289 ();
 FILLCELL_X32 FILLER_234_321 ();
 FILLCELL_X32 FILLER_234_353 ();
 FILLCELL_X32 FILLER_234_385 ();
 FILLCELL_X32 FILLER_234_417 ();
 FILLCELL_X32 FILLER_234_449 ();
 FILLCELL_X32 FILLER_234_481 ();
 FILLCELL_X32 FILLER_234_513 ();
 FILLCELL_X32 FILLER_234_545 ();
 FILLCELL_X32 FILLER_234_577 ();
 FILLCELL_X16 FILLER_234_609 ();
 FILLCELL_X4 FILLER_234_625 ();
 FILLCELL_X2 FILLER_234_629 ();
 FILLCELL_X32 FILLER_234_632 ();
 FILLCELL_X32 FILLER_234_664 ();
 FILLCELL_X32 FILLER_234_696 ();
 FILLCELL_X32 FILLER_234_728 ();
 FILLCELL_X32 FILLER_234_760 ();
 FILLCELL_X32 FILLER_234_792 ();
 FILLCELL_X32 FILLER_234_824 ();
 FILLCELL_X32 FILLER_234_856 ();
 FILLCELL_X32 FILLER_234_888 ();
 FILLCELL_X32 FILLER_234_920 ();
 FILLCELL_X32 FILLER_234_952 ();
 FILLCELL_X32 FILLER_234_984 ();
 FILLCELL_X32 FILLER_234_1016 ();
 FILLCELL_X32 FILLER_234_1048 ();
 FILLCELL_X32 FILLER_234_1080 ();
 FILLCELL_X32 FILLER_234_1112 ();
 FILLCELL_X32 FILLER_234_1144 ();
 FILLCELL_X32 FILLER_234_1176 ();
 FILLCELL_X32 FILLER_234_1208 ();
 FILLCELL_X32 FILLER_234_1240 ();
 FILLCELL_X32 FILLER_234_1272 ();
 FILLCELL_X32 FILLER_234_1304 ();
 FILLCELL_X32 FILLER_234_1336 ();
 FILLCELL_X32 FILLER_234_1368 ();
 FILLCELL_X32 FILLER_234_1400 ();
 FILLCELL_X32 FILLER_234_1432 ();
 FILLCELL_X32 FILLER_234_1464 ();
 FILLCELL_X32 FILLER_234_1496 ();
 FILLCELL_X32 FILLER_234_1528 ();
 FILLCELL_X32 FILLER_234_1560 ();
 FILLCELL_X32 FILLER_234_1592 ();
 FILLCELL_X32 FILLER_234_1624 ();
 FILLCELL_X32 FILLER_234_1656 ();
 FILLCELL_X32 FILLER_234_1688 ();
 FILLCELL_X32 FILLER_234_1720 ();
 FILLCELL_X4 FILLER_234_1752 ();
 FILLCELL_X32 FILLER_235_1 ();
 FILLCELL_X32 FILLER_235_33 ();
 FILLCELL_X32 FILLER_235_65 ();
 FILLCELL_X32 FILLER_235_97 ();
 FILLCELL_X32 FILLER_235_129 ();
 FILLCELL_X32 FILLER_235_161 ();
 FILLCELL_X32 FILLER_235_193 ();
 FILLCELL_X32 FILLER_235_225 ();
 FILLCELL_X32 FILLER_235_257 ();
 FILLCELL_X32 FILLER_235_289 ();
 FILLCELL_X32 FILLER_235_321 ();
 FILLCELL_X32 FILLER_235_353 ();
 FILLCELL_X32 FILLER_235_385 ();
 FILLCELL_X32 FILLER_235_417 ();
 FILLCELL_X32 FILLER_235_449 ();
 FILLCELL_X32 FILLER_235_481 ();
 FILLCELL_X32 FILLER_235_513 ();
 FILLCELL_X32 FILLER_235_545 ();
 FILLCELL_X32 FILLER_235_577 ();
 FILLCELL_X32 FILLER_235_609 ();
 FILLCELL_X32 FILLER_235_641 ();
 FILLCELL_X32 FILLER_235_673 ();
 FILLCELL_X32 FILLER_235_705 ();
 FILLCELL_X32 FILLER_235_737 ();
 FILLCELL_X32 FILLER_235_769 ();
 FILLCELL_X32 FILLER_235_801 ();
 FILLCELL_X32 FILLER_235_833 ();
 FILLCELL_X32 FILLER_235_865 ();
 FILLCELL_X32 FILLER_235_897 ();
 FILLCELL_X32 FILLER_235_929 ();
 FILLCELL_X32 FILLER_235_961 ();
 FILLCELL_X32 FILLER_235_993 ();
 FILLCELL_X32 FILLER_235_1025 ();
 FILLCELL_X32 FILLER_235_1057 ();
 FILLCELL_X32 FILLER_235_1089 ();
 FILLCELL_X32 FILLER_235_1121 ();
 FILLCELL_X32 FILLER_235_1153 ();
 FILLCELL_X32 FILLER_235_1185 ();
 FILLCELL_X32 FILLER_235_1217 ();
 FILLCELL_X8 FILLER_235_1249 ();
 FILLCELL_X4 FILLER_235_1257 ();
 FILLCELL_X2 FILLER_235_1261 ();
 FILLCELL_X32 FILLER_235_1264 ();
 FILLCELL_X32 FILLER_235_1296 ();
 FILLCELL_X32 FILLER_235_1328 ();
 FILLCELL_X32 FILLER_235_1360 ();
 FILLCELL_X32 FILLER_235_1392 ();
 FILLCELL_X32 FILLER_235_1424 ();
 FILLCELL_X32 FILLER_235_1456 ();
 FILLCELL_X32 FILLER_235_1488 ();
 FILLCELL_X32 FILLER_235_1520 ();
 FILLCELL_X32 FILLER_235_1552 ();
 FILLCELL_X32 FILLER_235_1584 ();
 FILLCELL_X32 FILLER_235_1616 ();
 FILLCELL_X32 FILLER_235_1648 ();
 FILLCELL_X32 FILLER_235_1680 ();
 FILLCELL_X32 FILLER_235_1712 ();
 FILLCELL_X8 FILLER_235_1744 ();
 FILLCELL_X4 FILLER_235_1752 ();
 FILLCELL_X4 FILLER_236_1 ();
 FILLCELL_X32 FILLER_236_8 ();
 FILLCELL_X32 FILLER_236_40 ();
 FILLCELL_X32 FILLER_236_72 ();
 FILLCELL_X32 FILLER_236_104 ();
 FILLCELL_X32 FILLER_236_136 ();
 FILLCELL_X32 FILLER_236_168 ();
 FILLCELL_X32 FILLER_236_200 ();
 FILLCELL_X32 FILLER_236_232 ();
 FILLCELL_X32 FILLER_236_264 ();
 FILLCELL_X32 FILLER_236_296 ();
 FILLCELL_X32 FILLER_236_328 ();
 FILLCELL_X32 FILLER_236_360 ();
 FILLCELL_X32 FILLER_236_392 ();
 FILLCELL_X32 FILLER_236_424 ();
 FILLCELL_X32 FILLER_236_456 ();
 FILLCELL_X32 FILLER_236_488 ();
 FILLCELL_X32 FILLER_236_520 ();
 FILLCELL_X32 FILLER_236_552 ();
 FILLCELL_X32 FILLER_236_584 ();
 FILLCELL_X8 FILLER_236_616 ();
 FILLCELL_X4 FILLER_236_624 ();
 FILLCELL_X2 FILLER_236_628 ();
 FILLCELL_X1 FILLER_236_630 ();
 FILLCELL_X32 FILLER_236_632 ();
 FILLCELL_X32 FILLER_236_664 ();
 FILLCELL_X32 FILLER_236_696 ();
 FILLCELL_X32 FILLER_236_728 ();
 FILLCELL_X32 FILLER_236_760 ();
 FILLCELL_X32 FILLER_236_792 ();
 FILLCELL_X32 FILLER_236_824 ();
 FILLCELL_X32 FILLER_236_856 ();
 FILLCELL_X32 FILLER_236_888 ();
 FILLCELL_X32 FILLER_236_920 ();
 FILLCELL_X32 FILLER_236_952 ();
 FILLCELL_X32 FILLER_236_984 ();
 FILLCELL_X32 FILLER_236_1016 ();
 FILLCELL_X32 FILLER_236_1048 ();
 FILLCELL_X32 FILLER_236_1080 ();
 FILLCELL_X32 FILLER_236_1112 ();
 FILLCELL_X32 FILLER_236_1144 ();
 FILLCELL_X32 FILLER_236_1176 ();
 FILLCELL_X32 FILLER_236_1208 ();
 FILLCELL_X32 FILLER_236_1240 ();
 FILLCELL_X32 FILLER_236_1272 ();
 FILLCELL_X32 FILLER_236_1304 ();
 FILLCELL_X32 FILLER_236_1336 ();
 FILLCELL_X32 FILLER_236_1368 ();
 FILLCELL_X32 FILLER_236_1400 ();
 FILLCELL_X32 FILLER_236_1432 ();
 FILLCELL_X32 FILLER_236_1464 ();
 FILLCELL_X32 FILLER_236_1496 ();
 FILLCELL_X32 FILLER_236_1528 ();
 FILLCELL_X32 FILLER_236_1560 ();
 FILLCELL_X32 FILLER_236_1592 ();
 FILLCELL_X32 FILLER_236_1624 ();
 FILLCELL_X32 FILLER_236_1656 ();
 FILLCELL_X32 FILLER_236_1688 ();
 FILLCELL_X32 FILLER_236_1720 ();
 FILLCELL_X4 FILLER_236_1752 ();
 FILLCELL_X8 FILLER_237_1 ();
 FILLCELL_X32 FILLER_237_12 ();
 FILLCELL_X32 FILLER_237_44 ();
 FILLCELL_X4 FILLER_237_76 ();
 FILLCELL_X32 FILLER_237_83 ();
 FILLCELL_X32 FILLER_237_115 ();
 FILLCELL_X2 FILLER_237_147 ();
 FILLCELL_X1 FILLER_237_149 ();
 FILLCELL_X32 FILLER_237_153 ();
 FILLCELL_X32 FILLER_237_185 ();
 FILLCELL_X4 FILLER_237_217 ();
 FILLCELL_X32 FILLER_237_224 ();
 FILLCELL_X32 FILLER_237_256 ();
 FILLCELL_X4 FILLER_237_288 ();
 FILLCELL_X32 FILLER_237_295 ();
 FILLCELL_X32 FILLER_237_327 ();
 FILLCELL_X4 FILLER_237_359 ();
 FILLCELL_X32 FILLER_237_366 ();
 FILLCELL_X32 FILLER_237_398 ();
 FILLCELL_X2 FILLER_237_430 ();
 FILLCELL_X1 FILLER_237_432 ();
 FILLCELL_X32 FILLER_237_436 ();
 FILLCELL_X32 FILLER_237_468 ();
 FILLCELL_X4 FILLER_237_500 ();
 FILLCELL_X32 FILLER_237_507 ();
 FILLCELL_X32 FILLER_237_539 ();
 FILLCELL_X4 FILLER_237_571 ();
 FILLCELL_X32 FILLER_237_582 ();
 FILLCELL_X16 FILLER_237_614 ();
 FILLCELL_X1 FILLER_237_630 ();
 FILLCELL_X8 FILLER_237_632 ();
 FILLCELL_X4 FILLER_237_640 ();
 FILLCELL_X2 FILLER_237_644 ();
 FILLCELL_X32 FILLER_237_653 ();
 FILLCELL_X16 FILLER_237_685 ();
 FILLCELL_X8 FILLER_237_701 ();
 FILLCELL_X4 FILLER_237_709 ();
 FILLCELL_X2 FILLER_237_713 ();
 FILLCELL_X1 FILLER_237_715 ();
 FILLCELL_X32 FILLER_237_719 ();
 FILLCELL_X32 FILLER_237_751 ();
 FILLCELL_X4 FILLER_237_783 ();
 FILLCELL_X32 FILLER_237_794 ();
 FILLCELL_X32 FILLER_237_826 ();
 FILLCELL_X32 FILLER_237_861 ();
 FILLCELL_X32 FILLER_237_893 ();
 FILLCELL_X2 FILLER_237_925 ();
 FILLCELL_X1 FILLER_237_927 ();
 FILLCELL_X32 FILLER_237_931 ();
 FILLCELL_X32 FILLER_237_963 ();
 FILLCELL_X4 FILLER_237_995 ();
 FILLCELL_X32 FILLER_237_1006 ();
 FILLCELL_X32 FILLER_237_1038 ();
 FILLCELL_X32 FILLER_237_1077 ();
 FILLCELL_X32 FILLER_237_1109 ();
 FILLCELL_X32 FILLER_237_1144 ();
 FILLCELL_X32 FILLER_237_1176 ();
 FILLCELL_X2 FILLER_237_1208 ();
 FILLCELL_X1 FILLER_237_1210 ();
 FILLCELL_X32 FILLER_237_1214 ();
 FILLCELL_X16 FILLER_237_1246 ();
 FILLCELL_X16 FILLER_237_1263 ();
 FILLCELL_X2 FILLER_237_1279 ();
 FILLCELL_X1 FILLER_237_1281 ();
 FILLCELL_X32 FILLER_237_1285 ();
 FILLCELL_X32 FILLER_237_1317 ();
 FILLCELL_X4 FILLER_237_1349 ();
 FILLCELL_X32 FILLER_237_1356 ();
 FILLCELL_X32 FILLER_237_1388 ();
 FILLCELL_X4 FILLER_237_1420 ();
 FILLCELL_X32 FILLER_237_1427 ();
 FILLCELL_X32 FILLER_237_1459 ();
 FILLCELL_X2 FILLER_237_1491 ();
 FILLCELL_X1 FILLER_237_1493 ();
 FILLCELL_X32 FILLER_237_1497 ();
 FILLCELL_X32 FILLER_237_1529 ();
 FILLCELL_X4 FILLER_237_1561 ();
 FILLCELL_X32 FILLER_237_1568 ();
 FILLCELL_X32 FILLER_237_1600 ();
 FILLCELL_X4 FILLER_237_1632 ();
 FILLCELL_X32 FILLER_237_1639 ();
 FILLCELL_X32 FILLER_237_1671 ();
 FILLCELL_X4 FILLER_237_1703 ();
 FILLCELL_X32 FILLER_237_1714 ();
 FILLCELL_X2 FILLER_237_1746 ();
 FILLCELL_X1 FILLER_237_1748 ();
 FILLCELL_X4 FILLER_237_1752 ();
 assign init_done = curr_state[1];
 assign valid_out = valid_reg_out;
endmodule
