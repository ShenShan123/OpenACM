module sram_multiplier_system (clk,
    init_done,
    init_enable,
    pe_ce,
    rst_n,
    valid_out,
    data_in,
    data_out);
 input clk;
 output init_done;
 input init_enable;
 input pe_ce;
 input rst_n;
 output valid_out;
 input [7:0] data_in;
 output [15:0] data_out;

 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire \u_multiplier/_0345_ ;
 wire \u_multiplier/_0346_ ;
 wire \u_multiplier/_0347_ ;
 wire \u_multiplier/_0348_ ;
 wire \u_multiplier/_0349_ ;
 wire \u_multiplier/_0350_ ;
 wire \u_multiplier/_0351_ ;
 wire \u_multiplier/_0352_ ;
 wire \u_multiplier/_0353_ ;
 wire \u_multiplier/_0354_ ;
 wire \u_multiplier/_0355_ ;
 wire \u_multiplier/_0392_ ;
 wire \u_multiplier/_0393_ ;
 wire \u_multiplier/_0394_ ;
 wire \u_multiplier/_0395_ ;
 wire \u_multiplier/_0396_ ;
 wire \u_multiplier/_0397_ ;
 wire \u_multiplier/_0398_ ;
 wire \u_multiplier/_0399_ ;
 wire \u_multiplier/_0400_ ;
 wire \u_multiplier/_0401_ ;
 wire \u_multiplier/_0402_ ;
 wire \u_multiplier/_0403_ ;
 wire \u_multiplier/_0404_ ;
 wire \u_multiplier/_0405_ ;
 wire \u_multiplier/_0406_ ;
 wire \u_multiplier/_0407_ ;
 wire \u_multiplier/_0408_ ;
 wire \u_multiplier/_0409_ ;
 wire \u_multiplier/_0410_ ;
 wire \u_multiplier/_0411_ ;
 wire \u_multiplier/_0412_ ;
 wire \u_multiplier/_0413_ ;
 wire \u_multiplier/_0414_ ;
 wire \u_multiplier/_0415_ ;
 wire \u_multiplier/_0416_ ;
 wire \u_multiplier/_0417_ ;
 wire \u_multiplier/_0418_ ;
 wire \u_multiplier/_0419_ ;
 wire \u_multiplier/_0420_ ;
 wire \u_multiplier/_0421_ ;
 wire \u_multiplier/_0422_ ;
 wire \u_multiplier/_0423_ ;
 wire \u_multiplier/_0424_ ;
 wire \u_multiplier/_0425_ ;
 wire \u_multiplier/_0426_ ;
 wire \u_multiplier/_0427_ ;
 wire \u_multiplier/_0428_ ;
 wire \u_multiplier/_0429_ ;
 wire \u_multiplier/_0430_ ;
 wire \u_multiplier/_0431_ ;
 wire \u_multiplier/_0432_ ;
 wire \u_multiplier/_0433_ ;
 wire \u_multiplier/_0434_ ;
 wire \u_multiplier/_0435_ ;
 wire \u_multiplier/_0436_ ;
 wire \u_multiplier/_0437_ ;
 wire \u_multiplier/_0438_ ;
 wire \u_multiplier/_0439_ ;
 wire \u_multiplier/_0440_ ;
 wire \u_multiplier/_0441_ ;
 wire \u_multiplier/_0442_ ;
 wire \u_multiplier/_0443_ ;
 wire \u_multiplier/_0444_ ;
 wire \u_multiplier/_0445_ ;
 wire \u_multiplier/_0446_ ;
 wire \u_multiplier/_0447_ ;
 wire \u_multiplier/_0448_ ;
 wire \u_multiplier/_0449_ ;
 wire \u_multiplier/_0450_ ;
 wire \u_multiplier/_0451_ ;
 wire \u_multiplier/_0452_ ;
 wire \u_multiplier/_0453_ ;
 wire \u_multiplier/_0454_ ;
 wire \u_multiplier/_0455_ ;
 wire \u_multiplier/_0456_ ;
 wire \u_multiplier/_0457_ ;
 wire \u_multiplier/_0458_ ;
 wire \u_multiplier/_0459_ ;
 wire \u_multiplier/_0460_ ;
 wire \u_multiplier/_0461_ ;
 wire \u_multiplier/_0462_ ;
 wire \u_multiplier/_0463_ ;
 wire \u_multiplier/_0464_ ;
 wire \u_multiplier/_0465_ ;
 wire \u_multiplier/_0466_ ;
 wire \u_multiplier/_0467_ ;
 wire \u_multiplier/_0468_ ;
 wire \u_multiplier/_0469_ ;
 wire \u_multiplier/_0470_ ;
 wire \u_multiplier/_0471_ ;
 wire \u_multiplier/_0472_ ;
 wire \u_multiplier/_0473_ ;
 wire \u_multiplier/_0474_ ;
 wire \u_multiplier/_0475_ ;
 wire \u_multiplier/_0476_ ;
 wire \u_multiplier/_0477_ ;
 wire \u_multiplier/_0478_ ;
 wire \u_multiplier/_0479_ ;
 wire \u_multiplier/_0480_ ;
 wire \u_multiplier/_0481_ ;
 wire \u_multiplier/_0482_ ;
 wire \u_multiplier/_0483_ ;
 wire \u_multiplier/_0484_ ;
 wire \u_multiplier/_0485_ ;
 wire \u_multiplier/_0486_ ;
 wire \u_multiplier/_0487_ ;
 wire \u_multiplier/_0488_ ;
 wire \u_multiplier/_0489_ ;
 wire \u_multiplier/_0490_ ;
 wire \u_multiplier/_0491_ ;
 wire \u_multiplier/_0492_ ;
 wire \u_multiplier/_0493_ ;
 wire \u_multiplier/_0494_ ;
 wire \u_multiplier/_0495_ ;
 wire \u_multiplier/_0496_ ;
 wire \u_multiplier/_0497_ ;
 wire \u_multiplier/_0498_ ;
 wire \u_multiplier/_0499_ ;
 wire \u_multiplier/_0500_ ;
 wire \u_multiplier/_0501_ ;
 wire \u_multiplier/_0502_ ;
 wire \u_multiplier/_0503_ ;
 wire \u_multiplier/_0504_ ;
 wire \u_multiplier/_0505_ ;
 wire \u_multiplier/_0506_ ;
 wire \u_multiplier/_0507_ ;
 wire \u_multiplier/_0508_ ;
 wire \u_multiplier/_0509_ ;
 wire \u_multiplier/_0510_ ;
 wire \u_multiplier/_0511_ ;
 wire \u_multiplier/_0512_ ;
 wire \u_multiplier/_0513_ ;
 wire \u_multiplier/_0514_ ;
 wire \u_multiplier/_0515_ ;
 wire \u_multiplier/_0516_ ;
 wire \u_multiplier/_0517_ ;
 wire \u_multiplier/_0518_ ;
 wire \u_multiplier/_0519_ ;
 wire \u_multiplier/_0520_ ;
 wire \u_multiplier/_0521_ ;
 wire \u_multiplier/_0522_ ;
 wire \u_multiplier/_0523_ ;
 wire \u_multiplier/_0524_ ;
 wire \u_multiplier/_0525_ ;
 wire \u_multiplier/_0526_ ;
 wire \u_multiplier/_0527_ ;
 wire \u_multiplier/_0528_ ;
 wire \u_multiplier/_0529_ ;
 wire \u_multiplier/_0530_ ;
 wire \u_multiplier/_0531_ ;
 wire \u_multiplier/_0532_ ;
 wire \u_multiplier/_0533_ ;
 wire \u_multiplier/_0534_ ;
 wire \u_multiplier/_0535_ ;
 wire \u_multiplier/_0536_ ;
 wire \u_multiplier/_0537_ ;
 wire \u_multiplier/_0538_ ;
 wire \u_multiplier/_0539_ ;
 wire \u_multiplier/_0540_ ;
 wire \u_multiplier/_0541_ ;
 wire \u_multiplier/_0542_ ;
 wire \u_multiplier/_0543_ ;
 wire \u_multiplier/_0544_ ;
 wire \u_multiplier/_0545_ ;
 wire \u_multiplier/_0546_ ;
 wire \u_multiplier/_0547_ ;
 wire \u_multiplier/_0548_ ;
 wire \u_multiplier/_0549_ ;
 wire \u_multiplier/_0550_ ;
 wire \u_multiplier/_0551_ ;
 wire \u_multiplier/_0552_ ;
 wire \u_multiplier/_0553_ ;
 wire \u_multiplier/_0554_ ;
 wire \u_multiplier/_0555_ ;
 wire \u_multiplier/_0556_ ;
 wire \u_multiplier/_0557_ ;
 wire \u_multiplier/_0558_ ;
 wire \u_multiplier/_0559_ ;
 wire \u_multiplier/_0560_ ;
 wire \u_multiplier/_0561_ ;
 wire \u_multiplier/_0562_ ;
 wire \u_multiplier/_0563_ ;
 wire \u_multiplier/_0564_ ;
 wire \u_multiplier/_0565_ ;
 wire \u_multiplier/_0566_ ;
 wire \u_multiplier/_0567_ ;
 wire \u_multiplier/_0568_ ;
 wire \u_multiplier/_0569_ ;
 wire \u_multiplier/_0570_ ;
 wire \u_multiplier/_0571_ ;
 wire \u_multiplier/_0572_ ;
 wire \u_multiplier/_0573_ ;
 wire \u_multiplier/_0574_ ;
 wire \u_multiplier/_0575_ ;
 wire \u_multiplier/_0576_ ;
 wire \u_multiplier/_0577_ ;
 wire \u_multiplier/_0578_ ;
 wire \u_multiplier/_0579_ ;
 wire \u_multiplier/_0580_ ;
 wire \u_multiplier/_0581_ ;
 wire \u_multiplier/_0582_ ;
 wire \u_multiplier/_0583_ ;
 wire \u_multiplier/_0584_ ;
 wire \u_multiplier/_0585_ ;
 wire \u_multiplier/_0586_ ;
 wire \u_multiplier/_0587_ ;
 wire \u_multiplier/_0588_ ;
 wire \u_multiplier/_0589_ ;
 wire \u_multiplier/_0590_ ;
 wire \u_multiplier/_0591_ ;
 wire \u_multiplier/_0592_ ;
 wire \u_multiplier/_0593_ ;
 wire \u_multiplier/_0594_ ;
 wire \u_multiplier/_0595_ ;
 wire \u_multiplier/_0596_ ;
 wire \u_multiplier/_0597_ ;
 wire \u_multiplier/_0598_ ;
 wire \u_multiplier/_0599_ ;
 wire \u_multiplier/_0600_ ;
 wire \u_multiplier/_0601_ ;
 wire \u_multiplier/_0602_ ;
 wire \u_multiplier/_0603_ ;
 wire \u_multiplier/_0604_ ;
 wire \u_multiplier/_0605_ ;
 wire \u_multiplier/_0606_ ;
 wire \u_multiplier/_0607_ ;
 wire \u_multiplier/_0608_ ;
 wire \u_multiplier/_0609_ ;
 wire \u_multiplier/_0610_ ;
 wire \u_multiplier/_0611_ ;
 wire \u_multiplier/_0612_ ;
 wire \u_multiplier/_0613_ ;
 wire \u_multiplier/_0614_ ;
 wire \u_multiplier/_0615_ ;
 wire \u_multiplier/_0616_ ;
 wire \u_multiplier/_0617_ ;
 wire \u_multiplier/_0618_ ;
 wire \u_multiplier/_0619_ ;
 wire \u_multiplier/_0620_ ;
 wire \u_multiplier/_0621_ ;
 wire \u_multiplier/_0622_ ;
 wire \u_multiplier/_0623_ ;
 wire \u_multiplier/_0624_ ;
 wire \u_multiplier/_0625_ ;
 wire \u_multiplier/_0626_ ;
 wire \u_multiplier/_0627_ ;
 wire \u_multiplier/_0628_ ;
 wire \u_multiplier/_0629_ ;
 wire \u_multiplier/_0630_ ;
 wire \u_multiplier/_0631_ ;
 wire \u_multiplier/_0632_ ;
 wire \u_multiplier/_0633_ ;
 wire \u_multiplier/_0634_ ;
 wire \u_multiplier/_0635_ ;
 wire \u_multiplier/_0636_ ;
 wire \u_multiplier/_0637_ ;
 wire \u_multiplier/_0638_ ;
 wire \u_multiplier/_0639_ ;
 wire \u_multiplier/_0640_ ;
 wire \u_multiplier/_0641_ ;
 wire \u_multiplier/_0642_ ;
 wire \u_multiplier/_0643_ ;
 wire \u_multiplier/_0644_ ;
 wire \u_multiplier/_0645_ ;
 wire \u_multiplier/_0646_ ;
 wire \u_multiplier/_0647_ ;
 wire \u_multiplier/_0648_ ;
 wire \u_multiplier/_0649_ ;
 wire \u_multiplier/_0650_ ;
 wire \u_multiplier/_0651_ ;
 wire \u_multiplier/_0652_ ;
 wire \u_multiplier/_0653_ ;
 wire \u_multiplier/_0654_ ;
 wire \u_multiplier/_0655_ ;
 wire \u_multiplier/_0656_ ;
 wire \u_multiplier/_0657_ ;
 wire \u_multiplier/_0658_ ;
 wire \u_multiplier/_0659_ ;
 wire \u_multiplier/_0660_ ;
 wire \u_multiplier/_0661_ ;
 wire \u_multiplier/_0662_ ;
 wire \u_multiplier/_0663_ ;
 wire \u_multiplier/_0664_ ;
 wire \u_multiplier/_0665_ ;
 wire \u_multiplier/_0666_ ;
 wire \u_multiplier/_0667_ ;
 wire \u_multiplier/_0668_ ;
 wire \u_multiplier/_0669_ ;
 wire \u_multiplier/_0670_ ;
 wire \u_multiplier/_0671_ ;
 wire \u_multiplier/_0672_ ;
 wire \u_multiplier/_0673_ ;
 wire \u_multiplier/_0674_ ;
 wire \u_multiplier/_0675_ ;
 wire \u_multiplier/_0676_ ;
 wire \u_multiplier/_0677_ ;
 wire \u_multiplier/_0678_ ;
 wire \u_multiplier/_0679_ ;
 wire \u_multiplier/_0680_ ;
 wire \u_multiplier/_0681_ ;
 wire \u_multiplier/_0682_ ;
 wire \u_multiplier/_0683_ ;
 wire \u_multiplier/_0684_ ;
 wire \u_multiplier/_0685_ ;
 wire \u_multiplier/_0686_ ;
 wire \u_multiplier/_0687_ ;
 wire \u_multiplier/_0688_ ;
 wire \u_multiplier/_0689_ ;
 wire \u_multiplier/_0690_ ;
 wire \u_multiplier/_0691_ ;
 wire \u_multiplier/_0692_ ;
 wire \u_multiplier/_0693_ ;
 wire \u_multiplier/_0694_ ;
 wire \u_multiplier/_0695_ ;
 wire \u_multiplier/_0696_ ;
 wire \u_multiplier/_0697_ ;
 wire \u_multiplier/_0698_ ;
 wire \u_multiplier/_0699_ ;
 wire \u_multiplier/_0700_ ;
 wire \u_multiplier/_0701_ ;
 wire \u_multiplier/_0702_ ;
 wire \u_multiplier/_0703_ ;
 wire \u_multiplier/_0704_ ;
 wire \u_multiplier/_0705_ ;
 wire \u_multiplier/_0706_ ;
 wire \u_multiplier/_0707_ ;
 wire \u_multiplier/_0708_ ;
 wire \u_multiplier/_0709_ ;
 wire \u_multiplier/_0710_ ;
 wire \u_multiplier/_0711_ ;
 wire \u_multiplier/_0712_ ;
 wire \u_multiplier/_0713_ ;
 wire \u_multiplier/_0714_ ;
 wire \u_multiplier/_0715_ ;
 wire \u_multiplier/_0716_ ;
 wire \u_multiplier/_0717_ ;
 wire \u_multiplier/_0718_ ;
 wire \u_multiplier/_0719_ ;
 wire \u_multiplier/_0720_ ;
 wire \u_multiplier/_0721_ ;
 wire \u_multiplier/_0722_ ;
 wire \u_multiplier/_0723_ ;
 wire net30;
 wire \u_multiplier/zero_x ;
 wire \u_multiplier/zero_y ;
 wire \u_multiplier/LODx/_12_ ;
 wire \u_multiplier/LODx/_13_ ;
 wire \u_multiplier/LODx/Middle/_3_ ;
 wire \u_multiplier/LODx/lod2_0/_09_ ;
 wire \u_multiplier/LODx/lod2_0/_10_ ;
 wire \u_multiplier/LODx/lod2_0/_11_ ;
 wire \u_multiplier/LODx/lod2_1/_09_ ;
 wire \u_multiplier/LODx/lod2_1/_10_ ;
 wire \u_multiplier/LODx/lod2_1/_11_ ;
 wire \u_multiplier/LODy/_12_ ;
 wire \u_multiplier/LODy/_13_ ;
 wire \u_multiplier/LODy/Middle/_3_ ;
 wire \u_multiplier/LODy/lod2_0/_09_ ;
 wire \u_multiplier/LODy/lod2_0/_10_ ;
 wire \u_multiplier/LODy/lod2_0/_11_ ;
 wire \u_multiplier/LODy/lod2_1/_09_ ;
 wire \u_multiplier/LODy/lod2_1/_10_ ;
 wire \u_multiplier/LODy/lod2_1/_11_ ;
 wire \u_multiplier/NOD/_11_ ;
 wire \u_multiplier/NOD/_12_ ;
 wire \u_multiplier/NOD/_13_ ;
 wire net31;
 wire \u_multiplier/NOD/nod_basic_unit15/_5_ ;
 wire \u_multiplier/NOD/nod_cels[2].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[2].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[2].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[2].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[3].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[3].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[3].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[3].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[4].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[4].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[4].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[4].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/NOD/nod_cels[5].Nod_bits/_02_ ;
 wire \u_multiplier/NOD/nod_cels[5].Nod_bits/_03_ ;
 wire \u_multiplier/NOD/nod_cels[5].Nod_bits/tmp1 ;
 wire \u_multiplier/NOD/nod_cels[5].Nod_bits/nod_basic_unit/_5_ ;
 wire \u_multiplier/dec/_34_ ;
 wire \u_multiplier/dec/_35_ ;
 wire \u_multiplier/dec/_36_ ;
 wire \u_multiplier/dec/_37_ ;
 wire \u_multiplier/dec/_38_ ;
 wire \u_multiplier/dec/_39_ ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire valid_reg_out;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire [3:0] addr_ptr;
 wire [2:0] curr_state;
 wire [7:0] data_in_reg;
 wire [3:0] init_count;
 wire [15:0] product;
 wire [7:0] sram_rdata;
 wire [7:0] sram_rdata_reg;
 wire [2:0] \u_multiplier/K ;
 wire [1:0] \u_multiplier/LODx/select ;
 wire [7:0] \u_multiplier/LODx/z ;
 wire [1:0] \u_multiplier/LODy/select ;
 wire [7:0] \u_multiplier/LODy/z ;
 wire [4:0] \u_multiplier/NOD/t_in ;
 wire [7:0] \u_multiplier/NOD_Q1 ;
 wire [2:0] \u_multiplier/code_x ;
 wire [2:0] \u_multiplier/code_y ;
 wire [15:0] \u_multiplier/dec_out ;
 wire [7:0] \u_multiplier/kx ;
 wire [7:0] \u_multiplier/ky ;

 INV_X2 _281_ (.A(net11),
    .ZN(_165_));
 INV_X4 _282_ (.A(net10),
    .ZN(_134_));
 INV_X1 _283_ (.A(init_count[2]),
    .ZN(_166_));
 INV_X1 _284_ (.A(addr_ptr[0]),
    .ZN(_167_));
 INV_X1 _285_ (.A(addr_ptr[3]),
    .ZN(_168_));
 NAND2_X2 _286_ (.A1(net11),
    .A2(net82),
    .ZN(_135_));
 NAND2_X1 _287_ (.A1(init_count[3]),
    .A2(init_count[2]),
    .ZN(_169_));
 NAND2_X1 _288_ (.A1(init_count[1]),
    .A2(init_count[0]),
    .ZN(_170_));
 NAND4_X4 _289_ (.A1(init_count[1]),
    .A2(init_count[0]),
    .A3(init_count[3]),
    .A4(init_count[2]),
    .ZN(_171_));
 NOR2_X1 _290_ (.A1(_134_),
    .A2(_171_),
    .ZN(_172_));
 NAND3_X1 _291_ (.A1(net11),
    .A2(net10),
    .A3(net9),
    .ZN(_173_));
 OAI22_X1 _292_ (.A1(_135_),
    .A2(_172_),
    .B1(_173_),
    .B2(net57),
    .ZN(_133_));
 OR2_X1 _293_ (.A1(_165_),
    .A2(net85),
    .ZN(_174_));
 AND2_X1 _294_ (.A1(_173_),
    .A2(_174_),
    .ZN(_131_));
 AND2_X4 _295_ (.A1(net11),
    .A2(net12),
    .ZN(_130_));
 NOR3_X1 _296_ (.A1(_134_),
    .A2(_135_),
    .A3(_171_),
    .ZN(_175_));
 OR2_X1 _297_ (.A1(_130_),
    .A2(_175_),
    .ZN(_132_));
 AND2_X1 _298_ (.A1(net11),
    .A2(sram_rdata[0]),
    .ZN(_122_));
 AND2_X1 _299_ (.A1(net11),
    .A2(sram_rdata[1]),
    .ZN(_123_));
 AND2_X1 _300_ (.A1(net11),
    .A2(sram_rdata[2]),
    .ZN(_124_));
 AND2_X1 _301_ (.A1(net11),
    .A2(sram_rdata[3]),
    .ZN(_125_));
 AND2_X1 _302_ (.A1(net11),
    .A2(sram_rdata[4]),
    .ZN(_126_));
 AND2_X1 _303_ (.A1(net11),
    .A2(sram_rdata[5]),
    .ZN(_127_));
 AND2_X1 _304_ (.A1(net11),
    .A2(sram_rdata[6]),
    .ZN(_128_));
 AND2_X1 _305_ (.A1(net11),
    .A2(sram_rdata[7]),
    .ZN(_129_));
 AND2_X1 _306_ (.A1(product[0]),
    .A2(_130_),
    .ZN(_102_));
 AND2_X1 _307_ (.A1(product[1]),
    .A2(_130_),
    .ZN(_109_));
 AND2_X1 _308_ (.A1(product[2]),
    .A2(_130_),
    .ZN(_110_));
 AND2_X1 _309_ (.A1(product[3]),
    .A2(_130_),
    .ZN(_111_));
 AND2_X1 _310_ (.A1(product[4]),
    .A2(_130_),
    .ZN(_112_));
 AND2_X1 _311_ (.A1(product[5]),
    .A2(_130_),
    .ZN(_113_));
 AND2_X1 _312_ (.A1(product[6]),
    .A2(_130_),
    .ZN(_114_));
 AND2_X1 _313_ (.A1(product[7]),
    .A2(_130_),
    .ZN(_115_));
 AND2_X1 _314_ (.A1(product[8]),
    .A2(_130_),
    .ZN(_116_));
 AND2_X1 _315_ (.A1(product[9]),
    .A2(_130_),
    .ZN(_117_));
 AND2_X1 _316_ (.A1(product[10]),
    .A2(_130_),
    .ZN(_103_));
 AND2_X1 _317_ (.A1(product[11]),
    .A2(_130_),
    .ZN(_104_));
 AND2_X1 _318_ (.A1(product[12]),
    .A2(_130_),
    .ZN(_105_));
 AND2_X1 _319_ (.A1(product[13]),
    .A2(_130_),
    .ZN(_106_));
 AND2_X1 _320_ (.A1(product[14]),
    .A2(_130_),
    .ZN(_107_));
 AND2_X1 _321_ (.A1(product[15]),
    .A2(_130_),
    .ZN(_108_));
 AND2_X1 _322_ (.A1(net11),
    .A2(net1),
    .ZN(_094_));
 AND2_X1 _323_ (.A1(net11),
    .A2(net2),
    .ZN(_095_));
 AND2_X1 _324_ (.A1(net11),
    .A2(net3),
    .ZN(_096_));
 AND2_X1 _325_ (.A1(net11),
    .A2(net4),
    .ZN(_097_));
 AND2_X1 _326_ (.A1(net11),
    .A2(net5),
    .ZN(_098_));
 AND2_X1 _327_ (.A1(net11),
    .A2(net6),
    .ZN(_099_));
 AND2_X1 _328_ (.A1(net11),
    .A2(net7),
    .ZN(_100_));
 AND2_X1 _329_ (.A1(net11),
    .A2(net8),
    .ZN(_101_));
 OAI21_X1 _330_ (.A(init_count[0]),
    .B1(_269_),
    .B2(_169_),
    .ZN(_176_));
 AOI221_X2 _331_ (.A(_134_),
    .B1(init_count[0]),
    .B2(net12),
    .C1(_176_),
    .C2(curr_state[2]),
    .ZN(_177_));
 AOI211_X1 _332_ (.A(_165_),
    .B(_177_),
    .C1(net61),
    .C2(_134_),
    .ZN(_118_));
 NAND3_X1 _333_ (.A1(init_count[1]),
    .A2(init_count[0]),
    .A3(_169_),
    .ZN(_178_));
 AOI21_X1 _334_ (.A(_134_),
    .B1(init_count[1]),
    .B2(net12),
    .ZN(_179_));
 OAI211_X1 _335_ (.A(curr_state[2]),
    .B(_178_),
    .C1(init_count[1]),
    .C2(init_count[0]),
    .ZN(_180_));
 AOI221_X1 _336_ (.A(_165_),
    .B1(_134_),
    .B2(net79),
    .C1(_179_),
    .C2(_180_),
    .ZN(_119_));
 OR2_X1 _337_ (.A1(init_count[3]),
    .A2(_166_),
    .ZN(_181_));
 NAND2_X1 _338_ (.A1(_166_),
    .A2(_170_),
    .ZN(_182_));
 OAI211_X1 _339_ (.A(curr_state[2]),
    .B(_182_),
    .C1(_181_),
    .C2(_170_),
    .ZN(_183_));
 AOI21_X1 _340_ (.A(_134_),
    .B1(init_count[2]),
    .B2(net12),
    .ZN(_184_));
 AOI221_X1 _341_ (.A(_165_),
    .B1(_134_),
    .B2(net72),
    .C1(_183_),
    .C2(_184_),
    .ZN(_120_));
 NAND2_X1 _342_ (.A1(init_count[3]),
    .A2(net12),
    .ZN(_185_));
 OAI21_X1 _343_ (.A(net76),
    .B1(_170_),
    .B2(net71),
    .ZN(_186_));
 OAI21_X1 _344_ (.A(_186_),
    .B1(curr_state[2]),
    .B2(_134_),
    .ZN(_187_));
 AOI221_X1 _345_ (.A(_165_),
    .B1(_134_),
    .B2(net39),
    .C1(_185_),
    .C2(_187_),
    .ZN(_121_));
 NAND3_X1 _346_ (.A1(curr_state[2]),
    .A2(net63),
    .A3(_171_),
    .ZN(_188_));
 AOI21_X1 _347_ (.A(_134_),
    .B1(net12),
    .B2(_167_),
    .ZN(_189_));
 AOI221_X1 _348_ (.A(_165_),
    .B1(_134_),
    .B2(net40),
    .C1(net64),
    .C2(_189_),
    .ZN(_090_));
 AOI21_X2 _349_ (.A(net12),
    .B1(_171_),
    .B2(curr_state[2]),
    .ZN(_190_));
 NAND2_X1 _350_ (.A1(addr_ptr[0]),
    .A2(addr_ptr[1]),
    .ZN(_191_));
 XNOR2_X1 _351_ (.A(addr_ptr[0]),
    .B(addr_ptr[1]),
    .ZN(_192_));
 OAI21_X1 _352_ (.A(net10),
    .B1(_190_),
    .B2(_192_),
    .ZN(_193_));
 AOI21_X1 _353_ (.A(_165_),
    .B1(_134_),
    .B2(net47),
    .ZN(_194_));
 AND2_X1 _354_ (.A1(_193_),
    .A2(net48),
    .ZN(_091_));
 XOR2_X1 _355_ (.A(addr_ptr[2]),
    .B(_191_),
    .Z(_195_));
 OAI21_X1 _356_ (.A(net10),
    .B1(_190_),
    .B2(_195_),
    .ZN(_196_));
 AOI21_X1 _357_ (.A(_165_),
    .B1(_134_),
    .B2(net49),
    .ZN(_197_));
 AND2_X1 _358_ (.A1(_196_),
    .A2(net50),
    .ZN(_092_));
 AOI21_X1 _359_ (.A(_168_),
    .B1(_171_),
    .B2(curr_state[2]),
    .ZN(_198_));
 NAND4_X1 _360_ (.A1(net10),
    .A2(addr_ptr[0]),
    .A3(addr_ptr[1]),
    .A4(addr_ptr[2]),
    .ZN(_199_));
 OR2_X1 _361_ (.A1(_198_),
    .A2(_199_),
    .ZN(_200_));
 OAI21_X1 _362_ (.A(net11),
    .B1(net53),
    .B2(_199_),
    .ZN(_201_));
 AOI221_X1 _363_ (.A(net54),
    .B1(_200_),
    .B2(net34),
    .C1(net10),
    .C2(_190_),
    .ZN(_093_));
 DFF_X1 _364_ (.D(_102_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net13),
    .QN(_228_));
 DFF_X1 _365_ (.D(_109_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net20),
    .QN(_229_));
 DFF_X1 _366_ (.D(_110_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net21),
    .QN(_230_));
 DFF_X1 _367_ (.D(_111_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net22),
    .QN(_231_));
 DFF_X1 _368_ (.D(_112_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net23),
    .QN(_232_));
 DFF_X2 _369_ (.D(_113_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net24),
    .QN(_233_));
 DFF_X1 _370_ (.D(_114_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net25),
    .QN(_234_));
 DFF_X1 _371_ (.D(_115_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net26),
    .QN(_235_));
 DFF_X1 _372_ (.D(_116_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net27),
    .QN(_236_));
 DFF_X2 _373_ (.D(_117_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net28),
    .QN(_237_));
 DFF_X1 _374_ (.D(_103_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net14),
    .QN(_238_));
 DFF_X1 _375_ (.D(_104_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net15),
    .QN(_239_));
 DFF_X1 _376_ (.D(_105_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net16),
    .QN(_240_));
 DFF_X1 _377_ (.D(_106_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net17),
    .QN(_241_));
 DFF_X1 _378_ (.D(_107_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net18),
    .QN(_242_));
 DFF_X1 _379_ (.D(_108_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net19),
    .QN(_243_));
 DFF_X1 _380_ (.D(_131_),
    .CK(clknet_2_1__leaf_clk),
    .Q(curr_state[0]),
    .QN(_244_));
 DFF_X2 _381_ (.D(_132_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net12),
    .QN(_245_));
 DFF_X2 _382_ (.D(net58),
    .CK(clknet_2_1__leaf_clk),
    .Q(curr_state[2]),
    .QN(_246_));
 DFF_X2 _383_ (.D(_094_),
    .CK(clknet_2_0__leaf_clk),
    .Q(data_in_reg[0]),
    .QN(_247_));
 DFF_X2 _384_ (.D(_095_),
    .CK(clknet_2_2__leaf_clk),
    .Q(data_in_reg[1]),
    .QN(_248_));
 DFF_X2 _385_ (.D(_096_),
    .CK(clknet_2_2__leaf_clk),
    .Q(data_in_reg[2]),
    .QN(_249_));
 DFF_X2 _386_ (.D(_097_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\u_multiplier/LODx/z [3]),
    .QN(_250_));
 DFF_X2 _387_ (.D(_098_),
    .CK(clknet_2_2__leaf_clk),
    .Q(data_in_reg[4]),
    .QN(_251_));
 DFF_X2 _388_ (.D(_099_),
    .CK(clknet_2_2__leaf_clk),
    .Q(data_in_reg[5]),
    .QN(_252_));
 DFF_X2 _389_ (.D(_100_),
    .CK(clknet_2_0__leaf_clk),
    .Q(data_in_reg[6]),
    .QN(_253_));
 DFF_X2 _390_ (.D(_101_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\u_multiplier/LODx/z [7]),
    .QN(_254_));
 DFF_X2 _391_ (.D(_122_),
    .CK(clknet_2_0__leaf_clk),
    .Q(sram_rdata_reg[0]),
    .QN(_255_));
 DFF_X2 _392_ (.D(_123_),
    .CK(clknet_2_0__leaf_clk),
    .Q(sram_rdata_reg[1]),
    .QN(_256_));
 DFF_X2 _393_ (.D(_124_),
    .CK(clknet_2_0__leaf_clk),
    .Q(sram_rdata_reg[2]),
    .QN(_257_));
 DFF_X2 _394_ (.D(_125_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\u_multiplier/LODy/z [3]),
    .QN(_258_));
 DFF_X2 _395_ (.D(_126_),
    .CK(clknet_2_2__leaf_clk),
    .Q(sram_rdata_reg[4]),
    .QN(_259_));
 DFF_X2 _396_ (.D(_127_),
    .CK(clknet_2_2__leaf_clk),
    .Q(sram_rdata_reg[5]),
    .QN(_260_));
 DFF_X2 _397_ (.D(_128_),
    .CK(clknet_2_2__leaf_clk),
    .Q(sram_rdata_reg[6]),
    .QN(_261_));
 DFF_X2 _398_ (.D(_129_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\u_multiplier/LODy/z [7]),
    .QN(_262_));
 DFF_X1 _399_ (.D(_130_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net29),
    .QN(_263_));
 DFF_X2 _400_ (.D(_090_),
    .CK(clknet_2_1__leaf_clk),
    .Q(addr_ptr[0]),
    .QN(_264_));
 DFF_X1 _401_ (.D(_091_),
    .CK(clknet_2_1__leaf_clk),
    .Q(addr_ptr[1]),
    .QN(_265_));
 DFF_X1 _402_ (.D(_092_),
    .CK(clknet_2_1__leaf_clk),
    .Q(addr_ptr[2]),
    .QN(_266_));
 DFF_X1 _403_ (.D(net55),
    .CK(clknet_2_1__leaf_clk),
    .Q(addr_ptr[3]),
    .QN(_267_));
 DFF_X2 _404_ (.D(net62),
    .CK(clknet_2_1__leaf_clk),
    .Q(init_count[0]),
    .QN(_268_));
 DFF_X2 _405_ (.D(net80),
    .CK(clknet_2_1__leaf_clk),
    .Q(init_count[1]),
    .QN(_269_));
 DFF_X2 _406_ (.D(net73),
    .CK(clknet_2_1__leaf_clk),
    .Q(init_count[2]),
    .QN(_270_));
 DFF_X2 _407_ (.D(net77),
    .CK(clknet_2_1__leaf_clk),
    .Q(init_count[3]),
    .QN(_271_));
 SRAM_6T_CORE_16x8_MC_TB sram_inst (.ce_in(_134_),
    .we_in(_135_),
    .clk(clknet_2_0__leaf_clk),
    .addr_in({net68,
    net70,
    net66,
    net75}),
    .rd_out({sram_rdata[7],
    sram_rdata[6],
    sram_rdata[5],
    sram_rdata[4],
    sram_rdata[3],
    sram_rdata[2],
    sram_rdata[1],
    sram_rdata[0]}),
    .wd_in({net42,
    net59,
    net43,
    net44,
    net52,
    net51,
    net46,
    net45}));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_0/_09_  (.A1(\u_multiplier/LODx/z [1]),
    .A2(\u_multiplier/LODx/select [0]),
    .ZN(\u_multiplier/kx [1]));
 AND2_X1 \u_multiplier/LODx/Inst_MUX214_0/_10_  (.A1(\u_multiplier/LODx/select [0]),
    .A2(\u_multiplier/LODx/z [0]),
    .ZN(\u_multiplier/kx [0]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_0/_11_  (.A1(\u_multiplier/LODx/select [0]),
    .A2(\u_multiplier/LODx/z [3]),
    .ZN(\u_multiplier/kx [3]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_0/_12_  (.A1(\u_multiplier/LODx/select [0]),
    .A2(\u_multiplier/LODx/z [2]),
    .ZN(\u_multiplier/kx [2]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_1/_09_  (.A1(\u_multiplier/LODx/z [5]),
    .A2(\u_multiplier/LODx/select [1]),
    .ZN(\u_multiplier/kx [5]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_1/_10_  (.A1(\u_multiplier/LODx/select [1]),
    .A2(\u_multiplier/LODx/z [4]),
    .ZN(\u_multiplier/kx [4]));
 AND2_X1 \u_multiplier/LODx/Inst_MUX214_1/_11_  (.A1(\u_multiplier/LODx/select [1]),
    .A2(\u_multiplier/LODx/z [7]),
    .ZN(\u_multiplier/kx [7]));
 AND2_X2 \u_multiplier/LODx/Inst_MUX214_1/_12_  (.A1(\u_multiplier/LODx/select [1]),
    .A2(\u_multiplier/LODx/z [6]),
    .ZN(\u_multiplier/kx [6]));
 INV_X1 \u_multiplier/LODx/Middle/_4_  (.A(\u_multiplier/LODx/_12_ ),
    .ZN(\u_multiplier/LODx/Middle/_3_ ));
 NOR2_X1 \u_multiplier/LODx/Middle/_5_  (.A1(\u_multiplier/LODx/Middle/_3_ ),
    .A2(\u_multiplier/LODx/select [1]),
    .ZN(\u_multiplier/LODx/select [0]));
 OR4_X1 \u_multiplier/LODx/_15_  (.A1(data_in_reg[2]),
    .A2(\u_multiplier/LODx/z [3]),
    .A3(data_in_reg[0]),
    .A4(data_in_reg[1]),
    .ZN(\u_multiplier/LODx/_12_ ));
 OR4_X2 \u_multiplier/LODx/_16_  (.A1(data_in_reg[6]),
    .A2(\u_multiplier/LODx/z [7]),
    .A3(data_in_reg[4]),
    .A4(data_in_reg[5]),
    .ZN(\u_multiplier/LODx/select [1]));
 NOR2_X2 \u_multiplier/LODx/_17_  (.A1(\u_multiplier/LODx/_12_ ),
    .A2(\u_multiplier/LODx/select [1]),
    .ZN(\u_multiplier/zero_x ));
 INV_X1 \u_multiplier/LODx/lod2_0/_12_  (.A(data_in_reg[2]),
    .ZN(\u_multiplier/LODx/lod2_0/_10_ ));
 INV_X1 \u_multiplier/LODx/lod2_0/_13_  (.A(data_in_reg[1]),
    .ZN(\u_multiplier/LODx/lod2_0/_11_ ));
 INV_X1 \u_multiplier/LODx/lod2_0/_14_  (.A(data_in_reg[0]),
    .ZN(\u_multiplier/LODx/lod2_0/_09_ ));
 NOR2_X1 \u_multiplier/LODx/lod2_0/_15_  (.A1(\u_multiplier/LODx/lod2_0/_10_ ),
    .A2(\u_multiplier/LODx/z [3]),
    .ZN(\u_multiplier/LODx/z [2]));
 NOR3_X1 \u_multiplier/LODx/lod2_0/_16_  (.A1(data_in_reg[2]),
    .A2(\u_multiplier/LODx/z [3]),
    .A3(\u_multiplier/LODx/lod2_0/_11_ ),
    .ZN(\u_multiplier/LODx/z [1]));
 NOR4_X1 \u_multiplier/LODx/lod2_0/_17_  (.A1(data_in_reg[2]),
    .A2(\u_multiplier/LODx/z [3]),
    .A3(data_in_reg[1]),
    .A4(\u_multiplier/LODx/lod2_0/_09_ ),
    .ZN(\u_multiplier/LODx/z [0]));
 INV_X1 \u_multiplier/LODx/lod2_1/_12_  (.A(data_in_reg[6]),
    .ZN(\u_multiplier/LODx/lod2_1/_10_ ));
 INV_X1 \u_multiplier/LODx/lod2_1/_13_  (.A(data_in_reg[5]),
    .ZN(\u_multiplier/LODx/lod2_1/_11_ ));
 INV_X1 \u_multiplier/LODx/lod2_1/_14_  (.A(data_in_reg[4]),
    .ZN(\u_multiplier/LODx/lod2_1/_09_ ));
 NOR2_X1 \u_multiplier/LODx/lod2_1/_15_  (.A1(\u_multiplier/LODx/lod2_1/_10_ ),
    .A2(\u_multiplier/LODx/z [7]),
    .ZN(\u_multiplier/LODx/z [6]));
 NOR3_X1 \u_multiplier/LODx/lod2_1/_16_  (.A1(data_in_reg[6]),
    .A2(\u_multiplier/LODx/z [7]),
    .A3(\u_multiplier/LODx/lod2_1/_11_ ),
    .ZN(\u_multiplier/LODx/z [5]));
 NOR4_X1 \u_multiplier/LODx/lod2_1/_17_  (.A1(data_in_reg[6]),
    .A2(\u_multiplier/LODx/z [7]),
    .A3(data_in_reg[5]),
    .A4(\u_multiplier/LODx/lod2_1/_09_ ),
    .ZN(\u_multiplier/LODx/z [4]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_0/_09_  (.A1(\u_multiplier/LODy/z [1]),
    .A2(\u_multiplier/LODy/select [0]),
    .ZN(\u_multiplier/ky [1]));
 AND2_X1 \u_multiplier/LODy/Inst_MUX214_0/_10_  (.A1(\u_multiplier/LODy/select [0]),
    .A2(\u_multiplier/LODy/z [0]),
    .ZN(\u_multiplier/ky [0]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_0/_11_  (.A1(\u_multiplier/LODy/select [0]),
    .A2(\u_multiplier/LODy/z [3]),
    .ZN(\u_multiplier/ky [3]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_0/_12_  (.A1(\u_multiplier/LODy/select [0]),
    .A2(\u_multiplier/LODy/z [2]),
    .ZN(\u_multiplier/ky [2]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_1/_09_  (.A1(\u_multiplier/LODy/z [5]),
    .A2(\u_multiplier/LODy/select [1]),
    .ZN(\u_multiplier/ky [5]));
 AND2_X1 \u_multiplier/LODy/Inst_MUX214_1/_10_  (.A1(\u_multiplier/LODy/select [1]),
    .A2(\u_multiplier/LODy/z [4]),
    .ZN(\u_multiplier/ky [4]));
 AND2_X1 \u_multiplier/LODy/Inst_MUX214_1/_11_  (.A1(\u_multiplier/LODy/select [1]),
    .A2(\u_multiplier/LODy/z [7]),
    .ZN(\u_multiplier/ky [7]));
 AND2_X2 \u_multiplier/LODy/Inst_MUX214_1/_12_  (.A1(\u_multiplier/LODy/select [1]),
    .A2(\u_multiplier/LODy/z [6]),
    .ZN(\u_multiplier/ky [6]));
 INV_X1 \u_multiplier/LODy/Middle/_4_  (.A(\u_multiplier/LODy/_12_ ),
    .ZN(\u_multiplier/LODy/Middle/_3_ ));
 NOR2_X1 \u_multiplier/LODy/Middle/_5_  (.A1(\u_multiplier/LODy/Middle/_3_ ),
    .A2(\u_multiplier/LODy/select [1]),
    .ZN(\u_multiplier/LODy/select [0]));
 OR4_X1 \u_multiplier/LODy/_15_  (.A1(sram_rdata_reg[2]),
    .A2(\u_multiplier/LODy/z [3]),
    .A3(sram_rdata_reg[0]),
    .A4(sram_rdata_reg[1]),
    .ZN(\u_multiplier/LODy/_12_ ));
 OR4_X2 \u_multiplier/LODy/_16_  (.A1(sram_rdata_reg[6]),
    .A2(\u_multiplier/LODy/z [7]),
    .A3(sram_rdata_reg[4]),
    .A4(sram_rdata_reg[5]),
    .ZN(\u_multiplier/LODy/select [1]));
 NOR2_X2 \u_multiplier/LODy/_17_  (.A1(\u_multiplier/LODy/_12_ ),
    .A2(\u_multiplier/LODy/select [1]),
    .ZN(\u_multiplier/zero_y ));
 INV_X1 \u_multiplier/LODy/lod2_0/_12_  (.A(sram_rdata_reg[2]),
    .ZN(\u_multiplier/LODy/lod2_0/_10_ ));
 INV_X1 \u_multiplier/LODy/lod2_0/_13_  (.A(sram_rdata_reg[1]),
    .ZN(\u_multiplier/LODy/lod2_0/_11_ ));
 INV_X1 \u_multiplier/LODy/lod2_0/_14_  (.A(sram_rdata_reg[0]),
    .ZN(\u_multiplier/LODy/lod2_0/_09_ ));
 NOR2_X1 \u_multiplier/LODy/lod2_0/_15_  (.A1(\u_multiplier/LODy/lod2_0/_10_ ),
    .A2(\u_multiplier/LODy/z [3]),
    .ZN(\u_multiplier/LODy/z [2]));
 NOR3_X1 \u_multiplier/LODy/lod2_0/_16_  (.A1(sram_rdata_reg[2]),
    .A2(\u_multiplier/LODy/z [3]),
    .A3(\u_multiplier/LODy/lod2_0/_11_ ),
    .ZN(\u_multiplier/LODy/z [1]));
 NOR4_X1 \u_multiplier/LODy/lod2_0/_17_  (.A1(sram_rdata_reg[2]),
    .A2(\u_multiplier/LODy/z [3]),
    .A3(sram_rdata_reg[1]),
    .A4(\u_multiplier/LODy/lod2_0/_09_ ),
    .ZN(\u_multiplier/LODy/z [0]));
 INV_X1 \u_multiplier/LODy/lod2_1/_12_  (.A(sram_rdata_reg[6]),
    .ZN(\u_multiplier/LODy/lod2_1/_10_ ));
 INV_X1 \u_multiplier/LODy/lod2_1/_13_  (.A(sram_rdata_reg[5]),
    .ZN(\u_multiplier/LODy/lod2_1/_11_ ));
 INV_X1 \u_multiplier/LODy/lod2_1/_14_  (.A(sram_rdata_reg[4]),
    .ZN(\u_multiplier/LODy/lod2_1/_09_ ));
 NOR2_X1 \u_multiplier/LODy/lod2_1/_15_  (.A1(\u_multiplier/LODy/lod2_1/_10_ ),
    .A2(\u_multiplier/LODy/z [7]),
    .ZN(\u_multiplier/LODy/z [6]));
 NOR3_X1 \u_multiplier/LODy/lod2_1/_16_  (.A1(sram_rdata_reg[6]),
    .A2(\u_multiplier/LODy/z [7]),
    .A3(\u_multiplier/LODy/lod2_1/_11_ ),
    .ZN(\u_multiplier/LODy/z [5]));
 NOR4_X1 \u_multiplier/LODy/lod2_1/_17_  (.A1(sram_rdata_reg[6]),
    .A2(\u_multiplier/LODy/z [7]),
    .A3(sram_rdata_reg[5]),
    .A4(\u_multiplier/LODy/lod2_1/_09_ ),
    .ZN(\u_multiplier/LODy/z [4]));
 INV_X1 \u_multiplier/NOD/_15_  (.A(\u_multiplier/NOD/t_in [1]),
    .ZN(\u_multiplier/NOD/_11_ ));
 INV_X1 \u_multiplier/NOD/_16_  (.A(\u_multiplier/_0346_ ),
    .ZN(\u_multiplier/NOD/_12_ ));
 INV_X1 \u_multiplier/NOD/_17_  (.A(\u_multiplier/_0345_ ),
    .ZN(\u_multiplier/NOD/_13_ ));
 AND2_X1 \u_multiplier/NOD/_18_  (.A1(\u_multiplier/_0350_ ),
    .A2(\u_multiplier/_0351_ ),
    .ZN(\u_multiplier/NOD_Q1 [7]));
 NOR4_X2 \u_multiplier/NOD/_19_  (.A1(\u_multiplier/_0347_ ),
    .A2(\u_multiplier/NOD/_11_ ),
    .A3(\u_multiplier/NOD/_12_ ),
    .A4(\u_multiplier/_0345_ ),
    .ZN(\u_multiplier/NOD_Q1 [1]));
 NOR4_X1 \u_multiplier/NOD/_20_  (.A1(\u_multiplier/_0347_ ),
    .A2(\u_multiplier/NOD/_11_ ),
    .A3(\u_multiplier/_0346_ ),
    .A4(\u_multiplier/NOD/_13_ ),
    .ZN(\u_multiplier/NOD_Q1 [0]));
 AOI21_X1 \u_multiplier/NOD/nod_basic_unit15/_7_  (.A(\u_multiplier/_0351_ ),
    .B1(\u_multiplier/_0349_ ),
    .B2(\u_multiplier/_0350_ ),
    .ZN(\u_multiplier/NOD/nod_basic_unit15/_5_ ));
 AOI21_X2 \u_multiplier/NOD/nod_basic_unit15/_8_  (.A(\u_multiplier/NOD/nod_basic_unit15/_5_ ),
    .B1(\u_multiplier/_0351_ ),
    .B2(\u_multiplier/_0350_ ),
    .ZN(\u_multiplier/NOD_Q1 [6]));
 INV_X1 \u_multiplier/NOD/nod_cels[2].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [2]),
    .ZN(\u_multiplier/NOD/nod_cels[2].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[2].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[2].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[2].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[2].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[2].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0348_ ),
    .ZN(\u_multiplier/NOD/t_in [1]));
 NOR3_X1 \u_multiplier/NOD/nod_cels[2].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[2].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0348_ ),
    .A3(\u_multiplier/NOD/nod_cels[2].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [2]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[2].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_0347_ ),
    .B1(\u_multiplier/_0345_ ),
    .B2(\u_multiplier/_0346_ ),
    .ZN(\u_multiplier/NOD/nod_cels[2].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[2].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[2].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_0347_ ),
    .B2(\u_multiplier/_0346_ ),
    .ZN(\u_multiplier/NOD/nod_cels[2].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[3].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [3]),
    .ZN(\u_multiplier/NOD/nod_cels[3].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[3].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[3].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[3].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[3].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[3].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0349_ ),
    .ZN(\u_multiplier/NOD/t_in [2]));
 NOR3_X2 \u_multiplier/NOD/nod_cels[3].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[3].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0349_ ),
    .A3(\u_multiplier/NOD/nod_cels[3].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [3]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[3].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_0348_ ),
    .B1(\u_multiplier/_0346_ ),
    .B2(\u_multiplier/_0347_ ),
    .ZN(\u_multiplier/NOD/nod_cels[3].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[3].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[3].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_0348_ ),
    .B2(\u_multiplier/_0347_ ),
    .ZN(\u_multiplier/NOD/nod_cels[3].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[4].Nod_bits/_07_  (.A(\u_multiplier/NOD/t_in [4]),
    .ZN(\u_multiplier/NOD/nod_cels[4].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[4].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[4].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[4].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[4].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[4].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0350_ ),
    .ZN(\u_multiplier/NOD/t_in [3]));
 NOR3_X1 \u_multiplier/NOD/nod_cels[4].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[4].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0350_ ),
    .A3(\u_multiplier/NOD/nod_cels[4].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [4]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[4].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_0349_ ),
    .B1(\u_multiplier/_0347_ ),
    .B2(\u_multiplier/_0348_ ),
    .ZN(\u_multiplier/NOD/nod_cels[4].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[4].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[4].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_0349_ ),
    .B2(\u_multiplier/_0348_ ),
    .ZN(\u_multiplier/NOD/nod_cels[4].Nod_bits/tmp1 ));
 INV_X1 \u_multiplier/NOD/nod_cels[5].Nod_bits/_07_  (.A(net30),
    .ZN(\u_multiplier/NOD/nod_cels[5].Nod_bits/_02_ ));
 INV_X1 \u_multiplier/NOD/nod_cels[5].Nod_bits/_08_  (.A(\u_multiplier/NOD/nod_cels[5].Nod_bits/tmp1 ),
    .ZN(\u_multiplier/NOD/nod_cels[5].Nod_bits/_03_ ));
 NOR2_X1 \u_multiplier/NOD/nod_cels[5].Nod_bits/_09_  (.A1(\u_multiplier/NOD/nod_cels[5].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0351_ ),
    .ZN(\u_multiplier/NOD/t_in [4]));
 NOR3_X2 \u_multiplier/NOD/nod_cels[5].Nod_bits/_10_  (.A1(\u_multiplier/NOD/nod_cels[5].Nod_bits/_02_ ),
    .A2(\u_multiplier/_0351_ ),
    .A3(\u_multiplier/NOD/nod_cels[5].Nod_bits/_03_ ),
    .ZN(\u_multiplier/NOD_Q1 [5]));
 AOI21_X1 \u_multiplier/NOD/nod_cels[5].Nod_bits/nod_basic_unit/_7_  (.A(\u_multiplier/_0350_ ),
    .B1(\u_multiplier/_0348_ ),
    .B2(\u_multiplier/_0349_ ),
    .ZN(\u_multiplier/NOD/nod_cels[5].Nod_bits/nod_basic_unit/_5_ ));
 AOI21_X1 \u_multiplier/NOD/nod_cels[5].Nod_bits/nod_basic_unit/_8_  (.A(\u_multiplier/NOD/nod_cels[5].Nod_bits/nod_basic_unit/_5_ ),
    .B1(\u_multiplier/_0350_ ),
    .B2(\u_multiplier/_0349_ ),
    .ZN(\u_multiplier/NOD/nod_cels[5].Nod_bits/tmp1 ));
 OR4_X4 \u_multiplier/PE/code0/_7_  (.A1(\u_multiplier/NOD_Q1 [5]),
    .A2(\u_multiplier/NOD_Q1 [1]),
    .A3(\u_multiplier/NOD_Q1 [7]),
    .A4(\u_multiplier/NOD_Q1 [3]),
    .ZN(\u_multiplier/K [0]));
 OR4_X4 \u_multiplier/PE/code1/_7_  (.A1(\u_multiplier/NOD_Q1 [6]),
    .A2(\u_multiplier/NOD_Q1 [2]),
    .A3(\u_multiplier/NOD_Q1 [7]),
    .A4(\u_multiplier/NOD_Q1 [3]),
    .ZN(\u_multiplier/K [1]));
 OR4_X4 \u_multiplier/PE/code2/_7_  (.A1(\u_multiplier/NOD_Q1 [6]),
    .A2(\u_multiplier/NOD_Q1 [4]),
    .A3(\u_multiplier/NOD_Q1 [7]),
    .A4(\u_multiplier/NOD_Q1 [5]),
    .ZN(\u_multiplier/K [2]));
 OR4_X4 \u_multiplier/PEx/code0/_7_  (.A1(\u_multiplier/kx [5]),
    .A2(\u_multiplier/kx [1]),
    .A3(\u_multiplier/kx [7]),
    .A4(\u_multiplier/kx [3]),
    .ZN(\u_multiplier/code_x [0]));
 OR4_X4 \u_multiplier/PEx/code1/_7_  (.A1(\u_multiplier/kx [6]),
    .A2(\u_multiplier/kx [2]),
    .A3(\u_multiplier/kx [7]),
    .A4(\u_multiplier/kx [3]),
    .ZN(\u_multiplier/code_x [1]));
 OR4_X4 \u_multiplier/PEx/code2/_7_  (.A1(\u_multiplier/kx [6]),
    .A2(\u_multiplier/kx [4]),
    .A3(\u_multiplier/kx [7]),
    .A4(\u_multiplier/kx [5]),
    .ZN(\u_multiplier/code_x [2]));
 OR4_X4 \u_multiplier/PEy/code0/_7_  (.A1(\u_multiplier/ky [5]),
    .A2(\u_multiplier/ky [1]),
    .A3(\u_multiplier/ky [7]),
    .A4(\u_multiplier/ky [3]),
    .ZN(\u_multiplier/code_y [0]));
 OR4_X4 \u_multiplier/PEy/code1/_7_  (.A1(\u_multiplier/ky [6]),
    .A2(\u_multiplier/ky [2]),
    .A3(\u_multiplier/ky [7]),
    .A4(\u_multiplier/ky [3]),
    .ZN(\u_multiplier/code_y [1]));
 OR4_X4 \u_multiplier/PEy/code2/_7_  (.A1(\u_multiplier/ky [6]),
    .A2(\u_multiplier/ky [4]),
    .A3(\u_multiplier/ky [7]),
    .A4(\u_multiplier/ky [5]),
    .ZN(\u_multiplier/code_y [2]));
 INV_X1 \u_multiplier/_0756_  (.A(\u_multiplier/code_y [2]),
    .ZN(\u_multiplier/_0707_ ));
 INV_X1 \u_multiplier/_0757_  (.A(\u_multiplier/code_x [2]),
    .ZN(\u_multiplier/_0708_ ));
 INV_X2 \u_multiplier/_0758_  (.A(\u_multiplier/K [0]),
    .ZN(\u_multiplier/_0709_ ));
 INV_X2 \u_multiplier/_0759_  (.A(\u_multiplier/K [1]),
    .ZN(\u_multiplier/_0710_ ));
 INV_X4 \u_multiplier/_0760_  (.A(\u_multiplier/K [2]),
    .ZN(\u_multiplier/_0711_ ));
 INV_X1 \u_multiplier/_0761_  (.A(\u_multiplier/dec_out [12]),
    .ZN(\u_multiplier/_0712_ ));
 INV_X1 \u_multiplier/_0762_  (.A(\u_multiplier/dec_out [15]),
    .ZN(\u_multiplier/_0713_ ));
 XNOR2_X2 \u_multiplier/_0763_  (.A(\u_multiplier/ky [0]),
    .B(sram_rdata_reg[0]),
    .ZN(\u_multiplier/_0714_ ));
 XOR2_X2 \u_multiplier/_0764_  (.A(\u_multiplier/ky [0]),
    .B(sram_rdata_reg[0]),
    .Z(\u_multiplier/_0715_ ));
 XOR2_X2 \u_multiplier/_0765_  (.A(\u_multiplier/kx [6]),
    .B(data_in_reg[6]),
    .Z(\u_multiplier/_0716_ ));
 XNOR2_X2 \u_multiplier/_0766_  (.A(\u_multiplier/kx [6]),
    .B(data_in_reg[6]),
    .ZN(\u_multiplier/_0717_ ));
 XOR2_X2 \u_multiplier/_0767_  (.A(\u_multiplier/ky [6]),
    .B(sram_rdata_reg[6]),
    .Z(\u_multiplier/_0718_ ));
 XNOR2_X2 \u_multiplier/_0768_  (.A(\u_multiplier/ky [6]),
    .B(sram_rdata_reg[6]),
    .ZN(\u_multiplier/_0719_ ));
 NOR2_X2 \u_multiplier/_0769_  (.A1(\u_multiplier/_0716_ ),
    .A2(\u_multiplier/_0719_ ),
    .ZN(\u_multiplier/_0720_ ));
 XOR2_X2 \u_multiplier/_0770_  (.A(\u_multiplier/ky [1]),
    .B(sram_rdata_reg[1]),
    .Z(\u_multiplier/_0721_ ));
 XNOR2_X2 \u_multiplier/_0771_  (.A(\u_multiplier/ky [1]),
    .B(sram_rdata_reg[1]),
    .ZN(\u_multiplier/_0722_ ));
 XNOR2_X2 \u_multiplier/_0772_  (.A(\u_multiplier/kx [1]),
    .B(data_in_reg[1]),
    .ZN(\u_multiplier/_0723_ ));
 XOR2_X2 \u_multiplier/_0773_  (.A(\u_multiplier/kx [1]),
    .B(data_in_reg[1]),
    .Z(\u_multiplier/_0392_ ));
 XNOR2_X2 \u_multiplier/_0774_  (.A(\u_multiplier/kx [0]),
    .B(data_in_reg[0]),
    .ZN(\u_multiplier/_0393_ ));
 XOR2_X2 \u_multiplier/_0775_  (.A(\u_multiplier/kx [0]),
    .B(data_in_reg[0]),
    .Z(\u_multiplier/_0394_ ));
 AOI211_X1 \u_multiplier/_0776_  (.A(\u_multiplier/_0715_ ),
    .B(\u_multiplier/_0393_ ),
    .C1(\u_multiplier/_0723_ ),
    .C2(\u_multiplier/_0721_ ),
    .ZN(\u_multiplier/_0395_ ));
 OAI211_X1 \u_multiplier/_0777_  (.A(\u_multiplier/_0714_ ),
    .B(\u_multiplier/_0394_ ),
    .C1(\u_multiplier/_0392_ ),
    .C2(\u_multiplier/_0722_ ),
    .ZN(\u_multiplier/_0396_ ));
 XOR2_X2 \u_multiplier/_0778_  (.A(\u_multiplier/ky [2]),
    .B(sram_rdata_reg[2]),
    .Z(\u_multiplier/_0397_ ));
 XNOR2_X2 \u_multiplier/_0779_  (.A(\u_multiplier/ky [2]),
    .B(sram_rdata_reg[2]),
    .ZN(\u_multiplier/_0398_ ));
 XNOR2_X2 \u_multiplier/_0780_  (.A(\u_multiplier/kx [2]),
    .B(data_in_reg[2]),
    .ZN(\u_multiplier/_0399_ ));
 XOR2_X2 \u_multiplier/_0781_  (.A(\u_multiplier/kx [2]),
    .B(data_in_reg[2]),
    .Z(\u_multiplier/_0400_ ));
 AOI22_X1 \u_multiplier/_0782_  (.A1(\u_multiplier/_0722_ ),
    .A2(\u_multiplier/_0392_ ),
    .B1(\u_multiplier/_0398_ ),
    .B2(\u_multiplier/_0400_ ),
    .ZN(\u_multiplier/_0401_ ));
 OAI22_X1 \u_multiplier/_0783_  (.A1(\u_multiplier/_0721_ ),
    .A2(\u_multiplier/_0723_ ),
    .B1(\u_multiplier/_0397_ ),
    .B2(\u_multiplier/_0399_ ),
    .ZN(\u_multiplier/_0402_ ));
 XOR2_X2 \u_multiplier/_0784_  (.A(\u_multiplier/ky [3]),
    .B(\u_multiplier/LODy/z [3]),
    .Z(\u_multiplier/_0403_ ));
 XNOR2_X2 \u_multiplier/_0785_  (.A(\u_multiplier/kx [3]),
    .B(\u_multiplier/LODx/z [3]),
    .ZN(\u_multiplier/_0404_ ));
 XOR2_X2 \u_multiplier/_0786_  (.A(\u_multiplier/kx [3]),
    .B(\u_multiplier/LODx/z [3]),
    .Z(\u_multiplier/_0405_ ));
 AOI22_X1 \u_multiplier/_0787_  (.A1(\u_multiplier/_0397_ ),
    .A2(\u_multiplier/_0399_ ),
    .B1(\u_multiplier/_0403_ ),
    .B2(\u_multiplier/_0404_ ),
    .ZN(\u_multiplier/_0406_ ));
 AOI222_X2 \u_multiplier/_0788_  (.A1(\u_multiplier/_0397_ ),
    .A2(\u_multiplier/_0399_ ),
    .B1(\u_multiplier/_0403_ ),
    .B2(\u_multiplier/_0404_ ),
    .C1(\u_multiplier/_0401_ ),
    .C2(\u_multiplier/_0396_ ),
    .ZN(\u_multiplier/_0407_ ));
 OAI21_X1 \u_multiplier/_0789_  (.A(\u_multiplier/_0406_ ),
    .B1(\u_multiplier/_0402_ ),
    .B2(\u_multiplier/_0395_ ),
    .ZN(\u_multiplier/_0408_ ));
 XOR2_X2 \u_multiplier/_0790_  (.A(\u_multiplier/ky [4]),
    .B(sram_rdata_reg[4]),
    .Z(\u_multiplier/_0409_ ));
 XNOR2_X2 \u_multiplier/_0791_  (.A(\u_multiplier/kx [4]),
    .B(data_in_reg[4]),
    .ZN(\u_multiplier/_0410_ ));
 XOR2_X2 \u_multiplier/_0792_  (.A(\u_multiplier/kx [4]),
    .B(data_in_reg[4]),
    .Z(\u_multiplier/_0411_ ));
 OAI22_X2 \u_multiplier/_0793_  (.A1(\u_multiplier/_0403_ ),
    .A2(\u_multiplier/_0404_ ),
    .B1(\u_multiplier/_0409_ ),
    .B2(\u_multiplier/_0410_ ),
    .ZN(\u_multiplier/_0412_ ));
 INV_X1 \u_multiplier/_0794_  (.A(\u_multiplier/_0412_ ),
    .ZN(\u_multiplier/_0413_ ));
 XOR2_X2 \u_multiplier/_0795_  (.A(\u_multiplier/kx [5]),
    .B(data_in_reg[5]),
    .Z(\u_multiplier/_0414_ ));
 XNOR2_X2 \u_multiplier/_0796_  (.A(\u_multiplier/ky [5]),
    .B(sram_rdata_reg[5]),
    .ZN(\u_multiplier/_0415_ ));
 XOR2_X2 \u_multiplier/_0797_  (.A(\u_multiplier/ky [5]),
    .B(sram_rdata_reg[5]),
    .Z(\u_multiplier/_0416_ ));
 NOR2_X1 \u_multiplier/_0798_  (.A1(\u_multiplier/_0414_ ),
    .A2(\u_multiplier/_0415_ ),
    .ZN(\u_multiplier/_0417_ ));
 NAND2_X1 \u_multiplier/_0799_  (.A1(\u_multiplier/_0409_ ),
    .A2(\u_multiplier/_0410_ ),
    .ZN(\u_multiplier/_0418_ ));
 AOI221_X2 \u_multiplier/_0800_  (.A(\u_multiplier/_0417_ ),
    .B1(\u_multiplier/_0410_ ),
    .B2(\u_multiplier/_0409_ ),
    .C1(\u_multiplier/_0408_ ),
    .C2(\u_multiplier/_0413_ ),
    .ZN(\u_multiplier/_0419_ ));
 OAI221_X2 \u_multiplier/_0801_  (.A(\u_multiplier/_0418_ ),
    .B1(\u_multiplier/_0415_ ),
    .B2(\u_multiplier/_0414_ ),
    .C1(\u_multiplier/_0407_ ),
    .C2(\u_multiplier/_0412_ ),
    .ZN(\u_multiplier/_0420_ ));
 NAND2_X1 \u_multiplier/_0802_  (.A1(\u_multiplier/_0414_ ),
    .A2(\u_multiplier/_0415_ ),
    .ZN(\u_multiplier/_0421_ ));
 AOI22_X4 \u_multiplier/_0803_  (.A1(\u_multiplier/_0716_ ),
    .A2(\u_multiplier/_0719_ ),
    .B1(\u_multiplier/_0414_ ),
    .B2(\u_multiplier/_0415_ ),
    .ZN(\u_multiplier/_0422_ ));
 OAI21_X2 \u_multiplier/_0804_  (.A(\u_multiplier/_0421_ ),
    .B1(\u_multiplier/_0718_ ),
    .B2(\u_multiplier/_0717_ ),
    .ZN(\u_multiplier/_0423_ ));
 AOI21_X4 \u_multiplier/_0805_  (.A(\u_multiplier/_0720_ ),
    .B1(\u_multiplier/_0420_ ),
    .B2(\u_multiplier/_0422_ ),
    .ZN(\u_multiplier/_0424_ ));
 OAI22_X4 \u_multiplier/_0806_  (.A1(\u_multiplier/_0716_ ),
    .A2(\u_multiplier/_0719_ ),
    .B1(\u_multiplier/_0419_ ),
    .B2(\u_multiplier/_0423_ ),
    .ZN(\u_multiplier/_0425_ ));
 MUX2_X1 \u_multiplier/_0807_  (.A(\u_multiplier/_0715_ ),
    .B(\u_multiplier/_0394_ ),
    .S(\u_multiplier/_0424_ ),
    .Z(\u_multiplier/_0345_ ));
 MUX2_X2 \u_multiplier/_0808_  (.A(\u_multiplier/_0721_ ),
    .B(\u_multiplier/_0392_ ),
    .S(\u_multiplier/_0424_ ),
    .Z(\u_multiplier/_0346_ ));
 MUX2_X2 \u_multiplier/_0809_  (.A(\u_multiplier/_0397_ ),
    .B(\u_multiplier/_0400_ ),
    .S(\u_multiplier/_0424_ ),
    .Z(\u_multiplier/_0347_ ));
 MUX2_X2 \u_multiplier/_0810_  (.A(\u_multiplier/_0403_ ),
    .B(\u_multiplier/_0405_ ),
    .S(\u_multiplier/_0424_ ),
    .Z(\u_multiplier/_0348_ ));
 MUX2_X2 \u_multiplier/_0811_  (.A(\u_multiplier/_0409_ ),
    .B(\u_multiplier/_0411_ ),
    .S(\u_multiplier/_0424_ ),
    .Z(\u_multiplier/_0349_ ));
 MUX2_X2 \u_multiplier/_0812_  (.A(\u_multiplier/_0414_ ),
    .B(\u_multiplier/_0416_ ),
    .S(\u_multiplier/_0425_ ),
    .Z(\u_multiplier/_0350_ ));
 NAND2_X2 \u_multiplier/_0813_  (.A1(\u_multiplier/_0717_ ),
    .A2(\u_multiplier/_0719_ ),
    .ZN(\u_multiplier/_0351_ ));
 MUX2_X2 \u_multiplier/_0814_  (.A(\u_multiplier/_0714_ ),
    .B(\u_multiplier/_0393_ ),
    .S(\u_multiplier/_0425_ ),
    .Z(\u_multiplier/_0426_ ));
 NOR3_X1 \u_multiplier/_0815_  (.A1(\u_multiplier/K [0]),
    .A2(\u_multiplier/K [1]),
    .A3(\u_multiplier/_0426_ ),
    .ZN(\u_multiplier/_0427_ ));
 NOR4_X2 \u_multiplier/_0816_  (.A1(\u_multiplier/K [0]),
    .A2(\u_multiplier/K [1]),
    .A3(\u_multiplier/K [2]),
    .A4(\u_multiplier/_0426_ ),
    .ZN(\u_multiplier/_0428_ ));
 NOR2_X1 \u_multiplier/_0817_  (.A1(\u_multiplier/code_x [0]),
    .A2(\u_multiplier/_0714_ ),
    .ZN(\u_multiplier/_0429_ ));
 NOR3_X1 \u_multiplier/_0818_  (.A1(\u_multiplier/code_x [0]),
    .A2(\u_multiplier/code_x [1]),
    .A3(\u_multiplier/_0714_ ),
    .ZN(\u_multiplier/_0430_ ));
 AND2_X1 \u_multiplier/_0819_  (.A1(\u_multiplier/_0708_ ),
    .A2(\u_multiplier/_0430_ ),
    .ZN(\u_multiplier/_0431_ ));
 NOR2_X1 \u_multiplier/_0820_  (.A1(\u_multiplier/code_y [0]),
    .A2(\u_multiplier/_0393_ ),
    .ZN(\u_multiplier/_0432_ ));
 OR3_X1 \u_multiplier/_0821_  (.A1(\u_multiplier/code_y [0]),
    .A2(\u_multiplier/code_y [1]),
    .A3(\u_multiplier/_0393_ ),
    .ZN(\u_multiplier/_0433_ ));
 NOR2_X1 \u_multiplier/_0822_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_0433_ ),
    .ZN(\u_multiplier/_0434_ ));
 NAND2_X1 \u_multiplier/_0823_  (.A1(\u_multiplier/_0431_ ),
    .A2(\u_multiplier/_0434_ ),
    .ZN(\u_multiplier/_0435_ ));
 XOR2_X1 \u_multiplier/_0824_  (.A(\u_multiplier/_0431_ ),
    .B(\u_multiplier/_0434_ ),
    .Z(\u_multiplier/_0436_ ));
 OR3_X1 \u_multiplier/_0825_  (.A1(\u_multiplier/dec_out [0]),
    .A2(\u_multiplier/_0428_ ),
    .A3(\u_multiplier/_0436_ ),
    .ZN(\u_multiplier/_0437_ ));
 OAI21_X1 \u_multiplier/_0826_  (.A(\u_multiplier/_0436_ ),
    .B1(\u_multiplier/_0428_ ),
    .B2(\u_multiplier/dec_out [0]),
    .ZN(\u_multiplier/_0438_ ));
 NOR2_X4 \u_multiplier/_0827_  (.A1(\u_multiplier/zero_y ),
    .A2(\u_multiplier/zero_x ),
    .ZN(\u_multiplier/_0439_ ));
 OR2_X2 \u_multiplier/_0828_  (.A1(\u_multiplier/zero_y ),
    .A2(\u_multiplier/zero_x ),
    .ZN(\u_multiplier/_0440_ ));
 AND3_X1 \u_multiplier/_0829_  (.A1(\u_multiplier/_0437_ ),
    .A2(\u_multiplier/_0438_ ),
    .A3(\u_multiplier/_0439_ ),
    .ZN(product[0]));
 NAND2_X1 \u_multiplier/_0830_  (.A1(\u_multiplier/_0435_ ),
    .A2(\u_multiplier/_0438_ ),
    .ZN(\u_multiplier/_0441_ ));
 AOI211_X2 \u_multiplier/_0831_  (.A(\u_multiplier/_0720_ ),
    .B(\u_multiplier/_0722_ ),
    .C1(\u_multiplier/_0420_ ),
    .C2(\u_multiplier/_0422_ ),
    .ZN(\u_multiplier/_0442_ ));
 AOI211_X2 \u_multiplier/_0832_  (.A(\u_multiplier/K [0]),
    .B(\u_multiplier/_0442_ ),
    .C1(\u_multiplier/_0425_ ),
    .C2(\u_multiplier/_0392_ ),
    .ZN(\u_multiplier/_0443_ ));
 AOI21_X1 \u_multiplier/_0833_  (.A(\u_multiplier/_0443_ ),
    .B1(\u_multiplier/_0426_ ),
    .B2(\u_multiplier/K [0]),
    .ZN(\u_multiplier/_0444_ ));
 AOI211_X2 \u_multiplier/_0834_  (.A(\u_multiplier/K [1]),
    .B(\u_multiplier/_0443_ ),
    .C1(\u_multiplier/_0426_ ),
    .C2(\u_multiplier/K [0]),
    .ZN(\u_multiplier/_0445_ ));
 AOI21_X4 \u_multiplier/_0835_  (.A(\u_multiplier/dec_out [1]),
    .B1(\u_multiplier/_0445_ ),
    .B2(\u_multiplier/_0711_ ),
    .ZN(\u_multiplier/_0446_ ));
 MUX2_X1 \u_multiplier/_0836_  (.A(\u_multiplier/_0722_ ),
    .B(\u_multiplier/_0714_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_0447_ ));
 OR2_X1 \u_multiplier/_0837_  (.A1(\u_multiplier/code_x [1]),
    .A2(\u_multiplier/_0447_ ),
    .ZN(\u_multiplier/_0448_ ));
 MUX2_X1 \u_multiplier/_0838_  (.A(\u_multiplier/_0723_ ),
    .B(\u_multiplier/_0393_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_0449_ ));
 OR2_X1 \u_multiplier/_0839_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_0449_ ),
    .ZN(\u_multiplier/_0450_ ));
 OAI22_X1 \u_multiplier/_0840_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_0448_ ),
    .B1(\u_multiplier/_0450_ ),
    .B2(\u_multiplier/code_y [2]),
    .ZN(\u_multiplier/_0451_ ));
 OR4_X1 \u_multiplier/_0841_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/code_x [2]),
    .A3(\u_multiplier/_0448_ ),
    .A4(\u_multiplier/_0450_ ),
    .ZN(\u_multiplier/_0452_ ));
 NAND2_X1 \u_multiplier/_0842_  (.A1(\u_multiplier/_0451_ ),
    .A2(\u_multiplier/_0452_ ),
    .ZN(\u_multiplier/_0453_ ));
 XOR2_X2 \u_multiplier/_0843_  (.A(\u_multiplier/_0446_ ),
    .B(\u_multiplier/_0453_ ),
    .Z(\u_multiplier/_0454_ ));
 NAND2_X2 \u_multiplier/_0844_  (.A1(\u_multiplier/_0441_ ),
    .A2(\u_multiplier/_0454_ ),
    .ZN(\u_multiplier/_0455_ ));
 OAI21_X1 \u_multiplier/_0845_  (.A(\u_multiplier/_0439_ ),
    .B1(\u_multiplier/_0441_ ),
    .B2(\u_multiplier/_0454_ ),
    .ZN(\u_multiplier/_0456_ ));
 AOI21_X1 \u_multiplier/_0846_  (.A(\u_multiplier/_0456_ ),
    .B1(\u_multiplier/_0454_ ),
    .B2(\u_multiplier/_0441_ ),
    .ZN(product[1]));
 OAI21_X2 \u_multiplier/_0847_  (.A(\u_multiplier/_0452_ ),
    .B1(\u_multiplier/_0453_ ),
    .B2(\u_multiplier/_0446_ ),
    .ZN(\u_multiplier/_0457_ ));
 AOI211_X2 \u_multiplier/_0848_  (.A(\u_multiplier/_0720_ ),
    .B(\u_multiplier/_0398_ ),
    .C1(\u_multiplier/_0420_ ),
    .C2(\u_multiplier/_0422_ ),
    .ZN(\u_multiplier/_0458_ ));
 MUX2_X1 \u_multiplier/_0849_  (.A(\u_multiplier/_0397_ ),
    .B(\u_multiplier/_0400_ ),
    .S(\u_multiplier/_0425_ ),
    .Z(\u_multiplier/_0459_ ));
 AOI211_X2 \u_multiplier/_0850_  (.A(\u_multiplier/_0709_ ),
    .B(\u_multiplier/_0442_ ),
    .C1(\u_multiplier/_0425_ ),
    .C2(\u_multiplier/_0392_ ),
    .ZN(\u_multiplier/_0460_ ));
 AOI211_X2 \u_multiplier/_0851_  (.A(\u_multiplier/K [0]),
    .B(\u_multiplier/_0458_ ),
    .C1(\u_multiplier/_0425_ ),
    .C2(\u_multiplier/_0400_ ),
    .ZN(\u_multiplier/_0461_ ));
 OAI21_X1 \u_multiplier/_0852_  (.A(\u_multiplier/K [1]),
    .B1(\u_multiplier/_0426_ ),
    .B2(\u_multiplier/K [0]),
    .ZN(\u_multiplier/_0462_ ));
 OAI21_X1 \u_multiplier/_0853_  (.A(\u_multiplier/_0710_ ),
    .B1(\u_multiplier/_0460_ ),
    .B2(\u_multiplier/_0461_ ),
    .ZN(\u_multiplier/_0463_ ));
 AND3_X1 \u_multiplier/_0854_  (.A1(\u_multiplier/_0711_ ),
    .A2(\u_multiplier/_0462_ ),
    .A3(\u_multiplier/_0463_ ),
    .ZN(\u_multiplier/_0464_ ));
 MUX2_X1 \u_multiplier/_0855_  (.A(\u_multiplier/_0398_ ),
    .B(\u_multiplier/_0722_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_0465_ ));
 NOR2_X1 \u_multiplier/_0856_  (.A1(\u_multiplier/code_x [1]),
    .A2(\u_multiplier/_0465_ ),
    .ZN(\u_multiplier/_0466_ ));
 AOI21_X2 \u_multiplier/_0857_  (.A(\u_multiplier/_0466_ ),
    .B1(\u_multiplier/_0429_ ),
    .B2(\u_multiplier/code_x [1]),
    .ZN(\u_multiplier/_0467_ ));
 NOR2_X1 \u_multiplier/_0858_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_0467_ ),
    .ZN(\u_multiplier/_0468_ ));
 MUX2_X1 \u_multiplier/_0859_  (.A(\u_multiplier/_0399_ ),
    .B(\u_multiplier/_0723_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_0469_ ));
 NOR2_X1 \u_multiplier/_0860_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_0469_ ),
    .ZN(\u_multiplier/_0470_ ));
 AOI21_X2 \u_multiplier/_0861_  (.A(\u_multiplier/_0470_ ),
    .B1(\u_multiplier/_0432_ ),
    .B2(\u_multiplier/code_y [1]),
    .ZN(\u_multiplier/_0471_ ));
 NOR2_X1 \u_multiplier/_0862_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_0471_ ),
    .ZN(\u_multiplier/_0472_ ));
 NAND2_X1 \u_multiplier/_0863_  (.A1(\u_multiplier/_0468_ ),
    .A2(\u_multiplier/_0472_ ),
    .ZN(\u_multiplier/_0473_ ));
 XOR2_X2 \u_multiplier/_0864_  (.A(\u_multiplier/_0468_ ),
    .B(\u_multiplier/_0472_ ),
    .Z(\u_multiplier/_0474_ ));
 OAI21_X2 \u_multiplier/_0865_  (.A(\u_multiplier/_0474_ ),
    .B1(\u_multiplier/_0464_ ),
    .B2(\u_multiplier/dec_out [2]),
    .ZN(\u_multiplier/_0475_ ));
 OR3_X1 \u_multiplier/_0866_  (.A1(\u_multiplier/dec_out [2]),
    .A2(\u_multiplier/_0464_ ),
    .A3(\u_multiplier/_0474_ ),
    .ZN(\u_multiplier/_0476_ ));
 AND2_X1 \u_multiplier/_0867_  (.A1(\u_multiplier/_0475_ ),
    .A2(\u_multiplier/_0476_ ),
    .ZN(\u_multiplier/_0477_ ));
 NAND3_X1 \u_multiplier/_0868_  (.A1(\u_multiplier/_0457_ ),
    .A2(\u_multiplier/_0475_ ),
    .A3(\u_multiplier/_0476_ ),
    .ZN(\u_multiplier/_0478_ ));
 AOI21_X1 \u_multiplier/_0869_  (.A(\u_multiplier/_0457_ ),
    .B1(\u_multiplier/_0475_ ),
    .B2(\u_multiplier/_0476_ ),
    .ZN(\u_multiplier/_0479_ ));
 XNOR2_X1 \u_multiplier/_0870_  (.A(\u_multiplier/_0457_ ),
    .B(\u_multiplier/_0477_ ),
    .ZN(\u_multiplier/_0480_ ));
 OAI21_X1 \u_multiplier/_0871_  (.A(\u_multiplier/_0439_ ),
    .B1(\u_multiplier/_0455_ ),
    .B2(\u_multiplier/_0480_ ),
    .ZN(\u_multiplier/_0481_ ));
 AOI21_X2 \u_multiplier/_0872_  (.A(\u_multiplier/_0481_ ),
    .B1(\u_multiplier/_0480_ ),
    .B2(\u_multiplier/_0455_ ),
    .ZN(product[2]));
 OAI21_X2 \u_multiplier/_0873_  (.A(\u_multiplier/_0478_ ),
    .B1(\u_multiplier/_0479_ ),
    .B2(\u_multiplier/_0455_ ),
    .ZN(\u_multiplier/_0482_ ));
 NAND2_X1 \u_multiplier/_0874_  (.A1(\u_multiplier/_0473_ ),
    .A2(\u_multiplier/_0475_ ),
    .ZN(\u_multiplier/_0483_ ));
 MUX2_X1 \u_multiplier/_0875_  (.A(\u_multiplier/_0403_ ),
    .B(\u_multiplier/_0405_ ),
    .S(\u_multiplier/_0425_ ),
    .Z(\u_multiplier/_0484_ ));
 MUX2_X1 \u_multiplier/_0876_  (.A(\u_multiplier/_0459_ ),
    .B(\u_multiplier/_0484_ ),
    .S(\u_multiplier/_0709_ ),
    .Z(\u_multiplier/_0485_ ));
 MUX2_X1 \u_multiplier/_0877_  (.A(\u_multiplier/_0444_ ),
    .B(\u_multiplier/_0485_ ),
    .S(\u_multiplier/_0710_ ),
    .Z(\u_multiplier/_0486_ ));
 AOI21_X2 \u_multiplier/_0878_  (.A(\u_multiplier/dec_out [3]),
    .B1(\u_multiplier/_0486_ ),
    .B2(\u_multiplier/_0711_ ),
    .ZN(\u_multiplier/_0487_ ));
 MUX2_X1 \u_multiplier/_0879_  (.A(\u_multiplier/_0403_ ),
    .B(\u_multiplier/_0397_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_0488_ ));
 NAND2_X1 \u_multiplier/_0880_  (.A1(\u_multiplier/code_x [1]),
    .A2(\u_multiplier/_0447_ ),
    .ZN(\u_multiplier/_0489_ ));
 OAI21_X2 \u_multiplier/_0881_  (.A(\u_multiplier/_0489_ ),
    .B1(\u_multiplier/_0488_ ),
    .B2(\u_multiplier/code_x [1]),
    .ZN(\u_multiplier/_0490_ ));
 NOR2_X2 \u_multiplier/_0882_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_0490_ ),
    .ZN(\u_multiplier/_0491_ ));
 MUX2_X1 \u_multiplier/_0883_  (.A(\u_multiplier/_0404_ ),
    .B(\u_multiplier/_0399_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_0492_ ));
 MUX2_X1 \u_multiplier/_0884_  (.A(\u_multiplier/_0492_ ),
    .B(\u_multiplier/_0449_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_0493_ ));
 NOR2_X2 \u_multiplier/_0885_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_0493_ ),
    .ZN(\u_multiplier/_0494_ ));
 XNOR2_X2 \u_multiplier/_0886_  (.A(\u_multiplier/_0491_ ),
    .B(\u_multiplier/_0494_ ),
    .ZN(\u_multiplier/_0495_ ));
 NOR2_X1 \u_multiplier/_0887_  (.A1(\u_multiplier/_0487_ ),
    .A2(\u_multiplier/_0495_ ),
    .ZN(\u_multiplier/_0496_ ));
 XOR2_X2 \u_multiplier/_0888_  (.A(\u_multiplier/_0487_ ),
    .B(\u_multiplier/_0495_ ),
    .Z(\u_multiplier/_0497_ ));
 AND2_X1 \u_multiplier/_0889_  (.A1(\u_multiplier/_0483_ ),
    .A2(\u_multiplier/_0497_ ),
    .ZN(\u_multiplier/_0498_ ));
 XOR2_X2 \u_multiplier/_0890_  (.A(\u_multiplier/_0483_ ),
    .B(\u_multiplier/_0497_ ),
    .Z(\u_multiplier/_0499_ ));
 NAND2_X1 \u_multiplier/_0891_  (.A1(\u_multiplier/_0482_ ),
    .A2(\u_multiplier/_0499_ ),
    .ZN(\u_multiplier/_0500_ ));
 OR2_X1 \u_multiplier/_0892_  (.A1(\u_multiplier/_0482_ ),
    .A2(\u_multiplier/_0499_ ),
    .ZN(\u_multiplier/_0501_ ));
 NAND3_X1 \u_multiplier/_0893_  (.A1(\u_multiplier/_0439_ ),
    .A2(\u_multiplier/_0500_ ),
    .A3(\u_multiplier/_0501_ ),
    .ZN(\u_multiplier/_0502_ ));
 INV_X1 \u_multiplier/_0894_  (.A(\u_multiplier/_0502_ ),
    .ZN(product[3]));
 AOI21_X2 \u_multiplier/_0895_  (.A(\u_multiplier/_0498_ ),
    .B1(\u_multiplier/_0499_ ),
    .B2(\u_multiplier/_0482_ ),
    .ZN(\u_multiplier/_0503_ ));
 AOI21_X2 \u_multiplier/_0896_  (.A(\u_multiplier/_0496_ ),
    .B1(\u_multiplier/_0494_ ),
    .B2(\u_multiplier/_0491_ ),
    .ZN(\u_multiplier/_0504_ ));
 MUX2_X1 \u_multiplier/_0897_  (.A(\u_multiplier/_0409_ ),
    .B(\u_multiplier/_0411_ ),
    .S(\u_multiplier/_0425_ ),
    .Z(\u_multiplier/_0505_ ));
 MUX2_X1 \u_multiplier/_0898_  (.A(\u_multiplier/_0484_ ),
    .B(\u_multiplier/_0505_ ),
    .S(\u_multiplier/_0709_ ),
    .Z(\u_multiplier/_0506_ ));
 NAND2_X1 \u_multiplier/_0899_  (.A1(\u_multiplier/_0710_ ),
    .A2(\u_multiplier/_0506_ ),
    .ZN(\u_multiplier/_0507_ ));
 OR3_X1 \u_multiplier/_0900_  (.A1(\u_multiplier/_0710_ ),
    .A2(\u_multiplier/_0460_ ),
    .A3(\u_multiplier/_0461_ ),
    .ZN(\u_multiplier/_0508_ ));
 AND2_X1 \u_multiplier/_0901_  (.A1(\u_multiplier/_0507_ ),
    .A2(\u_multiplier/_0508_ ),
    .ZN(\u_multiplier/_0509_ ));
 AOI21_X1 \u_multiplier/_0902_  (.A(\u_multiplier/dec_out [4]),
    .B1(\u_multiplier/_0427_ ),
    .B2(\u_multiplier/K [2]),
    .ZN(\u_multiplier/_0510_ ));
 OAI21_X2 \u_multiplier/_0903_  (.A(\u_multiplier/_0510_ ),
    .B1(\u_multiplier/_0509_ ),
    .B2(\u_multiplier/K [2]),
    .ZN(\u_multiplier/_0511_ ));
 MUX2_X1 \u_multiplier/_0904_  (.A(\u_multiplier/_0409_ ),
    .B(\u_multiplier/_0403_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_0512_ ));
 NOR2_X1 \u_multiplier/_0905_  (.A1(\u_multiplier/code_x [1]),
    .A2(\u_multiplier/_0512_ ),
    .ZN(\u_multiplier/_0513_ ));
 AOI21_X2 \u_multiplier/_0906_  (.A(\u_multiplier/_0513_ ),
    .B1(\u_multiplier/_0465_ ),
    .B2(\u_multiplier/code_x [1]),
    .ZN(\u_multiplier/_0514_ ));
 MUX2_X1 \u_multiplier/_0907_  (.A(\u_multiplier/_0430_ ),
    .B(\u_multiplier/_0514_ ),
    .S(\u_multiplier/_0708_ ),
    .Z(\u_multiplier/_0515_ ));
 MUX2_X1 \u_multiplier/_0908_  (.A(\u_multiplier/_0411_ ),
    .B(\u_multiplier/_0405_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_0516_ ));
 NOR2_X1 \u_multiplier/_0909_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_0516_ ),
    .ZN(\u_multiplier/_0517_ ));
 AOI21_X2 \u_multiplier/_0910_  (.A(\u_multiplier/_0517_ ),
    .B1(\u_multiplier/_0469_ ),
    .B2(\u_multiplier/code_y [1]),
    .ZN(\u_multiplier/_0518_ ));
 NOR2_X1 \u_multiplier/_0911_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_0518_ ),
    .ZN(\u_multiplier/_0519_ ));
 AOI21_X2 \u_multiplier/_0912_  (.A(\u_multiplier/_0519_ ),
    .B1(\u_multiplier/_0433_ ),
    .B2(\u_multiplier/code_y [2]),
    .ZN(\u_multiplier/_0520_ ));
 NAND2_X1 \u_multiplier/_0913_  (.A1(\u_multiplier/_0515_ ),
    .A2(\u_multiplier/_0520_ ),
    .ZN(\u_multiplier/_0521_ ));
 XOR2_X2 \u_multiplier/_0914_  (.A(\u_multiplier/_0515_ ),
    .B(\u_multiplier/_0520_ ),
    .Z(\u_multiplier/_0522_ ));
 NAND2_X1 \u_multiplier/_0915_  (.A1(\u_multiplier/_0511_ ),
    .A2(\u_multiplier/_0522_ ),
    .ZN(\u_multiplier/_0523_ ));
 XNOR2_X2 \u_multiplier/_0916_  (.A(\u_multiplier/_0511_ ),
    .B(\u_multiplier/_0522_ ),
    .ZN(\u_multiplier/_0524_ ));
 OR2_X1 \u_multiplier/_0917_  (.A1(\u_multiplier/_0504_ ),
    .A2(\u_multiplier/_0524_ ),
    .ZN(\u_multiplier/_0525_ ));
 XNOR2_X2 \u_multiplier/_0918_  (.A(\u_multiplier/_0504_ ),
    .B(\u_multiplier/_0524_ ),
    .ZN(\u_multiplier/_0526_ ));
 AOI21_X1 \u_multiplier/_0919_  (.A(\u_multiplier/_0440_ ),
    .B1(\u_multiplier/_0503_ ),
    .B2(\u_multiplier/_0526_ ),
    .ZN(\u_multiplier/_0527_ ));
 OAI21_X1 \u_multiplier/_0920_  (.A(\u_multiplier/_0527_ ),
    .B1(\u_multiplier/_0526_ ),
    .B2(\u_multiplier/_0503_ ),
    .ZN(\u_multiplier/_0528_ ));
 INV_X1 \u_multiplier/_0921_  (.A(\u_multiplier/_0528_ ),
    .ZN(product[4]));
 OAI21_X2 \u_multiplier/_0922_  (.A(\u_multiplier/_0525_ ),
    .B1(\u_multiplier/_0526_ ),
    .B2(\u_multiplier/_0503_ ),
    .ZN(\u_multiplier/_0529_ ));
 MUX2_X1 \u_multiplier/_0923_  (.A(\u_multiplier/_0414_ ),
    .B(\u_multiplier/_0416_ ),
    .S(\u_multiplier/_0424_ ),
    .Z(\u_multiplier/_0530_ ));
 MUX2_X1 \u_multiplier/_0924_  (.A(\u_multiplier/_0505_ ),
    .B(\u_multiplier/_0530_ ),
    .S(\u_multiplier/_0709_ ),
    .Z(\u_multiplier/_0531_ ));
 MUX2_X1 \u_multiplier/_0925_  (.A(\u_multiplier/_0485_ ),
    .B(\u_multiplier/_0531_ ),
    .S(\u_multiplier/_0710_ ),
    .Z(\u_multiplier/_0532_ ));
 INV_X1 \u_multiplier/_0926_  (.A(\u_multiplier/_0532_ ),
    .ZN(\u_multiplier/_0533_ ));
 AOI21_X1 \u_multiplier/_0927_  (.A(\u_multiplier/dec_out [5]),
    .B1(\u_multiplier/_0445_ ),
    .B2(\u_multiplier/K [2]),
    .ZN(\u_multiplier/_0534_ ));
 OAI21_X2 \u_multiplier/_0928_  (.A(\u_multiplier/_0534_ ),
    .B1(\u_multiplier/_0533_ ),
    .B2(\u_multiplier/K [2]),
    .ZN(\u_multiplier/_0535_ ));
 INV_X1 \u_multiplier/_0929_  (.A(\u_multiplier/_0535_ ),
    .ZN(\u_multiplier/_0536_ ));
 MUX2_X1 \u_multiplier/_0930_  (.A(\u_multiplier/_0416_ ),
    .B(\u_multiplier/_0409_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_0537_ ));
 MUX2_X1 \u_multiplier/_0931_  (.A(\u_multiplier/_0537_ ),
    .B(\u_multiplier/_0488_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_0538_ ));
 NOR2_X1 \u_multiplier/_0932_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_0538_ ),
    .ZN(\u_multiplier/_0539_ ));
 AOI21_X2 \u_multiplier/_0933_  (.A(\u_multiplier/_0539_ ),
    .B1(\u_multiplier/_0448_ ),
    .B2(\u_multiplier/code_x [2]),
    .ZN(\u_multiplier/_0540_ ));
 MUX2_X1 \u_multiplier/_0934_  (.A(\u_multiplier/_0414_ ),
    .B(\u_multiplier/_0411_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_0541_ ));
 NOR2_X1 \u_multiplier/_0935_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_0541_ ),
    .ZN(\u_multiplier/_0542_ ));
 AOI21_X2 \u_multiplier/_0936_  (.A(\u_multiplier/_0542_ ),
    .B1(\u_multiplier/_0492_ ),
    .B2(\u_multiplier/code_y [1]),
    .ZN(\u_multiplier/_0543_ ));
 NOR2_X1 \u_multiplier/_0937_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_0543_ ),
    .ZN(\u_multiplier/_0544_ ));
 AOI21_X2 \u_multiplier/_0938_  (.A(\u_multiplier/_0544_ ),
    .B1(\u_multiplier/_0450_ ),
    .B2(\u_multiplier/code_y [2]),
    .ZN(\u_multiplier/_0545_ ));
 XNOR2_X2 \u_multiplier/_0939_  (.A(\u_multiplier/_0540_ ),
    .B(\u_multiplier/_0545_ ),
    .ZN(\u_multiplier/_0546_ ));
 NOR2_X1 \u_multiplier/_0940_  (.A1(\u_multiplier/_0536_ ),
    .A2(\u_multiplier/_0546_ ),
    .ZN(\u_multiplier/_0547_ ));
 XOR2_X2 \u_multiplier/_0941_  (.A(\u_multiplier/_0535_ ),
    .B(\u_multiplier/_0546_ ),
    .Z(\u_multiplier/_0548_ ));
 AOI21_X2 \u_multiplier/_0942_  (.A(\u_multiplier/_0548_ ),
    .B1(\u_multiplier/_0523_ ),
    .B2(\u_multiplier/_0521_ ),
    .ZN(\u_multiplier/_0549_ ));
 AND3_X1 \u_multiplier/_0943_  (.A1(\u_multiplier/_0521_ ),
    .A2(\u_multiplier/_0523_ ),
    .A3(\u_multiplier/_0548_ ),
    .ZN(\u_multiplier/_0550_ ));
 NOR2_X2 \u_multiplier/_0944_  (.A1(\u_multiplier/_0549_ ),
    .A2(\u_multiplier/_0550_ ),
    .ZN(\u_multiplier/_0551_ ));
 OAI21_X1 \u_multiplier/_0945_  (.A(\u_multiplier/_0439_ ),
    .B1(\u_multiplier/_0529_ ),
    .B2(\u_multiplier/_0551_ ),
    .ZN(\u_multiplier/_0552_ ));
 AOI21_X1 \u_multiplier/_0946_  (.A(\u_multiplier/_0552_ ),
    .B1(\u_multiplier/_0551_ ),
    .B2(\u_multiplier/_0529_ ),
    .ZN(product[5]));
 AOI21_X2 \u_multiplier/_0947_  (.A(\u_multiplier/_0549_ ),
    .B1(\u_multiplier/_0551_ ),
    .B2(\u_multiplier/_0529_ ),
    .ZN(\u_multiplier/_0553_ ));
 AOI21_X2 \u_multiplier/_0948_  (.A(\u_multiplier/_0547_ ),
    .B1(\u_multiplier/_0545_ ),
    .B2(\u_multiplier/_0540_ ),
    .ZN(\u_multiplier/_0554_ ));
 NOR2_X1 \u_multiplier/_0949_  (.A1(\u_multiplier/_0717_ ),
    .A2(\u_multiplier/_0719_ ),
    .ZN(\u_multiplier/_0555_ ));
 MUX2_X1 \u_multiplier/_0950_  (.A(\u_multiplier/_0530_ ),
    .B(\u_multiplier/_0555_ ),
    .S(\u_multiplier/_0709_ ),
    .Z(\u_multiplier/_0556_ ));
 MUX2_X1 \u_multiplier/_0951_  (.A(\u_multiplier/_0506_ ),
    .B(\u_multiplier/_0556_ ),
    .S(\u_multiplier/_0710_ ),
    .Z(\u_multiplier/_0557_ ));
 AND3_X1 \u_multiplier/_0952_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/_0462_ ),
    .A3(\u_multiplier/_0463_ ),
    .ZN(\u_multiplier/_0558_ ));
 AOI211_X2 \u_multiplier/_0953_  (.A(\u_multiplier/dec_out [6]),
    .B(\u_multiplier/_0558_ ),
    .C1(\u_multiplier/_0557_ ),
    .C2(\u_multiplier/_0711_ ),
    .ZN(\u_multiplier/_0559_ ));
 MUX2_X1 \u_multiplier/_0954_  (.A(\u_multiplier/_0718_ ),
    .B(\u_multiplier/_0416_ ),
    .S(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_0560_ ));
 MUX2_X1 \u_multiplier/_0955_  (.A(\u_multiplier/_0560_ ),
    .B(\u_multiplier/_0512_ ),
    .S(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_0561_ ));
 NOR2_X1 \u_multiplier/_0956_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_0561_ ),
    .ZN(\u_multiplier/_0562_ ));
 AOI21_X1 \u_multiplier/_0957_  (.A(\u_multiplier/_0562_ ),
    .B1(\u_multiplier/_0467_ ),
    .B2(\u_multiplier/code_x [2]),
    .ZN(\u_multiplier/_0563_ ));
 MUX2_X1 \u_multiplier/_0958_  (.A(\u_multiplier/_0716_ ),
    .B(\u_multiplier/_0414_ ),
    .S(\u_multiplier/code_y [0]),
    .Z(\u_multiplier/_0564_ ));
 MUX2_X1 \u_multiplier/_0959_  (.A(\u_multiplier/_0564_ ),
    .B(\u_multiplier/_0516_ ),
    .S(\u_multiplier/code_y [1]),
    .Z(\u_multiplier/_0565_ ));
 NAND2_X1 \u_multiplier/_0960_  (.A1(\u_multiplier/_0707_ ),
    .A2(\u_multiplier/_0565_ ),
    .ZN(\u_multiplier/_0566_ ));
 OAI21_X1 \u_multiplier/_0961_  (.A(\u_multiplier/_0566_ ),
    .B1(\u_multiplier/_0471_ ),
    .B2(\u_multiplier/_0707_ ),
    .ZN(\u_multiplier/_0567_ ));
 NAND2_X1 \u_multiplier/_0962_  (.A1(\u_multiplier/_0563_ ),
    .A2(\u_multiplier/_0567_ ),
    .ZN(\u_multiplier/_0568_ ));
 XOR2_X1 \u_multiplier/_0963_  (.A(\u_multiplier/_0563_ ),
    .B(\u_multiplier/_0567_ ),
    .Z(\u_multiplier/_0569_ ));
 INV_X1 \u_multiplier/_0964_  (.A(\u_multiplier/_0569_ ),
    .ZN(\u_multiplier/_0570_ ));
 XNOR2_X2 \u_multiplier/_0965_  (.A(\u_multiplier/_0559_ ),
    .B(\u_multiplier/_0570_ ),
    .ZN(\u_multiplier/_0571_ ));
 OR2_X1 \u_multiplier/_0966_  (.A1(\u_multiplier/_0554_ ),
    .A2(\u_multiplier/_0571_ ),
    .ZN(\u_multiplier/_0572_ ));
 XNOR2_X2 \u_multiplier/_0967_  (.A(\u_multiplier/_0554_ ),
    .B(\u_multiplier/_0571_ ),
    .ZN(\u_multiplier/_0573_ ));
 OAI21_X1 \u_multiplier/_0968_  (.A(\u_multiplier/_0439_ ),
    .B1(\u_multiplier/_0553_ ),
    .B2(\u_multiplier/_0573_ ),
    .ZN(\u_multiplier/_0574_ ));
 AOI21_X1 \u_multiplier/_0969_  (.A(\u_multiplier/_0574_ ),
    .B1(\u_multiplier/_0573_ ),
    .B2(\u_multiplier/_0553_ ),
    .ZN(product[6]));
 OAI21_X2 \u_multiplier/_0970_  (.A(\u_multiplier/_0572_ ),
    .B1(\u_multiplier/_0573_ ),
    .B2(\u_multiplier/_0553_ ),
    .ZN(\u_multiplier/_0575_ ));
 OAI21_X1 \u_multiplier/_0971_  (.A(\u_multiplier/_0568_ ),
    .B1(\u_multiplier/_0570_ ),
    .B2(\u_multiplier/_0559_ ),
    .ZN(\u_multiplier/_0576_ ));
 NOR3_X1 \u_multiplier/_0972_  (.A1(\u_multiplier/_0709_ ),
    .A2(\u_multiplier/_0717_ ),
    .A3(\u_multiplier/_0719_ ),
    .ZN(\u_multiplier/_0577_ ));
 MUX2_X1 \u_multiplier/_0973_  (.A(\u_multiplier/_0531_ ),
    .B(\u_multiplier/_0577_ ),
    .S(\u_multiplier/_0710_ ),
    .Z(\u_multiplier/_0578_ ));
 AND2_X1 \u_multiplier/_0974_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/_0486_ ),
    .ZN(\u_multiplier/_0579_ ));
 AOI211_X2 \u_multiplier/_0975_  (.A(\u_multiplier/dec_out [7]),
    .B(\u_multiplier/_0579_ ),
    .C1(\u_multiplier/_0578_ ),
    .C2(\u_multiplier/_0711_ ),
    .ZN(\u_multiplier/_0580_ ));
 INV_X1 \u_multiplier/_0976_  (.A(\u_multiplier/_0580_ ),
    .ZN(\u_multiplier/_0581_ ));
 NAND2_X1 \u_multiplier/_0977_  (.A1(\u_multiplier/code_x [0]),
    .A2(\u_multiplier/_0718_ ),
    .ZN(\u_multiplier/_0582_ ));
 NAND2_X1 \u_multiplier/_0978_  (.A1(\u_multiplier/code_x [1]),
    .A2(\u_multiplier/_0537_ ),
    .ZN(\u_multiplier/_0583_ ));
 OAI21_X2 \u_multiplier/_0979_  (.A(\u_multiplier/_0583_ ),
    .B1(\u_multiplier/_0582_ ),
    .B2(\u_multiplier/code_x [1]),
    .ZN(\u_multiplier/_0584_ ));
 NAND2_X1 \u_multiplier/_0980_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_0490_ ),
    .ZN(\u_multiplier/_0585_ ));
 OAI21_X2 \u_multiplier/_0981_  (.A(\u_multiplier/_0585_ ),
    .B1(\u_multiplier/_0584_ ),
    .B2(\u_multiplier/code_x [2]),
    .ZN(\u_multiplier/_0586_ ));
 NAND2_X1 \u_multiplier/_0982_  (.A1(\u_multiplier/code_y [0]),
    .A2(\u_multiplier/_0716_ ),
    .ZN(\u_multiplier/_0587_ ));
 NAND2_X1 \u_multiplier/_0983_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_0541_ ),
    .ZN(\u_multiplier/_0588_ ));
 OAI21_X2 \u_multiplier/_0984_  (.A(\u_multiplier/_0588_ ),
    .B1(\u_multiplier/_0587_ ),
    .B2(\u_multiplier/code_y [1]),
    .ZN(\u_multiplier/_0589_ ));
 NAND2_X1 \u_multiplier/_0985_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_0493_ ),
    .ZN(\u_multiplier/_0590_ ));
 OAI21_X2 \u_multiplier/_0986_  (.A(\u_multiplier/_0590_ ),
    .B1(\u_multiplier/_0589_ ),
    .B2(\u_multiplier/code_y [2]),
    .ZN(\u_multiplier/_0591_ ));
 XOR2_X2 \u_multiplier/_0987_  (.A(\u_multiplier/_0586_ ),
    .B(\u_multiplier/_0591_ ),
    .Z(\u_multiplier/_0592_ ));
 NAND2_X1 \u_multiplier/_0988_  (.A1(\u_multiplier/_0581_ ),
    .A2(\u_multiplier/_0592_ ),
    .ZN(\u_multiplier/_0593_ ));
 XNOR2_X1 \u_multiplier/_0989_  (.A(\u_multiplier/_0580_ ),
    .B(\u_multiplier/_0592_ ),
    .ZN(\u_multiplier/_0594_ ));
 AND2_X1 \u_multiplier/_0990_  (.A1(\u_multiplier/_0576_ ),
    .A2(\u_multiplier/_0594_ ),
    .ZN(\u_multiplier/_0595_ ));
 XNOR2_X1 \u_multiplier/_0991_  (.A(\u_multiplier/_0576_ ),
    .B(\u_multiplier/_0594_ ),
    .ZN(\u_multiplier/_0596_ ));
 INV_X1 \u_multiplier/_0992_  (.A(\u_multiplier/_0596_ ),
    .ZN(\u_multiplier/_0597_ ));
 OAI21_X1 \u_multiplier/_0993_  (.A(\u_multiplier/_0439_ ),
    .B1(\u_multiplier/_0575_ ),
    .B2(\u_multiplier/_0597_ ),
    .ZN(\u_multiplier/_0598_ ));
 AOI21_X1 \u_multiplier/_0994_  (.A(\u_multiplier/_0598_ ),
    .B1(\u_multiplier/_0597_ ),
    .B2(\u_multiplier/_0575_ ),
    .ZN(product[7]));
 AOI21_X2 \u_multiplier/_0995_  (.A(\u_multiplier/_0595_ ),
    .B1(\u_multiplier/_0597_ ),
    .B2(\u_multiplier/_0575_ ),
    .ZN(\u_multiplier/_0599_ ));
 OAI21_X1 \u_multiplier/_0996_  (.A(\u_multiplier/_0593_ ),
    .B1(\u_multiplier/_0591_ ),
    .B2(\u_multiplier/_0586_ ),
    .ZN(\u_multiplier/_0600_ ));
 NAND2_X1 \u_multiplier/_0997_  (.A1(\u_multiplier/K [1]),
    .A2(\u_multiplier/_0556_ ),
    .ZN(\u_multiplier/_0601_ ));
 NOR2_X1 \u_multiplier/_0998_  (.A1(\u_multiplier/K [2]),
    .A2(\u_multiplier/_0601_ ),
    .ZN(\u_multiplier/_0602_ ));
 NOR2_X1 \u_multiplier/_0999_  (.A1(\u_multiplier/dec_out [8]),
    .A2(\u_multiplier/_0602_ ),
    .ZN(\u_multiplier/_0603_ ));
 OAI21_X2 \u_multiplier/_1000_  (.A(\u_multiplier/_0603_ ),
    .B1(\u_multiplier/_0509_ ),
    .B2(\u_multiplier/_0711_ ),
    .ZN(\u_multiplier/_0604_ ));
 AND2_X1 \u_multiplier/_1001_  (.A1(\u_multiplier/code_x [1]),
    .A2(\u_multiplier/_0560_ ),
    .ZN(\u_multiplier/_0605_ ));
 OR2_X1 \u_multiplier/_1002_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_0605_ ),
    .ZN(\u_multiplier/_0606_ ));
 OAI21_X2 \u_multiplier/_1003_  (.A(\u_multiplier/_0606_ ),
    .B1(\u_multiplier/_0514_ ),
    .B2(\u_multiplier/_0708_ ),
    .ZN(\u_multiplier/_0607_ ));
 AND2_X1 \u_multiplier/_1004_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/_0564_ ),
    .ZN(\u_multiplier/_0608_ ));
 OR2_X1 \u_multiplier/_1005_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_0608_ ),
    .ZN(\u_multiplier/_0609_ ));
 OAI21_X2 \u_multiplier/_1006_  (.A(\u_multiplier/_0609_ ),
    .B1(\u_multiplier/_0518_ ),
    .B2(\u_multiplier/_0707_ ),
    .ZN(\u_multiplier/_0610_ ));
 NOR2_X1 \u_multiplier/_1007_  (.A1(\u_multiplier/_0607_ ),
    .A2(\u_multiplier/_0610_ ),
    .ZN(\u_multiplier/_0611_ ));
 XOR2_X2 \u_multiplier/_1008_  (.A(\u_multiplier/_0607_ ),
    .B(\u_multiplier/_0610_ ),
    .Z(\u_multiplier/_0612_ ));
 XNOR2_X1 \u_multiplier/_1009_  (.A(\u_multiplier/_0604_ ),
    .B(\u_multiplier/_0612_ ),
    .ZN(\u_multiplier/_0613_ ));
 INV_X1 \u_multiplier/_1010_  (.A(\u_multiplier/_0613_ ),
    .ZN(\u_multiplier/_0614_ ));
 NAND2_X1 \u_multiplier/_1011_  (.A1(\u_multiplier/_0600_ ),
    .A2(\u_multiplier/_0614_ ),
    .ZN(\u_multiplier/_0615_ ));
 XNOR2_X1 \u_multiplier/_1012_  (.A(\u_multiplier/_0600_ ),
    .B(\u_multiplier/_0613_ ),
    .ZN(\u_multiplier/_0616_ ));
 INV_X1 \u_multiplier/_1013_  (.A(\u_multiplier/_0616_ ),
    .ZN(\u_multiplier/_0617_ ));
 OAI21_X1 \u_multiplier/_1014_  (.A(\u_multiplier/_0439_ ),
    .B1(\u_multiplier/_0599_ ),
    .B2(\u_multiplier/_0617_ ),
    .ZN(\u_multiplier/_0618_ ));
 AOI21_X2 \u_multiplier/_1015_  (.A(\u_multiplier/_0618_ ),
    .B1(\u_multiplier/_0617_ ),
    .B2(\u_multiplier/_0599_ ),
    .ZN(product[8]));
 OAI21_X2 \u_multiplier/_1016_  (.A(\u_multiplier/_0615_ ),
    .B1(\u_multiplier/_0617_ ),
    .B2(\u_multiplier/_0599_ ),
    .ZN(\u_multiplier/_0619_ ));
 AOI21_X2 \u_multiplier/_1017_  (.A(\u_multiplier/_0611_ ),
    .B1(\u_multiplier/_0612_ ),
    .B2(\u_multiplier/_0604_ ),
    .ZN(\u_multiplier/_0620_ ));
 NOR2_X1 \u_multiplier/_1018_  (.A1(\u_multiplier/_0711_ ),
    .A2(\u_multiplier/_0533_ ),
    .ZN(\u_multiplier/_0621_ ));
 AND2_X1 \u_multiplier/_1019_  (.A1(\u_multiplier/K [1]),
    .A2(\u_multiplier/_0577_ ),
    .ZN(\u_multiplier/_0622_ ));
 AOI211_X2 \u_multiplier/_1020_  (.A(\u_multiplier/dec_out [9]),
    .B(\u_multiplier/_0621_ ),
    .C1(\u_multiplier/_0622_ ),
    .C2(\u_multiplier/_0711_ ),
    .ZN(\u_multiplier/_0623_ ));
 INV_X1 \u_multiplier/_1021_  (.A(\u_multiplier/_0623_ ),
    .ZN(\u_multiplier/_0624_ ));
 AND3_X1 \u_multiplier/_1022_  (.A1(\u_multiplier/code_x [0]),
    .A2(\u_multiplier/code_x [1]),
    .A3(\u_multiplier/_0718_ ),
    .ZN(\u_multiplier/_0625_ ));
 OR2_X1 \u_multiplier/_1023_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_0625_ ),
    .ZN(\u_multiplier/_0626_ ));
 OAI21_X2 \u_multiplier/_1024_  (.A(\u_multiplier/_0626_ ),
    .B1(\u_multiplier/_0538_ ),
    .B2(\u_multiplier/_0708_ ),
    .ZN(\u_multiplier/_0627_ ));
 AND3_X1 \u_multiplier/_1025_  (.A1(\u_multiplier/code_y [0]),
    .A2(\u_multiplier/code_y [1]),
    .A3(\u_multiplier/_0716_ ),
    .ZN(\u_multiplier/_0628_ ));
 OR2_X1 \u_multiplier/_1026_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_0628_ ),
    .ZN(\u_multiplier/_0629_ ));
 OAI21_X2 \u_multiplier/_1027_  (.A(\u_multiplier/_0629_ ),
    .B1(\u_multiplier/_0543_ ),
    .B2(\u_multiplier/_0707_ ),
    .ZN(\u_multiplier/_0630_ ));
 NOR2_X1 \u_multiplier/_1028_  (.A1(\u_multiplier/_0627_ ),
    .A2(\u_multiplier/_0630_ ),
    .ZN(\u_multiplier/_0631_ ));
 XOR2_X2 \u_multiplier/_1029_  (.A(\u_multiplier/_0627_ ),
    .B(\u_multiplier/_0630_ ),
    .Z(\u_multiplier/_0632_ ));
 XNOR2_X1 \u_multiplier/_1030_  (.A(\u_multiplier/_0623_ ),
    .B(\u_multiplier/_0632_ ),
    .ZN(\u_multiplier/_0633_ ));
 INV_X1 \u_multiplier/_1031_  (.A(\u_multiplier/_0633_ ),
    .ZN(\u_multiplier/_0634_ ));
 NOR2_X1 \u_multiplier/_1032_  (.A1(\u_multiplier/_0620_ ),
    .A2(\u_multiplier/_0634_ ),
    .ZN(\u_multiplier/_0635_ ));
 XOR2_X1 \u_multiplier/_1033_  (.A(\u_multiplier/_0620_ ),
    .B(\u_multiplier/_0633_ ),
    .Z(\u_multiplier/_0636_ ));
 INV_X1 \u_multiplier/_1034_  (.A(\u_multiplier/_0636_ ),
    .ZN(\u_multiplier/_0637_ ));
 OAI21_X1 \u_multiplier/_1035_  (.A(\u_multiplier/_0439_ ),
    .B1(\u_multiplier/_0619_ ),
    .B2(\u_multiplier/_0637_ ),
    .ZN(\u_multiplier/_0638_ ));
 AOI21_X1 \u_multiplier/_1036_  (.A(\u_multiplier/_0638_ ),
    .B1(\u_multiplier/_0637_ ),
    .B2(\u_multiplier/_0619_ ),
    .ZN(product[9]));
 AOI21_X2 \u_multiplier/_1037_  (.A(\u_multiplier/_0635_ ),
    .B1(\u_multiplier/_0637_ ),
    .B2(\u_multiplier/_0619_ ),
    .ZN(\u_multiplier/_0639_ ));
 AOI21_X1 \u_multiplier/_1038_  (.A(\u_multiplier/_0631_ ),
    .B1(\u_multiplier/_0632_ ),
    .B2(\u_multiplier/_0624_ ),
    .ZN(\u_multiplier/_0640_ ));
 AOI21_X2 \u_multiplier/_1039_  (.A(\u_multiplier/dec_out [10]),
    .B1(\u_multiplier/_0557_ ),
    .B2(\u_multiplier/K [2]),
    .ZN(\u_multiplier/_0641_ ));
 NAND2_X1 \u_multiplier/_1040_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_0561_ ),
    .ZN(\u_multiplier/_0642_ ));
 NAND2_X1 \u_multiplier/_1041_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_0565_ ),
    .ZN(\u_multiplier/_0643_ ));
 OR2_X1 \u_multiplier/_1042_  (.A1(\u_multiplier/_0642_ ),
    .A2(\u_multiplier/_0643_ ),
    .ZN(\u_multiplier/_0644_ ));
 XOR2_X1 \u_multiplier/_1043_  (.A(\u_multiplier/_0642_ ),
    .B(\u_multiplier/_0643_ ),
    .Z(\u_multiplier/_0645_ ));
 INV_X1 \u_multiplier/_1044_  (.A(\u_multiplier/_0645_ ),
    .ZN(\u_multiplier/_0646_ ));
 XNOR2_X1 \u_multiplier/_1045_  (.A(\u_multiplier/_0641_ ),
    .B(\u_multiplier/_0646_ ),
    .ZN(\u_multiplier/_0647_ ));
 OR2_X1 \u_multiplier/_1046_  (.A1(\u_multiplier/_0640_ ),
    .A2(\u_multiplier/_0647_ ),
    .ZN(\u_multiplier/_0648_ ));
 XOR2_X1 \u_multiplier/_1047_  (.A(\u_multiplier/_0640_ ),
    .B(\u_multiplier/_0647_ ),
    .Z(\u_multiplier/_0649_ ));
 INV_X1 \u_multiplier/_1048_  (.A(\u_multiplier/_0649_ ),
    .ZN(\u_multiplier/_0650_ ));
 NOR2_X1 \u_multiplier/_1049_  (.A1(\u_multiplier/_0639_ ),
    .A2(\u_multiplier/_0650_ ),
    .ZN(\u_multiplier/_0651_ ));
 AND2_X1 \u_multiplier/_1050_  (.A1(\u_multiplier/_0639_ ),
    .A2(\u_multiplier/_0650_ ),
    .ZN(\u_multiplier/_0652_ ));
 NOR3_X1 \u_multiplier/_1051_  (.A1(\u_multiplier/_0440_ ),
    .A2(\u_multiplier/_0651_ ),
    .A3(\u_multiplier/_0652_ ),
    .ZN(product[10]));
 OAI21_X2 \u_multiplier/_1052_  (.A(\u_multiplier/_0648_ ),
    .B1(\u_multiplier/_0650_ ),
    .B2(\u_multiplier/_0639_ ),
    .ZN(\u_multiplier/_0653_ ));
 OAI21_X2 \u_multiplier/_1053_  (.A(\u_multiplier/_0644_ ),
    .B1(\u_multiplier/_0646_ ),
    .B2(\u_multiplier/_0641_ ),
    .ZN(\u_multiplier/_0654_ ));
 INV_X1 \u_multiplier/_1054_  (.A(\u_multiplier/_0654_ ),
    .ZN(\u_multiplier/_0655_ ));
 AOI21_X2 \u_multiplier/_1055_  (.A(\u_multiplier/dec_out [11]),
    .B1(\u_multiplier/_0578_ ),
    .B2(\u_multiplier/K [2]),
    .ZN(\u_multiplier/_0656_ ));
 NAND2_X1 \u_multiplier/_1056_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_0584_ ),
    .ZN(\u_multiplier/_0657_ ));
 NAND2_X2 \u_multiplier/_1057_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/_0589_ ),
    .ZN(\u_multiplier/_0658_ ));
 XNOR2_X2 \u_multiplier/_1058_  (.A(\u_multiplier/_0657_ ),
    .B(\u_multiplier/_0658_ ),
    .ZN(\u_multiplier/_0659_ ));
 OR2_X1 \u_multiplier/_1059_  (.A1(\u_multiplier/_0656_ ),
    .A2(\u_multiplier/_0659_ ),
    .ZN(\u_multiplier/_0660_ ));
 XNOR2_X2 \u_multiplier/_1060_  (.A(\u_multiplier/_0656_ ),
    .B(\u_multiplier/_0659_ ),
    .ZN(\u_multiplier/_0661_ ));
 NOR2_X1 \u_multiplier/_1061_  (.A1(\u_multiplier/_0655_ ),
    .A2(\u_multiplier/_0661_ ),
    .ZN(\u_multiplier/_0662_ ));
 XNOR2_X2 \u_multiplier/_1062_  (.A(\u_multiplier/_0654_ ),
    .B(\u_multiplier/_0661_ ),
    .ZN(\u_multiplier/_0663_ ));
 OAI21_X1 \u_multiplier/_1063_  (.A(\u_multiplier/_0439_ ),
    .B1(\u_multiplier/_0653_ ),
    .B2(\u_multiplier/_0663_ ),
    .ZN(\u_multiplier/_0664_ ));
 AOI21_X1 \u_multiplier/_1064_  (.A(\u_multiplier/_0664_ ),
    .B1(\u_multiplier/_0663_ ),
    .B2(\u_multiplier/_0653_ ),
    .ZN(product[11]));
 AOI21_X2 \u_multiplier/_1065_  (.A(\u_multiplier/_0662_ ),
    .B1(\u_multiplier/_0663_ ),
    .B2(\u_multiplier/_0653_ ),
    .ZN(\u_multiplier/_0665_ ));
 OAI21_X2 \u_multiplier/_1066_  (.A(\u_multiplier/_0660_ ),
    .B1(\u_multiplier/_0658_ ),
    .B2(\u_multiplier/_0657_ ),
    .ZN(\u_multiplier/_0666_ ));
 OAI21_X2 \u_multiplier/_1067_  (.A(\u_multiplier/_0712_ ),
    .B1(\u_multiplier/_0601_ ),
    .B2(\u_multiplier/_0711_ ),
    .ZN(\u_multiplier/_0667_ ));
 AND4_X1 \u_multiplier/_1068_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/code_x [2]),
    .A3(\u_multiplier/_0605_ ),
    .A4(\u_multiplier/_0608_ ),
    .ZN(\u_multiplier/_0668_ ));
 AOI22_X1 \u_multiplier/_1069_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_0605_ ),
    .B1(\u_multiplier/_0608_ ),
    .B2(\u_multiplier/code_y [2]),
    .ZN(\u_multiplier/_0669_ ));
 NOR2_X1 \u_multiplier/_1070_  (.A1(\u_multiplier/_0668_ ),
    .A2(\u_multiplier/_0669_ ),
    .ZN(\u_multiplier/_0670_ ));
 XNOR2_X1 \u_multiplier/_1071_  (.A(\u_multiplier/_0667_ ),
    .B(\u_multiplier/_0670_ ),
    .ZN(\u_multiplier/_0671_ ));
 INV_X1 \u_multiplier/_1072_  (.A(\u_multiplier/_0671_ ),
    .ZN(\u_multiplier/_0672_ ));
 NAND2_X1 \u_multiplier/_1073_  (.A1(\u_multiplier/_0666_ ),
    .A2(\u_multiplier/_0672_ ),
    .ZN(\u_multiplier/_0673_ ));
 XNOR2_X2 \u_multiplier/_1074_  (.A(\u_multiplier/_0666_ ),
    .B(\u_multiplier/_0672_ ),
    .ZN(\u_multiplier/_0674_ ));
 AOI21_X1 \u_multiplier/_1075_  (.A(\u_multiplier/_0440_ ),
    .B1(\u_multiplier/_0665_ ),
    .B2(\u_multiplier/_0674_ ),
    .ZN(\u_multiplier/_0675_ ));
 OAI21_X1 \u_multiplier/_1076_  (.A(\u_multiplier/_0675_ ),
    .B1(\u_multiplier/_0674_ ),
    .B2(\u_multiplier/_0665_ ),
    .ZN(\u_multiplier/_0676_ ));
 INV_X1 \u_multiplier/_1077_  (.A(\u_multiplier/_0676_ ),
    .ZN(product[12]));
 OAI21_X2 \u_multiplier/_1078_  (.A(\u_multiplier/_0673_ ),
    .B1(\u_multiplier/_0674_ ),
    .B2(\u_multiplier/_0665_ ),
    .ZN(\u_multiplier/_0677_ ));
 AOI21_X2 \u_multiplier/_1079_  (.A(\u_multiplier/_0668_ ),
    .B1(\u_multiplier/_0670_ ),
    .B2(\u_multiplier/_0667_ ),
    .ZN(\u_multiplier/_0678_ ));
 INV_X1 \u_multiplier/_1080_  (.A(\u_multiplier/_0678_ ),
    .ZN(\u_multiplier/_0679_ ));
 AOI21_X2 \u_multiplier/_1081_  (.A(\u_multiplier/dec_out [13]),
    .B1(\u_multiplier/_0622_ ),
    .B2(\u_multiplier/K [2]),
    .ZN(\u_multiplier/_0680_ ));
 INV_X1 \u_multiplier/_1082_  (.A(\u_multiplier/_0680_ ),
    .ZN(\u_multiplier/_0681_ ));
 AND4_X1 \u_multiplier/_1083_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/code_x [2]),
    .A3(\u_multiplier/_0625_ ),
    .A4(\u_multiplier/_0628_ ),
    .ZN(\u_multiplier/_0682_ ));
 AOI22_X2 \u_multiplier/_1084_  (.A1(\u_multiplier/code_x [2]),
    .A2(\u_multiplier/_0625_ ),
    .B1(\u_multiplier/_0628_ ),
    .B2(\u_multiplier/code_y [2]),
    .ZN(\u_multiplier/_0683_ ));
 NOR2_X2 \u_multiplier/_1085_  (.A1(\u_multiplier/_0682_ ),
    .A2(\u_multiplier/_0683_ ),
    .ZN(\u_multiplier/_0684_ ));
 XNOR2_X2 \u_multiplier/_1086_  (.A(\u_multiplier/_0680_ ),
    .B(\u_multiplier/_0684_ ),
    .ZN(\u_multiplier/_0685_ ));
 NAND2_X1 \u_multiplier/_1087_  (.A1(\u_multiplier/_0679_ ),
    .A2(\u_multiplier/_0685_ ),
    .ZN(\u_multiplier/_0686_ ));
 INV_X1 \u_multiplier/_1088_  (.A(\u_multiplier/_0686_ ),
    .ZN(\u_multiplier/_0687_ ));
 XNOR2_X2 \u_multiplier/_1089_  (.A(\u_multiplier/_0678_ ),
    .B(\u_multiplier/_0685_ ),
    .ZN(\u_multiplier/_0688_ ));
 OAI21_X1 \u_multiplier/_1090_  (.A(\u_multiplier/_0439_ ),
    .B1(\u_multiplier/_0677_ ),
    .B2(\u_multiplier/_0688_ ),
    .ZN(\u_multiplier/_0689_ ));
 AOI21_X1 \u_multiplier/_1091_  (.A(\u_multiplier/_0689_ ),
    .B1(\u_multiplier/_0688_ ),
    .B2(\u_multiplier/_0677_ ),
    .ZN(product[13]));
 AOI21_X2 \u_multiplier/_1092_  (.A(\u_multiplier/_0687_ ),
    .B1(\u_multiplier/_0688_ ),
    .B2(\u_multiplier/_0677_ ),
    .ZN(\u_multiplier/_0690_ ));
 AOI21_X2 \u_multiplier/_1093_  (.A(\u_multiplier/_0682_ ),
    .B1(\u_multiplier/_0684_ ),
    .B2(\u_multiplier/_0681_ ),
    .ZN(\u_multiplier/_0691_ ));
 INV_X1 \u_multiplier/_1094_  (.A(\u_multiplier/_0691_ ),
    .ZN(\u_multiplier/_0692_ ));
 NAND2_X1 \u_multiplier/_1095_  (.A1(\u_multiplier/dec_out [14]),
    .A2(\u_multiplier/_0692_ ),
    .ZN(\u_multiplier/_0693_ ));
 XOR2_X2 \u_multiplier/_1096_  (.A(\u_multiplier/dec_out [14]),
    .B(\u_multiplier/_0691_ ),
    .Z(\u_multiplier/_0694_ ));
 OR2_X1 \u_multiplier/_1097_  (.A1(\u_multiplier/_0690_ ),
    .A2(\u_multiplier/_0694_ ),
    .ZN(\u_multiplier/_0695_ ));
 NAND2_X1 \u_multiplier/_1098_  (.A1(\u_multiplier/_0439_ ),
    .A2(\u_multiplier/_0695_ ),
    .ZN(\u_multiplier/_0696_ ));
 AOI21_X4 \u_multiplier/_1099_  (.A(\u_multiplier/_0696_ ),
    .B1(\u_multiplier/_0694_ ),
    .B2(\u_multiplier/_0690_ ),
    .ZN(product[14]));
 AOI21_X1 \u_multiplier/_1100_  (.A(\u_multiplier/_0713_ ),
    .B1(\u_multiplier/_0693_ ),
    .B2(\u_multiplier/_0695_ ),
    .ZN(\u_multiplier/_0697_ ));
 AND3_X1 \u_multiplier/_1101_  (.A1(\u_multiplier/_0713_ ),
    .A2(\u_multiplier/_0693_ ),
    .A3(\u_multiplier/_0695_ ),
    .ZN(\u_multiplier/_0698_ ));
 NOR3_X1 \u_multiplier/_1102_  (.A1(\u_multiplier/_0440_ ),
    .A2(\u_multiplier/_0697_ ),
    .A3(\u_multiplier/_0698_ ),
    .ZN(product[15]));
 NAND2_X1 \u_multiplier/_1103_  (.A1(\u_multiplier/code_y [2]),
    .A2(\u_multiplier/code_x [2]),
    .ZN(\u_multiplier/_0699_ ));
 NAND2_X1 \u_multiplier/_1104_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/code_x [1]),
    .ZN(\u_multiplier/_0700_ ));
 NAND2_X1 \u_multiplier/_1105_  (.A1(\u_multiplier/code_y [0]),
    .A2(\u_multiplier/code_x [0]),
    .ZN(\u_multiplier/_0701_ ));
 NOR2_X1 \u_multiplier/_1106_  (.A1(\u_multiplier/code_y [1]),
    .A2(\u_multiplier/code_x [1]),
    .ZN(\u_multiplier/_0702_ ));
 XOR2_X2 \u_multiplier/_1107_  (.A(\u_multiplier/code_y [1]),
    .B(\u_multiplier/code_x [1]),
    .Z(\u_multiplier/_0703_ ));
 OAI21_X2 \u_multiplier/_1108_  (.A(\u_multiplier/_0700_ ),
    .B1(\u_multiplier/_0701_ ),
    .B2(\u_multiplier/_0702_ ),
    .ZN(\u_multiplier/_0704_ ));
 INV_X1 \u_multiplier/_1109_  (.A(\u_multiplier/_0704_ ),
    .ZN(\u_multiplier/_0705_ ));
 XNOR2_X2 \u_multiplier/_1110_  (.A(\u_multiplier/code_y [2]),
    .B(\u_multiplier/code_x [2]),
    .ZN(\u_multiplier/_0706_ ));
 OAI21_X4 \u_multiplier/_1111_  (.A(\u_multiplier/_0699_ ),
    .B1(\u_multiplier/_0705_ ),
    .B2(\u_multiplier/_0706_ ),
    .ZN(\u_multiplier/_0355_ ));
 XNOR2_X2 \u_multiplier/_1112_  (.A(\u_multiplier/_0701_ ),
    .B(\u_multiplier/_0703_ ),
    .ZN(\u_multiplier/_0353_ ));
 XNOR2_X2 \u_multiplier/_1113_  (.A(\u_multiplier/_0704_ ),
    .B(\u_multiplier/_0706_ ),
    .ZN(\u_multiplier/_0354_ ));
 XOR2_X2 \u_multiplier/_1114_  (.A(\u_multiplier/code_y [0]),
    .B(\u_multiplier/code_x [0]),
    .Z(\u_multiplier/_0352_ ));
 INV_X2 \u_multiplier/dec/_40_  (.A(\u_multiplier/_0355_ ),
    .ZN(\u_multiplier/dec/_34_ ));
 INV_X1 \u_multiplier/dec/_41_  (.A(\u_multiplier/_0352_ ),
    .ZN(\u_multiplier/dec/_35_ ));
 INV_X2 \u_multiplier/dec/_42_  (.A(\u_multiplier/_0353_ ),
    .ZN(\u_multiplier/dec/_36_ ));
 INV_X2 \u_multiplier/dec/_43_  (.A(\u_multiplier/_0354_ ),
    .ZN(\u_multiplier/dec/_37_ ));
 NOR4_X1 \u_multiplier/dec/_44_  (.A1(\u_multiplier/_0355_ ),
    .A2(\u_multiplier/_0352_ ),
    .A3(\u_multiplier/_0353_ ),
    .A4(\u_multiplier/_0354_ ),
    .ZN(\u_multiplier/dec_out [0]));
 NOR4_X2 \u_multiplier/dec/_45_  (.A1(\u_multiplier/_0355_ ),
    .A2(\u_multiplier/dec/_35_ ),
    .A3(\u_multiplier/_0353_ ),
    .A4(\u_multiplier/_0354_ ),
    .ZN(\u_multiplier/dec_out [1]));
 NOR4_X2 \u_multiplier/dec/_46_  (.A1(\u_multiplier/_0355_ ),
    .A2(\u_multiplier/_0352_ ),
    .A3(\u_multiplier/dec/_36_ ),
    .A4(\u_multiplier/_0354_ ),
    .ZN(\u_multiplier/dec_out [2]));
 NAND2_X1 \u_multiplier/dec/_47_  (.A1(\u_multiplier/_0352_ ),
    .A2(\u_multiplier/_0353_ ),
    .ZN(\u_multiplier/dec/_38_ ));
 NOR3_X1 \u_multiplier/dec/_48_  (.A1(\u_multiplier/_0355_ ),
    .A2(\u_multiplier/_0354_ ),
    .A3(\u_multiplier/dec/_38_ ),
    .ZN(\u_multiplier/dec_out [3]));
 NOR4_X1 \u_multiplier/dec/_49_  (.A1(\u_multiplier/_0355_ ),
    .A2(\u_multiplier/_0352_ ),
    .A3(\u_multiplier/_0353_ ),
    .A4(\u_multiplier/dec/_37_ ),
    .ZN(\u_multiplier/dec_out [4]));
 NOR4_X1 \u_multiplier/dec/_50_  (.A1(\u_multiplier/_0355_ ),
    .A2(\u_multiplier/dec/_35_ ),
    .A3(\u_multiplier/_0353_ ),
    .A4(\u_multiplier/dec/_37_ ),
    .ZN(\u_multiplier/dec_out [5]));
 NOR4_X1 \u_multiplier/dec/_51_  (.A1(\u_multiplier/_0355_ ),
    .A2(\u_multiplier/_0352_ ),
    .A3(\u_multiplier/dec/_36_ ),
    .A4(\u_multiplier/dec/_37_ ),
    .ZN(\u_multiplier/dec_out [6]));
 NAND3_X1 \u_multiplier/dec/_52_  (.A1(\u_multiplier/_0352_ ),
    .A2(\u_multiplier/_0353_ ),
    .A3(\u_multiplier/_0354_ ),
    .ZN(\u_multiplier/dec/_39_ ));
 NOR2_X1 \u_multiplier/dec/_53_  (.A1(\u_multiplier/_0355_ ),
    .A2(\u_multiplier/dec/_39_ ),
    .ZN(\u_multiplier/dec_out [7]));
 NOR4_X1 \u_multiplier/dec/_54_  (.A1(\u_multiplier/dec/_34_ ),
    .A2(\u_multiplier/_0352_ ),
    .A3(\u_multiplier/_0353_ ),
    .A4(\u_multiplier/_0354_ ),
    .ZN(\u_multiplier/dec_out [8]));
 NOR4_X1 \u_multiplier/dec/_55_  (.A1(\u_multiplier/dec/_34_ ),
    .A2(\u_multiplier/dec/_35_ ),
    .A3(\u_multiplier/_0353_ ),
    .A4(\u_multiplier/_0354_ ),
    .ZN(\u_multiplier/dec_out [9]));
 NOR4_X2 \u_multiplier/dec/_56_  (.A1(\u_multiplier/dec/_34_ ),
    .A2(\u_multiplier/_0352_ ),
    .A3(\u_multiplier/dec/_36_ ),
    .A4(\u_multiplier/_0354_ ),
    .ZN(\u_multiplier/dec_out [10]));
 NOR3_X1 \u_multiplier/dec/_57_  (.A1(\u_multiplier/dec/_34_ ),
    .A2(\u_multiplier/_0354_ ),
    .A3(\u_multiplier/dec/_38_ ),
    .ZN(\u_multiplier/dec_out [11]));
 NOR4_X1 \u_multiplier/dec/_58_  (.A1(\u_multiplier/dec/_34_ ),
    .A2(\u_multiplier/_0352_ ),
    .A3(\u_multiplier/_0353_ ),
    .A4(\u_multiplier/dec/_37_ ),
    .ZN(\u_multiplier/dec_out [12]));
 NOR4_X1 \u_multiplier/dec/_59_  (.A1(\u_multiplier/dec/_34_ ),
    .A2(\u_multiplier/dec/_35_ ),
    .A3(\u_multiplier/_0353_ ),
    .A4(\u_multiplier/dec/_37_ ),
    .ZN(\u_multiplier/dec_out [13]));
 NOR4_X4 \u_multiplier/dec/_60_  (.A1(\u_multiplier/dec/_34_ ),
    .A2(\u_multiplier/_0352_ ),
    .A3(\u_multiplier/dec/_36_ ),
    .A4(\u_multiplier/dec/_37_ ),
    .ZN(\u_multiplier/dec_out [14]));
 NOR2_X1 \u_multiplier/dec/_61_  (.A1(\u_multiplier/dec/_34_ ),
    .A2(\u_multiplier/dec/_39_ ),
    .ZN(\u_multiplier/dec_out [15]));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_2_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_2_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_2_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_2_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_2_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_2_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_2_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_2_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_2_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_2_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_2_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_2_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_2_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_2_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_2_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_2_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_2_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_2_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_2_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_2_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_2_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_2_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_2_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_2_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_2_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_2_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_2_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_2_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_2_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_2_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_2_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_2_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_2_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_2_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_2_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_2_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_2_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_2_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_2_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_2_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_2_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_2_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_2_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_2_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_2_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_2_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_2_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_2_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_2_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_2_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_2_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_2_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_2_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_2_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_2_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_2_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_2_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_2_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_2_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_2_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_2_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_2_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_2_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_2_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_2_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_2_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_2_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_2_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_2_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_2_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_2_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_2_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_2_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_2_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_1_Left_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_1_Left_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_1_Left_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_1_Left_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_1_Left_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_1_Left_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_1_Left_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_1_Left_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_1_Left_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_1_Left_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_1_Left_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_1_Left_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_1_Left_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_1_Left_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_1_Left_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_1_Left_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_1_Left_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_1_Left_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_1_Left_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_1_Left_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_1_Left_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_1_Left_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_1_Left_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_1_Left_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_1_Left_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_1_Left_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_1_Left_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_1_Left_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_1_Left_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_1_Left_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_1_Left_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_1_Left_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_1_Left_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_1_Left_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_1_Left_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_1_Left_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_1_Left_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_1_Left_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_1_Left_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_1_Left_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_1_Left_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_1_Left_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_1_Left_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_1_Left_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_1_Left_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_1_Left_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_1_Left_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_1_Left_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_1_Left_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_1_Left_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_1_Left_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_1_Left_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_1_Left_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_1_Left_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_1_Left_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_1_Left_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_1_Left_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_1_Left_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_1_Left_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_1_Left_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_1_Left_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_1_Left_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_1_Left_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_1_Left_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_1_Left_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_1_Left_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_1_Left_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_1_Left_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_1_Left_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_1_Left_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_1_Left_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_1_Left_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_1_Left_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Left_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Left_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Left_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Left_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Left_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Left_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Left_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Left_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Left_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Left_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_1_Left_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_2_Left_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_2_Left_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_2_Left_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_2_Left_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_2_Left_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_2_Left_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_2_Left_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_2_Left_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_2_Left_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_2_Left_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_2_Left_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_2_Left_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_2_Left_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_2_Left_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_2_Left_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_2_Left_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_2_Left_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_2_Left_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_2_Left_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_2_Left_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_2_Left_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_2_Left_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_2_Left_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_2_Left_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_2_Left_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_2_Left_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_2_Left_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_2_Left_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_2_Left_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_2_Left_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_2_Left_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_2_Left_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_2_Left_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_2_Left_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_2_Left_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_2_Left_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_2_Left_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_2_Left_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_2_Left_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_2_Left_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_2_Left_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_2_Left_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_2_Left_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_2_Left_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_2_Left_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_2_Left_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_2_Left_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_2_Left_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_2_Left_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_2_Left_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_2_Left_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_2_Left_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_2_Left_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_2_Left_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_2_Left_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_2_Left_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_2_Left_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_2_Left_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_2_Left_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_2_Left_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_2_Left_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_2_Left_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_2_Left_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_2_Left_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_2_Left_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_2_Left_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_2_Left_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_2_Left_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_2_Left_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_2_Left_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_2_Left_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_2_Left_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_2_Left_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_2_Left_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_1_Right_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_1_Right_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_1_Right_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_1_Right_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_1_Right_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_1_Right_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_1_Right_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_1_Right_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_1_Right_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_1_Right_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_1_Right_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_1_Right_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_1_Right_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_1_Right_265 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_1_Right_266 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_1_Right_267 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_1_Right_268 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_1_Right_269 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_1_Right_270 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_1_Right_271 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_1_Right_272 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_1_Right_273 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_1_Right_274 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_1_Right_275 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_1_Right_276 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_1_Right_277 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_1_Right_278 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_1_Right_279 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_1_Right_280 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_1_Right_281 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_1_Right_282 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_1_Right_283 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_1_Right_284 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_1_Right_285 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_1_Right_286 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_1_Right_287 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_1_Right_288 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_1_Right_289 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_1_Right_290 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_1_Right_291 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_1_Right_292 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_1_Right_293 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_1_Right_294 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_1_Right_295 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_1_Right_296 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_1_Right_297 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_1_Right_298 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_1_Right_299 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_1_Right_300 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_1_Right_301 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_1_Right_302 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_1_Right_303 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_1_Right_304 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_1_Right_305 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_1_Right_306 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_1_Right_307 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_1_Right_308 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_1_Right_309 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_1_Right_310 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_1_Right_311 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_1_Right_312 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_1_Right_313 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_1_Right_314 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_1_Right_315 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_1_Right_316 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_1_Right_317 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_1_Right_318 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_1_Right_319 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_1_Right_320 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_1_Right_321 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_1_Right_322 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_1_Right_323 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_1_Right_324 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_1_Right_325 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_326 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_327 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_328 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_79_329 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_330 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_331 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_332 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_333 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_334 ();
 LOGIC1_X1 \u_multiplier/NOD/nod_cels[5].Nod_bits/_07__30  (.Z(net30));
 CLKBUF_X1 hold31 (.A(net56),
    .Z(net31));
 BUF_X2 input1 (.A(data_in[0]),
    .Z(net1));
 BUF_X1 input2 (.A(data_in[1]),
    .Z(net2));
 BUF_X1 input3 (.A(data_in[2]),
    .Z(net3));
 CLKBUF_X2 input4 (.A(data_in[3]),
    .Z(net4));
 CLKBUF_X2 input5 (.A(data_in[4]),
    .Z(net5));
 BUF_X1 input6 (.A(data_in[5]),
    .Z(net6));
 BUF_X2 input7 (.A(data_in[6]),
    .Z(net7));
 BUF_X1 input8 (.A(data_in[7]),
    .Z(net8));
 BUF_X2 input9 (.A(init_enable),
    .Z(net9));
 BUF_X2 input10 (.A(pe_ce),
    .Z(net10));
 BUF_X8 input11 (.A(rst_n),
    .Z(net11));
 BUF_X1 output12 (.A(net12),
    .Z(curr_state[1]));
 BUF_X1 output13 (.A(net13),
    .Z(data_out[0]));
 BUF_X1 output14 (.A(net14),
    .Z(data_out[10]));
 BUF_X1 output15 (.A(net15),
    .Z(data_out[11]));
 BUF_X1 output16 (.A(net16),
    .Z(data_out[12]));
 BUF_X1 output17 (.A(net17),
    .Z(data_out[13]));
 BUF_X1 output18 (.A(net18),
    .Z(data_out[14]));
 BUF_X1 output19 (.A(net19),
    .Z(data_out[15]));
 BUF_X1 output20 (.A(net20),
    .Z(data_out[1]));
 BUF_X1 output21 (.A(net21),
    .Z(data_out[2]));
 BUF_X1 output22 (.A(net22),
    .Z(data_out[3]));
 BUF_X1 output23 (.A(net23),
    .Z(data_out[4]));
 BUF_X1 output24 (.A(net24),
    .Z(data_out[5]));
 BUF_X1 output25 (.A(net25),
    .Z(data_out[6]));
 BUF_X1 output26 (.A(net26),
    .Z(data_out[7]));
 BUF_X1 output27 (.A(net27),
    .Z(data_out[8]));
 BUF_X1 output28 (.A(net28),
    .Z(data_out[9]));
 BUF_X1 output29 (.A(net29),
    .Z(valid_reg_out));
 CLKBUF_X1 hold32 (.A(net60),
    .Z(net32));
 CLKBUF_X1 hold33 (.A(net67),
    .Z(net33));
 CLKBUF_X1 hold34 (.A(net53),
    .Z(net34));
 CLKBUF_X1 hold35 (.A(net65),
    .Z(net35));
 CLKBUF_X1 hold36 (.A(net69),
    .Z(net36));
 CLKBUF_X1 hold37 (.A(net71),
    .Z(net37));
 CLKBUF_X1 hold38 (.A(net78),
    .Z(net38));
 CLKBUF_X1 hold39 (.A(net76),
    .Z(net39));
 CLKBUF_X1 hold40 (.A(net63),
    .Z(net40));
 CLKBUF_X1 hold41 (.A(net74),
    .Z(net41));
 CLKBUF_X1 hold42 (.A(net81),
    .Z(net42));
 CLKBUF_X1 hold43 (.A(net83),
    .Z(net43));
 CLKBUF_X1 hold44 (.A(net84),
    .Z(net44));
 CLKBUF_X1 hold45 (.A(net86),
    .Z(net45));
 CLKBUF_X1 hold46 (.A(net87),
    .Z(net46));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 CLKBUF_X3 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 CLKBUF_X3 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 CLKBUF_X3 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 INV_X2 clkload0 (.A(clknet_2_0__leaf_clk));
 CLKBUF_X1 clkload1 (.A(clknet_2_2__leaf_clk));
 INV_X1 clkload2 (.A(clknet_2_3__leaf_clk));
 CLKBUF_X1 hold1 (.A(_265_),
    .Z(net47));
 CLKBUF_X1 hold2 (.A(_194_),
    .Z(net48));
 CLKBUF_X1 hold3 (.A(_266_),
    .Z(net49));
 CLKBUF_X1 hold4 (.A(_197_),
    .Z(net50));
 CLKBUF_X1 hold5 (.A(net89),
    .Z(net51));
 CLKBUF_X1 hold6 (.A(net88),
    .Z(net52));
 CLKBUF_X1 hold7 (.A(_267_),
    .Z(net53));
 CLKBUF_X1 hold8 (.A(_201_),
    .Z(net54));
 CLKBUF_X1 hold9 (.A(_093_),
    .Z(net55));
 CLKBUF_X1 hold10 (.A(_244_),
    .Z(net56));
 CLKBUF_X1 hold11 (.A(net31),
    .Z(net57));
 CLKBUF_X1 hold12 (.A(_133_),
    .Z(net58));
 CLKBUF_X1 hold13 (.A(net90),
    .Z(net59));
 CLKBUF_X1 hold14 (.A(_268_),
    .Z(net60));
 CLKBUF_X1 hold15 (.A(net32),
    .Z(net61));
 CLKBUF_X1 hold16 (.A(_118_),
    .Z(net62));
 CLKBUF_X1 hold17 (.A(_264_),
    .Z(net63));
 CLKBUF_X1 hold18 (.A(_188_),
    .Z(net64));
 CLKBUF_X1 hold19 (.A(addr_ptr[1]),
    .Z(net65));
 CLKBUF_X1 hold20 (.A(net35),
    .Z(net66));
 CLKBUF_X1 hold21 (.A(addr_ptr[3]),
    .Z(net67));
 CLKBUF_X1 hold22 (.A(net33),
    .Z(net68));
 CLKBUF_X1 hold23 (.A(addr_ptr[2]),
    .Z(net69));
 CLKBUF_X1 hold24 (.A(net36),
    .Z(net70));
 CLKBUF_X1 hold25 (.A(_270_),
    .Z(net71));
 CLKBUF_X1 hold26 (.A(net37),
    .Z(net72));
 CLKBUF_X1 hold27 (.A(_120_),
    .Z(net73));
 CLKBUF_X1 hold28 (.A(addr_ptr[0]),
    .Z(net74));
 CLKBUF_X1 hold29 (.A(net41),
    .Z(net75));
 CLKBUF_X1 hold30 (.A(_271_),
    .Z(net76));
 CLKBUF_X1 hold47 (.A(_121_),
    .Z(net77));
 CLKBUF_X1 hold48 (.A(_269_),
    .Z(net78));
 CLKBUF_X1 hold49 (.A(net38),
    .Z(net79));
 CLKBUF_X1 hold50 (.A(_119_),
    .Z(net80));
 CLKBUF_X1 hold51 (.A(\u_multiplier/LODx/z [7]),
    .Z(net81));
 CLKBUF_X1 hold52 (.A(curr_state[2]),
    .Z(net82));
 CLKBUF_X1 hold53 (.A(data_in_reg[5]),
    .Z(net83));
 CLKBUF_X1 hold54 (.A(data_in_reg[4]),
    .Z(net84));
 CLKBUF_X1 hold55 (.A(curr_state[0]),
    .Z(net85));
 CLKBUF_X1 hold56 (.A(data_in_reg[0]),
    .Z(net86));
 CLKBUF_X1 hold57 (.A(data_in_reg[1]),
    .Z(net87));
 CLKBUF_X1 hold58 (.A(\u_multiplier/LODx/z [3]),
    .Z(net88));
 CLKBUF_X1 hold59 (.A(data_in_reg[2]),
    .Z(net89));
 CLKBUF_X1 hold60 (.A(data_in_reg[6]),
    .Z(net90));
 assign init_done = curr_state[1];
 assign valid_out = valid_reg_out;
endmodule
