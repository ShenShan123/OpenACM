module sram_multiplier_system (clk,
    init_done,
    init_enable,
    pe_ce,
    rst_n,
    valid_out,
    data_in,
    data_out);
 input clk;
 output init_done;
 input init_enable;
 input pe_ce;
 input rst_n;
 output valid_out;
 input [31:0] data_in;
 output [63:0] data_out;

 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net161;
 wire net163;
 wire \u_multiplier/pp1_0 ;
 wire \u_multiplier/pp1_62 ;
 wire net132;
 wire \u_multiplier/pp2_0 ;
 wire \u_multiplier/pp2_62 ;
 wire net140;
 wire \u_multiplier/pp3_0 ;
 wire \u_multiplier/pp3_62 ;
 wire net147;
 wire \u_multiplier/Final_add/Cout ;
 wire \u_multiplier/Final_add/c1 ;
 wire \u_multiplier/Final_add/cla1/c1 ;
 wire \u_multiplier/Final_add/cla1/cla1/c1 ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/c1 ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_25_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_26_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_27_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_28_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_29_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_30_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_31_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_32_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_33_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_34_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_35_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_36_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_37_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_38_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_39_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_25_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_26_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_27_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_28_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_29_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_30_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_31_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_32_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_33_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_34_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_35_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_36_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_37_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_38_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_39_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/c1 ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_25_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_26_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_27_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_28_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_29_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_30_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_31_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_32_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_33_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_34_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_35_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_36_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_37_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_38_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_39_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_25_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_26_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_27_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_28_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_29_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_30_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_31_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_32_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_33_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_34_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_35_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_36_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_37_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_38_ ;
 wire \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_39_ ;
 wire \u_multiplier/Final_add/cla1/cla2/c1 ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/c1 ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_25_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_26_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_27_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_28_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_29_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_30_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_31_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_32_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_33_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_34_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_35_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_36_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_37_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_38_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_39_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_25_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_26_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_27_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_28_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_29_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_30_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_31_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_32_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_33_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_34_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_35_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_36_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_37_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_38_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_39_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/c1 ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_25_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_26_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_27_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_28_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_29_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_30_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_31_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_32_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_33_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_34_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_35_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_36_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_37_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_38_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_39_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_25_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_26_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_27_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_28_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_29_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_30_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_31_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_32_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_33_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_34_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_35_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_36_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_37_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_38_ ;
 wire \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_39_ ;
 wire \u_multiplier/Final_add/cla2/c1 ;
 wire \u_multiplier/Final_add/cla2/cla1/c1 ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/c1 ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_25_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_26_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_27_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_28_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_29_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_30_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_31_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_32_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_33_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_34_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_35_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_36_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_37_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_38_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_39_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_25_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_26_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_27_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_28_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_29_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_30_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_31_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_32_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_33_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_34_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_35_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_36_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_37_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_38_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_39_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/c1 ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_25_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_26_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_27_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_28_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_29_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_30_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_31_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_32_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_33_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_34_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_35_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_36_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_37_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_38_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_39_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_25_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_26_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_27_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_28_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_29_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_30_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_31_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_32_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_33_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_34_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_35_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_36_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_37_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_38_ ;
 wire \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_39_ ;
 wire \u_multiplier/Final_add/cla2/cla2/c1 ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/c1 ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_25_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_26_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_27_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_28_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_29_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_30_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_31_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_32_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_33_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_34_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_35_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_36_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_37_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_38_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_39_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_25_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_26_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_27_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_28_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_29_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_30_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_31_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_32_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_33_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_34_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_35_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_36_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_37_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_38_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_39_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/c1 ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_25_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_26_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_27_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_28_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_29_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_30_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_31_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_32_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_33_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_34_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_35_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_36_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_37_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_38_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_39_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_25_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_26_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_27_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_28_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_29_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_30_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_31_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_32_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_33_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_34_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_35_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_36_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_37_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_38_ ;
 wire \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_39_ ;
 wire \u_multiplier/STAGE1/_0607_ ;
 wire \u_multiplier/STAGE1/_0608_ ;
 wire \u_multiplier/STAGE1/_0609_ ;
 wire \u_multiplier/STAGE1/_0610_ ;
 wire \u_multiplier/STAGE1/_0611_ ;
 wire \u_multiplier/STAGE1/_0612_ ;
 wire \u_multiplier/STAGE1/_0613_ ;
 wire \u_multiplier/STAGE1/_0614_ ;
 wire \u_multiplier/STAGE1/_0615_ ;
 wire \u_multiplier/STAGE1/_0616_ ;
 wire \u_multiplier/STAGE1/_0617_ ;
 wire \u_multiplier/STAGE1/_0618_ ;
 wire \u_multiplier/STAGE1/_0619_ ;
 wire \u_multiplier/STAGE1/_0620_ ;
 wire \u_multiplier/STAGE1/_0621_ ;
 wire \u_multiplier/STAGE1/_0622_ ;
 wire \u_multiplier/STAGE1/_0623_ ;
 wire \u_multiplier/STAGE1/_0624_ ;
 wire \u_multiplier/STAGE1/_0625_ ;
 wire \u_multiplier/STAGE1/_0626_ ;
 wire \u_multiplier/STAGE1/_0627_ ;
 wire \u_multiplier/STAGE1/_0628_ ;
 wire \u_multiplier/STAGE1/_0629_ ;
 wire \u_multiplier/STAGE1/_0630_ ;
 wire \u_multiplier/STAGE1/_0631_ ;
 wire \u_multiplier/STAGE1/_0632_ ;
 wire \u_multiplier/STAGE1/_0633_ ;
 wire \u_multiplier/STAGE1/_0634_ ;
 wire \u_multiplier/STAGE1/_0635_ ;
 wire \u_multiplier/STAGE1/_0636_ ;
 wire \u_multiplier/STAGE1/_0637_ ;
 wire \u_multiplier/STAGE1/_0638_ ;
 wire \u_multiplier/STAGE1/_0639_ ;
 wire \u_multiplier/STAGE1/_0640_ ;
 wire \u_multiplier/STAGE1/_0641_ ;
 wire \u_multiplier/STAGE1/_0642_ ;
 wire \u_multiplier/STAGE1/_0643_ ;
 wire \u_multiplier/STAGE1/_0644_ ;
 wire \u_multiplier/STAGE1/_0645_ ;
 wire \u_multiplier/STAGE1/_0646_ ;
 wire \u_multiplier/STAGE1/_0647_ ;
 wire \u_multiplier/STAGE1/_0648_ ;
 wire \u_multiplier/STAGE1/_0649_ ;
 wire \u_multiplier/STAGE1/_0650_ ;
 wire \u_multiplier/STAGE1/_0651_ ;
 wire \u_multiplier/STAGE1/_0652_ ;
 wire \u_multiplier/STAGE1/_0653_ ;
 wire \u_multiplier/STAGE1/_0654_ ;
 wire \u_multiplier/STAGE1/_0655_ ;
 wire \u_multiplier/STAGE1/_0656_ ;
 wire \u_multiplier/STAGE1/_0657_ ;
 wire \u_multiplier/STAGE1/_0658_ ;
 wire \u_multiplier/STAGE1/_0659_ ;
 wire \u_multiplier/STAGE1/_0660_ ;
 wire \u_multiplier/STAGE1/_0661_ ;
 wire \u_multiplier/STAGE1/_0662_ ;
 wire \u_multiplier/STAGE1/_0663_ ;
 wire \u_multiplier/STAGE1/_0664_ ;
 wire \u_multiplier/STAGE1/_0665_ ;
 wire \u_multiplier/STAGE1/_0666_ ;
 wire \u_multiplier/STAGE1/_0667_ ;
 wire \u_multiplier/STAGE1/_0668_ ;
 wire \u_multiplier/STAGE1/_0669_ ;
 wire \u_multiplier/STAGE1/_0670_ ;
 wire \u_multiplier/STAGE1/_0671_ ;
 wire \u_multiplier/STAGE1/_0672_ ;
 wire \u_multiplier/STAGE1/_0673_ ;
 wire \u_multiplier/STAGE1/_0674_ ;
 wire \u_multiplier/STAGE1/_0675_ ;
 wire \u_multiplier/STAGE1/_0676_ ;
 wire \u_multiplier/STAGE1/_0677_ ;
 wire \u_multiplier/STAGE1/_0678_ ;
 wire \u_multiplier/STAGE1/_0679_ ;
 wire \u_multiplier/STAGE1/_0680_ ;
 wire \u_multiplier/STAGE1/_0681_ ;
 wire \u_multiplier/STAGE1/_0682_ ;
 wire \u_multiplier/STAGE1/_0683_ ;
 wire \u_multiplier/STAGE1/_0684_ ;
 wire \u_multiplier/STAGE1/_0685_ ;
 wire \u_multiplier/STAGE1/_0686_ ;
 wire \u_multiplier/STAGE1/_0687_ ;
 wire \u_multiplier/STAGE1/_0688_ ;
 wire \u_multiplier/STAGE1/_0689_ ;
 wire \u_multiplier/STAGE1/_0690_ ;
 wire \u_multiplier/STAGE1/_0691_ ;
 wire \u_multiplier/STAGE1/_0692_ ;
 wire \u_multiplier/STAGE1/_0693_ ;
 wire \u_multiplier/STAGE1/_0694_ ;
 wire \u_multiplier/STAGE1/_0695_ ;
 wire \u_multiplier/STAGE1/_0696_ ;
 wire \u_multiplier/STAGE1/_0697_ ;
 wire \u_multiplier/STAGE1/_0698_ ;
 wire \u_multiplier/STAGE1/_0699_ ;
 wire \u_multiplier/STAGE1/_0700_ ;
 wire \u_multiplier/STAGE1/_0701_ ;
 wire \u_multiplier/STAGE1/_0702_ ;
 wire \u_multiplier/STAGE1/_0703_ ;
 wire \u_multiplier/STAGE1/_0704_ ;
 wire \u_multiplier/STAGE1/_0705_ ;
 wire \u_multiplier/STAGE1/_0706_ ;
 wire \u_multiplier/STAGE1/_0707_ ;
 wire \u_multiplier/STAGE1/_0708_ ;
 wire \u_multiplier/STAGE1/_0709_ ;
 wire \u_multiplier/STAGE1/_0710_ ;
 wire \u_multiplier/STAGE1/_0711_ ;
 wire \u_multiplier/STAGE1/_0712_ ;
 wire \u_multiplier/STAGE1/_0713_ ;
 wire \u_multiplier/STAGE1/_0714_ ;
 wire \u_multiplier/STAGE1/_0715_ ;
 wire \u_multiplier/STAGE1/_0716_ ;
 wire \u_multiplier/STAGE1/_0717_ ;
 wire \u_multiplier/STAGE1/_0718_ ;
 wire \u_multiplier/STAGE1/_0719_ ;
 wire \u_multiplier/STAGE1/_0720_ ;
 wire \u_multiplier/STAGE1/_0721_ ;
 wire \u_multiplier/STAGE1/_0722_ ;
 wire \u_multiplier/STAGE1/_0723_ ;
 wire \u_multiplier/STAGE1/_0724_ ;
 wire \u_multiplier/STAGE1/_0725_ ;
 wire \u_multiplier/STAGE1/_0726_ ;
 wire \u_multiplier/STAGE1/_0727_ ;
 wire \u_multiplier/STAGE1/_0728_ ;
 wire \u_multiplier/STAGE1/_0729_ ;
 wire \u_multiplier/STAGE1/_0730_ ;
 wire \u_multiplier/STAGE1/_0731_ ;
 wire \u_multiplier/STAGE1/_0732_ ;
 wire \u_multiplier/STAGE1/_0733_ ;
 wire \u_multiplier/STAGE1/_0734_ ;
 wire \u_multiplier/STAGE1/_0735_ ;
 wire \u_multiplier/STAGE1/_0736_ ;
 wire \u_multiplier/STAGE1/_0737_ ;
 wire \u_multiplier/STAGE1/_0738_ ;
 wire \u_multiplier/STAGE1/_0739_ ;
 wire \u_multiplier/STAGE1/_0740_ ;
 wire \u_multiplier/STAGE1/_0741_ ;
 wire \u_multiplier/STAGE1/_0742_ ;
 wire \u_multiplier/STAGE1/_0743_ ;
 wire \u_multiplier/STAGE1/_0744_ ;
 wire \u_multiplier/STAGE1/_0745_ ;
 wire \u_multiplier/STAGE1/_0746_ ;
 wire \u_multiplier/STAGE1/_0747_ ;
 wire \u_multiplier/STAGE1/_0748_ ;
 wire \u_multiplier/STAGE1/_0749_ ;
 wire \u_multiplier/STAGE1/_0750_ ;
 wire \u_multiplier/STAGE1/_0751_ ;
 wire \u_multiplier/STAGE1/_0752_ ;
 wire \u_multiplier/STAGE1/_0753_ ;
 wire \u_multiplier/STAGE1/_0754_ ;
 wire \u_multiplier/STAGE1/_0755_ ;
 wire \u_multiplier/STAGE1/_0756_ ;
 wire \u_multiplier/STAGE1/_0757_ ;
 wire \u_multiplier/STAGE1/_0758_ ;
 wire \u_multiplier/STAGE1/_0759_ ;
 wire \u_multiplier/STAGE1/_0760_ ;
 wire \u_multiplier/STAGE1/_0761_ ;
 wire \u_multiplier/STAGE1/_0762_ ;
 wire \u_multiplier/STAGE1/_0763_ ;
 wire \u_multiplier/STAGE1/_0764_ ;
 wire \u_multiplier/STAGE1/_0765_ ;
 wire \u_multiplier/STAGE1/_0766_ ;
 wire \u_multiplier/STAGE1/_0767_ ;
 wire \u_multiplier/STAGE1/_0768_ ;
 wire \u_multiplier/STAGE1/_0769_ ;
 wire \u_multiplier/STAGE1/_0770_ ;
 wire \u_multiplier/STAGE1/_0771_ ;
 wire \u_multiplier/STAGE1/_0772_ ;
 wire \u_multiplier/STAGE1/_0773_ ;
 wire \u_multiplier/STAGE1/_0774_ ;
 wire \u_multiplier/STAGE1/_0775_ ;
 wire \u_multiplier/STAGE1/_0776_ ;
 wire \u_multiplier/STAGE1/_0777_ ;
 wire \u_multiplier/STAGE1/_0778_ ;
 wire \u_multiplier/STAGE1/_0779_ ;
 wire \u_multiplier/STAGE1/_0780_ ;
 wire \u_multiplier/STAGE1/_0781_ ;
 wire \u_multiplier/STAGE1/_0782_ ;
 wire \u_multiplier/STAGE1/_0783_ ;
 wire \u_multiplier/STAGE1/_0784_ ;
 wire \u_multiplier/STAGE1/_0785_ ;
 wire \u_multiplier/STAGE1/_0786_ ;
 wire \u_multiplier/STAGE1/_0787_ ;
 wire \u_multiplier/STAGE1/_0788_ ;
 wire \u_multiplier/STAGE1/_0789_ ;
 wire \u_multiplier/STAGE1/_0790_ ;
 wire \u_multiplier/STAGE1/_0791_ ;
 wire \u_multiplier/STAGE1/_0792_ ;
 wire \u_multiplier/STAGE1/_0793_ ;
 wire \u_multiplier/STAGE1/_0794_ ;
 wire \u_multiplier/STAGE1/_0795_ ;
 wire \u_multiplier/STAGE1/_0796_ ;
 wire \u_multiplier/STAGE1/_0797_ ;
 wire \u_multiplier/STAGE1/_0798_ ;
 wire \u_multiplier/STAGE1/_0799_ ;
 wire \u_multiplier/STAGE1/_0800_ ;
 wire \u_multiplier/STAGE1/_0801_ ;
 wire \u_multiplier/STAGE1/_0802_ ;
 wire \u_multiplier/STAGE1/_0803_ ;
 wire \u_multiplier/STAGE1/_0804_ ;
 wire \u_multiplier/STAGE1/_0805_ ;
 wire \u_multiplier/STAGE1/_0806_ ;
 wire \u_multiplier/STAGE1/_0807_ ;
 wire \u_multiplier/STAGE1/_0808_ ;
 wire \u_multiplier/STAGE1/_0809_ ;
 wire \u_multiplier/STAGE1/_0810_ ;
 wire \u_multiplier/STAGE1/_0811_ ;
 wire \u_multiplier/STAGE1/_0812_ ;
 wire \u_multiplier/STAGE1/_0813_ ;
 wire \u_multiplier/STAGE1/_0814_ ;
 wire \u_multiplier/STAGE1/_0815_ ;
 wire \u_multiplier/STAGE1/_0816_ ;
 wire \u_multiplier/STAGE1/_0817_ ;
 wire \u_multiplier/STAGE1/_0818_ ;
 wire \u_multiplier/STAGE1/_0819_ ;
 wire \u_multiplier/STAGE1/_0820_ ;
 wire \u_multiplier/STAGE1/_0821_ ;
 wire \u_multiplier/STAGE1/_0822_ ;
 wire \u_multiplier/STAGE1/_0823_ ;
 wire \u_multiplier/STAGE1/_0824_ ;
 wire \u_multiplier/STAGE1/_0825_ ;
 wire \u_multiplier/STAGE1/_0826_ ;
 wire \u_multiplier/STAGE1/_0827_ ;
 wire \u_multiplier/STAGE1/_0828_ ;
 wire \u_multiplier/STAGE1/_0829_ ;
 wire \u_multiplier/STAGE1/_0830_ ;
 wire \u_multiplier/STAGE1/_0831_ ;
 wire \u_multiplier/STAGE1/_0832_ ;
 wire \u_multiplier/STAGE1/_0833_ ;
 wire \u_multiplier/STAGE1/_0834_ ;
 wire \u_multiplier/STAGE1/_0835_ ;
 wire \u_multiplier/STAGE1/_0836_ ;
 wire \u_multiplier/STAGE1/_0837_ ;
 wire \u_multiplier/STAGE1/_0838_ ;
 wire \u_multiplier/STAGE1/_0839_ ;
 wire \u_multiplier/STAGE1/_0840_ ;
 wire \u_multiplier/STAGE1/_0841_ ;
 wire \u_multiplier/STAGE1/_0842_ ;
 wire \u_multiplier/STAGE1/_0843_ ;
 wire \u_multiplier/STAGE1/_0844_ ;
 wire \u_multiplier/STAGE1/_0845_ ;
 wire \u_multiplier/STAGE1/_0846_ ;
 wire \u_multiplier/STAGE1/_0847_ ;
 wire \u_multiplier/STAGE1/_0848_ ;
 wire \u_multiplier/STAGE1/_0849_ ;
 wire \u_multiplier/STAGE1/_0850_ ;
 wire \u_multiplier/STAGE1/_0851_ ;
 wire \u_multiplier/STAGE1/_0852_ ;
 wire \u_multiplier/STAGE1/_0853_ ;
 wire \u_multiplier/STAGE1/_0854_ ;
 wire \u_multiplier/STAGE1/_0855_ ;
 wire \u_multiplier/STAGE1/_0856_ ;
 wire \u_multiplier/STAGE1/_0857_ ;
 wire \u_multiplier/STAGE1/_0858_ ;
 wire \u_multiplier/STAGE1/_0859_ ;
 wire \u_multiplier/STAGE1/_0860_ ;
 wire \u_multiplier/STAGE1/_0861_ ;
 wire \u_multiplier/STAGE1/_0862_ ;
 wire \u_multiplier/STAGE1/_0863_ ;
 wire \u_multiplier/STAGE1/_0864_ ;
 wire \u_multiplier/STAGE1/_0865_ ;
 wire \u_multiplier/STAGE1/_0866_ ;
 wire \u_multiplier/STAGE1/_0867_ ;
 wire \u_multiplier/STAGE1/_0868_ ;
 wire \u_multiplier/STAGE1/_0869_ ;
 wire \u_multiplier/STAGE1/_0870_ ;
 wire \u_multiplier/STAGE1/_0871_ ;
 wire \u_multiplier/STAGE1/_0872_ ;
 wire \u_multiplier/STAGE1/_0873_ ;
 wire \u_multiplier/STAGE1/_0874_ ;
 wire \u_multiplier/STAGE1/_0875_ ;
 wire \u_multiplier/STAGE1/_0876_ ;
 wire \u_multiplier/STAGE1/_0877_ ;
 wire \u_multiplier/STAGE1/_0878_ ;
 wire \u_multiplier/STAGE1/_0879_ ;
 wire \u_multiplier/STAGE1/_0880_ ;
 wire \u_multiplier/STAGE1/_0881_ ;
 wire \u_multiplier/STAGE1/_0882_ ;
 wire \u_multiplier/STAGE1/_0883_ ;
 wire \u_multiplier/STAGE1/_0884_ ;
 wire \u_multiplier/STAGE1/_0885_ ;
 wire \u_multiplier/STAGE1/_0886_ ;
 wire \u_multiplier/STAGE1/_0887_ ;
 wire \u_multiplier/STAGE1/_0888_ ;
 wire \u_multiplier/STAGE1/_0889_ ;
 wire \u_multiplier/STAGE1/_0890_ ;
 wire \u_multiplier/STAGE1/_0891_ ;
 wire \u_multiplier/STAGE1/_0892_ ;
 wire \u_multiplier/STAGE1/_0893_ ;
 wire \u_multiplier/STAGE1/_0894_ ;
 wire \u_multiplier/STAGE1/_0895_ ;
 wire \u_multiplier/STAGE1/_0896_ ;
 wire \u_multiplier/STAGE1/_0897_ ;
 wire \u_multiplier/STAGE1/_0898_ ;
 wire \u_multiplier/STAGE1/_0899_ ;
 wire \u_multiplier/STAGE1/_0900_ ;
 wire \u_multiplier/STAGE1/_0901_ ;
 wire \u_multiplier/STAGE1/_0902_ ;
 wire \u_multiplier/STAGE1/_0903_ ;
 wire \u_multiplier/STAGE1/_0904_ ;
 wire \u_multiplier/STAGE1/_0905_ ;
 wire \u_multiplier/STAGE1/_0906_ ;
 wire \u_multiplier/STAGE1/_0907_ ;
 wire \u_multiplier/STAGE1/_0908_ ;
 wire \u_multiplier/STAGE1/_0909_ ;
 wire \u_multiplier/STAGE1/_0910_ ;
 wire \u_multiplier/STAGE1/_0911_ ;
 wire \u_multiplier/STAGE1/_0912_ ;
 wire \u_multiplier/STAGE1/_0913_ ;
 wire \u_multiplier/STAGE1/_0914_ ;
 wire \u_multiplier/STAGE1/_0915_ ;
 wire \u_multiplier/STAGE1/_0916_ ;
 wire \u_multiplier/STAGE1/_0917_ ;
 wire \u_multiplier/STAGE1/_0918_ ;
 wire \u_multiplier/STAGE1/_0919_ ;
 wire \u_multiplier/STAGE1/_0920_ ;
 wire \u_multiplier/STAGE1/_0921_ ;
 wire \u_multiplier/STAGE1/_0922_ ;
 wire \u_multiplier/STAGE1/_0923_ ;
 wire \u_multiplier/STAGE1/_0924_ ;
 wire \u_multiplier/STAGE1/_0925_ ;
 wire \u_multiplier/STAGE1/_0926_ ;
 wire \u_multiplier/STAGE1/_0927_ ;
 wire \u_multiplier/STAGE1/_0928_ ;
 wire \u_multiplier/STAGE1/_0929_ ;
 wire \u_multiplier/STAGE1/_0930_ ;
 wire \u_multiplier/STAGE1/_0931_ ;
 wire \u_multiplier/STAGE1/_0932_ ;
 wire \u_multiplier/STAGE1/_0933_ ;
 wire \u_multiplier/STAGE1/_0934_ ;
 wire \u_multiplier/STAGE1/_0935_ ;
 wire \u_multiplier/STAGE1/_0936_ ;
 wire \u_multiplier/STAGE1/_0937_ ;
 wire \u_multiplier/STAGE1/_0938_ ;
 wire \u_multiplier/STAGE1/_0939_ ;
 wire \u_multiplier/STAGE1/_0940_ ;
 wire \u_multiplier/STAGE1/_0941_ ;
 wire \u_multiplier/STAGE1/_0942_ ;
 wire \u_multiplier/STAGE1/_0943_ ;
 wire \u_multiplier/STAGE1/_0944_ ;
 wire \u_multiplier/STAGE1/_0945_ ;
 wire \u_multiplier/STAGE1/_0946_ ;
 wire \u_multiplier/STAGE1/_0947_ ;
 wire \u_multiplier/STAGE1/_0948_ ;
 wire \u_multiplier/STAGE1/_0949_ ;
 wire \u_multiplier/STAGE1/_0950_ ;
 wire \u_multiplier/STAGE1/_0951_ ;
 wire \u_multiplier/STAGE1/_0952_ ;
 wire \u_multiplier/STAGE1/_0953_ ;
 wire \u_multiplier/STAGE1/_0954_ ;
 wire \u_multiplier/STAGE1/_0955_ ;
 wire \u_multiplier/STAGE1/_0956_ ;
 wire \u_multiplier/STAGE1/_0957_ ;
 wire \u_multiplier/STAGE1/_0958_ ;
 wire \u_multiplier/STAGE1/_0959_ ;
 wire \u_multiplier/STAGE1/_0960_ ;
 wire \u_multiplier/STAGE1/_0961_ ;
 wire \u_multiplier/STAGE1/_0962_ ;
 wire \u_multiplier/STAGE1/_0963_ ;
 wire \u_multiplier/STAGE1/_0964_ ;
 wire \u_multiplier/STAGE1/_0965_ ;
 wire \u_multiplier/STAGE1/_0966_ ;
 wire \u_multiplier/STAGE1/_0967_ ;
 wire \u_multiplier/STAGE1/_0968_ ;
 wire \u_multiplier/STAGE1/_0969_ ;
 wire \u_multiplier/STAGE1/_0970_ ;
 wire \u_multiplier/STAGE1/_0971_ ;
 wire \u_multiplier/STAGE1/_0972_ ;
 wire \u_multiplier/STAGE1/_0973_ ;
 wire \u_multiplier/STAGE1/_0974_ ;
 wire \u_multiplier/STAGE1/_0975_ ;
 wire \u_multiplier/STAGE1/_0976_ ;
 wire \u_multiplier/STAGE1/_0977_ ;
 wire \u_multiplier/STAGE1/_0978_ ;
 wire \u_multiplier/STAGE1/_0979_ ;
 wire \u_multiplier/STAGE1/_0980_ ;
 wire \u_multiplier/STAGE1/_0981_ ;
 wire \u_multiplier/STAGE1/_0982_ ;
 wire \u_multiplier/STAGE1/_0983_ ;
 wire \u_multiplier/STAGE1/_0984_ ;
 wire \u_multiplier/STAGE1/_0985_ ;
 wire \u_multiplier/STAGE1/_0986_ ;
 wire \u_multiplier/STAGE1/_0987_ ;
 wire \u_multiplier/STAGE1/_0988_ ;
 wire \u_multiplier/STAGE1/_0989_ ;
 wire \u_multiplier/STAGE1/_0990_ ;
 wire \u_multiplier/STAGE1/_0991_ ;
 wire \u_multiplier/STAGE1/_0992_ ;
 wire \u_multiplier/STAGE1/_0993_ ;
 wire \u_multiplier/STAGE1/_0994_ ;
 wire \u_multiplier/STAGE1/_0995_ ;
 wire \u_multiplier/STAGE1/_0996_ ;
 wire \u_multiplier/STAGE1/_0997_ ;
 wire \u_multiplier/STAGE1/_0998_ ;
 wire \u_multiplier/STAGE1/_0999_ ;
 wire \u_multiplier/STAGE1/_1000_ ;
 wire \u_multiplier/STAGE1/_1001_ ;
 wire \u_multiplier/STAGE1/_1002_ ;
 wire \u_multiplier/STAGE1/_1003_ ;
 wire \u_multiplier/STAGE1/_1004_ ;
 wire \u_multiplier/STAGE1/_1005_ ;
 wire \u_multiplier/STAGE1/_1006_ ;
 wire \u_multiplier/STAGE1/_1007_ ;
 wire \u_multiplier/STAGE1/_1008_ ;
 wire \u_multiplier/STAGE1/_1009_ ;
 wire \u_multiplier/STAGE1/_1010_ ;
 wire \u_multiplier/STAGE1/_1011_ ;
 wire \u_multiplier/STAGE1/_1012_ ;
 wire \u_multiplier/STAGE1/_1013_ ;
 wire \u_multiplier/STAGE1/_1014_ ;
 wire \u_multiplier/STAGE1/_1015_ ;
 wire \u_multiplier/STAGE1/_1016_ ;
 wire \u_multiplier/STAGE1/_1017_ ;
 wire \u_multiplier/STAGE1/_1018_ ;
 wire \u_multiplier/STAGE1/_1019_ ;
 wire \u_multiplier/STAGE1/_1020_ ;
 wire \u_multiplier/STAGE1/_1021_ ;
 wire \u_multiplier/STAGE1/_1022_ ;
 wire \u_multiplier/STAGE1/_1023_ ;
 wire \u_multiplier/STAGE1/_1024_ ;
 wire \u_multiplier/STAGE1/_1025_ ;
 wire \u_multiplier/STAGE1/_1026_ ;
 wire \u_multiplier/STAGE1/_1027_ ;
 wire \u_multiplier/STAGE1/_1028_ ;
 wire \u_multiplier/STAGE1/_1029_ ;
 wire \u_multiplier/STAGE1/_1030_ ;
 wire \u_multiplier/STAGE1/_1031_ ;
 wire \u_multiplier/STAGE1/_1032_ ;
 wire \u_multiplier/STAGE1/_1033_ ;
 wire \u_multiplier/STAGE1/_1034_ ;
 wire \u_multiplier/STAGE1/_1035_ ;
 wire \u_multiplier/STAGE1/_1036_ ;
 wire \u_multiplier/STAGE1/_1037_ ;
 wire \u_multiplier/STAGE1/_1038_ ;
 wire \u_multiplier/STAGE1/_1039_ ;
 wire \u_multiplier/STAGE1/_1040_ ;
 wire \u_multiplier/STAGE1/_1041_ ;
 wire \u_multiplier/STAGE1/_1042_ ;
 wire \u_multiplier/STAGE1/_1043_ ;
 wire \u_multiplier/STAGE1/_1044_ ;
 wire \u_multiplier/STAGE1/_1045_ ;
 wire \u_multiplier/STAGE1/_1046_ ;
 wire \u_multiplier/STAGE1/_1047_ ;
 wire \u_multiplier/STAGE1/_1048_ ;
 wire \u_multiplier/STAGE1/_1049_ ;
 wire \u_multiplier/STAGE1/_1050_ ;
 wire \u_multiplier/STAGE1/_1051_ ;
 wire \u_multiplier/STAGE1/_1052_ ;
 wire \u_multiplier/STAGE1/_1053_ ;
 wire \u_multiplier/STAGE1/_1054_ ;
 wire \u_multiplier/STAGE1/_1055_ ;
 wire \u_multiplier/STAGE1/_1056_ ;
 wire \u_multiplier/STAGE1/_1057_ ;
 wire \u_multiplier/STAGE1/_1058_ ;
 wire \u_multiplier/STAGE1/_1059_ ;
 wire \u_multiplier/STAGE1/_1060_ ;
 wire \u_multiplier/STAGE1/_1061_ ;
 wire \u_multiplier/STAGE1/_1062_ ;
 wire \u_multiplier/STAGE1/_1063_ ;
 wire \u_multiplier/STAGE1/_1064_ ;
 wire \u_multiplier/STAGE1/_1065_ ;
 wire \u_multiplier/STAGE1/_1066_ ;
 wire \u_multiplier/STAGE1/_1067_ ;
 wire \u_multiplier/STAGE1/_1068_ ;
 wire \u_multiplier/STAGE1/_1069_ ;
 wire \u_multiplier/STAGE1/_1070_ ;
 wire \u_multiplier/STAGE1/_1071_ ;
 wire \u_multiplier/STAGE1/_1072_ ;
 wire \u_multiplier/STAGE1/_1073_ ;
 wire \u_multiplier/STAGE1/_1074_ ;
 wire \u_multiplier/STAGE1/_1075_ ;
 wire \u_multiplier/STAGE1/_1076_ ;
 wire \u_multiplier/STAGE1/_1077_ ;
 wire \u_multiplier/STAGE1/_1078_ ;
 wire \u_multiplier/STAGE1/_1079_ ;
 wire \u_multiplier/STAGE1/_1080_ ;
 wire \u_multiplier/STAGE1/_1081_ ;
 wire \u_multiplier/STAGE1/_1082_ ;
 wire \u_multiplier/STAGE1/_1083_ ;
 wire \u_multiplier/STAGE1/_1084_ ;
 wire \u_multiplier/STAGE1/_1085_ ;
 wire \u_multiplier/STAGE1/_1086_ ;
 wire \u_multiplier/STAGE1/_1087_ ;
 wire \u_multiplier/STAGE1/_1088_ ;
 wire \u_multiplier/STAGE1/_1089_ ;
 wire \u_multiplier/STAGE1/_1090_ ;
 wire \u_multiplier/STAGE1/_1091_ ;
 wire \u_multiplier/STAGE1/_1092_ ;
 wire \u_multiplier/STAGE1/_1093_ ;
 wire \u_multiplier/STAGE1/_1094_ ;
 wire \u_multiplier/STAGE1/_1095_ ;
 wire \u_multiplier/STAGE1/_1096_ ;
 wire \u_multiplier/STAGE1/_1097_ ;
 wire \u_multiplier/STAGE1/_1098_ ;
 wire \u_multiplier/STAGE1/_1099_ ;
 wire \u_multiplier/STAGE1/_1100_ ;
 wire \u_multiplier/STAGE1/_1101_ ;
 wire \u_multiplier/STAGE1/_1102_ ;
 wire \u_multiplier/STAGE1/_1103_ ;
 wire \u_multiplier/STAGE1/_1104_ ;
 wire \u_multiplier/STAGE1/_1105_ ;
 wire \u_multiplier/STAGE1/_1106_ ;
 wire \u_multiplier/STAGE1/_1107_ ;
 wire \u_multiplier/STAGE1/_1108_ ;
 wire \u_multiplier/STAGE1/_1109_ ;
 wire \u_multiplier/STAGE1/_1110_ ;
 wire \u_multiplier/STAGE1/_1111_ ;
 wire \u_multiplier/STAGE1/_1112_ ;
 wire \u_multiplier/STAGE1/_1113_ ;
 wire \u_multiplier/STAGE1/_1114_ ;
 wire \u_multiplier/STAGE1/_1115_ ;
 wire \u_multiplier/STAGE1/_1116_ ;
 wire \u_multiplier/STAGE1/_1117_ ;
 wire \u_multiplier/STAGE1/_1118_ ;
 wire \u_multiplier/STAGE1/_1119_ ;
 wire \u_multiplier/STAGE1/_1120_ ;
 wire \u_multiplier/STAGE1/_1121_ ;
 wire \u_multiplier/STAGE1/_1122_ ;
 wire \u_multiplier/STAGE1/_1123_ ;
 wire \u_multiplier/STAGE1/_1124_ ;
 wire \u_multiplier/STAGE1/_1125_ ;
 wire \u_multiplier/STAGE1/_1126_ ;
 wire \u_multiplier/STAGE1/_1127_ ;
 wire \u_multiplier/STAGE1/_1128_ ;
 wire \u_multiplier/STAGE1/_1129_ ;
 wire \u_multiplier/STAGE1/_1130_ ;
 wire \u_multiplier/STAGE1/_1131_ ;
 wire \u_multiplier/STAGE1/_1132_ ;
 wire \u_multiplier/STAGE1/_1133_ ;
 wire \u_multiplier/STAGE1/_1134_ ;
 wire \u_multiplier/STAGE1/_1135_ ;
 wire \u_multiplier/STAGE1/_1136_ ;
 wire \u_multiplier/STAGE1/_1137_ ;
 wire \u_multiplier/STAGE1/_1138_ ;
 wire \u_multiplier/STAGE1/_1139_ ;
 wire \u_multiplier/STAGE1/_1140_ ;
 wire \u_multiplier/STAGE1/_1141_ ;
 wire \u_multiplier/STAGE1/_1142_ ;
 wire \u_multiplier/STAGE1/_1143_ ;
 wire \u_multiplier/STAGE1/_1144_ ;
 wire \u_multiplier/STAGE1/_1145_ ;
 wire \u_multiplier/STAGE1/_1146_ ;
 wire \u_multiplier/STAGE1/_1147_ ;
 wire \u_multiplier/STAGE1/_1148_ ;
 wire \u_multiplier/STAGE1/_1149_ ;
 wire net133;
 wire \u_multiplier/STAGE1/pp1_17_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_18_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_19_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_19_e42_2_cout ;
 wire \u_multiplier/STAGE1/pp1_20_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_20_e42_2_cout ;
 wire \u_multiplier/STAGE1/pp1_21_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_21_e42_2_cout ;
 wire \u_multiplier/STAGE1/pp1_21_e42_3_cout ;
 wire \u_multiplier/STAGE1/pp1_22_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_22_e42_2_cout ;
 wire \u_multiplier/STAGE1/pp1_22_e42_3_cout ;
 wire \u_multiplier/STAGE1/pp1_23_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_23_e42_2_cout ;
 wire \u_multiplier/STAGE1/pp1_23_e42_3_cout ;
 wire \u_multiplier/STAGE1/pp1_23_e42_4_cout ;
 wire \u_multiplier/STAGE1/pp1_24_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_24_e42_2_cout ;
 wire \u_multiplier/STAGE1/pp1_24_e42_3_cout ;
 wire \u_multiplier/STAGE1/pp1_24_e42_4_cout ;
 wire \u_multiplier/STAGE1/pp1_25_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_25_e42_2_cout ;
 wire \u_multiplier/STAGE1/pp1_25_e42_3_cout ;
 wire \u_multiplier/STAGE1/pp1_25_e42_4_cout ;
 wire \u_multiplier/STAGE1/pp1_25_e42_5_cout ;
 wire \u_multiplier/STAGE1/pp1_26_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_26_e42_2_cout ;
 wire \u_multiplier/STAGE1/pp1_26_e42_3_cout ;
 wire \u_multiplier/STAGE1/pp1_26_e42_4_cout ;
 wire \u_multiplier/STAGE1/pp1_26_e42_5_cout ;
 wire \u_multiplier/STAGE1/pp1_27_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_27_e42_2_cout ;
 wire \u_multiplier/STAGE1/pp1_27_e42_3_cout ;
 wire \u_multiplier/STAGE1/pp1_27_e42_4_cout ;
 wire \u_multiplier/STAGE1/pp1_27_e42_5_cout ;
 wire \u_multiplier/STAGE1/pp1_27_e42_6_cout ;
 wire \u_multiplier/STAGE1/pp1_28_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_28_e42_2_cout ;
 wire \u_multiplier/STAGE1/pp1_28_e42_3_cout ;
 wire \u_multiplier/STAGE1/pp1_28_e42_4_cout ;
 wire \u_multiplier/STAGE1/pp1_28_e42_5_cout ;
 wire \u_multiplier/STAGE1/pp1_28_e42_6_cout ;
 wire \u_multiplier/STAGE1/pp1_29_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_29_e42_2_cout ;
 wire \u_multiplier/STAGE1/pp1_29_e42_3_cout ;
 wire \u_multiplier/STAGE1/pp1_29_e42_4_cout ;
 wire \u_multiplier/STAGE1/pp1_29_e42_5_cout ;
 wire \u_multiplier/STAGE1/pp1_29_e42_6_cout ;
 wire \u_multiplier/STAGE1/pp1_29_e42_7_cout ;
 wire \u_multiplier/STAGE1/pp1_30_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_30_e42_2_cout ;
 wire \u_multiplier/STAGE1/pp1_30_e42_3_cout ;
 wire \u_multiplier/STAGE1/pp1_30_e42_4_cout ;
 wire \u_multiplier/STAGE1/pp1_30_e42_5_cout ;
 wire \u_multiplier/STAGE1/pp1_30_e42_6_cout ;
 wire \u_multiplier/STAGE1/pp1_30_e42_7_cout ;
 wire \u_multiplier/STAGE1/pp1_31_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_31_e42_2_cout ;
 wire \u_multiplier/STAGE1/pp1_31_e42_3_cout ;
 wire \u_multiplier/STAGE1/pp1_31_e42_4_cout ;
 wire \u_multiplier/STAGE1/pp1_31_e42_5_cout ;
 wire \u_multiplier/STAGE1/pp1_31_e42_6_cout ;
 wire \u_multiplier/STAGE1/pp1_31_e42_7_cout ;
 wire \u_multiplier/STAGE1/pp1_31_e42_8_cout ;
 wire \u_multiplier/STAGE1/pp1_32_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_32_e42_2_cout ;
 wire \u_multiplier/STAGE1/pp1_32_e42_3_cout ;
 wire \u_multiplier/STAGE1/pp1_32_e42_4_cout ;
 wire \u_multiplier/STAGE1/pp1_32_e42_5_cout ;
 wire \u_multiplier/STAGE1/pp1_32_e42_6_cout ;
 wire \u_multiplier/STAGE1/pp1_32_e42_7_cout ;
 wire \u_multiplier/STAGE1/pp1_32_e42_8_cout ;
 wire \u_multiplier/STAGE1/pp1_33_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_33_e42_2_cout ;
 wire \u_multiplier/STAGE1/pp1_33_e42_3_cout ;
 wire \u_multiplier/STAGE1/pp1_33_e42_4_cout ;
 wire \u_multiplier/STAGE1/pp1_33_e42_5_cout ;
 wire \u_multiplier/STAGE1/pp1_33_e42_6_cout ;
 wire \u_multiplier/STAGE1/pp1_33_e42_7_cout ;
 wire \u_multiplier/STAGE1/pp1_34_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_34_e42_2_cout ;
 wire \u_multiplier/STAGE1/pp1_34_e42_3_cout ;
 wire \u_multiplier/STAGE1/pp1_34_e42_4_cout ;
 wire \u_multiplier/STAGE1/pp1_34_e42_5_cout ;
 wire \u_multiplier/STAGE1/pp1_34_e42_6_cout ;
 wire \u_multiplier/STAGE1/pp1_34_e42_7_cout ;
 wire \u_multiplier/STAGE1/pp1_35_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_35_e42_2_cout ;
 wire \u_multiplier/STAGE1/pp1_35_e42_3_cout ;
 wire \u_multiplier/STAGE1/pp1_35_e42_4_cout ;
 wire \u_multiplier/STAGE1/pp1_35_e42_5_cout ;
 wire \u_multiplier/STAGE1/pp1_35_e42_6_cout ;
 wire \u_multiplier/STAGE1/pp1_36_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_36_e42_2_cout ;
 wire \u_multiplier/STAGE1/pp1_36_e42_3_cout ;
 wire \u_multiplier/STAGE1/pp1_36_e42_4_cout ;
 wire \u_multiplier/STAGE1/pp1_36_e42_5_cout ;
 wire \u_multiplier/STAGE1/pp1_36_e42_6_cout ;
 wire \u_multiplier/STAGE1/pp1_37_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_37_e42_2_cout ;
 wire \u_multiplier/STAGE1/pp1_37_e42_3_cout ;
 wire \u_multiplier/STAGE1/pp1_37_e42_4_cout ;
 wire \u_multiplier/STAGE1/pp1_37_e42_5_cout ;
 wire \u_multiplier/STAGE1/pp1_38_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_38_e42_2_cout ;
 wire \u_multiplier/STAGE1/pp1_38_e42_3_cout ;
 wire \u_multiplier/STAGE1/pp1_38_e42_4_cout ;
 wire \u_multiplier/STAGE1/pp1_38_e42_5_cout ;
 wire \u_multiplier/STAGE1/pp1_39_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_39_e42_2_cout ;
 wire \u_multiplier/STAGE1/pp1_39_e42_3_cout ;
 wire \u_multiplier/STAGE1/pp1_39_e42_4_cout ;
 wire \u_multiplier/STAGE1/pp1_40_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_40_e42_2_cout ;
 wire \u_multiplier/STAGE1/pp1_40_e42_3_cout ;
 wire \u_multiplier/STAGE1/pp1_40_e42_4_cout ;
 wire \u_multiplier/STAGE1/pp1_41_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_41_e42_2_cout ;
 wire \u_multiplier/STAGE1/pp1_41_e42_3_cout ;
 wire \u_multiplier/STAGE1/pp1_42_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_42_e42_2_cout ;
 wire \u_multiplier/STAGE1/pp1_42_e42_3_cout ;
 wire \u_multiplier/STAGE1/pp1_43_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_43_e42_2_cout ;
 wire \u_multiplier/STAGE1/pp1_44_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_44_e42_2_cout ;
 wire \u_multiplier/STAGE1/pp1_45_e42_1_cout ;
 wire \u_multiplier/STAGE1/pp1_46_e42_1_cout ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_17_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_18_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_19_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_20_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_21_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_22_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_4/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_4/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_4/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_4/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_4/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_4/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_23_4/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_4/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_4/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_4/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_4/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_4/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_4/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_24_4/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_4/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_4/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_4/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_4/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_4/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_4/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_4/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_5/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_5/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_5/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_5/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_5/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_5/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_25_5/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_4/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_4/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_4/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_4/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_4/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_4/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_4/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_5/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_5/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_5/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_5/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_5/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_5/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_26_5/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_4/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_4/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_4/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_4/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_4/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_4/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_4/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_5/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_5/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_5/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_5/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_5/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_5/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_5/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_6/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_6/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_6/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_6/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_6/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_6/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_27_6/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_4/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_4/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_4/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_4/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_4/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_4/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_4/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_5/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_5/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_5/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_5/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_5/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_5/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_5/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_6/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_6/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_6/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_6/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_6/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_6/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_28_6/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_4/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_4/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_4/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_4/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_4/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_4/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_4/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_5/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_5/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_5/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_5/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_5/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_5/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_5/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_6/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_6/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_6/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_6/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_6/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_6/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_6/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_7/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_7/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_7/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_7/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_7/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_7/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_29_7/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_4/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_4/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_4/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_4/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_4/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_4/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_4/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_5/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_5/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_5/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_5/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_5/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_5/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_5/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_6/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_6/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_6/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_6/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_6/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_6/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_6/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_7/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_7/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_7/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_7/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_7/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_7/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_30_7/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_4/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_4/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_4/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_4/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_4/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_4/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_4/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_5/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_5/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_5/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_5/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_5/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_5/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_5/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_6/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_6/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_6/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_6/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_6/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_6/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_6/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_7/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_7/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_7/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_7/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_7/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_7/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_7/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_8/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_8/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_8/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_8/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_8/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_8/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_31_8/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_4/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_4/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_4/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_4/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_4/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_4/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_4/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_5/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_5/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_5/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_5/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_5/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_5/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_5/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_6/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_6/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_6/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_6/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_6/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_6/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_6/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_7/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_7/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_7/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_7/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_7/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_7/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_7/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_8/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_8/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_8/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_8/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_8/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_8/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_32_8/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_4/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_4/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_4/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_4/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_4/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_4/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_4/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_5/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_5/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_5/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_5/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_5/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_5/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_5/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_6/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_6/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_6/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_6/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_6/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_6/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_6/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_7/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_7/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_7/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_7/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_7/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_7/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_33_7/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_4/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_4/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_4/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_4/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_4/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_4/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_4/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_5/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_5/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_5/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_5/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_5/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_5/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_5/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_6/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_6/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_6/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_6/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_6/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_6/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_6/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_7/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_7/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_7/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_7/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_7/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_7/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_34_7/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_4/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_4/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_4/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_4/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_4/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_4/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_4/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_5/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_5/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_5/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_5/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_5/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_5/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_5/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_6/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_6/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_6/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_6/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_6/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_6/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_35_6/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_4/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_4/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_4/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_4/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_4/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_4/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_4/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_5/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_5/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_5/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_5/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_5/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_5/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_5/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_6/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_6/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_6/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_6/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_6/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_6/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_36_6/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_4/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_4/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_4/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_4/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_4/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_4/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_4/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_5/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_5/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_5/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_5/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_5/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_5/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_37_5/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_4/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_4/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_4/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_4/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_4/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_4/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_4/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_5/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_5/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_5/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_5/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_5/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_5/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_38_5/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_4/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_4/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_4/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_4/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_4/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_4/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_39_4/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_4/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_4/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_4/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_4/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_4/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_4/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_40_4/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_41_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_41_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_41_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_41_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_41_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_41_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_41_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_41_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_41_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_41_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_41_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_41_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_41_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_41_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_41_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_41_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_41_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_41_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_41_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_41_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_41_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_42_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_42_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_42_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_42_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_42_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_42_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_42_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_42_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_42_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_42_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_42_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_42_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_42_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_42_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_42_3/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_42_3/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_42_3/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_42_3/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_42_3/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_42_3/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_42_3/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_43_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_43_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_43_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_43_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_43_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_43_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_43_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_43_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_43_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_43_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_43_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_43_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_43_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_43_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_44_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_44_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_44_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_44_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_44_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_44_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_44_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_44_2/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_44_2/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_44_2/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_44_2/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_44_2/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_44_2/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_44_2/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_45_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_45_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_45_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_45_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_45_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_45_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_45_1/_17_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_46_1/_11_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_46_1/_12_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_46_1/_13_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_46_1/_14_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_46_1/_15_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_46_1/_16_ ;
 wire \u_multiplier/STAGE1/E_4_2_pp_46_1/_17_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_33_1/_08_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_33_1/_09_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_33_1/_10_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_33_1/_11_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_35_1/_08_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_35_1/_09_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_35_1/_10_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_35_1/_11_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_37_1/_08_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_37_1/_09_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_37_1/_10_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_37_1/_11_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_39_1/_08_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_39_1/_09_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_39_1/_10_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_39_1/_11_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_41_1/_08_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_41_1/_09_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_41_1/_10_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_41_1/_11_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_43_1/_08_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_43_1/_09_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_43_1/_10_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_43_1/_11_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_45_1/_08_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_45_1/_09_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_45_1/_10_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_45_1/_11_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_47_1/_08_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_47_1/_09_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_47_1/_10_ ;
 wire \u_multiplier/STAGE1/Full_adder_pp_47_1/_11_ ;
 wire \u_multiplier/STAGE2/pp2_10_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_11_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_11_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_12_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_12_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_13_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_13_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_13_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_14_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_14_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_14_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_15_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_15_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_15_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_15_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_16_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_16_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_16_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_16_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_17_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_17_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_17_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_17_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_18_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_18_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_18_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_18_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_19_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_19_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_19_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_19_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_20_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_20_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_20_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_20_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_21_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_21_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_21_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_21_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_22_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_22_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_22_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_22_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_23_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_23_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_23_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_23_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_24_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_24_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_24_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_24_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_25_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_25_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_25_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_25_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_26_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_26_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_26_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_26_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_27_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_27_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_27_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_27_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_28_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_28_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_28_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_28_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_29_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_29_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_29_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_29_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_30_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_30_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_30_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_30_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_31_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_31_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_31_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_31_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_32_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_32_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_32_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_32_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_33_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_33_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_33_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_33_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_34_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_34_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_34_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_34_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_35_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_35_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_35_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_35_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_36_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_36_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_36_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_36_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_37_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_37_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_37_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_37_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_38_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_38_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_38_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_38_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_39_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_39_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_39_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_39_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_40_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_40_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_40_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_40_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_41_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_41_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_41_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_41_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_42_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_42_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_42_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_42_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_43_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_43_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_43_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_43_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_44_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_44_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_44_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_44_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_45_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_45_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_45_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_45_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_46_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_46_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_46_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_46_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_47_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_47_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_47_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_47_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_48_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_48_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_48_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_48_e42_4_cout ;
 wire \u_multiplier/STAGE2/pp2_49_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_49_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_49_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_50_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_50_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_50_e42_3_cout ;
 wire \u_multiplier/STAGE2/pp2_51_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_51_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_52_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_52_e42_2_cout ;
 wire \u_multiplier/STAGE2/pp2_53_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_54_e42_1_cout ;
 wire \u_multiplier/STAGE2/pp2_9_e42_1_cout ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_10_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_10_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_10_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_10_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_10_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_10_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_10_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_11_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_11_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_11_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_11_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_11_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_11_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_11_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_11_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_11_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_11_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_11_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_11_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_11_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_11_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_12_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_12_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_12_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_12_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_12_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_12_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_12_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_12_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_12_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_12_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_12_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_12_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_12_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_12_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_13_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_13_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_13_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_13_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_13_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_13_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_13_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_13_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_13_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_13_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_13_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_13_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_13_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_13_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_13_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_13_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_13_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_13_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_13_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_13_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_13_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_14_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_14_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_14_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_14_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_14_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_14_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_14_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_14_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_14_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_14_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_14_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_14_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_14_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_14_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_14_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_14_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_14_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_14_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_14_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_14_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_14_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_15_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_16_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_17_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_18_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_19_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_20_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_21_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_22_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_23_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_24_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_25_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_26_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_27_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_28_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_29_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_30_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_31_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_32_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_33_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_34_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_35_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_36_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_37_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_38_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_39_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_40_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_41_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_42_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_43_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_44_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_45_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_46_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_47_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_4/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_4/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_4/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_4/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_4/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_4/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_48_4/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_49_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_49_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_49_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_49_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_49_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_49_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_49_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_49_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_49_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_49_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_49_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_49_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_49_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_49_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_49_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_49_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_49_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_49_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_49_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_49_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_49_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_50_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_50_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_50_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_50_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_50_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_50_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_50_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_50_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_50_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_50_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_50_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_50_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_50_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_50_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_50_3/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_50_3/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_50_3/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_50_3/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_50_3/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_50_3/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_50_3/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_51_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_51_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_51_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_51_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_51_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_51_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_51_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_51_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_51_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_51_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_51_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_51_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_51_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_51_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_52_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_52_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_52_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_52_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_52_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_52_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_52_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_52_2/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_52_2/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_52_2/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_52_2/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_52_2/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_52_2/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_52_2/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_53_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_53_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_53_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_53_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_53_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_53_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_53_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_54_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_54_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_54_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_54_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_54_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_54_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_54_1/_17_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_9_1/_11_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_9_1/_12_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_9_1/_13_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_9_1/_14_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_9_1/_15_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_9_1/_16_ ;
 wire \u_multiplier/STAGE2/E_4_2_pp2_9_1/_17_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp2_49_1/_08_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp2_49_1/_09_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp2_49_1/_10_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp2_49_1/_11_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp2_51_1/_08_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp2_51_1/_09_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp2_51_1/_10_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp2_51_1/_11_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp2_53_1/_08_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp2_53_1/_09_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp2_53_1/_10_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp2_53_1/_11_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp2_55_1/_08_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp2_55_1/_09_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp2_55_1/_10_ ;
 wire \u_multiplier/STAGE2/Full_adder_pp2_55_1/_11_ ;
 wire \u_multiplier/STAGE3/pp3_10_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_10_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_11_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_11_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_12_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_12_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_13_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_13_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_14_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_14_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_15_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_15_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_16_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_16_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_17_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_17_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_18_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_18_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_19_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_19_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_20_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_20_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_21_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_21_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_22_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_22_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_23_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_23_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_24_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_24_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_25_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_25_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_26_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_26_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_27_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_27_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_28_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_28_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_29_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_29_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_30_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_30_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_31_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_31_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_32_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_32_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_33_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_33_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_34_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_34_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_35_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_35_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_36_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_36_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_37_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_37_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_38_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_38_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_39_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_39_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_40_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_40_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_41_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_41_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_42_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_42_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_43_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_43_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_44_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_44_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_45_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_45_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_46_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_46_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_47_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_47_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_48_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_48_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_49_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_49_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_50_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_50_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_51_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_51_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_52_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_52_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_53_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_53_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_54_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_54_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_55_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_55_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_56_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_56_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_57_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_58_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_5_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_6_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_7_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_7_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_8_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_8_e42_2_cout ;
 wire \u_multiplier/STAGE3/pp3_9_e42_1_cout ;
 wire \u_multiplier/STAGE3/pp3_9_e42_2_cout ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_10_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_10_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_10_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_10_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_10_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_10_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_10_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_10_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_10_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_10_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_10_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_10_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_10_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_10_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_11_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_11_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_11_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_11_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_11_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_11_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_11_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_11_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_11_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_11_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_11_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_11_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_11_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_11_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_12_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_12_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_12_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_12_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_12_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_12_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_12_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_12_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_12_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_12_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_12_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_12_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_12_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_12_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_13_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_13_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_13_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_13_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_13_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_13_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_13_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_13_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_13_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_13_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_13_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_13_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_13_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_13_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_14_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_14_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_14_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_14_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_14_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_14_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_14_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_14_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_14_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_14_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_14_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_14_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_14_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_14_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_15_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_15_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_15_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_15_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_15_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_15_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_15_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_15_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_15_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_15_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_15_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_15_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_15_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_15_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_16_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_16_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_16_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_16_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_16_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_16_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_16_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_16_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_16_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_16_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_16_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_16_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_16_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_16_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_17_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_17_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_17_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_17_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_17_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_17_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_17_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_17_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_17_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_17_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_17_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_17_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_17_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_17_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_18_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_18_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_18_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_18_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_18_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_18_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_18_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_18_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_18_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_18_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_18_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_18_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_18_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_18_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_19_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_19_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_19_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_19_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_19_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_19_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_19_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_19_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_19_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_19_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_19_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_19_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_19_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_19_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_20_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_20_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_20_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_20_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_20_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_20_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_20_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_20_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_20_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_20_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_20_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_20_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_20_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_20_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_21_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_21_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_21_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_21_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_21_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_21_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_21_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_21_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_21_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_21_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_21_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_21_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_21_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_21_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_22_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_22_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_22_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_22_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_22_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_22_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_22_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_22_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_22_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_22_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_22_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_22_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_22_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_22_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_23_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_23_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_23_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_23_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_23_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_23_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_23_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_23_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_23_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_23_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_23_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_23_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_23_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_23_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_24_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_24_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_24_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_24_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_24_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_24_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_24_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_24_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_24_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_24_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_24_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_24_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_24_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_24_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_25_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_25_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_25_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_25_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_25_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_25_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_25_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_25_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_25_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_25_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_25_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_25_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_25_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_25_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_26_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_26_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_26_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_26_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_26_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_26_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_26_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_26_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_26_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_26_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_26_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_26_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_26_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_26_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_27_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_27_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_27_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_27_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_27_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_27_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_27_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_27_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_27_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_27_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_27_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_27_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_27_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_27_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_28_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_28_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_28_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_28_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_28_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_28_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_28_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_28_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_28_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_28_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_28_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_28_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_28_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_28_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_29_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_29_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_29_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_29_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_29_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_29_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_29_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_29_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_29_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_29_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_29_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_29_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_29_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_29_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_30_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_30_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_30_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_30_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_30_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_30_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_30_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_30_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_30_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_30_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_30_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_30_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_30_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_30_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_31_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_31_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_31_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_31_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_31_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_31_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_31_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_31_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_31_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_31_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_31_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_31_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_31_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_31_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_32_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_32_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_32_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_32_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_32_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_32_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_32_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_32_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_32_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_32_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_32_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_32_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_32_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_32_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_33_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_33_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_33_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_33_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_33_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_33_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_33_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_33_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_33_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_33_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_33_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_33_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_33_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_33_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_34_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_34_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_34_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_34_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_34_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_34_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_34_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_34_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_34_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_34_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_34_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_34_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_34_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_34_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_35_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_35_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_35_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_35_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_35_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_35_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_35_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_35_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_35_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_35_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_35_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_35_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_35_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_35_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_36_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_36_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_36_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_36_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_36_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_36_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_36_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_36_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_36_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_36_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_36_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_36_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_36_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_36_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_37_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_37_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_37_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_37_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_37_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_37_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_37_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_37_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_37_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_37_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_37_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_37_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_37_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_37_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_38_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_38_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_38_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_38_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_38_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_38_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_38_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_38_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_38_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_38_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_38_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_38_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_38_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_38_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_39_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_39_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_39_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_39_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_39_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_39_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_39_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_39_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_39_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_39_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_39_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_39_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_39_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_39_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_40_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_40_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_40_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_40_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_40_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_40_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_40_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_40_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_40_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_40_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_40_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_40_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_40_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_40_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_41_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_41_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_41_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_41_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_41_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_41_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_41_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_41_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_41_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_41_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_41_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_41_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_41_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_41_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_42_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_42_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_42_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_42_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_42_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_42_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_42_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_42_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_42_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_42_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_42_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_42_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_42_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_42_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_43_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_43_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_43_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_43_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_43_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_43_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_43_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_43_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_43_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_43_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_43_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_43_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_43_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_43_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_44_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_44_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_44_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_44_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_44_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_44_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_44_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_44_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_44_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_44_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_44_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_44_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_44_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_44_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_45_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_45_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_45_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_45_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_45_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_45_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_45_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_45_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_45_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_45_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_45_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_45_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_45_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_45_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_46_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_46_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_46_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_46_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_46_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_46_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_46_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_46_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_46_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_46_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_46_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_46_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_46_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_46_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_47_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_47_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_47_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_47_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_47_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_47_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_47_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_47_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_47_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_47_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_47_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_47_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_47_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_47_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_48_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_48_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_48_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_48_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_48_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_48_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_48_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_48_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_48_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_48_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_48_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_48_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_48_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_48_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_49_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_49_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_49_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_49_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_49_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_49_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_49_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_49_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_49_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_49_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_49_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_49_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_49_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_49_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_50_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_50_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_50_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_50_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_50_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_50_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_50_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_50_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_50_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_50_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_50_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_50_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_50_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_50_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_51_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_51_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_51_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_51_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_51_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_51_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_51_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_51_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_51_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_51_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_51_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_51_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_51_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_51_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_52_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_52_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_52_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_52_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_52_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_52_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_52_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_52_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_52_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_52_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_52_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_52_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_52_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_52_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_53_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_53_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_53_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_53_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_53_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_53_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_53_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_53_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_53_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_53_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_53_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_53_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_53_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_53_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_54_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_54_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_54_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_54_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_54_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_54_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_54_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_54_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_54_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_54_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_54_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_54_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_54_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_54_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_55_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_55_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_55_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_55_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_55_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_55_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_55_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_55_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_55_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_55_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_55_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_55_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_55_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_55_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_56_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_56_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_56_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_56_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_56_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_56_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_56_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_56_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_56_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_56_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_56_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_56_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_56_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_56_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_57_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_57_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_57_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_57_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_57_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_57_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_57_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_58_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_58_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_58_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_58_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_58_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_58_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_58_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_5_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_5_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_5_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_5_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_5_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_5_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_5_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_6_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_6_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_6_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_6_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_6_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_6_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_6_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_7_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_7_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_7_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_7_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_7_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_7_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_7_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_7_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_7_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_7_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_7_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_7_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_7_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_7_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_8_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_8_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_8_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_8_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_8_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_8_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_8_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_8_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_8_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_8_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_8_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_8_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_8_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_8_2/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_9_1/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_9_1/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_9_1/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_9_1/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_9_1/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_9_1/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_9_1/_17_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_9_2/_11_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_9_2/_12_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_9_2/_13_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_9_2/_14_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_9_2/_15_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_9_2/_16_ ;
 wire \u_multiplier/STAGE3/E_4_2_pp3_9_2/_17_ ;
 wire \u_multiplier/STAGE3/Full_adder_pp3_57_1/_08_ ;
 wire \u_multiplier/STAGE3/Full_adder_pp3_57_1/_09_ ;
 wire \u_multiplier/STAGE3/Full_adder_pp3_57_1/_10_ ;
 wire \u_multiplier/STAGE3/Full_adder_pp3_57_1/_11_ ;
 wire \u_multiplier/STAGE3/Full_adder_pp3_59_1/_08_ ;
 wire \u_multiplier/STAGE3/Full_adder_pp3_59_1/_09_ ;
 wire \u_multiplier/STAGE3/Full_adder_pp3_59_1/_10_ ;
 wire \u_multiplier/STAGE3/Full_adder_pp3_59_1/_11_ ;
 wire \u_multiplier/STAGE4/pp4_10_cout ;
 wire \u_multiplier/STAGE4/pp4_11_cout ;
 wire \u_multiplier/STAGE4/pp4_12_cout ;
 wire \u_multiplier/STAGE4/pp4_13_cout ;
 wire \u_multiplier/STAGE4/pp4_14_cout ;
 wire \u_multiplier/STAGE4/pp4_15_cout ;
 wire \u_multiplier/STAGE4/pp4_16_cout ;
 wire \u_multiplier/STAGE4/pp4_17_cout ;
 wire \u_multiplier/STAGE4/pp4_18_cout ;
 wire \u_multiplier/STAGE4/pp4_19_cout ;
 wire \u_multiplier/STAGE4/pp4_1_ha_c ;
 wire \u_multiplier/STAGE4/pp4_20_cout ;
 wire \u_multiplier/STAGE4/pp4_21_cout ;
 wire \u_multiplier/STAGE4/pp4_22_cout ;
 wire \u_multiplier/STAGE4/pp4_23_cout ;
 wire \u_multiplier/STAGE4/pp4_24_cout ;
 wire \u_multiplier/STAGE4/pp4_25_cout ;
 wire \u_multiplier/STAGE4/pp4_26_cout ;
 wire \u_multiplier/STAGE4/pp4_27_cout ;
 wire \u_multiplier/STAGE4/pp4_28_cout ;
 wire \u_multiplier/STAGE4/pp4_29_cout ;
 wire \u_multiplier/STAGE4/pp4_2_cout ;
 wire \u_multiplier/STAGE4/pp4_30_cout ;
 wire \u_multiplier/STAGE4/pp4_31_cout ;
 wire \u_multiplier/STAGE4/pp4_32_cout ;
 wire \u_multiplier/STAGE4/pp4_33_cout ;
 wire \u_multiplier/STAGE4/pp4_34_cout ;
 wire \u_multiplier/STAGE4/pp4_35_cout ;
 wire \u_multiplier/STAGE4/pp4_36_cout ;
 wire \u_multiplier/STAGE4/pp4_37_cout ;
 wire \u_multiplier/STAGE4/pp4_38_cout ;
 wire \u_multiplier/STAGE4/pp4_39_cout ;
 wire \u_multiplier/STAGE4/pp4_3_cout ;
 wire \u_multiplier/STAGE4/pp4_40_cout ;
 wire \u_multiplier/STAGE4/pp4_41_cout ;
 wire \u_multiplier/STAGE4/pp4_42_cout ;
 wire \u_multiplier/STAGE4/pp4_43_cout ;
 wire \u_multiplier/STAGE4/pp4_44_cout ;
 wire \u_multiplier/STAGE4/pp4_45_cout ;
 wire \u_multiplier/STAGE4/pp4_46_cout ;
 wire \u_multiplier/STAGE4/pp4_47_cout ;
 wire \u_multiplier/STAGE4/pp4_48_cout ;
 wire \u_multiplier/STAGE4/pp4_49_cout ;
 wire \u_multiplier/STAGE4/pp4_4_cout ;
 wire \u_multiplier/STAGE4/pp4_50_cout ;
 wire \u_multiplier/STAGE4/pp4_51_cout ;
 wire \u_multiplier/STAGE4/pp4_52_cout ;
 wire \u_multiplier/STAGE4/pp4_53_cout ;
 wire \u_multiplier/STAGE4/pp4_54_cout ;
 wire \u_multiplier/STAGE4/pp4_55_cout ;
 wire \u_multiplier/STAGE4/pp4_56_cout ;
 wire \u_multiplier/STAGE4/pp4_57_cout ;
 wire \u_multiplier/STAGE4/pp4_58_cout ;
 wire \u_multiplier/STAGE4/pp4_59_cout ;
 wire \u_multiplier/STAGE4/pp4_5_cout ;
 wire \u_multiplier/STAGE4/pp4_60_cout ;
 wire \u_multiplier/STAGE4/pp4_6_cout ;
 wire \u_multiplier/STAGE4/pp4_7_cout ;
 wire \u_multiplier/STAGE4/pp4_8_cout ;
 wire \u_multiplier/STAGE4/pp4_9_cout ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_10/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_10/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_10/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_10/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_10/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_10/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_10/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_11/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_11/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_11/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_11/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_11/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_11/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_11/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_12/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_12/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_12/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_12/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_12/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_12/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_12/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_13/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_13/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_13/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_13/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_13/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_13/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_13/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_14/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_14/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_14/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_14/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_14/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_14/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_14/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_15/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_15/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_15/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_15/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_15/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_15/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_15/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_16/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_16/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_16/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_16/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_16/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_16/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_16/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_17/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_17/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_17/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_17/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_17/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_17/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_17/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_18/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_18/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_18/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_18/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_18/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_18/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_18/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_19/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_19/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_19/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_19/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_19/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_19/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_19/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_2/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_2/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_2/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_2/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_2/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_2/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_2/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_20/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_20/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_20/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_20/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_20/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_20/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_20/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_21/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_21/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_21/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_21/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_21/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_21/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_21/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_22/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_22/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_22/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_22/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_22/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_22/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_22/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_23/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_23/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_23/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_23/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_23/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_23/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_23/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_24/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_24/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_24/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_24/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_24/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_24/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_24/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_25/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_25/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_25/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_25/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_25/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_25/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_25/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_26/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_26/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_26/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_26/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_26/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_26/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_26/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_27/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_27/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_27/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_27/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_27/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_27/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_27/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_28/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_28/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_28/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_28/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_28/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_28/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_28/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_29/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_29/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_29/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_29/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_29/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_29/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_29/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_3/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_3/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_3/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_3/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_3/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_3/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_3/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_30/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_30/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_30/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_30/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_30/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_30/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_30/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_31/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_31/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_31/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_31/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_31/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_31/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_31/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_32/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_32/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_32/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_32/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_32/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_32/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_32/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_33/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_33/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_33/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_33/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_33/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_33/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_33/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_34/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_34/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_34/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_34/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_34/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_34/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_34/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_35/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_35/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_35/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_35/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_35/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_35/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_35/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_36/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_36/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_36/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_36/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_36/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_36/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_36/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_37/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_37/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_37/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_37/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_37/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_37/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_37/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_38/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_38/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_38/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_38/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_38/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_38/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_38/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_39/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_39/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_39/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_39/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_39/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_39/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_39/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_4/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_4/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_4/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_4/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_4/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_4/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_4/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_40/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_40/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_40/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_40/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_40/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_40/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_40/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_41/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_41/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_41/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_41/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_41/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_41/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_41/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_42/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_42/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_42/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_42/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_42/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_42/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_42/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_43/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_43/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_43/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_43/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_43/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_43/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_43/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_44/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_44/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_44/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_44/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_44/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_44/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_44/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_45/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_45/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_45/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_45/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_45/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_45/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_45/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_46/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_46/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_46/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_46/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_46/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_46/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_46/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_47/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_47/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_47/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_47/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_47/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_47/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_47/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_48/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_48/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_48/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_48/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_48/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_48/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_48/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_49/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_49/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_49/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_49/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_49/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_49/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_49/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_5/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_5/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_5/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_5/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_5/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_5/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_5/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_50/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_50/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_50/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_50/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_50/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_50/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_50/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_51/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_51/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_51/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_51/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_51/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_51/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_51/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_52/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_52/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_52/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_52/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_52/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_52/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_52/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_53/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_53/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_53/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_53/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_53/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_53/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_53/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_54/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_54/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_54/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_54/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_54/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_54/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_54/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_55/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_55/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_55/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_55/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_55/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_55/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_55/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_56/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_56/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_56/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_56/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_56/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_56/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_56/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_57/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_57/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_57/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_57/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_57/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_57/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_57/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_58/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_58/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_58/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_58/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_58/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_58/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_58/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_59/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_59/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_59/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_59/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_59/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_59/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_59/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_6/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_6/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_6/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_6/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_6/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_6/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_6/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_60/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_60/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_60/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_60/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_60/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_60/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_60/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_7/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_7/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_7/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_7/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_7/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_7/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_7/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_8/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_8/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_8/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_8/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_8/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_8/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_8/_17_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_9/_11_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_9/_12_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_9/_13_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_9/_14_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_9/_15_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_9/_16_ ;
 wire \u_multiplier/STAGE4/E_4_2_pp4_9/_17_ ;
 wire \u_multiplier/STAGE4/Full_adder_pp4_61/_08_ ;
 wire \u_multiplier/STAGE4/Full_adder_pp4_61/_09_ ;
 wire \u_multiplier/STAGE4/Full_adder_pp4_61/_10_ ;
 wire \u_multiplier/STAGE4/Full_adder_pp4_61/_11_ ;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire valid_reg_out;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net162;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire clknet_0_clk;
 wire clknet_1_0_0_clk;
 wire clknet_1_1_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_4_0__leaf_clk;
 wire clknet_4_1__leaf_clk;
 wire clknet_4_2__leaf_clk;
 wire clknet_4_3__leaf_clk;
 wire clknet_4_4__leaf_clk;
 wire clknet_4_5__leaf_clk;
 wire clknet_4_6__leaf_clk;
 wire clknet_4_7__leaf_clk;
 wire clknet_4_8__leaf_clk;
 wire clknet_4_9__leaf_clk;
 wire clknet_4_10__leaf_clk;
 wire clknet_4_11__leaf_clk;
 wire clknet_4_12__leaf_clk;
 wire clknet_4_13__leaf_clk;
 wire clknet_4_14__leaf_clk;
 wire clknet_4_15__leaf_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire [5:0] addr_ptr;
 wire [2:0] curr_state;
 wire [31:0] data_in_reg;
 wire [5:0] init_count;
 wire [63:0] product;
 wire [31:0] sram_rdata;
 wire [31:0] sram_rdata_reg;
 wire [63:0] \u_multiplier/A ;
 wire [62:0] \u_multiplier/B ;
 wire [1:0] \u_multiplier/pp1_1 ;
 wire [10:0] \u_multiplier/pp1_10 ;
 wire [11:0] \u_multiplier/pp1_11 ;
 wire [12:0] \u_multiplier/pp1_12 ;
 wire [13:0] \u_multiplier/pp1_13 ;
 wire [14:0] \u_multiplier/pp1_14 ;
 wire [15:0] \u_multiplier/pp1_15 ;
 wire [15:0] \u_multiplier/pp1_16 ;
 wire [15:0] \u_multiplier/pp1_17 ;
 wire [15:0] \u_multiplier/pp1_18 ;
 wire [15:0] \u_multiplier/pp1_19 ;
 wire [2:0] \u_multiplier/pp1_2 ;
 wire [15:0] \u_multiplier/pp1_20 ;
 wire [15:0] \u_multiplier/pp1_21 ;
 wire [15:0] \u_multiplier/pp1_22 ;
 wire [15:0] \u_multiplier/pp1_23 ;
 wire [15:0] \u_multiplier/pp1_24 ;
 wire [15:0] \u_multiplier/pp1_25 ;
 wire [15:0] \u_multiplier/pp1_26 ;
 wire [15:0] \u_multiplier/pp1_27 ;
 wire [15:0] \u_multiplier/pp1_28 ;
 wire [15:0] \u_multiplier/pp1_29 ;
 wire [3:0] \u_multiplier/pp1_3 ;
 wire [15:0] \u_multiplier/pp1_30 ;
 wire [15:0] \u_multiplier/pp1_31 ;
 wire [15:0] \u_multiplier/pp1_32 ;
 wire [15:0] \u_multiplier/pp1_33 ;
 wire [15:0] \u_multiplier/pp1_34 ;
 wire [15:0] \u_multiplier/pp1_35 ;
 wire [15:0] \u_multiplier/pp1_36 ;
 wire [15:0] \u_multiplier/pp1_37 ;
 wire [15:0] \u_multiplier/pp1_38 ;
 wire [15:0] \u_multiplier/pp1_39 ;
 wire [4:0] \u_multiplier/pp1_4 ;
 wire [15:0] \u_multiplier/pp1_40 ;
 wire [15:0] \u_multiplier/pp1_41 ;
 wire [15:0] \u_multiplier/pp1_42 ;
 wire [15:0] \u_multiplier/pp1_43 ;
 wire [15:0] \u_multiplier/pp1_44 ;
 wire [15:0] \u_multiplier/pp1_45 ;
 wire [15:0] \u_multiplier/pp1_46 ;
 wire [15:0] \u_multiplier/pp1_47 ;
 wire [15:0] \u_multiplier/pp1_48 ;
 wire [13:0] \u_multiplier/pp1_49 ;
 wire [5:0] \u_multiplier/pp1_5 ;
 wire [12:0] \u_multiplier/pp1_50 ;
 wire [11:0] \u_multiplier/pp1_51 ;
 wire [10:0] \u_multiplier/pp1_52 ;
 wire [9:0] \u_multiplier/pp1_53 ;
 wire [8:0] \u_multiplier/pp1_54 ;
 wire [7:0] \u_multiplier/pp1_55 ;
 wire [6:0] \u_multiplier/pp1_56 ;
 wire [5:0] \u_multiplier/pp1_57 ;
 wire [4:0] \u_multiplier/pp1_58 ;
 wire [3:0] \u_multiplier/pp1_59 ;
 wire [6:0] \u_multiplier/pp1_6 ;
 wire [2:0] \u_multiplier/pp1_60 ;
 wire [1:0] \u_multiplier/pp1_61 ;
 wire [7:0] \u_multiplier/pp1_7 ;
 wire [8:0] \u_multiplier/pp1_8 ;
 wire [9:0] \u_multiplier/pp1_9 ;
 wire [1:0] \u_multiplier/pp2_1 ;
 wire [7:0] \u_multiplier/pp2_10 ;
 wire [7:0] \u_multiplier/pp2_11 ;
 wire [7:0] \u_multiplier/pp2_12 ;
 wire [7:0] \u_multiplier/pp2_13 ;
 wire [7:0] \u_multiplier/pp2_14 ;
 wire [7:0] \u_multiplier/pp2_15 ;
 wire [7:0] \u_multiplier/pp2_16 ;
 wire [7:0] \u_multiplier/pp2_17 ;
 wire [7:0] \u_multiplier/pp2_18 ;
 wire [7:0] \u_multiplier/pp2_19 ;
 wire [2:0] \u_multiplier/pp2_2 ;
 wire [7:0] \u_multiplier/pp2_20 ;
 wire [7:0] \u_multiplier/pp2_21 ;
 wire [7:0] \u_multiplier/pp2_22 ;
 wire [7:0] \u_multiplier/pp2_23 ;
 wire [7:0] \u_multiplier/pp2_24 ;
 wire [7:0] \u_multiplier/pp2_25 ;
 wire [7:0] \u_multiplier/pp2_26 ;
 wire [7:0] \u_multiplier/pp2_27 ;
 wire [7:0] \u_multiplier/pp2_28 ;
 wire [7:0] \u_multiplier/pp2_29 ;
 wire [3:0] \u_multiplier/pp2_3 ;
 wire [7:0] \u_multiplier/pp2_30 ;
 wire [7:0] \u_multiplier/pp2_31 ;
 wire [7:0] \u_multiplier/pp2_32 ;
 wire [7:0] \u_multiplier/pp2_33 ;
 wire [7:0] \u_multiplier/pp2_34 ;
 wire [7:0] \u_multiplier/pp2_35 ;
 wire [7:0] \u_multiplier/pp2_36 ;
 wire [7:0] \u_multiplier/pp2_37 ;
 wire [7:0] \u_multiplier/pp2_38 ;
 wire [7:0] \u_multiplier/pp2_39 ;
 wire [4:0] \u_multiplier/pp2_4 ;
 wire [7:0] \u_multiplier/pp2_40 ;
 wire [7:0] \u_multiplier/pp2_41 ;
 wire [7:0] \u_multiplier/pp2_42 ;
 wire [7:0] \u_multiplier/pp2_43 ;
 wire [7:0] \u_multiplier/pp2_44 ;
 wire [7:0] \u_multiplier/pp2_45 ;
 wire [7:0] \u_multiplier/pp2_46 ;
 wire [7:0] \u_multiplier/pp2_47 ;
 wire [7:0] \u_multiplier/pp2_48 ;
 wire [7:0] \u_multiplier/pp2_49 ;
 wire [5:0] \u_multiplier/pp2_5 ;
 wire [7:0] \u_multiplier/pp2_50 ;
 wire [7:0] \u_multiplier/pp2_51 ;
 wire [7:0] \u_multiplier/pp2_52 ;
 wire [7:0] \u_multiplier/pp2_53 ;
 wire [7:0] \u_multiplier/pp2_54 ;
 wire [7:0] \u_multiplier/pp2_55 ;
 wire [7:0] \u_multiplier/pp2_56 ;
 wire [5:0] \u_multiplier/pp2_57 ;
 wire [4:0] \u_multiplier/pp2_58 ;
 wire [3:0] \u_multiplier/pp2_59 ;
 wire [6:0] \u_multiplier/pp2_6 ;
 wire [2:0] \u_multiplier/pp2_60 ;
 wire [1:0] \u_multiplier/pp2_61 ;
 wire [7:0] \u_multiplier/pp2_7 ;
 wire [7:0] \u_multiplier/pp2_8 ;
 wire [7:0] \u_multiplier/pp2_9 ;
 wire [1:0] \u_multiplier/pp3_1 ;
 wire [3:0] \u_multiplier/pp3_10 ;
 wire [3:0] \u_multiplier/pp3_11 ;
 wire [3:0] \u_multiplier/pp3_12 ;
 wire [3:0] \u_multiplier/pp3_13 ;
 wire [3:0] \u_multiplier/pp3_14 ;
 wire [3:0] \u_multiplier/pp3_15 ;
 wire [3:0] \u_multiplier/pp3_16 ;
 wire [3:0] \u_multiplier/pp3_17 ;
 wire [3:0] \u_multiplier/pp3_18 ;
 wire [3:0] \u_multiplier/pp3_19 ;
 wire [2:0] \u_multiplier/pp3_2 ;
 wire [3:0] \u_multiplier/pp3_20 ;
 wire [3:0] \u_multiplier/pp3_21 ;
 wire [3:0] \u_multiplier/pp3_22 ;
 wire [3:0] \u_multiplier/pp3_23 ;
 wire [3:0] \u_multiplier/pp3_24 ;
 wire [3:0] \u_multiplier/pp3_25 ;
 wire [3:0] \u_multiplier/pp3_26 ;
 wire [3:0] \u_multiplier/pp3_27 ;
 wire [3:0] \u_multiplier/pp3_28 ;
 wire [3:0] \u_multiplier/pp3_29 ;
 wire [3:0] \u_multiplier/pp3_3 ;
 wire [3:0] \u_multiplier/pp3_30 ;
 wire [3:0] \u_multiplier/pp3_31 ;
 wire [3:0] \u_multiplier/pp3_32 ;
 wire [3:0] \u_multiplier/pp3_33 ;
 wire [3:0] \u_multiplier/pp3_34 ;
 wire [3:0] \u_multiplier/pp3_35 ;
 wire [3:0] \u_multiplier/pp3_36 ;
 wire [3:0] \u_multiplier/pp3_37 ;
 wire [3:0] \u_multiplier/pp3_38 ;
 wire [3:0] \u_multiplier/pp3_39 ;
 wire [3:0] \u_multiplier/pp3_4 ;
 wire [3:0] \u_multiplier/pp3_40 ;
 wire [3:0] \u_multiplier/pp3_41 ;
 wire [3:0] \u_multiplier/pp3_42 ;
 wire [3:0] \u_multiplier/pp3_43 ;
 wire [3:0] \u_multiplier/pp3_44 ;
 wire [3:0] \u_multiplier/pp3_45 ;
 wire [3:0] \u_multiplier/pp3_46 ;
 wire [3:0] \u_multiplier/pp3_47 ;
 wire [3:0] \u_multiplier/pp3_48 ;
 wire [3:0] \u_multiplier/pp3_49 ;
 wire [3:0] \u_multiplier/pp3_5 ;
 wire [3:0] \u_multiplier/pp3_50 ;
 wire [3:0] \u_multiplier/pp3_51 ;
 wire [3:0] \u_multiplier/pp3_52 ;
 wire [3:0] \u_multiplier/pp3_53 ;
 wire [3:0] \u_multiplier/pp3_54 ;
 wire [3:0] \u_multiplier/pp3_55 ;
 wire [3:0] \u_multiplier/pp3_56 ;
 wire [3:0] \u_multiplier/pp3_57 ;
 wire [3:0] \u_multiplier/pp3_58 ;
 wire [3:0] \u_multiplier/pp3_59 ;
 wire [3:0] \u_multiplier/pp3_6 ;
 wire [3:0] \u_multiplier/pp3_60 ;
 wire [1:0] \u_multiplier/pp3_61 ;
 wire [3:0] \u_multiplier/pp3_7 ;
 wire [3:0] \u_multiplier/pp3_8 ;
 wire [3:0] \u_multiplier/pp3_9 ;

 INV_X2 _0675_ (.A(net12),
    .ZN(_0370_));
 INV_X2 _0676_ (.A(net46),
    .ZN(_0307_));
 INV_X1 _0677_ (.A(init_count[5]),
    .ZN(_0371_));
 INV_X1 _0678_ (.A(curr_state[2]),
    .ZN(_0372_));
 INV_X1 _0679_ (.A(net48),
    .ZN(_0373_));
 INV_X1 _0680_ (.A(net180),
    .ZN(_0374_));
 NOR2_X4 _0681_ (.A1(_0370_),
    .A2(_0373_),
    .ZN(_0303_));
 NAND2_X2 _0682_ (.A1(net12),
    .A2(net220),
    .ZN(_0308_));
 NAND2_X1 _0683_ (.A1(init_count[1]),
    .A2(init_count[0]),
    .ZN(_0375_));
 AND4_X2 _0684_ (.A1(init_count[1]),
    .A2(init_count[0]),
    .A3(init_count[3]),
    .A4(init_count[2]),
    .ZN(_0376_));
 INV_X1 _0685_ (.A(_0376_),
    .ZN(_0377_));
 AND2_X1 _0686_ (.A1(init_count[5]),
    .A2(init_count[4]),
    .ZN(_0378_));
 AND3_X1 _0687_ (.A1(net46),
    .A2(_0376_),
    .A3(_0378_),
    .ZN(_0379_));
 NOR2_X2 _0688_ (.A1(_0370_),
    .A2(_0307_),
    .ZN(_0380_));
 NAND2_X2 _0689_ (.A1(net12),
    .A2(net46),
    .ZN(_0381_));
 AND3_X1 _0690_ (.A1(curr_state[2]),
    .A2(_0376_),
    .A3(_0378_),
    .ZN(_0382_));
 NAND2_X1 _0691_ (.A1(_0380_),
    .A2(_0382_),
    .ZN(_0383_));
 OAI21_X1 _0692_ (.A(_0383_),
    .B1(_0373_),
    .B2(_0370_),
    .ZN(_0305_));
 NAND3_X1 _0693_ (.A1(net45),
    .A2(net200),
    .A3(_0380_),
    .ZN(_0384_));
 OAI21_X1 _0694_ (.A(net201),
    .B1(_0379_),
    .B2(_0308_),
    .ZN(_0306_));
 AOI22_X1 _0695_ (.A1(net12),
    .A2(net163),
    .B1(_0380_),
    .B2(net45),
    .ZN(_0304_));
 AND2_X1 _0696_ (.A1(net11),
    .A2(sram_rdata[0]),
    .ZN(_0271_));
 AND2_X1 _0697_ (.A1(net11),
    .A2(sram_rdata[1]),
    .ZN(_0282_));
 AND2_X1 _0698_ (.A1(net11),
    .A2(sram_rdata[2]),
    .ZN(_0293_));
 AND2_X1 _0699_ (.A1(net11),
    .A2(sram_rdata[3]),
    .ZN(_0296_));
 AND2_X1 _0700_ (.A1(net11),
    .A2(sram_rdata[4]),
    .ZN(_0297_));
 AND2_X1 _0701_ (.A1(net11),
    .A2(sram_rdata[5]),
    .ZN(_0298_));
 AND2_X1 _0702_ (.A1(net11),
    .A2(sram_rdata[6]),
    .ZN(_0299_));
 AND2_X1 _0703_ (.A1(net11),
    .A2(sram_rdata[7]),
    .ZN(_0300_));
 AND2_X1 _0704_ (.A1(net11),
    .A2(sram_rdata[8]),
    .ZN(_0301_));
 AND2_X1 _0705_ (.A1(net11),
    .A2(sram_rdata[9]),
    .ZN(_0302_));
 AND2_X1 _0706_ (.A1(net11),
    .A2(sram_rdata[10]),
    .ZN(_0272_));
 AND2_X1 _0707_ (.A1(net11),
    .A2(sram_rdata[11]),
    .ZN(_0273_));
 AND2_X1 _0708_ (.A1(net11),
    .A2(sram_rdata[12]),
    .ZN(_0274_));
 AND2_X1 _0709_ (.A1(net11),
    .A2(sram_rdata[13]),
    .ZN(_0275_));
 AND2_X1 _0710_ (.A1(net11),
    .A2(sram_rdata[14]),
    .ZN(_0276_));
 AND2_X1 _0711_ (.A1(net11),
    .A2(sram_rdata[15]),
    .ZN(_0277_));
 AND2_X1 _0712_ (.A1(net11),
    .A2(sram_rdata[16]),
    .ZN(_0278_));
 AND2_X1 _0713_ (.A1(net11),
    .A2(sram_rdata[17]),
    .ZN(_0279_));
 AND2_X1 _0714_ (.A1(net11),
    .A2(sram_rdata[18]),
    .ZN(_0280_));
 AND2_X1 _0715_ (.A1(net11),
    .A2(sram_rdata[19]),
    .ZN(_0281_));
 AND2_X1 _0716_ (.A1(net11),
    .A2(sram_rdata[20]),
    .ZN(_0283_));
 AND2_X1 _0717_ (.A1(net11),
    .A2(sram_rdata[21]),
    .ZN(_0284_));
 AND2_X1 _0718_ (.A1(net11),
    .A2(sram_rdata[22]),
    .ZN(_0285_));
 AND2_X1 _0719_ (.A1(net11),
    .A2(sram_rdata[23]),
    .ZN(_0286_));
 AND2_X1 _0720_ (.A1(net11),
    .A2(sram_rdata[24]),
    .ZN(_0287_));
 AND2_X1 _0721_ (.A1(net11),
    .A2(sram_rdata[25]),
    .ZN(_0288_));
 AND2_X1 _0722_ (.A1(net11),
    .A2(sram_rdata[26]),
    .ZN(_0289_));
 AND2_X1 _0723_ (.A1(net11),
    .A2(sram_rdata[27]),
    .ZN(_0290_));
 AND2_X1 _0724_ (.A1(net11),
    .A2(sram_rdata[28]),
    .ZN(_0291_));
 AND2_X1 _0725_ (.A1(net11),
    .A2(sram_rdata[29]),
    .ZN(_0292_));
 AND2_X1 _0726_ (.A1(net11),
    .A2(sram_rdata[30]),
    .ZN(_0294_));
 AND2_X1 _0727_ (.A1(net11),
    .A2(sram_rdata[31]),
    .ZN(_0295_));
 AND2_X1 _0728_ (.A1(product[0]),
    .A2(net9),
    .ZN(_0201_));
 AND2_X1 _0729_ (.A1(product[1]),
    .A2(net9),
    .ZN(_0212_));
 AND2_X1 _0730_ (.A1(product[2]),
    .A2(net9),
    .ZN(_0223_));
 AND2_X1 _0731_ (.A1(product[3]),
    .A2(net9),
    .ZN(_0234_));
 AND2_X1 _0732_ (.A1(product[4]),
    .A2(_0303_),
    .ZN(_0245_));
 AND2_X1 _0733_ (.A1(product[5]),
    .A2(net9),
    .ZN(_0256_));
 AND2_X1 _0734_ (.A1(product[6]),
    .A2(net10),
    .ZN(_0261_));
 AND2_X1 _0735_ (.A1(product[7]),
    .A2(net10),
    .ZN(_0262_));
 AND2_X1 _0736_ (.A1(product[8]),
    .A2(_0303_),
    .ZN(_0263_));
 AND2_X1 _0737_ (.A1(product[9]),
    .A2(net10),
    .ZN(_0264_));
 AND2_X1 _0738_ (.A1(product[10]),
    .A2(net9),
    .ZN(_0202_));
 AND2_X1 _0739_ (.A1(product[11]),
    .A2(net10),
    .ZN(_0203_));
 AND2_X1 _0740_ (.A1(product[12]),
    .A2(net9),
    .ZN(_0204_));
 AND2_X1 _0741_ (.A1(product[13]),
    .A2(net9),
    .ZN(_0205_));
 AND2_X1 _0742_ (.A1(product[14]),
    .A2(net9),
    .ZN(_0206_));
 AND2_X1 _0743_ (.A1(product[15]),
    .A2(net9),
    .ZN(_0207_));
 AND2_X1 _0744_ (.A1(product[16]),
    .A2(net9),
    .ZN(_0208_));
 AND2_X1 _0745_ (.A1(product[17]),
    .A2(net9),
    .ZN(_0209_));
 AND2_X1 _0746_ (.A1(product[18]),
    .A2(net10),
    .ZN(_0210_));
 AND2_X1 _0747_ (.A1(product[19]),
    .A2(_0303_),
    .ZN(_0211_));
 AND2_X1 _0748_ (.A1(product[20]),
    .A2(net9),
    .ZN(_0213_));
 AND2_X1 _0749_ (.A1(product[21]),
    .A2(net9),
    .ZN(_0214_));
 AND2_X1 _0750_ (.A1(product[22]),
    .A2(_0303_),
    .ZN(_0215_));
 AND2_X1 _0751_ (.A1(product[23]),
    .A2(net10),
    .ZN(_0216_));
 AND2_X1 _0752_ (.A1(product[24]),
    .A2(net9),
    .ZN(_0217_));
 AND2_X1 _0753_ (.A1(product[25]),
    .A2(_0303_),
    .ZN(_0218_));
 AND2_X1 _0754_ (.A1(product[26]),
    .A2(_0303_),
    .ZN(_0219_));
 AND2_X1 _0755_ (.A1(product[27]),
    .A2(_0303_),
    .ZN(_0220_));
 AND2_X1 _0756_ (.A1(product[28]),
    .A2(_0303_),
    .ZN(_0221_));
 AND2_X1 _0757_ (.A1(product[29]),
    .A2(net9),
    .ZN(_0222_));
 AND2_X1 _0758_ (.A1(product[30]),
    .A2(_0303_),
    .ZN(_0224_));
 AND2_X1 _0759_ (.A1(product[31]),
    .A2(net10),
    .ZN(_0225_));
 AND2_X1 _0760_ (.A1(product[32]),
    .A2(net9),
    .ZN(_0226_));
 AND2_X1 _0761_ (.A1(product[33]),
    .A2(net9),
    .ZN(_0227_));
 AND2_X1 _0762_ (.A1(product[34]),
    .A2(net9),
    .ZN(_0228_));
 AND2_X1 _0763_ (.A1(product[35]),
    .A2(net9),
    .ZN(_0229_));
 AND2_X1 _0764_ (.A1(product[36]),
    .A2(_0303_),
    .ZN(_0230_));
 AND2_X1 _0765_ (.A1(product[37]),
    .A2(_0303_),
    .ZN(_0231_));
 AND2_X1 _0766_ (.A1(product[38]),
    .A2(net9),
    .ZN(_0232_));
 AND2_X1 _0767_ (.A1(product[39]),
    .A2(net10),
    .ZN(_0233_));
 AND2_X1 _0768_ (.A1(product[40]),
    .A2(net9),
    .ZN(_0235_));
 AND2_X1 _0769_ (.A1(product[41]),
    .A2(net9),
    .ZN(_0236_));
 AND2_X1 _0770_ (.A1(product[42]),
    .A2(net9),
    .ZN(_0237_));
 AND2_X1 _0771_ (.A1(product[43]),
    .A2(net10),
    .ZN(_0238_));
 AND2_X1 _0772_ (.A1(product[44]),
    .A2(_0303_),
    .ZN(_0239_));
 AND2_X1 _0773_ (.A1(product[45]),
    .A2(net9),
    .ZN(_0240_));
 AND2_X1 _0774_ (.A1(product[46]),
    .A2(_0303_),
    .ZN(_0241_));
 AND2_X1 _0775_ (.A1(product[47]),
    .A2(_0303_),
    .ZN(_0242_));
 AND2_X1 _0776_ (.A1(product[48]),
    .A2(_0303_),
    .ZN(_0243_));
 AND2_X1 _0777_ (.A1(product[49]),
    .A2(net10),
    .ZN(_0244_));
 AND2_X1 _0778_ (.A1(product[50]),
    .A2(_0303_),
    .ZN(_0246_));
 AND2_X1 _0779_ (.A1(product[51]),
    .A2(_0303_),
    .ZN(_0247_));
 AND2_X1 _0780_ (.A1(product[52]),
    .A2(_0303_),
    .ZN(_0248_));
 AND2_X1 _0781_ (.A1(product[53]),
    .A2(net9),
    .ZN(_0249_));
 AND2_X1 _0782_ (.A1(product[54]),
    .A2(net10),
    .ZN(_0250_));
 AND2_X1 _0783_ (.A1(product[55]),
    .A2(net9),
    .ZN(_0251_));
 AND2_X1 _0784_ (.A1(product[56]),
    .A2(net9),
    .ZN(_0252_));
 AND2_X1 _0785_ (.A1(product[57]),
    .A2(net9),
    .ZN(_0253_));
 AND2_X1 _0786_ (.A1(product[58]),
    .A2(net10),
    .ZN(_0254_));
 AND2_X1 _0787_ (.A1(product[59]),
    .A2(net9),
    .ZN(_0255_));
 AND2_X1 _0788_ (.A1(product[60]),
    .A2(net9),
    .ZN(_0257_));
 AND2_X1 _0789_ (.A1(product[61]),
    .A2(_0303_),
    .ZN(_0258_));
 AND2_X1 _0790_ (.A1(product[62]),
    .A2(net9),
    .ZN(_0259_));
 AND2_X1 _0791_ (.A1(product[63]),
    .A2(net9),
    .ZN(_0260_));
 AND2_X1 _0792_ (.A1(net11),
    .A2(net13),
    .ZN(_0169_));
 AND2_X1 _0793_ (.A1(net12),
    .A2(net24),
    .ZN(_0180_));
 AND2_X1 _0794_ (.A1(net12),
    .A2(net35),
    .ZN(_0191_));
 AND2_X1 _0795_ (.A1(net11),
    .A2(net38),
    .ZN(_0194_));
 AND2_X1 _0796_ (.A1(net11),
    .A2(net39),
    .ZN(_0195_));
 AND2_X1 _0797_ (.A1(net11),
    .A2(net40),
    .ZN(_0196_));
 AND2_X1 _0798_ (.A1(net12),
    .A2(net41),
    .ZN(_0197_));
 AND2_X1 _0799_ (.A1(net12),
    .A2(net42),
    .ZN(_0198_));
 AND2_X1 _0800_ (.A1(net11),
    .A2(net43),
    .ZN(_0199_));
 AND2_X1 _0801_ (.A1(net11),
    .A2(net44),
    .ZN(_0200_));
 AND2_X1 _0802_ (.A1(net11),
    .A2(net14),
    .ZN(_0170_));
 AND2_X1 _0803_ (.A1(net12),
    .A2(net15),
    .ZN(_0171_));
 AND2_X1 _0804_ (.A1(net12),
    .A2(net16),
    .ZN(_0172_));
 AND2_X1 _0805_ (.A1(net47),
    .A2(net17),
    .ZN(_0173_));
 AND2_X1 _0806_ (.A1(net11),
    .A2(net18),
    .ZN(_0174_));
 AND2_X1 _0807_ (.A1(net12),
    .A2(net19),
    .ZN(_0175_));
 AND2_X1 _0808_ (.A1(net12),
    .A2(net20),
    .ZN(_0176_));
 AND2_X1 _0809_ (.A1(net47),
    .A2(net21),
    .ZN(_0177_));
 AND2_X1 _0810_ (.A1(net12),
    .A2(net22),
    .ZN(_0178_));
 AND2_X1 _0811_ (.A1(net12),
    .A2(net23),
    .ZN(_0179_));
 AND2_X1 _0812_ (.A1(net12),
    .A2(net25),
    .ZN(_0181_));
 AND2_X1 _0813_ (.A1(net12),
    .A2(net26),
    .ZN(_0182_));
 AND2_X1 _0814_ (.A1(net11),
    .A2(net27),
    .ZN(_0183_));
 AND2_X1 _0815_ (.A1(net11),
    .A2(net28),
    .ZN(_0184_));
 AND2_X1 _0816_ (.A1(net12),
    .A2(net29),
    .ZN(_0185_));
 AND2_X1 _0817_ (.A1(net12),
    .A2(net30),
    .ZN(_0186_));
 AND2_X1 _0818_ (.A1(net47),
    .A2(net31),
    .ZN(_0187_));
 AND2_X1 _0819_ (.A1(net12),
    .A2(net32),
    .ZN(_0188_));
 AND2_X1 _0820_ (.A1(net12),
    .A2(net33),
    .ZN(_0189_));
 AND2_X1 _0821_ (.A1(net12),
    .A2(net34),
    .ZN(_0190_));
 AND2_X1 _0822_ (.A1(net12),
    .A2(net36),
    .ZN(_0192_));
 AND2_X1 _0823_ (.A1(net11),
    .A2(net37),
    .ZN(_0193_));
 NAND2_X2 _0824_ (.A1(net12),
    .A2(_0307_),
    .ZN(_0385_));
 OAI21_X1 _0825_ (.A(net12),
    .B1(_0307_),
    .B2(_0382_),
    .ZN(_0386_));
 AOI21_X4 _0826_ (.A(_0372_),
    .B1(_0376_),
    .B2(_0378_),
    .ZN(_0387_));
 AOI22_X1 _0827_ (.A1(init_count[0]),
    .A2(net48),
    .B1(net184),
    .B2(_0387_),
    .ZN(_0388_));
 OAI22_X1 _0828_ (.A1(net185),
    .A2(_0386_),
    .B1(_0388_),
    .B2(_0381_),
    .ZN(_0265_));
 AOI21_X1 _0829_ (.A(net48),
    .B1(_0375_),
    .B2(curr_state[2]),
    .ZN(_0389_));
 INV_X1 _0830_ (.A(_0389_),
    .ZN(_0390_));
 AOI21_X1 _0831_ (.A(init_count[1]),
    .B1(init_count[0]),
    .B2(curr_state[2]),
    .ZN(_0391_));
 OR3_X1 _0832_ (.A1(_0381_),
    .A2(_0389_),
    .A3(_0391_),
    .ZN(_0392_));
 OAI211_X1 _0833_ (.A(_0383_),
    .B(_0392_),
    .C1(_0385_),
    .C2(net199),
    .ZN(_0266_));
 NOR3_X1 _0834_ (.A1(init_count[2]),
    .A2(_0372_),
    .A3(_0375_),
    .ZN(_0393_));
 AOI211_X1 _0835_ (.A(_0382_),
    .B(_0393_),
    .C1(_0390_),
    .C2(init_count[2]),
    .ZN(_0394_));
 OAI22_X1 _0836_ (.A1(net193),
    .A2(_0385_),
    .B1(_0394_),
    .B2(_0381_),
    .ZN(_0267_));
 NOR2_X1 _0837_ (.A1(_0658_),
    .A2(_0375_),
    .ZN(_0395_));
 XOR2_X2 _0838_ (.A(init_count[3]),
    .B(_0395_),
    .Z(_0396_));
 AOI221_X2 _0839_ (.A(_0382_),
    .B1(_0396_),
    .B2(curr_state[2]),
    .C1(net48),
    .C2(init_count[3]),
    .ZN(_0397_));
 OAI22_X1 _0840_ (.A1(net204),
    .A2(_0385_),
    .B1(_0397_),
    .B2(_0381_),
    .ZN(_0268_));
 NAND3_X1 _0841_ (.A1(_0371_),
    .A2(init_count[4]),
    .A3(_0376_),
    .ZN(_0398_));
 OAI21_X1 _0842_ (.A(curr_state[2]),
    .B1(_0376_),
    .B2(init_count[4]),
    .ZN(_0399_));
 INV_X1 _0843_ (.A(_0399_),
    .ZN(_0400_));
 AOI22_X1 _0844_ (.A1(net234),
    .A2(net48),
    .B1(_0398_),
    .B2(_0400_),
    .ZN(_0401_));
 OAI22_X1 _0845_ (.A1(net196),
    .A2(_0385_),
    .B1(_0401_),
    .B2(_0381_),
    .ZN(_0269_));
 OAI21_X1 _0846_ (.A(net189),
    .B1(_0377_),
    .B2(_0660_),
    .ZN(_0402_));
 AOI22_X1 _0847_ (.A1(net233),
    .A2(net48),
    .B1(_0402_),
    .B2(curr_state[2]),
    .ZN(_0403_));
 OAI22_X1 _0848_ (.A1(net190),
    .A2(_0385_),
    .B1(_0403_),
    .B2(_0381_),
    .ZN(_0270_));
 NOR2_X1 _0849_ (.A1(_0373_),
    .A2(addr_ptr[0]),
    .ZN(_0404_));
 AOI21_X1 _0850_ (.A(_0404_),
    .B1(_0387_),
    .B2(net208),
    .ZN(_0405_));
 OAI22_X1 _0851_ (.A1(net176),
    .A2(_0385_),
    .B1(net209),
    .B2(_0381_),
    .ZN(_0163_));
 NAND2_X1 _0852_ (.A1(addr_ptr[0]),
    .A2(addr_ptr[1]),
    .ZN(_0406_));
 XOR2_X1 _0853_ (.A(addr_ptr[0]),
    .B(addr_ptr[1]),
    .Z(_0407_));
 OAI211_X1 _0854_ (.A(_0380_),
    .B(_0407_),
    .C1(_0387_),
    .C2(net48),
    .ZN(_0408_));
 OAI21_X1 _0855_ (.A(_0408_),
    .B1(_0385_),
    .B2(net2),
    .ZN(_0164_));
 AND4_X1 _0856_ (.A1(addr_ptr[0]),
    .A2(addr_ptr[1]),
    .A3(addr_ptr[3]),
    .A4(addr_ptr[2]),
    .ZN(_0409_));
 NAND3_X1 _0857_ (.A1(net187),
    .A2(net182),
    .A3(_0409_),
    .ZN(_0410_));
 AOI21_X2 _0858_ (.A(_0387_),
    .B1(_0410_),
    .B2(net48),
    .ZN(_0411_));
 AOI21_X1 _0859_ (.A(_0381_),
    .B1(_0406_),
    .B2(net213),
    .ZN(_0412_));
 OAI21_X1 _0860_ (.A(_0412_),
    .B1(_0406_),
    .B2(net213),
    .ZN(_0413_));
 OAI22_X1 _0861_ (.A1(net214),
    .A2(_0385_),
    .B1(_0411_),
    .B2(_0413_),
    .ZN(_0165_));
 NOR3_X1 _0862_ (.A1(_0307_),
    .A2(net213),
    .A3(_0406_),
    .ZN(_0414_));
 OAI21_X1 _0863_ (.A(net12),
    .B1(_0374_),
    .B2(_0414_),
    .ZN(_0415_));
 AOI221_X1 _0864_ (.A(_0415_),
    .B1(_0414_),
    .B2(_0374_),
    .C1(net46),
    .C2(_0411_),
    .ZN(_0166_));
 NAND2_X1 _0865_ (.A1(net46),
    .A2(_0409_),
    .ZN(_0416_));
 OR2_X1 _0866_ (.A1(_0654_),
    .A2(_0416_),
    .ZN(_0417_));
 XNOR2_X1 _0867_ (.A(net206),
    .B(_0416_),
    .ZN(_0418_));
 AOI211_X1 _0868_ (.A(_0370_),
    .B(net207),
    .C1(_0411_),
    .C2(net46),
    .ZN(_0167_));
 XNOR2_X1 _0869_ (.A(net7),
    .B(_0417_),
    .ZN(_0419_));
 AOI211_X1 _0870_ (.A(_0370_),
    .B(net8),
    .C1(_0411_),
    .C2(net46),
    .ZN(_0168_));
 DFF_X1 _0871_ (.D(net164),
    .CK(clknet_4_7__leaf_clk),
    .Q(curr_state[0]),
    .QN(_0518_));
 DFF_X2 _0872_ (.D(_0305_),
    .CK(clknet_4_7__leaf_clk),
    .Q(net48),
    .QN(_0519_));
 DFF_X2 _0873_ (.D(net202),
    .CK(clknet_4_6__leaf_clk),
    .Q(curr_state[2]),
    .QN(_0520_));
 DFF_X2 _0874_ (.D(_0201_),
    .CK(clknet_4_9__leaf_clk),
    .Q(net49),
    .QN(_0521_));
 DFF_X2 _0875_ (.D(_0212_),
    .CK(clknet_4_9__leaf_clk),
    .Q(net60),
    .QN(_0522_));
 DFF_X2 _0876_ (.D(_0223_),
    .CK(clknet_4_9__leaf_clk),
    .Q(net71),
    .QN(_0523_));
 DFF_X2 _0877_ (.D(_0234_),
    .CK(clknet_4_9__leaf_clk),
    .Q(net82),
    .QN(_0524_));
 DFF_X1 _0878_ (.D(_0245_),
    .CK(clknet_4_3__leaf_clk),
    .Q(net93),
    .QN(_0525_));
 DFF_X2 _0879_ (.D(_0256_),
    .CK(clknet_4_9__leaf_clk),
    .Q(net104),
    .QN(_0526_));
 DFF_X2 _0880_ (.D(_0261_),
    .CK(clknet_4_15__leaf_clk),
    .Q(net109),
    .QN(_0527_));
 DFF_X2 _0881_ (.D(_0262_),
    .CK(clknet_4_15__leaf_clk),
    .Q(net110),
    .QN(_0528_));
 DFF_X2 _0882_ (.D(_0263_),
    .CK(clknet_4_12__leaf_clk),
    .Q(net111),
    .QN(_0529_));
 DFF_X2 _0883_ (.D(_0264_),
    .CK(clknet_4_14__leaf_clk),
    .Q(net112),
    .QN(_0530_));
 DFF_X2 _0884_ (.D(_0202_),
    .CK(clknet_4_14__leaf_clk),
    .Q(net50),
    .QN(_0531_));
 DFF_X2 _0885_ (.D(_0203_),
    .CK(clknet_4_14__leaf_clk),
    .Q(net51),
    .QN(_0532_));
 DFF_X2 _0886_ (.D(_0204_),
    .CK(clknet_4_14__leaf_clk),
    .Q(net52),
    .QN(_0533_));
 DFF_X2 _0887_ (.D(_0205_),
    .CK(clknet_4_14__leaf_clk),
    .Q(net53),
    .QN(_0534_));
 DFF_X1 _0888_ (.D(_0206_),
    .CK(clknet_4_12__leaf_clk),
    .Q(net54),
    .QN(_0535_));
 DFF_X2 _0889_ (.D(_0207_),
    .CK(clknet_4_14__leaf_clk),
    .Q(net55),
    .QN(_0536_));
 DFF_X2 _0890_ (.D(_0208_),
    .CK(clknet_4_2__leaf_clk),
    .Q(net56),
    .QN(_0537_));
 DFF_X2 _0891_ (.D(_0209_),
    .CK(clknet_4_10__leaf_clk),
    .Q(net57),
    .QN(_0538_));
 DFF_X2 _0892_ (.D(_0210_),
    .CK(clknet_4_1__leaf_clk),
    .Q(net58),
    .QN(_0539_));
 DFF_X2 _0893_ (.D(_0211_),
    .CK(clknet_4_4__leaf_clk),
    .Q(net59),
    .QN(_0540_));
 DFF_X2 _0894_ (.D(_0213_),
    .CK(clknet_4_11__leaf_clk),
    .Q(net61),
    .QN(_0541_));
 DFF_X2 _0895_ (.D(_0214_),
    .CK(clknet_4_11__leaf_clk),
    .Q(net62),
    .QN(_0542_));
 DFF_X2 _0896_ (.D(_0215_),
    .CK(clknet_4_6__leaf_clk),
    .Q(net63),
    .QN(_0543_));
 DFF_X1 _0897_ (.D(_0216_),
    .CK(clknet_4_4__leaf_clk),
    .Q(net64),
    .QN(_0544_));
 DFF_X2 _0898_ (.D(_0217_),
    .CK(clknet_4_11__leaf_clk),
    .Q(net65),
    .QN(_0545_));
 DFF_X1 _0899_ (.D(_0218_),
    .CK(clknet_4_5__leaf_clk),
    .Q(net66),
    .QN(_0546_));
 DFF_X2 _0900_ (.D(_0219_),
    .CK(clknet_4_5__leaf_clk),
    .Q(net67),
    .QN(_0547_));
 DFF_X2 _0901_ (.D(_0220_),
    .CK(clknet_4_5__leaf_clk),
    .Q(net68),
    .QN(_0548_));
 DFF_X2 _0902_ (.D(_0221_),
    .CK(clknet_4_4__leaf_clk),
    .Q(net69),
    .QN(_0549_));
 DFF_X2 _0903_ (.D(_0222_),
    .CK(clknet_4_9__leaf_clk),
    .Q(net70),
    .QN(_0550_));
 DFF_X1 _0904_ (.D(_0224_),
    .CK(clknet_4_1__leaf_clk),
    .Q(net72),
    .QN(_0551_));
 DFF_X2 _0905_ (.D(_0225_),
    .CK(clknet_4_1__leaf_clk),
    .Q(net73),
    .QN(_0552_));
 DFF_X1 _0906_ (.D(_0226_),
    .CK(clknet_4_3__leaf_clk),
    .Q(net74),
    .QN(_0553_));
 DFF_X2 _0907_ (.D(_0227_),
    .CK(clknet_4_12__leaf_clk),
    .Q(net75),
    .QN(_0554_));
 DFF_X2 _0908_ (.D(_0228_),
    .CK(clknet_4_8__leaf_clk),
    .Q(net76),
    .QN(_0555_));
 DFF_X2 _0909_ (.D(_0229_),
    .CK(clknet_4_8__leaf_clk),
    .Q(net77),
    .QN(_0556_));
 DFF_X2 _0910_ (.D(_0230_),
    .CK(clknet_4_12__leaf_clk),
    .Q(net78),
    .QN(_0557_));
 DFF_X2 _0911_ (.D(_0231_),
    .CK(clknet_4_12__leaf_clk),
    .Q(net79),
    .QN(_0558_));
 DFF_X2 _0912_ (.D(_0232_),
    .CK(clknet_4_8__leaf_clk),
    .Q(net80),
    .QN(_0559_));
 DFF_X2 _0913_ (.D(_0233_),
    .CK(clknet_4_10__leaf_clk),
    .Q(net81),
    .QN(_0560_));
 DFF_X2 _0914_ (.D(_0235_),
    .CK(clknet_4_8__leaf_clk),
    .Q(net83),
    .QN(_0561_));
 DFF_X2 _0915_ (.D(_0236_),
    .CK(clknet_4_8__leaf_clk),
    .Q(net84),
    .QN(_0562_));
 DFF_X2 _0916_ (.D(_0237_),
    .CK(clknet_4_8__leaf_clk),
    .Q(net85),
    .QN(_0563_));
 DFF_X2 _0917_ (.D(_0238_),
    .CK(clknet_4_2__leaf_clk),
    .Q(net86),
    .QN(_0564_));
 DFF_X2 _0918_ (.D(_0239_),
    .CK(clknet_4_2__leaf_clk),
    .Q(net87),
    .QN(_0565_));
 DFF_X2 _0919_ (.D(_0240_),
    .CK(clknet_4_2__leaf_clk),
    .Q(net88),
    .QN(_0566_));
 DFF_X1 _0920_ (.D(_0241_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net89),
    .QN(_0567_));
 DFF_X2 _0921_ (.D(_0242_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net90),
    .QN(_0568_));
 DFF_X2 _0922_ (.D(_0243_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net91),
    .QN(_0569_));
 DFF_X2 _0923_ (.D(_0244_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net92),
    .QN(_0570_));
 DFF_X2 _0924_ (.D(_0246_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net94),
    .QN(_0571_));
 DFF_X1 _0925_ (.D(_0247_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net95),
    .QN(_0572_));
 DFF_X1 _0926_ (.D(_0248_),
    .CK(clknet_4_0__leaf_clk),
    .Q(net96),
    .QN(_0573_));
 DFF_X2 _0927_ (.D(_0249_),
    .CK(clknet_4_2__leaf_clk),
    .Q(net97),
    .QN(_0574_));
 DFF_X2 _0928_ (.D(_0250_),
    .CK(clknet_4_12__leaf_clk),
    .Q(net98),
    .QN(_0575_));
 DFF_X1 _0929_ (.D(_0251_),
    .CK(clknet_4_14__leaf_clk),
    .Q(net99),
    .QN(_0576_));
 DFF_X2 _0930_ (.D(_0252_),
    .CK(clknet_4_10__leaf_clk),
    .Q(net100),
    .QN(_0577_));
 DFF_X1 _0931_ (.D(_0253_),
    .CK(clknet_4_10__leaf_clk),
    .Q(net101),
    .QN(_0578_));
 DFF_X2 _0932_ (.D(_0254_),
    .CK(clknet_4_10__leaf_clk),
    .Q(net102),
    .QN(_0579_));
 DFF_X2 _0933_ (.D(_0255_),
    .CK(clknet_4_11__leaf_clk),
    .Q(net103),
    .QN(_0580_));
 DFF_X2 _0934_ (.D(_0257_),
    .CK(clknet_4_11__leaf_clk),
    .Q(net105),
    .QN(_0581_));
 DFF_X2 _0935_ (.D(_0258_),
    .CK(clknet_4_15__leaf_clk),
    .Q(net106),
    .QN(_0582_));
 DFF_X2 _0936_ (.D(_0259_),
    .CK(clknet_4_11__leaf_clk),
    .Q(net107),
    .QN(_0583_));
 DFF_X1 _0937_ (.D(_0260_),
    .CK(clknet_4_9__leaf_clk),
    .Q(net108),
    .QN(_0584_));
 DFF_X2 _0938_ (.D(_0169_),
    .CK(clknet_4_14__leaf_clk),
    .Q(data_in_reg[0]),
    .QN(_0585_));
 DFF_X2 _0939_ (.D(_0180_),
    .CK(clknet_4_1__leaf_clk),
    .Q(data_in_reg[1]),
    .QN(_0586_));
 DFF_X2 _0940_ (.D(_0191_),
    .CK(clknet_4_9__leaf_clk),
    .Q(data_in_reg[2]),
    .QN(_0587_));
 DFF_X2 _0941_ (.D(_0194_),
    .CK(clknet_4_10__leaf_clk),
    .Q(data_in_reg[3]),
    .QN(_0588_));
 DFF_X2 _0942_ (.D(_0195_),
    .CK(clknet_4_0__leaf_clk),
    .Q(data_in_reg[4]),
    .QN(_0589_));
 DFF_X2 _0943_ (.D(_0196_),
    .CK(clknet_4_10__leaf_clk),
    .Q(data_in_reg[5]),
    .QN(_0590_));
 DFF_X2 _0944_ (.D(_0197_),
    .CK(clknet_4_12__leaf_clk),
    .Q(data_in_reg[6]),
    .QN(_0591_));
 DFF_X2 _0945_ (.D(_0198_),
    .CK(clknet_4_4__leaf_clk),
    .Q(data_in_reg[7]),
    .QN(_0592_));
 DFF_X2 _0946_ (.D(_0199_),
    .CK(clknet_4_10__leaf_clk),
    .Q(data_in_reg[8]),
    .QN(_0593_));
 DFF_X2 _0947_ (.D(_0200_),
    .CK(clknet_4_1__leaf_clk),
    .Q(data_in_reg[9]),
    .QN(_0594_));
 DFF_X2 _0948_ (.D(_0170_),
    .CK(clknet_4_10__leaf_clk),
    .Q(data_in_reg[10]),
    .QN(_0595_));
 DFF_X2 _0949_ (.D(_0171_),
    .CK(clknet_4_4__leaf_clk),
    .Q(data_in_reg[11]),
    .QN(_0596_));
 DFF_X2 _0950_ (.D(_0172_),
    .CK(clknet_4_14__leaf_clk),
    .Q(data_in_reg[12]),
    .QN(_0597_));
 DFF_X2 _0951_ (.D(_0173_),
    .CK(clknet_4_1__leaf_clk),
    .Q(data_in_reg[13]),
    .QN(_0598_));
 DFF_X2 _0952_ (.D(_0174_),
    .CK(clknet_4_10__leaf_clk),
    .Q(data_in_reg[14]),
    .QN(_0599_));
 DFF_X2 _0953_ (.D(_0175_),
    .CK(clknet_4_10__leaf_clk),
    .Q(data_in_reg[15]),
    .QN(_0600_));
 DFF_X2 _0954_ (.D(_0176_),
    .CK(clknet_4_1__leaf_clk),
    .Q(data_in_reg[16]),
    .QN(_0601_));
 DFF_X2 _0955_ (.D(_0177_),
    .CK(clknet_4_1__leaf_clk),
    .Q(data_in_reg[17]),
    .QN(_0602_));
 DFF_X2 _0956_ (.D(_0178_),
    .CK(clknet_4_2__leaf_clk),
    .Q(data_in_reg[18]),
    .QN(_0603_));
 DFF_X2 _0957_ (.D(_0179_),
    .CK(clknet_4_5__leaf_clk),
    .Q(data_in_reg[19]),
    .QN(_0604_));
 DFF_X2 _0958_ (.D(_0181_),
    .CK(clknet_4_5__leaf_clk),
    .Q(data_in_reg[20]),
    .QN(_0605_));
 DFF_X2 _0959_ (.D(_0182_),
    .CK(clknet_4_5__leaf_clk),
    .Q(data_in_reg[21]),
    .QN(_0606_));
 DFF_X2 _0960_ (.D(_0183_),
    .CK(clknet_4_10__leaf_clk),
    .Q(data_in_reg[22]),
    .QN(_0607_));
 DFF_X2 _0961_ (.D(_0184_),
    .CK(clknet_4_2__leaf_clk),
    .Q(data_in_reg[23]),
    .QN(_0608_));
 DFF_X2 _0962_ (.D(_0185_),
    .CK(clknet_4_10__leaf_clk),
    .Q(data_in_reg[24]),
    .QN(_0609_));
 DFF_X2 _0963_ (.D(_0186_),
    .CK(clknet_4_0__leaf_clk),
    .Q(data_in_reg[25]),
    .QN(_0610_));
 DFF_X2 _0964_ (.D(_0187_),
    .CK(clknet_4_3__leaf_clk),
    .Q(data_in_reg[26]),
    .QN(_0611_));
 DFF_X2 _0965_ (.D(_0188_),
    .CK(clknet_4_0__leaf_clk),
    .Q(data_in_reg[27]),
    .QN(_0612_));
 DFF_X2 _0966_ (.D(_0189_),
    .CK(clknet_4_14__leaf_clk),
    .Q(data_in_reg[28]),
    .QN(_0613_));
 DFF_X2 _0967_ (.D(_0190_),
    .CK(clknet_4_14__leaf_clk),
    .Q(data_in_reg[29]),
    .QN(_0614_));
 DFF_X2 _0968_ (.D(_0192_),
    .CK(clknet_4_0__leaf_clk),
    .Q(data_in_reg[30]),
    .QN(_0615_));
 DFF_X2 _0969_ (.D(_0193_),
    .CK(clknet_4_11__leaf_clk),
    .Q(data_in_reg[31]),
    .QN(_0616_));
 DFF_X2 _0970_ (.D(_0271_),
    .CK(clknet_4_3__leaf_clk),
    .Q(sram_rdata_reg[0]),
    .QN(_0617_));
 DFF_X2 _0971_ (.D(_0282_),
    .CK(clknet_4_12__leaf_clk),
    .Q(sram_rdata_reg[1]),
    .QN(_0618_));
 DFF_X2 _0972_ (.D(_0293_),
    .CK(clknet_4_12__leaf_clk),
    .Q(sram_rdata_reg[2]),
    .QN(_0619_));
 DFF_X2 _0973_ (.D(_0296_),
    .CK(clknet_4_12__leaf_clk),
    .Q(sram_rdata_reg[3]),
    .QN(_0620_));
 DFF_X2 _0974_ (.D(_0297_),
    .CK(clknet_4_12__leaf_clk),
    .Q(sram_rdata_reg[4]),
    .QN(_0621_));
 DFF_X2 _0975_ (.D(_0298_),
    .CK(clknet_4_12__leaf_clk),
    .Q(sram_rdata_reg[5]),
    .QN(_0622_));
 DFF_X2 _0976_ (.D(_0299_),
    .CK(clknet_4_12__leaf_clk),
    .Q(sram_rdata_reg[6]),
    .QN(_0623_));
 DFF_X2 _0977_ (.D(_0300_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[7]),
    .QN(_0624_));
 DFF_X2 _0978_ (.D(_0301_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[8]),
    .QN(_0625_));
 DFF_X2 _0979_ (.D(_0302_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[9]),
    .QN(_0626_));
 DFF_X2 _0980_ (.D(_0272_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[10]),
    .QN(_0627_));
 DFF_X2 _0981_ (.D(_0273_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[11]),
    .QN(_0628_));
 DFF_X2 _0982_ (.D(_0274_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[12]),
    .QN(_0629_));
 DFF_X2 _0983_ (.D(_0275_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[13]),
    .QN(_0630_));
 DFF_X2 _0984_ (.D(_0276_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[14]),
    .QN(_0631_));
 DFF_X2 _0985_ (.D(_0277_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[15]),
    .QN(_0632_));
 DFF_X2 _0986_ (.D(_0278_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[16]),
    .QN(_0633_));
 DFF_X2 _0987_ (.D(_0279_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[17]),
    .QN(_0634_));
 DFF_X2 _0988_ (.D(_0280_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[18]),
    .QN(_0635_));
 DFF_X2 _0989_ (.D(_0281_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[19]),
    .QN(_0636_));
 DFF_X2 _0990_ (.D(_0283_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[20]),
    .QN(_0637_));
 DFF_X2 _0991_ (.D(_0284_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[21]),
    .QN(_0638_));
 DFF_X2 _0992_ (.D(_0285_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[22]),
    .QN(_0639_));
 DFF_X2 _0993_ (.D(_0286_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[23]),
    .QN(_0640_));
 DFF_X2 _0994_ (.D(_0287_),
    .CK(clknet_4_13__leaf_clk),
    .Q(sram_rdata_reg[24]),
    .QN(_0641_));
 DFF_X2 _0995_ (.D(_0288_),
    .CK(clknet_4_15__leaf_clk),
    .Q(sram_rdata_reg[25]),
    .QN(_0642_));
 DFF_X2 _0996_ (.D(_0289_),
    .CK(clknet_4_15__leaf_clk),
    .Q(sram_rdata_reg[26]),
    .QN(_0643_));
 DFF_X2 _0997_ (.D(_0290_),
    .CK(clknet_4_15__leaf_clk),
    .Q(sram_rdata_reg[27]),
    .QN(_0644_));
 DFF_X2 _0998_ (.D(_0291_),
    .CK(clknet_4_15__leaf_clk),
    .Q(sram_rdata_reg[28]),
    .QN(_0645_));
 DFF_X2 _0999_ (.D(_0292_),
    .CK(clknet_4_15__leaf_clk),
    .Q(sram_rdata_reg[29]),
    .QN(_0646_));
 DFF_X2 _1000_ (.D(_0294_),
    .CK(clknet_4_15__leaf_clk),
    .Q(sram_rdata_reg[30]),
    .QN(_0647_));
 DFF_X2 _1001_ (.D(_0295_),
    .CK(clknet_4_15__leaf_clk),
    .Q(sram_rdata_reg[31]),
    .QN(_0648_));
 DFF_X2 _1002_ (.D(net9),
    .CK(clknet_4_11__leaf_clk),
    .Q(net113),
    .QN(_0649_));
 DFF_X2 _1003_ (.D(net210),
    .CK(clknet_4_7__leaf_clk),
    .Q(addr_ptr[0]),
    .QN(_0650_));
 DFF_X1 _1004_ (.D(_0164_),
    .CK(clknet_4_7__leaf_clk),
    .Q(addr_ptr[1]),
    .QN(_0651_));
 DFF_X1 _1005_ (.D(_0165_),
    .CK(clknet_4_7__leaf_clk),
    .Q(addr_ptr[2]),
    .QN(_0652_));
 DFF_X1 _1006_ (.D(_0166_),
    .CK(clknet_4_7__leaf_clk),
    .Q(addr_ptr[3]),
    .QN(_0653_));
 DFF_X1 _1007_ (.D(_0167_),
    .CK(clknet_4_7__leaf_clk),
    .Q(addr_ptr[4]),
    .QN(_0654_));
 DFF_X1 _1008_ (.D(net181),
    .CK(clknet_4_7__leaf_clk),
    .Q(addr_ptr[5]),
    .QN(_0655_));
 DFF_X1 _1009_ (.D(net186),
    .CK(clknet_4_6__leaf_clk),
    .Q(init_count[0]),
    .QN(_0656_));
 DFF_X1 _1010_ (.D(_0266_),
    .CK(clknet_4_6__leaf_clk),
    .Q(init_count[1]),
    .QN(_0657_));
 DFF_X1 _1011_ (.D(net194),
    .CK(clknet_4_6__leaf_clk),
    .Q(init_count[2]),
    .QN(_0658_));
 DFF_X2 _1012_ (.D(net205),
    .CK(clknet_4_6__leaf_clk),
    .Q(init_count[3]),
    .QN(_0659_));
 DFF_X1 _1013_ (.D(net197),
    .CK(clknet_4_6__leaf_clk),
    .Q(init_count[4]),
    .QN(_0660_));
 DFF_X1 _1014_ (.D(net191),
    .CK(clknet_4_6__leaf_clk),
    .Q(init_count[5]),
    .QN(_0661_));
 SRAM_6T_CORE_64x32_MC_TB sram_inst (.ce_in(_0307_),
    .we_in(_0308_),
    .clk(clknet_4_3__leaf_clk),
    .addr_in({net188,
    net183,
    net4,
    net6,
    net212,
    net179}),
    .rd_out({sram_rdata[31],
    sram_rdata[30],
    sram_rdata[29],
    sram_rdata[28],
    sram_rdata[27],
    sram_rdata[26],
    sram_rdata[25],
    sram_rdata[24],
    sram_rdata[23],
    sram_rdata[22],
    sram_rdata[21],
    sram_rdata[20],
    sram_rdata[19],
    sram_rdata[18],
    sram_rdata[17],
    sram_rdata[16],
    sram_rdata[15],
    sram_rdata[14],
    sram_rdata[13],
    sram_rdata[12],
    sram_rdata[11],
    sram_rdata[10],
    sram_rdata[9],
    sram_rdata[8],
    sram_rdata[7],
    sram_rdata[6],
    sram_rdata[5],
    sram_rdata[4],
    sram_rdata[3],
    sram_rdata[2],
    sram_rdata[1],
    sram_rdata[0]}),
    .wd_in({net224,
    data_in_reg[30],
    net231,
    net227,
    data_in_reg[27],
    data_in_reg[26],
    data_in_reg[25],
    net226,
    data_in_reg[23],
    net228,
    data_in_reg[21],
    data_in_reg[20],
    data_in_reg[19],
    net230,
    data_in_reg[17],
    data_in_reg[16],
    net218,
    net225,
    data_in_reg[13],
    net223,
    data_in_reg[11],
    net232,
    data_in_reg[9],
    data_in_reg[8],
    data_in_reg[7],
    net219,
    data_in_reg[5],
    data_in_reg[4],
    data_in_reg[3],
    net221,
    net229,
    net222}));
 AND2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_40_  (.A1(net147),
    .A2(\u_multiplier/pp3_0 ),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_25_ ));
 OR2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_41_  (.A1(net148),
    .A2(\u_multiplier/pp3_0 ),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_26_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_42_  (.A(net149),
    .B(\u_multiplier/pp3_0 ),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_27_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_43_  (.A(net161),
    .B(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_27_ ),
    .ZN(product[0]));
 AOI21_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_44_  (.A(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_25_ ),
    .B1(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_26_ ),
    .B2(net162),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_28_ ));
 NOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_45_  (.A1(net150),
    .A2(\u_multiplier/A [1]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_29_ ));
 NAND2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_46_  (.A1(net151),
    .A2(\u_multiplier/A [1]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_30_ ));
 XOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_47_  (.A(net152),
    .B(\u_multiplier/A [1]),
    .Z(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_31_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_48_  (.A(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_28_ ),
    .B(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_31_ ),
    .ZN(product[1]));
 OAI21_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_49_  (.A(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_30_ ),
    .B1(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_29_ ),
    .B2(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_28_ ),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_32_ ));
 AND2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_50_  (.A1(net153),
    .A2(\u_multiplier/A [2]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_33_ ));
 OR2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_51_  (.A1(net154),
    .A2(\u_multiplier/A [2]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_34_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_52_  (.A(net155),
    .B(\u_multiplier/A [2]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_35_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_53_  (.A(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_32_ ),
    .B(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_35_ ),
    .ZN(product[2]));
 AOI21_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_54_  (.A(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_33_ ),
    .B1(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_34_ ),
    .B2(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_32_ ),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_36_ ));
 NOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_55_  (.A1(\u_multiplier/B [3]),
    .A2(\u_multiplier/A [3]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_37_ ));
 NAND2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_56_  (.A1(\u_multiplier/B [3]),
    .A2(\u_multiplier/A [3]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_38_ ));
 XOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_57_  (.A(\u_multiplier/B [3]),
    .B(\u_multiplier/A [3]),
    .Z(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_39_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_58_  (.A(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_36_ ),
    .B(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_39_ ),
    .ZN(product[3]));
 OAI21_X2 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_59_  (.A(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_38_ ),
    .B1(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_37_ ),
    .B2(\u_multiplier/Final_add/cla1/cla1/cla1/cla1/_36_ ),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla1/c1 ));
 AND2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_40_  (.A1(\u_multiplier/B [4]),
    .A2(\u_multiplier/A [4]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_25_ ));
 OR2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_41_  (.A1(\u_multiplier/B [4]),
    .A2(\u_multiplier/A [4]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_26_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_42_  (.A(\u_multiplier/B [4]),
    .B(\u_multiplier/A [4]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_27_ ));
 XNOR2_X2 \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_43_  (.A(\u_multiplier/Final_add/cla1/cla1/cla1/c1 ),
    .B(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_27_ ),
    .ZN(product[4]));
 AOI21_X2 \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_44_  (.A(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_25_ ),
    .B1(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_26_ ),
    .B2(\u_multiplier/Final_add/cla1/cla1/cla1/c1 ),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_28_ ));
 NOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_45_  (.A1(\u_multiplier/B [5]),
    .A2(\u_multiplier/A [5]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_29_ ));
 NAND2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_46_  (.A1(\u_multiplier/B [5]),
    .A2(\u_multiplier/A [5]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_30_ ));
 XOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_47_  (.A(\u_multiplier/B [5]),
    .B(\u_multiplier/A [5]),
    .Z(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_31_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_48_  (.A(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_28_ ),
    .B(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_31_ ),
    .ZN(product[5]));
 OAI21_X2 \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_49_  (.A(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_30_ ),
    .B1(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_29_ ),
    .B2(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_28_ ),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_32_ ));
 AND2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_50_  (.A1(\u_multiplier/B [6]),
    .A2(\u_multiplier/A [6]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_33_ ));
 OR2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_51_  (.A1(\u_multiplier/B [6]),
    .A2(\u_multiplier/A [6]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_34_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_52_  (.A(\u_multiplier/B [6]),
    .B(\u_multiplier/A [6]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_35_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_53_  (.A(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_32_ ),
    .B(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_35_ ),
    .ZN(product[6]));
 AOI21_X2 \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_54_  (.A(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_33_ ),
    .B1(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_34_ ),
    .B2(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_32_ ),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_36_ ));
 NOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_55_  (.A1(\u_multiplier/B [7]),
    .A2(\u_multiplier/A [7]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_37_ ));
 NAND2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_56_  (.A1(\u_multiplier/B [7]),
    .A2(\u_multiplier/A [7]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_38_ ));
 XOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_57_  (.A(\u_multiplier/B [7]),
    .B(\u_multiplier/A [7]),
    .Z(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_39_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_58_  (.A(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_36_ ),
    .B(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_39_ ),
    .ZN(product[7]));
 OAI21_X2 \u_multiplier/Final_add/cla1/cla1/cla1/cla2/_59_  (.A(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_38_ ),
    .B1(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_37_ ),
    .B2(\u_multiplier/Final_add/cla1/cla1/cla1/cla2/_36_ ),
    .ZN(\u_multiplier/Final_add/cla1/cla1/c1 ));
 AND2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_40_  (.A1(\u_multiplier/B [8]),
    .A2(\u_multiplier/A [8]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_25_ ));
 OR2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_41_  (.A1(\u_multiplier/B [8]),
    .A2(\u_multiplier/A [8]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_26_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_42_  (.A(\u_multiplier/B [8]),
    .B(\u_multiplier/A [8]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_27_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_43_  (.A(\u_multiplier/Final_add/cla1/cla1/c1 ),
    .B(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_27_ ),
    .ZN(product[8]));
 AOI21_X2 \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_44_  (.A(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_25_ ),
    .B1(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_26_ ),
    .B2(\u_multiplier/Final_add/cla1/cla1/c1 ),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_28_ ));
 NOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_45_  (.A1(\u_multiplier/B [9]),
    .A2(\u_multiplier/A [9]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_29_ ));
 NAND2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_46_  (.A1(\u_multiplier/B [9]),
    .A2(\u_multiplier/A [9]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_30_ ));
 XOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_47_  (.A(\u_multiplier/B [9]),
    .B(\u_multiplier/A [9]),
    .Z(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_31_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_48_  (.A(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_28_ ),
    .B(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_31_ ),
    .ZN(product[9]));
 OAI21_X2 \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_49_  (.A(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_30_ ),
    .B1(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_29_ ),
    .B2(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_28_ ),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_32_ ));
 AND2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_50_  (.A1(\u_multiplier/B [10]),
    .A2(\u_multiplier/A [10]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_33_ ));
 OR2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_51_  (.A1(\u_multiplier/B [10]),
    .A2(\u_multiplier/A [10]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_34_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_52_  (.A(\u_multiplier/B [10]),
    .B(\u_multiplier/A [10]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_35_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_53_  (.A(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_32_ ),
    .B(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_35_ ),
    .ZN(product[10]));
 AOI21_X2 \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_54_  (.A(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_33_ ),
    .B1(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_34_ ),
    .B2(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_32_ ),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_36_ ));
 NOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_55_  (.A1(\u_multiplier/B [11]),
    .A2(\u_multiplier/A [11]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_37_ ));
 NAND2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_56_  (.A1(\u_multiplier/B [11]),
    .A2(\u_multiplier/A [11]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_38_ ));
 XOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_57_  (.A(\u_multiplier/B [11]),
    .B(\u_multiplier/A [11]),
    .Z(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_39_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_58_  (.A(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_36_ ),
    .B(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_39_ ),
    .ZN(product[11]));
 OAI21_X2 \u_multiplier/Final_add/cla1/cla1/cla2/cla1/_59_  (.A(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_38_ ),
    .B1(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_37_ ),
    .B2(\u_multiplier/Final_add/cla1/cla1/cla2/cla1/_36_ ),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla2/c1 ));
 AND2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_40_  (.A1(\u_multiplier/B [12]),
    .A2(\u_multiplier/A [12]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_25_ ));
 OR2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_41_  (.A1(\u_multiplier/B [12]),
    .A2(\u_multiplier/A [12]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_26_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_42_  (.A(\u_multiplier/B [12]),
    .B(\u_multiplier/A [12]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_27_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_43_  (.A(\u_multiplier/Final_add/cla1/cla1/cla2/c1 ),
    .B(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_27_ ),
    .ZN(product[12]));
 AOI21_X2 \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_44_  (.A(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_25_ ),
    .B1(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_26_ ),
    .B2(\u_multiplier/Final_add/cla1/cla1/cla2/c1 ),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_28_ ));
 NOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_45_  (.A1(\u_multiplier/B [13]),
    .A2(\u_multiplier/A [13]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_29_ ));
 NAND2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_46_  (.A1(\u_multiplier/B [13]),
    .A2(\u_multiplier/A [13]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_30_ ));
 XOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_47_  (.A(\u_multiplier/B [13]),
    .B(\u_multiplier/A [13]),
    .Z(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_31_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_48_  (.A(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_28_ ),
    .B(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_31_ ),
    .ZN(product[13]));
 OAI21_X2 \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_49_  (.A(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_30_ ),
    .B1(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_29_ ),
    .B2(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_28_ ),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_32_ ));
 AND2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_50_  (.A1(\u_multiplier/B [14]),
    .A2(\u_multiplier/A [14]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_33_ ));
 OR2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_51_  (.A1(\u_multiplier/B [14]),
    .A2(\u_multiplier/A [14]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_34_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_52_  (.A(\u_multiplier/B [14]),
    .B(\u_multiplier/A [14]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_35_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_53_  (.A(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_32_ ),
    .B(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_35_ ),
    .ZN(product[14]));
 AOI21_X2 \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_54_  (.A(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_33_ ),
    .B1(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_34_ ),
    .B2(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_32_ ),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_36_ ));
 NOR2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_55_  (.A1(\u_multiplier/B [15]),
    .A2(\u_multiplier/A [15]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_37_ ));
 NAND2_X1 \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_56_  (.A1(\u_multiplier/B [15]),
    .A2(\u_multiplier/A [15]),
    .ZN(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_38_ ));
 XOR2_X2 \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_57_  (.A(\u_multiplier/B [15]),
    .B(\u_multiplier/A [15]),
    .Z(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_39_ ));
 XNOR2_X2 \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_58_  (.A(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_36_ ),
    .B(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_39_ ),
    .ZN(product[15]));
 OAI21_X2 \u_multiplier/Final_add/cla1/cla1/cla2/cla2/_59_  (.A(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_38_ ),
    .B1(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_37_ ),
    .B2(\u_multiplier/Final_add/cla1/cla1/cla2/cla2/_36_ ),
    .ZN(\u_multiplier/Final_add/cla1/c1 ));
 AND2_X1 \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_40_  (.A1(\u_multiplier/B [16]),
    .A2(\u_multiplier/A [16]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_25_ ));
 OR2_X1 \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_41_  (.A1(\u_multiplier/B [16]),
    .A2(\u_multiplier/A [16]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_26_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_42_  (.A(\u_multiplier/B [16]),
    .B(\u_multiplier/A [16]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_27_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_43_  (.A(\u_multiplier/Final_add/cla1/c1 ),
    .B(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_27_ ),
    .ZN(product[16]));
 AOI21_X2 \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_44_  (.A(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_25_ ),
    .B1(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_26_ ),
    .B2(\u_multiplier/Final_add/cla1/c1 ),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_28_ ));
 NOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_45_  (.A1(\u_multiplier/B [17]),
    .A2(\u_multiplier/A [17]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_29_ ));
 NAND2_X1 \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_46_  (.A1(\u_multiplier/B [17]),
    .A2(\u_multiplier/A [17]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_30_ ));
 XOR2_X2 \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_47_  (.A(\u_multiplier/B [17]),
    .B(\u_multiplier/A [17]),
    .Z(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_31_ ));
 XNOR2_X2 \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_48_  (.A(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_28_ ),
    .B(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_31_ ),
    .ZN(product[17]));
 OAI21_X2 \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_49_  (.A(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_30_ ),
    .B1(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_29_ ),
    .B2(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_28_ ),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_32_ ));
 AND2_X1 \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_50_  (.A1(\u_multiplier/B [18]),
    .A2(\u_multiplier/A [18]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_33_ ));
 OR2_X1 \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_51_  (.A1(\u_multiplier/B [18]),
    .A2(\u_multiplier/A [18]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_34_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_52_  (.A(\u_multiplier/B [18]),
    .B(\u_multiplier/A [18]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_35_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_53_  (.A(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_32_ ),
    .B(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_35_ ),
    .ZN(product[18]));
 AOI21_X2 \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_54_  (.A(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_33_ ),
    .B1(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_34_ ),
    .B2(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_32_ ),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_36_ ));
 NOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_55_  (.A1(\u_multiplier/B [19]),
    .A2(\u_multiplier/A [19]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_37_ ));
 NAND2_X1 \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_56_  (.A1(\u_multiplier/B [19]),
    .A2(\u_multiplier/A [19]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_38_ ));
 XOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_57_  (.A(\u_multiplier/B [19]),
    .B(\u_multiplier/A [19]),
    .Z(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_39_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_58_  (.A(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_36_ ),
    .B(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_39_ ),
    .ZN(product[19]));
 OAI21_X2 \u_multiplier/Final_add/cla1/cla2/cla1/cla1/_59_  (.A(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_38_ ),
    .B1(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_37_ ),
    .B2(\u_multiplier/Final_add/cla1/cla2/cla1/cla1/_36_ ),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla1/c1 ));
 AND2_X1 \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_40_  (.A1(\u_multiplier/B [20]),
    .A2(\u_multiplier/A [20]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_25_ ));
 OR2_X1 \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_41_  (.A1(\u_multiplier/B [20]),
    .A2(\u_multiplier/A [20]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_26_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_42_  (.A(\u_multiplier/B [20]),
    .B(\u_multiplier/A [20]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_27_ ));
 XNOR2_X2 \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_43_  (.A(\u_multiplier/Final_add/cla1/cla2/cla1/c1 ),
    .B(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_27_ ),
    .ZN(product[20]));
 AOI21_X2 \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_44_  (.A(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_25_ ),
    .B1(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_26_ ),
    .B2(\u_multiplier/Final_add/cla1/cla2/cla1/c1 ),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_28_ ));
 NOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_45_  (.A1(\u_multiplier/B [21]),
    .A2(\u_multiplier/A [21]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_29_ ));
 NAND2_X1 \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_46_  (.A1(\u_multiplier/B [21]),
    .A2(\u_multiplier/A [21]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_30_ ));
 XOR2_X2 \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_47_  (.A(\u_multiplier/B [21]),
    .B(\u_multiplier/A [21]),
    .Z(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_31_ ));
 XNOR2_X2 \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_48_  (.A(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_28_ ),
    .B(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_31_ ),
    .ZN(product[21]));
 OAI21_X2 \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_49_  (.A(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_30_ ),
    .B1(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_29_ ),
    .B2(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_28_ ),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_32_ ));
 AND2_X1 \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_50_  (.A1(\u_multiplier/B [22]),
    .A2(\u_multiplier/A [22]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_33_ ));
 OR2_X1 \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_51_  (.A1(\u_multiplier/B [22]),
    .A2(\u_multiplier/A [22]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_34_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_52_  (.A(\u_multiplier/B [22]),
    .B(\u_multiplier/A [22]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_35_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_53_  (.A(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_32_ ),
    .B(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_35_ ),
    .ZN(product[22]));
 AOI21_X2 \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_54_  (.A(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_33_ ),
    .B1(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_34_ ),
    .B2(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_32_ ),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_36_ ));
 NOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_55_  (.A1(\u_multiplier/B [23]),
    .A2(\u_multiplier/A [23]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_37_ ));
 NAND2_X1 \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_56_  (.A1(\u_multiplier/B [23]),
    .A2(\u_multiplier/A [23]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_38_ ));
 XOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_57_  (.A(\u_multiplier/B [23]),
    .B(\u_multiplier/A [23]),
    .Z(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_39_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_58_  (.A(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_36_ ),
    .B(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_39_ ),
    .ZN(product[23]));
 OAI21_X2 \u_multiplier/Final_add/cla1/cla2/cla1/cla2/_59_  (.A(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_38_ ),
    .B1(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_37_ ),
    .B2(\u_multiplier/Final_add/cla1/cla2/cla1/cla2/_36_ ),
    .ZN(\u_multiplier/Final_add/cla1/cla2/c1 ));
 AND2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_40_  (.A1(\u_multiplier/B [24]),
    .A2(\u_multiplier/A [24]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_25_ ));
 OR2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_41_  (.A1(\u_multiplier/B [24]),
    .A2(\u_multiplier/A [24]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_26_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_42_  (.A(\u_multiplier/B [24]),
    .B(\u_multiplier/A [24]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_27_ ));
 XNOR2_X2 \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_43_  (.A(\u_multiplier/Final_add/cla1/cla2/c1 ),
    .B(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_27_ ),
    .ZN(product[24]));
 AOI21_X2 \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_44_  (.A(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_25_ ),
    .B1(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_26_ ),
    .B2(\u_multiplier/Final_add/cla1/cla2/c1 ),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_28_ ));
 NOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_45_  (.A1(\u_multiplier/B [25]),
    .A2(\u_multiplier/A [25]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_29_ ));
 NAND2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_46_  (.A1(\u_multiplier/B [25]),
    .A2(\u_multiplier/A [25]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_30_ ));
 XOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_47_  (.A(\u_multiplier/B [25]),
    .B(\u_multiplier/A [25]),
    .Z(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_31_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_48_  (.A(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_28_ ),
    .B(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_31_ ),
    .ZN(product[25]));
 OAI21_X2 \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_49_  (.A(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_30_ ),
    .B1(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_29_ ),
    .B2(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_28_ ),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_32_ ));
 AND2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_50_  (.A1(\u_multiplier/B [26]),
    .A2(\u_multiplier/A [26]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_33_ ));
 OR2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_51_  (.A1(\u_multiplier/B [26]),
    .A2(\u_multiplier/A [26]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_34_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_52_  (.A(\u_multiplier/B [26]),
    .B(\u_multiplier/A [26]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_35_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_53_  (.A(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_32_ ),
    .B(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_35_ ),
    .ZN(product[26]));
 AOI21_X2 \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_54_  (.A(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_33_ ),
    .B1(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_34_ ),
    .B2(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_32_ ),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_36_ ));
 NOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_55_  (.A1(\u_multiplier/B [27]),
    .A2(\u_multiplier/A [27]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_37_ ));
 NAND2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_56_  (.A1(\u_multiplier/B [27]),
    .A2(\u_multiplier/A [27]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_38_ ));
 XOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_57_  (.A(\u_multiplier/B [27]),
    .B(\u_multiplier/A [27]),
    .Z(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_39_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_58_  (.A(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_36_ ),
    .B(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_39_ ),
    .ZN(product[27]));
 OAI21_X2 \u_multiplier/Final_add/cla1/cla2/cla2/cla1/_59_  (.A(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_38_ ),
    .B1(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_37_ ),
    .B2(\u_multiplier/Final_add/cla1/cla2/cla2/cla1/_36_ ),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla2/c1 ));
 AND2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_40_  (.A1(\u_multiplier/B [28]),
    .A2(\u_multiplier/A [28]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_25_ ));
 OR2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_41_  (.A1(\u_multiplier/B [28]),
    .A2(\u_multiplier/A [28]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_26_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_42_  (.A(\u_multiplier/B [28]),
    .B(\u_multiplier/A [28]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_27_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_43_  (.A(\u_multiplier/Final_add/cla1/cla2/cla2/c1 ),
    .B(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_27_ ),
    .ZN(product[28]));
 AOI21_X4 \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_44_  (.A(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_25_ ),
    .B1(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_26_ ),
    .B2(\u_multiplier/Final_add/cla1/cla2/cla2/c1 ),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_28_ ));
 NOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_45_  (.A1(\u_multiplier/B [29]),
    .A2(\u_multiplier/A [29]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_29_ ));
 NAND2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_46_  (.A1(\u_multiplier/B [29]),
    .A2(\u_multiplier/A [29]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_30_ ));
 XOR2_X2 \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_47_  (.A(\u_multiplier/B [29]),
    .B(\u_multiplier/A [29]),
    .Z(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_31_ ));
 XNOR2_X2 \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_48_  (.A(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_28_ ),
    .B(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_31_ ),
    .ZN(product[29]));
 OAI21_X2 \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_49_  (.A(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_30_ ),
    .B1(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_29_ ),
    .B2(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_28_ ),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_32_ ));
 AND2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_50_  (.A1(\u_multiplier/B [30]),
    .A2(\u_multiplier/A [30]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_33_ ));
 OR2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_51_  (.A1(\u_multiplier/B [30]),
    .A2(\u_multiplier/A [30]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_34_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_52_  (.A(\u_multiplier/B [30]),
    .B(\u_multiplier/A [30]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_35_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_53_  (.A(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_32_ ),
    .B(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_35_ ),
    .ZN(product[30]));
 AOI21_X4 \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_54_  (.A(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_33_ ),
    .B1(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_34_ ),
    .B2(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_32_ ),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_36_ ));
 NOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_55_  (.A1(\u_multiplier/B [31]),
    .A2(\u_multiplier/A [31]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_37_ ));
 NAND2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_56_  (.A1(\u_multiplier/B [31]),
    .A2(\u_multiplier/A [31]),
    .ZN(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_38_ ));
 XOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_57_  (.A(\u_multiplier/B [31]),
    .B(\u_multiplier/A [31]),
    .Z(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_39_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_58_  (.A(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_36_ ),
    .B(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_39_ ),
    .ZN(product[31]));
 OAI21_X4 \u_multiplier/Final_add/cla1/cla2/cla2/cla2/_59_  (.A(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_38_ ),
    .B1(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_37_ ),
    .B2(\u_multiplier/Final_add/cla1/cla2/cla2/cla2/_36_ ),
    .ZN(\u_multiplier/Final_add/c1 ));
 AND2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_40_  (.A1(\u_multiplier/B [32]),
    .A2(\u_multiplier/A [32]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_25_ ));
 OR2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_41_  (.A1(\u_multiplier/B [32]),
    .A2(\u_multiplier/A [32]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_26_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_42_  (.A(\u_multiplier/B [32]),
    .B(\u_multiplier/A [32]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_27_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_43_  (.A(\u_multiplier/Final_add/c1 ),
    .B(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_27_ ),
    .ZN(product[32]));
 AOI21_X4 \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_44_  (.A(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_25_ ),
    .B1(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_26_ ),
    .B2(\u_multiplier/Final_add/c1 ),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_28_ ));
 NOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_45_  (.A1(\u_multiplier/B [33]),
    .A2(\u_multiplier/A [33]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_29_ ));
 NAND2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_46_  (.A1(\u_multiplier/B [33]),
    .A2(\u_multiplier/A [33]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_30_ ));
 XOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_47_  (.A(\u_multiplier/B [33]),
    .B(\u_multiplier/A [33]),
    .Z(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_31_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_48_  (.A(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_28_ ),
    .B(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_31_ ),
    .ZN(product[33]));
 OAI21_X4 \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_49_  (.A(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_30_ ),
    .B1(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_29_ ),
    .B2(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_28_ ),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_32_ ));
 AND2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_50_  (.A1(\u_multiplier/B [34]),
    .A2(\u_multiplier/A [34]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_33_ ));
 OR2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_51_  (.A1(\u_multiplier/B [34]),
    .A2(\u_multiplier/A [34]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_34_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_52_  (.A(\u_multiplier/B [34]),
    .B(\u_multiplier/A [34]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_35_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_53_  (.A(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_32_ ),
    .B(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_35_ ),
    .ZN(product[34]));
 AOI21_X2 \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_54_  (.A(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_33_ ),
    .B1(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_34_ ),
    .B2(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_32_ ),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_36_ ));
 NOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_55_  (.A1(\u_multiplier/B [35]),
    .A2(\u_multiplier/A [35]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_37_ ));
 NAND2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_56_  (.A1(\u_multiplier/B [35]),
    .A2(\u_multiplier/A [35]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_38_ ));
 XOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_57_  (.A(\u_multiplier/B [35]),
    .B(\u_multiplier/A [35]),
    .Z(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_39_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_58_  (.A(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_36_ ),
    .B(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_39_ ),
    .ZN(product[35]));
 OAI21_X2 \u_multiplier/Final_add/cla2/cla1/cla1/cla1/_59_  (.A(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_38_ ),
    .B1(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_37_ ),
    .B2(\u_multiplier/Final_add/cla2/cla1/cla1/cla1/_36_ ),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla1/c1 ));
 AND2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_40_  (.A1(\u_multiplier/B [36]),
    .A2(\u_multiplier/A [36]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_25_ ));
 OR2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_41_  (.A1(\u_multiplier/B [36]),
    .A2(\u_multiplier/A [36]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_26_ ));
 XNOR2_X2 \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_42_  (.A(\u_multiplier/B [36]),
    .B(\u_multiplier/A [36]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_27_ ));
 XNOR2_X2 \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_43_  (.A(\u_multiplier/Final_add/cla2/cla1/cla1/c1 ),
    .B(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_27_ ),
    .ZN(product[36]));
 AOI21_X2 \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_44_  (.A(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_25_ ),
    .B1(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_26_ ),
    .B2(\u_multiplier/Final_add/cla2/cla1/cla1/c1 ),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_28_ ));
 NOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_45_  (.A1(\u_multiplier/B [37]),
    .A2(\u_multiplier/A [37]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_29_ ));
 NAND2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_46_  (.A1(\u_multiplier/B [37]),
    .A2(\u_multiplier/A [37]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_30_ ));
 XOR2_X2 \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_47_  (.A(\u_multiplier/B [37]),
    .B(\u_multiplier/A [37]),
    .Z(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_31_ ));
 XNOR2_X2 \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_48_  (.A(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_28_ ),
    .B(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_31_ ),
    .ZN(product[37]));
 OAI21_X2 \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_49_  (.A(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_30_ ),
    .B1(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_29_ ),
    .B2(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_28_ ),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_32_ ));
 AND2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_50_  (.A1(\u_multiplier/B [38]),
    .A2(\u_multiplier/A [38]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_33_ ));
 OR2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_51_  (.A1(\u_multiplier/B [38]),
    .A2(\u_multiplier/A [38]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_34_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_52_  (.A(\u_multiplier/B [38]),
    .B(\u_multiplier/A [38]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_35_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_53_  (.A(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_32_ ),
    .B(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_35_ ),
    .ZN(product[38]));
 AOI21_X2 \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_54_  (.A(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_33_ ),
    .B1(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_34_ ),
    .B2(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_32_ ),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_36_ ));
 NOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_55_  (.A1(\u_multiplier/B [39]),
    .A2(\u_multiplier/A [39]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_37_ ));
 NAND2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_56_  (.A1(\u_multiplier/B [39]),
    .A2(\u_multiplier/A [39]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_38_ ));
 XOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_57_  (.A(\u_multiplier/B [39]),
    .B(\u_multiplier/A [39]),
    .Z(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_39_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_58_  (.A(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_36_ ),
    .B(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_39_ ),
    .ZN(product[39]));
 OAI21_X2 \u_multiplier/Final_add/cla2/cla1/cla1/cla2/_59_  (.A(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_38_ ),
    .B1(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_37_ ),
    .B2(\u_multiplier/Final_add/cla2/cla1/cla1/cla2/_36_ ),
    .ZN(\u_multiplier/Final_add/cla2/cla1/c1 ));
 AND2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_40_  (.A1(\u_multiplier/B [40]),
    .A2(\u_multiplier/A [40]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_25_ ));
 OR2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_41_  (.A1(\u_multiplier/B [40]),
    .A2(\u_multiplier/A [40]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_26_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_42_  (.A(\u_multiplier/B [40]),
    .B(\u_multiplier/A [40]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_27_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_43_  (.A(\u_multiplier/Final_add/cla2/cla1/c1 ),
    .B(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_27_ ),
    .ZN(product[40]));
 AOI21_X2 \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_44_  (.A(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_25_ ),
    .B1(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_26_ ),
    .B2(\u_multiplier/Final_add/cla2/cla1/c1 ),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_28_ ));
 NOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_45_  (.A1(\u_multiplier/B [41]),
    .A2(\u_multiplier/A [41]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_29_ ));
 NAND2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_46_  (.A1(\u_multiplier/B [41]),
    .A2(\u_multiplier/A [41]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_30_ ));
 XOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_47_  (.A(\u_multiplier/B [41]),
    .B(\u_multiplier/A [41]),
    .Z(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_31_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_48_  (.A(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_28_ ),
    .B(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_31_ ),
    .ZN(product[41]));
 OAI21_X2 \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_49_  (.A(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_30_ ),
    .B1(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_29_ ),
    .B2(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_28_ ),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_32_ ));
 AND2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_50_  (.A1(\u_multiplier/B [42]),
    .A2(\u_multiplier/A [42]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_33_ ));
 OR2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_51_  (.A1(\u_multiplier/B [42]),
    .A2(\u_multiplier/A [42]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_34_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_52_  (.A(\u_multiplier/B [42]),
    .B(\u_multiplier/A [42]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_35_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_53_  (.A(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_32_ ),
    .B(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_35_ ),
    .ZN(product[42]));
 AOI21_X4 \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_54_  (.A(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_33_ ),
    .B1(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_34_ ),
    .B2(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_32_ ),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_36_ ));
 NOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_55_  (.A1(\u_multiplier/B [43]),
    .A2(\u_multiplier/A [43]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_37_ ));
 NAND2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_56_  (.A1(\u_multiplier/B [43]),
    .A2(\u_multiplier/A [43]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_38_ ));
 XOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_57_  (.A(\u_multiplier/B [43]),
    .B(\u_multiplier/A [43]),
    .Z(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_39_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_58_  (.A(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_36_ ),
    .B(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_39_ ),
    .ZN(product[43]));
 OAI21_X2 \u_multiplier/Final_add/cla2/cla1/cla2/cla1/_59_  (.A(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_38_ ),
    .B1(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_37_ ),
    .B2(\u_multiplier/Final_add/cla2/cla1/cla2/cla1/_36_ ),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla2/c1 ));
 AND2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_40_  (.A1(\u_multiplier/B [44]),
    .A2(\u_multiplier/A [44]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_25_ ));
 OR2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_41_  (.A1(\u_multiplier/B [44]),
    .A2(\u_multiplier/A [44]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_26_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_42_  (.A(\u_multiplier/B [44]),
    .B(\u_multiplier/A [44]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_27_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_43_  (.A(\u_multiplier/Final_add/cla2/cla1/cla2/c1 ),
    .B(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_27_ ),
    .ZN(product[44]));
 AOI21_X2 \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_44_  (.A(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_25_ ),
    .B1(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_26_ ),
    .B2(\u_multiplier/Final_add/cla2/cla1/cla2/c1 ),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_28_ ));
 NOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_45_  (.A1(\u_multiplier/B [45]),
    .A2(\u_multiplier/A [45]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_29_ ));
 NAND2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_46_  (.A1(\u_multiplier/B [45]),
    .A2(\u_multiplier/A [45]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_30_ ));
 XOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_47_  (.A(\u_multiplier/B [45]),
    .B(\u_multiplier/A [45]),
    .Z(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_31_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_48_  (.A(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_28_ ),
    .B(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_31_ ),
    .ZN(product[45]));
 OAI21_X2 \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_49_  (.A(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_30_ ),
    .B1(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_29_ ),
    .B2(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_28_ ),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_32_ ));
 AND2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_50_  (.A1(\u_multiplier/B [46]),
    .A2(\u_multiplier/A [46]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_33_ ));
 OR2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_51_  (.A1(\u_multiplier/B [46]),
    .A2(\u_multiplier/A [46]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_34_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_52_  (.A(\u_multiplier/B [46]),
    .B(\u_multiplier/A [46]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_35_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_53_  (.A(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_32_ ),
    .B(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_35_ ),
    .ZN(product[46]));
 AOI21_X2 \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_54_  (.A(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_33_ ),
    .B1(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_34_ ),
    .B2(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_32_ ),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_36_ ));
 NOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_55_  (.A1(\u_multiplier/B [47]),
    .A2(\u_multiplier/A [47]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_37_ ));
 NAND2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_56_  (.A1(\u_multiplier/B [47]),
    .A2(\u_multiplier/A [47]),
    .ZN(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_38_ ));
 XOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_57_  (.A(\u_multiplier/B [47]),
    .B(\u_multiplier/A [47]),
    .Z(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_39_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_58_  (.A(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_36_ ),
    .B(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_39_ ),
    .ZN(product[47]));
 OAI21_X2 \u_multiplier/Final_add/cla2/cla1/cla2/cla2/_59_  (.A(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_38_ ),
    .B1(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_37_ ),
    .B2(\u_multiplier/Final_add/cla2/cla1/cla2/cla2/_36_ ),
    .ZN(\u_multiplier/Final_add/cla2/c1 ));
 AND2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_40_  (.A1(\u_multiplier/B [48]),
    .A2(\u_multiplier/A [48]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_25_ ));
 OR2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_41_  (.A1(\u_multiplier/B [48]),
    .A2(\u_multiplier/A [48]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_26_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_42_  (.A(\u_multiplier/B [48]),
    .B(\u_multiplier/A [48]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_27_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_43_  (.A(\u_multiplier/Final_add/cla2/c1 ),
    .B(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_27_ ),
    .ZN(product[48]));
 AOI21_X2 \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_44_  (.A(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_25_ ),
    .B1(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_26_ ),
    .B2(\u_multiplier/Final_add/cla2/c1 ),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_28_ ));
 NOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_45_  (.A1(\u_multiplier/B [49]),
    .A2(\u_multiplier/A [49]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_29_ ));
 NAND2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_46_  (.A1(\u_multiplier/B [49]),
    .A2(\u_multiplier/A [49]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_30_ ));
 XOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_47_  (.A(\u_multiplier/B [49]),
    .B(\u_multiplier/A [49]),
    .Z(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_31_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_48_  (.A(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_28_ ),
    .B(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_31_ ),
    .ZN(product[49]));
 OAI21_X2 \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_49_  (.A(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_30_ ),
    .B1(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_29_ ),
    .B2(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_28_ ),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_32_ ));
 AND2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_50_  (.A1(\u_multiplier/B [50]),
    .A2(\u_multiplier/A [50]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_33_ ));
 OR2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_51_  (.A1(\u_multiplier/B [50]),
    .A2(\u_multiplier/A [50]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_34_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_52_  (.A(\u_multiplier/B [50]),
    .B(\u_multiplier/A [50]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_35_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_53_  (.A(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_32_ ),
    .B(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_35_ ),
    .ZN(product[50]));
 AOI21_X2 \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_54_  (.A(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_33_ ),
    .B1(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_34_ ),
    .B2(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_32_ ),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_36_ ));
 NOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_55_  (.A1(\u_multiplier/B [51]),
    .A2(\u_multiplier/A [51]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_37_ ));
 NAND2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_56_  (.A1(\u_multiplier/B [51]),
    .A2(\u_multiplier/A [51]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_38_ ));
 XOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_57_  (.A(\u_multiplier/B [51]),
    .B(\u_multiplier/A [51]),
    .Z(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_39_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_58_  (.A(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_36_ ),
    .B(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_39_ ),
    .ZN(product[51]));
 OAI21_X2 \u_multiplier/Final_add/cla2/cla2/cla1/cla1/_59_  (.A(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_38_ ),
    .B1(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_37_ ),
    .B2(\u_multiplier/Final_add/cla2/cla2/cla1/cla1/_36_ ),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla1/c1 ));
 AND2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_40_  (.A1(\u_multiplier/B [52]),
    .A2(\u_multiplier/A [52]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_25_ ));
 OR2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_41_  (.A1(\u_multiplier/B [52]),
    .A2(\u_multiplier/A [52]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_26_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_42_  (.A(\u_multiplier/B [52]),
    .B(\u_multiplier/A [52]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_27_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_43_  (.A(\u_multiplier/Final_add/cla2/cla2/cla1/c1 ),
    .B(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_27_ ),
    .ZN(product[52]));
 AOI21_X4 \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_44_  (.A(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_25_ ),
    .B1(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_26_ ),
    .B2(\u_multiplier/Final_add/cla2/cla2/cla1/c1 ),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_28_ ));
 NOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_45_  (.A1(\u_multiplier/B [53]),
    .A2(\u_multiplier/A [53]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_29_ ));
 NAND2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_46_  (.A1(\u_multiplier/B [53]),
    .A2(\u_multiplier/A [53]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_30_ ));
 XOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_47_  (.A(\u_multiplier/B [53]),
    .B(\u_multiplier/A [53]),
    .Z(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_31_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_48_  (.A(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_28_ ),
    .B(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_31_ ),
    .ZN(product[53]));
 OAI21_X4 \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_49_  (.A(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_30_ ),
    .B1(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_29_ ),
    .B2(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_28_ ),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_32_ ));
 AND2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_50_  (.A1(\u_multiplier/B [54]),
    .A2(\u_multiplier/A [54]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_33_ ));
 OR2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_51_  (.A1(\u_multiplier/B [54]),
    .A2(\u_multiplier/A [54]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_34_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_52_  (.A(\u_multiplier/B [54]),
    .B(\u_multiplier/A [54]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_35_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_53_  (.A(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_32_ ),
    .B(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_35_ ),
    .ZN(product[54]));
 AOI21_X4 \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_54_  (.A(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_33_ ),
    .B1(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_34_ ),
    .B2(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_32_ ),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_36_ ));
 NOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_55_  (.A1(\u_multiplier/B [55]),
    .A2(\u_multiplier/A [55]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_37_ ));
 NAND2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_56_  (.A1(\u_multiplier/B [55]),
    .A2(\u_multiplier/A [55]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_38_ ));
 XOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_57_  (.A(\u_multiplier/B [55]),
    .B(\u_multiplier/A [55]),
    .Z(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_39_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_58_  (.A(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_36_ ),
    .B(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_39_ ),
    .ZN(product[55]));
 OAI21_X4 \u_multiplier/Final_add/cla2/cla2/cla1/cla2/_59_  (.A(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_38_ ),
    .B1(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_37_ ),
    .B2(\u_multiplier/Final_add/cla2/cla2/cla1/cla2/_36_ ),
    .ZN(\u_multiplier/Final_add/cla2/cla2/c1 ));
 AND2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_40_  (.A1(\u_multiplier/B [56]),
    .A2(\u_multiplier/A [56]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_25_ ));
 OR2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_41_  (.A1(\u_multiplier/B [56]),
    .A2(\u_multiplier/A [56]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_26_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_42_  (.A(\u_multiplier/B [56]),
    .B(\u_multiplier/A [56]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_27_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_43_  (.A(\u_multiplier/Final_add/cla2/cla2/c1 ),
    .B(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_27_ ),
    .ZN(product[56]));
 AOI21_X2 \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_44_  (.A(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_25_ ),
    .B1(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_26_ ),
    .B2(\u_multiplier/Final_add/cla2/cla2/c1 ),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_28_ ));
 NOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_45_  (.A1(\u_multiplier/B [57]),
    .A2(\u_multiplier/A [57]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_29_ ));
 NAND2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_46_  (.A1(\u_multiplier/B [57]),
    .A2(\u_multiplier/A [57]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_30_ ));
 XOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_47_  (.A(\u_multiplier/B [57]),
    .B(\u_multiplier/A [57]),
    .Z(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_31_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_48_  (.A(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_28_ ),
    .B(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_31_ ),
    .ZN(product[57]));
 OAI21_X2 \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_49_  (.A(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_30_ ),
    .B1(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_29_ ),
    .B2(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_28_ ),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_32_ ));
 AND2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_50_  (.A1(\u_multiplier/B [58]),
    .A2(\u_multiplier/A [58]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_33_ ));
 OR2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_51_  (.A1(\u_multiplier/B [58]),
    .A2(\u_multiplier/A [58]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_34_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_52_  (.A(\u_multiplier/B [58]),
    .B(\u_multiplier/A [58]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_35_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_53_  (.A(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_32_ ),
    .B(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_35_ ),
    .ZN(product[58]));
 AOI21_X2 \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_54_  (.A(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_33_ ),
    .B1(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_34_ ),
    .B2(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_32_ ),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_36_ ));
 NOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_55_  (.A1(\u_multiplier/B [59]),
    .A2(\u_multiplier/A [59]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_37_ ));
 NAND2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_56_  (.A1(\u_multiplier/B [59]),
    .A2(\u_multiplier/A [59]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_38_ ));
 XOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_57_  (.A(\u_multiplier/B [59]),
    .B(\u_multiplier/A [59]),
    .Z(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_39_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_58_  (.A(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_36_ ),
    .B(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_39_ ),
    .ZN(product[59]));
 OAI21_X2 \u_multiplier/Final_add/cla2/cla2/cla2/cla1/_59_  (.A(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_38_ ),
    .B1(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_37_ ),
    .B2(\u_multiplier/Final_add/cla2/cla2/cla2/cla1/_36_ ),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla2/c1 ));
 AND2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_40_  (.A1(\u_multiplier/B [60]),
    .A2(\u_multiplier/A [60]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_25_ ));
 OR2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_41_  (.A1(\u_multiplier/B [60]),
    .A2(\u_multiplier/A [60]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_26_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_42_  (.A(\u_multiplier/B [60]),
    .B(\u_multiplier/A [60]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_27_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_43_  (.A(\u_multiplier/Final_add/cla2/cla2/cla2/c1 ),
    .B(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_27_ ),
    .ZN(product[60]));
 AOI21_X2 \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_44_  (.A(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_25_ ),
    .B1(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_26_ ),
    .B2(\u_multiplier/Final_add/cla2/cla2/cla2/c1 ),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_28_ ));
 NOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_45_  (.A1(\u_multiplier/B [61]),
    .A2(\u_multiplier/A [61]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_29_ ));
 NAND2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_46_  (.A1(\u_multiplier/B [61]),
    .A2(\u_multiplier/A [61]),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_30_ ));
 XOR2_X2 \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_47_  (.A(\u_multiplier/B [61]),
    .B(\u_multiplier/A [61]),
    .Z(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_31_ ));
 XNOR2_X2 \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_48_  (.A(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_28_ ),
    .B(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_31_ ),
    .ZN(product[61]));
 OAI21_X2 \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_49_  (.A(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_30_ ),
    .B1(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_29_ ),
    .B2(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_28_ ),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_32_ ));
 AND2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_50_  (.A1(\u_multiplier/B [62]),
    .A2(\u_multiplier/pp3_62 ),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_33_ ));
 OR2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_51_  (.A1(\u_multiplier/B [62]),
    .A2(\u_multiplier/pp3_62 ),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_34_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_52_  (.A(\u_multiplier/B [62]),
    .B(\u_multiplier/pp3_62 ),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_35_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_53_  (.A(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_32_ ),
    .B(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_35_ ),
    .ZN(product[62]));
 AOI21_X4 \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_54_  (.A(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_33_ ),
    .B1(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_34_ ),
    .B2(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_32_ ),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_36_ ));
 NOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_55_  (.A1(net156),
    .A2(net140),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_37_ ));
 NAND2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_56_  (.A1(net157),
    .A2(net141),
    .ZN(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_38_ ));
 XOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_57_  (.A(net158),
    .B(net142),
    .Z(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_39_ ));
 XNOR2_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_58_  (.A(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_36_ ),
    .B(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_39_ ),
    .ZN(product[63]));
 OAI21_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_59_  (.A(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_38_ ),
    .B1(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_37_ ),
    .B2(\u_multiplier/Final_add/cla2/cla2/cla2/cla2/_36_ ),
    .ZN(\u_multiplier/Final_add/Cout ));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_17_1/_18_  (.A(net114),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_1/_19_  (.A1(\u_multiplier/STAGE1/_0610_ ),
    .A2(\u_multiplier/STAGE1/_0609_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_1/_20_  (.A(\u_multiplier/STAGE1/_0610_ ),
    .B(\u_multiplier/STAGE1/_0609_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_17_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_1/_21_  (.A1(\u_multiplier/STAGE1/_0611_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_17_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_1/_22_  (.A(\u_multiplier/STAGE1/_0611_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_17_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_17_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_1/_23_  (.A1(\u_multiplier/STAGE1/_0612_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_17_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_1/_24_  (.A(\u_multiplier/STAGE1/_0612_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_17_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_17_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_17_1/_25_  (.A(net115),
    .B(\u_multiplier/STAGE1/E_4_2_pp_17_1/_16_ ),
    .ZN(\u_multiplier/pp1_17 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_17_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_17_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_17_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_17_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_17_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_17_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_17_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_17_1/_17_ ),
    .ZN(\u_multiplier/pp1_18 [2]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_18_1/_18_  (.A(\u_multiplier/STAGE1/pp1_17_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_18_1/_19_  (.A1(\u_multiplier/STAGE1/_0614_ ),
    .A2(\u_multiplier/STAGE1/_0613_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_1/_20_  (.A(\u_multiplier/STAGE1/_0614_ ),
    .B(\u_multiplier/STAGE1/_0613_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_18_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_18_1/_21_  (.A1(\u_multiplier/STAGE1/_0615_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_18_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_1/_22_  (.A(\u_multiplier/STAGE1/_0615_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_18_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_18_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_18_1/_23_  (.A1(\u_multiplier/STAGE1/_0616_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_18_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_1/_24_  (.A(\u_multiplier/STAGE1/_0616_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_18_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_18_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_18_1/_25_  (.A(\u_multiplier/STAGE1/pp1_17_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_18_1/_16_ ),
    .ZN(\u_multiplier/pp1_18 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_18_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_18_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_18_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_18_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_18_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_18_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_18_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_18_1/_17_ ),
    .ZN(\u_multiplier/pp1_19 [3]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_19_1/_18_  (.A(\u_multiplier/STAGE1/pp1_18_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_19_1/_19_  (.A1(\u_multiplier/STAGE1/_0620_ ),
    .A2(\u_multiplier/STAGE1/_0619_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_19_1/_20_  (.A(\u_multiplier/STAGE1/_0620_ ),
    .B(\u_multiplier/STAGE1/_0619_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_19_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_19_1/_21_  (.A1(\u_multiplier/STAGE1/_0621_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_19_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_19_1/_22_  (.A(\u_multiplier/STAGE1/_0621_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_19_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_19_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_19_1/_23_  (.A1(\u_multiplier/STAGE1/_0622_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_19_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_19_1/_24_  (.A(\u_multiplier/STAGE1/_0622_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_19_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_19_1/_25_  (.A(\u_multiplier/STAGE1/pp1_18_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_19_1/_16_ ),
    .ZN(\u_multiplier/pp1_19 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_19_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_19_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_19_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_19_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_19_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_19_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_19_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_19_1/_17_ ),
    .ZN(\u_multiplier/pp1_20 [4]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_19_2/_18_  (.A(net116),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_19_2/_19_  (.A1(\u_multiplier/STAGE1/_0624_ ),
    .A2(\u_multiplier/STAGE1/_0623_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_19_2/_20_  (.A(\u_multiplier/STAGE1/_0624_ ),
    .B(\u_multiplier/STAGE1/_0623_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_19_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_19_2/_21_  (.A1(\u_multiplier/STAGE1/_0625_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_19_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_19_2/_22_  (.A(\u_multiplier/STAGE1/_0625_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_19_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_19_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_19_2/_23_  (.A1(\u_multiplier/STAGE1/_0626_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_19_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_19_2/_24_  (.A(\u_multiplier/STAGE1/_0626_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_19_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_19_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_19_2/_25_  (.A(net117),
    .B(\u_multiplier/STAGE1/E_4_2_pp_19_2/_16_ ),
    .ZN(\u_multiplier/pp1_19 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_19_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_19_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_19_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_19_e42_2_cout ));
 OAI21_X1 \u_multiplier/STAGE1/E_4_2_pp_19_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_19_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_19_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_19_2/_17_ ),
    .ZN(\u_multiplier/pp1_20 [3]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_20_1/_18_  (.A(\u_multiplier/STAGE1/pp1_19_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_20_1/_19_  (.A1(\u_multiplier/STAGE1/_0628_ ),
    .A2(\u_multiplier/STAGE1/_0627_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_20_1/_20_  (.A(\u_multiplier/STAGE1/_0628_ ),
    .B(\u_multiplier/STAGE1/_0627_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_20_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_20_1/_21_  (.A1(\u_multiplier/STAGE1/_0629_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_20_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_20_1/_22_  (.A(\u_multiplier/STAGE1/_0629_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_20_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_20_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_20_1/_23_  (.A1(\u_multiplier/STAGE1/_0630_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_20_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_20_1/_24_  (.A(\u_multiplier/STAGE1/_0630_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_20_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_20_1/_25_  (.A(\u_multiplier/STAGE1/pp1_19_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_20_1/_16_ ),
    .ZN(\u_multiplier/pp1_20 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_20_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_20_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_20_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_20_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_20_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_20_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_20_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_20_1/_17_ ),
    .ZN(\u_multiplier/pp1_21 [5]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_20_2/_18_  (.A(\u_multiplier/STAGE1/pp1_19_e42_2_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_20_2/_19_  (.A1(\u_multiplier/STAGE1/_0632_ ),
    .A2(\u_multiplier/STAGE1/_0631_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_20_2/_20_  (.A(\u_multiplier/STAGE1/_0632_ ),
    .B(\u_multiplier/STAGE1/_0631_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_20_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_20_2/_21_  (.A1(\u_multiplier/STAGE1/_0633_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_20_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_20_2/_22_  (.A(\u_multiplier/STAGE1/_0633_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_20_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_20_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_20_2/_23_  (.A1(\u_multiplier/STAGE1/_0634_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_20_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_20_2/_24_  (.A(\u_multiplier/STAGE1/_0634_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_20_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_20_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_20_2/_25_  (.A(\u_multiplier/STAGE1/pp1_19_e42_2_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_20_2/_16_ ),
    .ZN(\u_multiplier/pp1_20 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_20_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_20_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_20_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_20_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_20_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_20_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_20_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_20_2/_17_ ),
    .ZN(\u_multiplier/pp1_21 [4]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_21_1/_18_  (.A(\u_multiplier/STAGE1/pp1_20_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_21_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_21_1/_19_  (.A1(\u_multiplier/STAGE1/_0638_ ),
    .A2(\u_multiplier/STAGE1/_0637_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_21_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_21_1/_20_  (.A(\u_multiplier/STAGE1/_0638_ ),
    .B(\u_multiplier/STAGE1/_0637_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_21_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_21_1/_21_  (.A1(\u_multiplier/STAGE1/_0639_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_21_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_21_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_21_1/_22_  (.A(\u_multiplier/STAGE1/_0639_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_21_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_21_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_21_1/_23_  (.A1(\u_multiplier/STAGE1/_0640_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_21_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_21_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_21_1/_24_  (.A(\u_multiplier/STAGE1/_0640_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_21_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_21_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_21_1/_25_  (.A(\u_multiplier/STAGE1/pp1_20_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_21_1/_16_ ),
    .ZN(\u_multiplier/pp1_21 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_21_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_21_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_21_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_21_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_21_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_21_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_21_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_21_1/_17_ ),
    .ZN(\u_multiplier/pp1_22 [6]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_21_2/_18_  (.A(\u_multiplier/STAGE1/pp1_20_e42_2_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_21_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_21_2/_19_  (.A1(\u_multiplier/STAGE1/_0642_ ),
    .A2(\u_multiplier/STAGE1/_0641_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_21_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_21_2/_20_  (.A(\u_multiplier/STAGE1/_0642_ ),
    .B(\u_multiplier/STAGE1/_0641_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_21_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_21_2/_21_  (.A1(\u_multiplier/STAGE1/_0643_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_21_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_21_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_21_2/_22_  (.A(\u_multiplier/STAGE1/_0643_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_21_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_21_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_21_2/_23_  (.A1(\u_multiplier/STAGE1/_0644_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_21_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_21_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_21_2/_24_  (.A(\u_multiplier/STAGE1/_0644_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_21_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_21_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_21_2/_25_  (.A(\u_multiplier/STAGE1/pp1_20_e42_2_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_21_2/_16_ ),
    .ZN(\u_multiplier/pp1_21 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_21_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_21_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_21_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_21_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_21_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_21_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_21_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_21_2/_17_ ),
    .ZN(\u_multiplier/pp1_22 [5]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_21_3/_18_  (.A(net118),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_21_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_21_3/_19_  (.A1(\u_multiplier/STAGE1/_0646_ ),
    .A2(\u_multiplier/STAGE1/_0645_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_21_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_21_3/_20_  (.A(\u_multiplier/STAGE1/_0646_ ),
    .B(\u_multiplier/STAGE1/_0645_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_21_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_21_3/_21_  (.A1(\u_multiplier/STAGE1/_0647_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_21_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_21_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_21_3/_22_  (.A(\u_multiplier/STAGE1/_0647_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_21_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_21_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_21_3/_23_  (.A1(\u_multiplier/STAGE1/_0648_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_21_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_21_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_21_3/_24_  (.A(\u_multiplier/STAGE1/_0648_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_21_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_21_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_21_3/_25_  (.A(net119),
    .B(\u_multiplier/STAGE1/E_4_2_pp_21_3/_16_ ),
    .ZN(\u_multiplier/pp1_21 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_21_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_21_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_21_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_21_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_21_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_21_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_21_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_21_3/_17_ ),
    .ZN(\u_multiplier/pp1_22 [4]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_22_1/_18_  (.A(\u_multiplier/STAGE1/pp1_21_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_22_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_22_1/_19_  (.A1(\u_multiplier/STAGE1/_0650_ ),
    .A2(\u_multiplier/STAGE1/_0649_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_22_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_22_1/_20_  (.A(\u_multiplier/STAGE1/_0650_ ),
    .B(\u_multiplier/STAGE1/_0649_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_22_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_22_1/_21_  (.A1(\u_multiplier/STAGE1/_0651_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_22_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_22_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_22_1/_22_  (.A(\u_multiplier/STAGE1/_0651_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_22_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_22_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_22_1/_23_  (.A1(\u_multiplier/STAGE1/_0652_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_22_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_22_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_22_1/_24_  (.A(\u_multiplier/STAGE1/_0652_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_22_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_22_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_22_1/_25_  (.A(\u_multiplier/STAGE1/pp1_21_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_22_1/_16_ ),
    .ZN(\u_multiplier/pp1_22 [3]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_22_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_22_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_22_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_22_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_22_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_22_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_22_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_22_1/_17_ ),
    .ZN(\u_multiplier/pp1_23 [7]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_22_2/_18_  (.A(\u_multiplier/STAGE1/pp1_21_e42_2_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_22_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_22_2/_19_  (.A1(\u_multiplier/STAGE1/_0654_ ),
    .A2(\u_multiplier/STAGE1/_0653_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_22_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_22_2/_20_  (.A(\u_multiplier/STAGE1/_0654_ ),
    .B(\u_multiplier/STAGE1/_0653_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_22_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_22_2/_21_  (.A1(\u_multiplier/STAGE1/_0655_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_22_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_22_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_22_2/_22_  (.A(\u_multiplier/STAGE1/_0655_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_22_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_22_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_22_2/_23_  (.A1(\u_multiplier/STAGE1/_0656_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_22_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_22_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_22_2/_24_  (.A(\u_multiplier/STAGE1/_0656_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_22_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_22_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_22_2/_25_  (.A(\u_multiplier/STAGE1/pp1_21_e42_2_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_22_2/_16_ ),
    .ZN(\u_multiplier/pp1_22 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_22_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_22_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_22_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_22_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_22_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_22_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_22_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_22_2/_17_ ),
    .ZN(\u_multiplier/pp1_23 [6]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_22_3/_18_  (.A(\u_multiplier/STAGE1/pp1_21_e42_3_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_22_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_22_3/_19_  (.A1(\u_multiplier/STAGE1/_0658_ ),
    .A2(\u_multiplier/STAGE1/_0657_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_22_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_22_3/_20_  (.A(\u_multiplier/STAGE1/_0658_ ),
    .B(\u_multiplier/STAGE1/_0657_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_22_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_22_3/_21_  (.A1(\u_multiplier/STAGE1/_0659_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_22_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_22_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_22_3/_22_  (.A(\u_multiplier/STAGE1/_0659_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_22_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_22_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_22_3/_23_  (.A1(\u_multiplier/STAGE1/_0660_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_22_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_22_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_22_3/_24_  (.A(\u_multiplier/STAGE1/_0660_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_22_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_22_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_22_3/_25_  (.A(\u_multiplier/STAGE1/pp1_21_e42_3_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_22_3/_16_ ),
    .ZN(\u_multiplier/pp1_22 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_22_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_22_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_22_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_22_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_22_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_22_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_22_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_22_3/_17_ ),
    .ZN(\u_multiplier/pp1_23 [5]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_23_1/_18_  (.A(\u_multiplier/STAGE1/pp1_22_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_23_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_23_1/_19_  (.A1(\u_multiplier/STAGE1/_0664_ ),
    .A2(\u_multiplier/STAGE1/_0663_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_23_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_23_1/_20_  (.A(\u_multiplier/STAGE1/_0664_ ),
    .B(\u_multiplier/STAGE1/_0663_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_23_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_23_1/_21_  (.A1(\u_multiplier/STAGE1/_0665_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_23_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_23_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_23_1/_22_  (.A(\u_multiplier/STAGE1/_0665_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_23_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_23_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_23_1/_23_  (.A1(\u_multiplier/STAGE1/_0666_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_23_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_23_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_23_1/_24_  (.A(\u_multiplier/STAGE1/_0666_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_23_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_23_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_23_1/_25_  (.A(\u_multiplier/STAGE1/pp1_22_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_23_1/_16_ ),
    .ZN(\u_multiplier/pp1_23 [3]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_23_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_23_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_23_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_23_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_23_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_23_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_23_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_23_1/_17_ ),
    .ZN(\u_multiplier/pp1_24 [8]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_23_2/_18_  (.A(\u_multiplier/STAGE1/pp1_22_e42_2_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_23_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_23_2/_19_  (.A1(\u_multiplier/STAGE1/_0668_ ),
    .A2(\u_multiplier/STAGE1/_0667_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_23_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_23_2/_20_  (.A(\u_multiplier/STAGE1/_0668_ ),
    .B(\u_multiplier/STAGE1/_0667_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_23_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_23_2/_21_  (.A1(\u_multiplier/STAGE1/_0669_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_23_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_23_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_23_2/_22_  (.A(\u_multiplier/STAGE1/_0669_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_23_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_23_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_23_2/_23_  (.A1(\u_multiplier/STAGE1/_0670_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_23_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_23_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_23_2/_24_  (.A(\u_multiplier/STAGE1/_0670_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_23_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_23_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_23_2/_25_  (.A(\u_multiplier/STAGE1/pp1_22_e42_2_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_23_2/_16_ ),
    .ZN(\u_multiplier/pp1_23 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_23_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_23_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_23_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_23_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_23_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_23_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_23_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_23_2/_17_ ),
    .ZN(\u_multiplier/pp1_24 [7]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_23_3/_18_  (.A(\u_multiplier/STAGE1/pp1_22_e42_3_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_23_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_23_3/_19_  (.A1(\u_multiplier/STAGE1/_0672_ ),
    .A2(\u_multiplier/STAGE1/_0671_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_23_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_23_3/_20_  (.A(\u_multiplier/STAGE1/_0672_ ),
    .B(\u_multiplier/STAGE1/_0671_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_23_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_23_3/_21_  (.A1(\u_multiplier/STAGE1/_0673_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_23_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_23_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_23_3/_22_  (.A(\u_multiplier/STAGE1/_0673_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_23_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_23_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_23_3/_23_  (.A1(\u_multiplier/STAGE1/_0674_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_23_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_23_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_23_3/_24_  (.A(\u_multiplier/STAGE1/_0674_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_23_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_23_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_23_3/_25_  (.A(\u_multiplier/STAGE1/pp1_22_e42_3_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_23_3/_16_ ),
    .ZN(\u_multiplier/pp1_23 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_23_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_23_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_23_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_23_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_23_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_23_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_23_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_23_3/_17_ ),
    .ZN(\u_multiplier/pp1_24 [6]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_23_4/_18_  (.A(net120),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_23_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_23_4/_19_  (.A1(\u_multiplier/STAGE1/_0676_ ),
    .A2(\u_multiplier/STAGE1/_0675_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_23_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_23_4/_20_  (.A(\u_multiplier/STAGE1/_0676_ ),
    .B(\u_multiplier/STAGE1/_0675_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_23_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_23_4/_21_  (.A1(\u_multiplier/STAGE1/_0677_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_23_4/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_23_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_23_4/_22_  (.A(\u_multiplier/STAGE1/_0677_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_23_4/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_23_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_23_4/_23_  (.A1(\u_multiplier/STAGE1/_0678_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_23_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_23_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_23_4/_24_  (.A(\u_multiplier/STAGE1/_0678_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_23_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_23_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_23_4/_25_  (.A(net121),
    .B(\u_multiplier/STAGE1/E_4_2_pp_23_4/_16_ ),
    .ZN(\u_multiplier/pp1_23 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_23_4/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_23_4/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_23_4/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_23_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_23_4/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_23_4/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_23_4/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_23_4/_17_ ),
    .ZN(\u_multiplier/pp1_24 [5]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_24_1/_18_  (.A(\u_multiplier/STAGE1/pp1_23_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_24_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_24_1/_19_  (.A1(\u_multiplier/STAGE1/_0680_ ),
    .A2(\u_multiplier/STAGE1/_0679_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_24_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_24_1/_20_  (.A(\u_multiplier/STAGE1/_0680_ ),
    .B(\u_multiplier/STAGE1/_0679_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_24_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_24_1/_21_  (.A1(\u_multiplier/STAGE1/_0681_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_24_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_24_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_24_1/_22_  (.A(\u_multiplier/STAGE1/_0681_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_24_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_24_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_24_1/_23_  (.A1(\u_multiplier/STAGE1/_0682_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_24_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_24_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_24_1/_24_  (.A(\u_multiplier/STAGE1/_0682_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_24_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_24_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_24_1/_25_  (.A(\u_multiplier/STAGE1/pp1_23_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_24_1/_16_ ),
    .ZN(\u_multiplier/pp1_24 [4]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_24_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_24_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_24_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_24_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_24_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_24_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_24_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_24_1/_17_ ),
    .ZN(\u_multiplier/pp1_25 [9]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_24_2/_18_  (.A(\u_multiplier/STAGE1/pp1_23_e42_2_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_24_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_24_2/_19_  (.A1(\u_multiplier/STAGE1/_0684_ ),
    .A2(\u_multiplier/STAGE1/_0683_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_24_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_24_2/_20_  (.A(\u_multiplier/STAGE1/_0684_ ),
    .B(\u_multiplier/STAGE1/_0683_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_24_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_24_2/_21_  (.A1(\u_multiplier/STAGE1/_0685_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_24_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_24_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_24_2/_22_  (.A(\u_multiplier/STAGE1/_0685_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_24_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_24_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_24_2/_23_  (.A1(\u_multiplier/STAGE1/_0686_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_24_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_24_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_24_2/_24_  (.A(\u_multiplier/STAGE1/_0686_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_24_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_24_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_24_2/_25_  (.A(\u_multiplier/STAGE1/pp1_23_e42_2_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_24_2/_16_ ),
    .ZN(\u_multiplier/pp1_24 [3]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_24_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_24_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_24_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_24_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_24_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_24_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_24_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_24_2/_17_ ),
    .ZN(\u_multiplier/pp1_25 [8]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_24_3/_18_  (.A(\u_multiplier/STAGE1/pp1_23_e42_3_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_24_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_24_3/_19_  (.A1(\u_multiplier/STAGE1/_0688_ ),
    .A2(\u_multiplier/STAGE1/_0687_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_24_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_24_3/_20_  (.A(\u_multiplier/STAGE1/_0688_ ),
    .B(\u_multiplier/STAGE1/_0687_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_24_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_24_3/_21_  (.A1(\u_multiplier/STAGE1/_0689_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_24_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_24_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_24_3/_22_  (.A(\u_multiplier/STAGE1/_0689_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_24_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_24_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_24_3/_23_  (.A1(\u_multiplier/STAGE1/_0690_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_24_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_24_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_24_3/_24_  (.A(\u_multiplier/STAGE1/_0690_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_24_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_24_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_24_3/_25_  (.A(\u_multiplier/STAGE1/pp1_23_e42_3_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_24_3/_16_ ),
    .ZN(\u_multiplier/pp1_24 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_24_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_24_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_24_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_24_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_24_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_24_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_24_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_24_3/_17_ ),
    .ZN(\u_multiplier/pp1_25 [7]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_24_4/_18_  (.A(\u_multiplier/STAGE1/pp1_23_e42_4_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_24_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_24_4/_19_  (.A1(\u_multiplier/STAGE1/_0692_ ),
    .A2(\u_multiplier/STAGE1/_0691_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_24_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_24_4/_20_  (.A(\u_multiplier/STAGE1/_0692_ ),
    .B(\u_multiplier/STAGE1/_0691_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_24_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_24_4/_21_  (.A1(\u_multiplier/STAGE1/_0693_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_24_4/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_24_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_24_4/_22_  (.A(\u_multiplier/STAGE1/_0693_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_24_4/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_24_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_24_4/_23_  (.A1(\u_multiplier/STAGE1/_0694_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_24_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_24_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_24_4/_24_  (.A(\u_multiplier/STAGE1/_0694_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_24_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_24_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_24_4/_25_  (.A(\u_multiplier/STAGE1/pp1_23_e42_4_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_24_4/_16_ ),
    .ZN(\u_multiplier/pp1_24 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_24_4/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_24_4/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_24_4/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_24_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_24_4/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_24_4/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_24_4/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_24_4/_17_ ),
    .ZN(\u_multiplier/pp1_25 [6]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_25_1/_18_  (.A(\u_multiplier/STAGE1/pp1_24_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_25_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_25_1/_19_  (.A1(\u_multiplier/STAGE1/_0698_ ),
    .A2(\u_multiplier/STAGE1/_0697_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_25_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_25_1/_20_  (.A(\u_multiplier/STAGE1/_0698_ ),
    .B(\u_multiplier/STAGE1/_0697_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_25_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_25_1/_21_  (.A1(\u_multiplier/STAGE1/_0699_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_25_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_25_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_25_1/_22_  (.A(\u_multiplier/STAGE1/_0699_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_25_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_25_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_25_1/_23_  (.A1(\u_multiplier/STAGE1/_0700_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_25_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_25_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_25_1/_24_  (.A(\u_multiplier/STAGE1/_0700_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_25_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_25_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_25_1/_25_  (.A(\u_multiplier/STAGE1/pp1_24_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_25_1/_16_ ),
    .ZN(\u_multiplier/pp1_25 [4]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_25_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_25_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_25_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_25_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_25_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_25_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_25_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_25_1/_17_ ),
    .ZN(\u_multiplier/pp1_26 [10]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_25_2/_18_  (.A(\u_multiplier/STAGE1/pp1_24_e42_2_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_25_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_25_2/_19_  (.A1(\u_multiplier/STAGE1/_0702_ ),
    .A2(\u_multiplier/STAGE1/_0701_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_25_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_25_2/_20_  (.A(\u_multiplier/STAGE1/_0702_ ),
    .B(\u_multiplier/STAGE1/_0701_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_25_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_25_2/_21_  (.A1(\u_multiplier/STAGE1/_0703_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_25_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_25_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_25_2/_22_  (.A(\u_multiplier/STAGE1/_0703_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_25_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_25_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_25_2/_23_  (.A1(\u_multiplier/STAGE1/_0704_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_25_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_25_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_25_2/_24_  (.A(\u_multiplier/STAGE1/_0704_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_25_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_25_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_25_2/_25_  (.A(\u_multiplier/STAGE1/pp1_24_e42_2_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_25_2/_16_ ),
    .ZN(\u_multiplier/pp1_25 [3]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_25_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_25_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_25_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_25_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_25_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_25_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_25_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_25_2/_17_ ),
    .ZN(\u_multiplier/pp1_26 [9]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_25_3/_18_  (.A(\u_multiplier/STAGE1/pp1_24_e42_3_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_25_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_25_3/_19_  (.A1(\u_multiplier/STAGE1/_0706_ ),
    .A2(\u_multiplier/STAGE1/_0705_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_25_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_25_3/_20_  (.A(\u_multiplier/STAGE1/_0706_ ),
    .B(\u_multiplier/STAGE1/_0705_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_25_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_25_3/_21_  (.A1(\u_multiplier/STAGE1/_0707_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_25_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_25_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_25_3/_22_  (.A(\u_multiplier/STAGE1/_0707_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_25_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_25_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_25_3/_23_  (.A1(\u_multiplier/STAGE1/_0708_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_25_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_25_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_25_3/_24_  (.A(\u_multiplier/STAGE1/_0708_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_25_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_25_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_25_3/_25_  (.A(\u_multiplier/STAGE1/pp1_24_e42_3_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_25_3/_16_ ),
    .ZN(\u_multiplier/pp1_25 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_25_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_25_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_25_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_25_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_25_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_25_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_25_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_25_3/_17_ ),
    .ZN(\u_multiplier/pp1_26 [8]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_25_4/_18_  (.A(\u_multiplier/STAGE1/pp1_24_e42_4_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_25_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_25_4/_19_  (.A1(\u_multiplier/STAGE1/_0710_ ),
    .A2(\u_multiplier/STAGE1/_0709_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_25_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_25_4/_20_  (.A(\u_multiplier/STAGE1/_0710_ ),
    .B(\u_multiplier/STAGE1/_0709_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_25_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_25_4/_21_  (.A1(\u_multiplier/STAGE1/_0711_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_25_4/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_25_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_25_4/_22_  (.A(\u_multiplier/STAGE1/_0711_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_25_4/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_25_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_25_4/_23_  (.A1(\u_multiplier/STAGE1/_0712_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_25_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_25_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_25_4/_24_  (.A(\u_multiplier/STAGE1/_0712_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_25_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_25_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_25_4/_25_  (.A(\u_multiplier/STAGE1/pp1_24_e42_4_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_25_4/_16_ ),
    .ZN(\u_multiplier/pp1_25 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_25_4/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_25_4/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_25_4/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_25_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_25_4/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_25_4/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_25_4/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_25_4/_17_ ),
    .ZN(\u_multiplier/pp1_26 [7]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_25_5/_18_  (.A(net122),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_25_5/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_25_5/_19_  (.A1(\u_multiplier/STAGE1/_0714_ ),
    .A2(\u_multiplier/STAGE1/_0713_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_25_5/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_25_5/_20_  (.A(\u_multiplier/STAGE1/_0714_ ),
    .B(\u_multiplier/STAGE1/_0713_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_25_5/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_25_5/_21_  (.A1(\u_multiplier/STAGE1/_0715_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_25_5/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_25_5/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_25_5/_22_  (.A(\u_multiplier/STAGE1/_0715_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_25_5/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_25_5/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_25_5/_23_  (.A1(\u_multiplier/STAGE1/_0716_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_25_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_25_5/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_25_5/_24_  (.A(\u_multiplier/STAGE1/_0716_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_25_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_25_5/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_25_5/_25_  (.A(net123),
    .B(\u_multiplier/STAGE1/E_4_2_pp_25_5/_16_ ),
    .ZN(\u_multiplier/pp1_25 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_25_5/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_25_5/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_25_5/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_25_e42_5_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_25_5/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_25_5/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_25_5/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_25_5/_17_ ),
    .ZN(\u_multiplier/pp1_26 [6]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_26_1/_18_  (.A(\u_multiplier/STAGE1/pp1_25_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_26_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_26_1/_19_  (.A1(\u_multiplier/STAGE1/_0718_ ),
    .A2(\u_multiplier/STAGE1/_0717_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_26_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_26_1/_20_  (.A(\u_multiplier/STAGE1/_0718_ ),
    .B(\u_multiplier/STAGE1/_0717_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_26_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_26_1/_21_  (.A1(\u_multiplier/STAGE1/_0719_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_26_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_26_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_26_1/_22_  (.A(\u_multiplier/STAGE1/_0719_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_26_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_26_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_26_1/_23_  (.A1(\u_multiplier/STAGE1/_0720_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_26_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_26_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_26_1/_24_  (.A(\u_multiplier/STAGE1/_0720_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_26_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_26_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_26_1/_25_  (.A(\u_multiplier/STAGE1/pp1_25_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_26_1/_16_ ),
    .ZN(\u_multiplier/pp1_26 [5]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_26_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_26_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_26_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_26_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE1/E_4_2_pp_26_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_26_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_26_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_26_1/_17_ ),
    .ZN(\u_multiplier/pp1_27 [11]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_26_2/_18_  (.A(\u_multiplier/STAGE1/pp1_25_e42_2_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_26_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_26_2/_19_  (.A1(\u_multiplier/STAGE1/_0722_ ),
    .A2(\u_multiplier/STAGE1/_0721_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_26_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_26_2/_20_  (.A(\u_multiplier/STAGE1/_0722_ ),
    .B(\u_multiplier/STAGE1/_0721_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_26_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_26_2/_21_  (.A1(\u_multiplier/STAGE1/_0723_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_26_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_26_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_26_2/_22_  (.A(\u_multiplier/STAGE1/_0723_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_26_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_26_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_26_2/_23_  (.A1(\u_multiplier/STAGE1/_0724_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_26_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_26_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_26_2/_24_  (.A(\u_multiplier/STAGE1/_0724_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_26_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_26_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_26_2/_25_  (.A(\u_multiplier/STAGE1/pp1_25_e42_2_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_26_2/_16_ ),
    .ZN(\u_multiplier/pp1_26 [4]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_26_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_26_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_26_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_26_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_26_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_26_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_26_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_26_2/_17_ ),
    .ZN(\u_multiplier/pp1_27 [10]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_26_3/_18_  (.A(\u_multiplier/STAGE1/pp1_25_e42_3_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_26_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_26_3/_19_  (.A1(\u_multiplier/STAGE1/_0726_ ),
    .A2(\u_multiplier/STAGE1/_0725_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_26_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_26_3/_20_  (.A(\u_multiplier/STAGE1/_0726_ ),
    .B(\u_multiplier/STAGE1/_0725_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_26_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_26_3/_21_  (.A1(\u_multiplier/STAGE1/_0727_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_26_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_26_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_26_3/_22_  (.A(\u_multiplier/STAGE1/_0727_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_26_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_26_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_26_3/_23_  (.A1(\u_multiplier/STAGE1/_0728_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_26_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_26_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_26_3/_24_  (.A(\u_multiplier/STAGE1/_0728_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_26_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_26_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_26_3/_25_  (.A(\u_multiplier/STAGE1/pp1_25_e42_3_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_26_3/_16_ ),
    .ZN(\u_multiplier/pp1_26 [3]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_26_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_26_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_26_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_26_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_26_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_26_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_26_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_26_3/_17_ ),
    .ZN(\u_multiplier/pp1_27 [9]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_26_4/_18_  (.A(\u_multiplier/STAGE1/pp1_25_e42_4_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_26_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_26_4/_19_  (.A1(\u_multiplier/STAGE1/_0730_ ),
    .A2(\u_multiplier/STAGE1/_0729_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_26_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_26_4/_20_  (.A(\u_multiplier/STAGE1/_0730_ ),
    .B(\u_multiplier/STAGE1/_0729_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_26_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_26_4/_21_  (.A1(\u_multiplier/STAGE1/_0731_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_26_4/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_26_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_26_4/_22_  (.A(\u_multiplier/STAGE1/_0731_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_26_4/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_26_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_26_4/_23_  (.A1(\u_multiplier/STAGE1/_0732_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_26_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_26_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_26_4/_24_  (.A(\u_multiplier/STAGE1/_0732_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_26_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_26_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_26_4/_25_  (.A(\u_multiplier/STAGE1/pp1_25_e42_4_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_26_4/_16_ ),
    .ZN(\u_multiplier/pp1_26 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_26_4/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_26_4/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_26_4/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_26_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_26_4/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_26_4/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_26_4/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_26_4/_17_ ),
    .ZN(\u_multiplier/pp1_27 [8]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_26_5/_18_  (.A(\u_multiplier/STAGE1/pp1_25_e42_5_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_26_5/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_26_5/_19_  (.A1(\u_multiplier/STAGE1/_0734_ ),
    .A2(\u_multiplier/STAGE1/_0733_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_26_5/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_26_5/_20_  (.A(\u_multiplier/STAGE1/_0734_ ),
    .B(\u_multiplier/STAGE1/_0733_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_26_5/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_26_5/_21_  (.A1(\u_multiplier/STAGE1/_0735_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_26_5/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_26_5/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_26_5/_22_  (.A(\u_multiplier/STAGE1/_0735_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_26_5/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_26_5/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_26_5/_23_  (.A1(\u_multiplier/STAGE1/_0736_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_26_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_26_5/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_26_5/_24_  (.A(\u_multiplier/STAGE1/_0736_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_26_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_26_5/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_26_5/_25_  (.A(\u_multiplier/STAGE1/pp1_25_e42_5_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_26_5/_16_ ),
    .ZN(\u_multiplier/pp1_26 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_26_5/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_26_5/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_26_5/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_26_e42_5_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_26_5/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_26_5/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_26_5/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_26_5/_17_ ),
    .ZN(\u_multiplier/pp1_27 [7]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_27_1/_18_  (.A(\u_multiplier/STAGE1/pp1_26_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_27_1/_19_  (.A1(\u_multiplier/STAGE1/_0740_ ),
    .A2(\u_multiplier/STAGE1/_0739_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_27_1/_20_  (.A(\u_multiplier/STAGE1/_0740_ ),
    .B(\u_multiplier/STAGE1/_0739_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_27_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_27_1/_21_  (.A1(\u_multiplier/STAGE1/_0741_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_27_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_27_1/_22_  (.A(\u_multiplier/STAGE1/_0741_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_27_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_27_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_27_1/_23_  (.A1(\u_multiplier/STAGE1/_0742_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_27_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_27_1/_24_  (.A(\u_multiplier/STAGE1/_0742_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_27_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_27_1/_25_  (.A(\u_multiplier/STAGE1/pp1_26_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_27_1/_16_ ),
    .ZN(\u_multiplier/pp1_27 [5]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_27_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_27_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_27_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_27_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_27_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_27_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_27_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_27_1/_17_ ),
    .ZN(\u_multiplier/pp1_28 [12]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_27_2/_18_  (.A(\u_multiplier/STAGE1/pp1_26_e42_2_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_27_2/_19_  (.A1(\u_multiplier/STAGE1/_0744_ ),
    .A2(\u_multiplier/STAGE1/_0743_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_27_2/_20_  (.A(\u_multiplier/STAGE1/_0744_ ),
    .B(\u_multiplier/STAGE1/_0743_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_27_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_27_2/_21_  (.A1(\u_multiplier/STAGE1/_0745_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_27_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_27_2/_22_  (.A(\u_multiplier/STAGE1/_0745_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_27_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_27_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_27_2/_23_  (.A1(\u_multiplier/STAGE1/_0746_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_27_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_27_2/_24_  (.A(\u_multiplier/STAGE1/_0746_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_27_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_27_2/_25_  (.A(\u_multiplier/STAGE1/pp1_26_e42_2_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_27_2/_16_ ),
    .ZN(\u_multiplier/pp1_27 [4]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_27_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_27_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_27_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_27_e42_2_cout ));
 OAI21_X1 \u_multiplier/STAGE1/E_4_2_pp_27_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_27_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_27_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_27_2/_17_ ),
    .ZN(\u_multiplier/pp1_28 [11]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_27_3/_18_  (.A(\u_multiplier/STAGE1/pp1_26_e42_3_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_27_3/_19_  (.A1(\u_multiplier/STAGE1/_0748_ ),
    .A2(\u_multiplier/STAGE1/_0747_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_27_3/_20_  (.A(\u_multiplier/STAGE1/_0748_ ),
    .B(\u_multiplier/STAGE1/_0747_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_27_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_27_3/_21_  (.A1(\u_multiplier/STAGE1/_0749_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_27_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_27_3/_22_  (.A(\u_multiplier/STAGE1/_0749_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_27_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_27_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_27_3/_23_  (.A1(\u_multiplier/STAGE1/_0750_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_27_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_27_3/_24_  (.A(\u_multiplier/STAGE1/_0750_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_27_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_27_3/_25_  (.A(\u_multiplier/STAGE1/pp1_26_e42_3_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_27_3/_16_ ),
    .ZN(\u_multiplier/pp1_27 [3]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_27_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_27_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_27_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_27_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_27_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_27_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_27_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_27_3/_17_ ),
    .ZN(\u_multiplier/pp1_28 [10]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_27_4/_18_  (.A(\u_multiplier/STAGE1/pp1_26_e42_4_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_27_4/_19_  (.A1(\u_multiplier/STAGE1/_0752_ ),
    .A2(\u_multiplier/STAGE1/_0751_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_27_4/_20_  (.A(\u_multiplier/STAGE1/_0752_ ),
    .B(\u_multiplier/STAGE1/_0751_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_27_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_27_4/_21_  (.A1(\u_multiplier/STAGE1/_0753_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_27_4/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_27_4/_22_  (.A(\u_multiplier/STAGE1/_0753_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_27_4/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_27_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_27_4/_23_  (.A1(\u_multiplier/STAGE1/_0754_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_27_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_27_4/_24_  (.A(\u_multiplier/STAGE1/_0754_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_27_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_27_4/_25_  (.A(\u_multiplier/STAGE1/pp1_26_e42_4_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_27_4/_16_ ),
    .ZN(\u_multiplier/pp1_27 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_27_4/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_27_4/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_27_4/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_27_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_27_4/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_27_4/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_27_4/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_27_4/_17_ ),
    .ZN(\u_multiplier/pp1_28 [9]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_27_5/_18_  (.A(\u_multiplier/STAGE1/pp1_26_e42_5_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_5/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_27_5/_19_  (.A1(\u_multiplier/STAGE1/_0756_ ),
    .A2(\u_multiplier/STAGE1/_0755_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_5/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_27_5/_20_  (.A(\u_multiplier/STAGE1/_0756_ ),
    .B(\u_multiplier/STAGE1/_0755_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_27_5/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_27_5/_21_  (.A1(\u_multiplier/STAGE1/_0757_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_27_5/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_5/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_27_5/_22_  (.A(\u_multiplier/STAGE1/_0757_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_27_5/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_27_5/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_27_5/_23_  (.A1(\u_multiplier/STAGE1/_0758_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_27_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_5/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_27_5/_24_  (.A(\u_multiplier/STAGE1/_0758_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_27_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_5/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_27_5/_25_  (.A(\u_multiplier/STAGE1/pp1_26_e42_5_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_27_5/_16_ ),
    .ZN(\u_multiplier/pp1_27 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_27_5/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_27_5/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_27_5/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_27_e42_5_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_27_5/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_27_5/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_27_5/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_27_5/_17_ ),
    .ZN(\u_multiplier/pp1_28 [8]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_27_6/_18_  (.A(net124),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_6/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_27_6/_19_  (.A1(\u_multiplier/STAGE1/_0760_ ),
    .A2(\u_multiplier/STAGE1/_0759_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_6/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_27_6/_20_  (.A(\u_multiplier/STAGE1/_0760_ ),
    .B(\u_multiplier/STAGE1/_0759_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_27_6/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_27_6/_21_  (.A1(\u_multiplier/STAGE1/_0761_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_27_6/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_6/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_27_6/_22_  (.A(\u_multiplier/STAGE1/_0761_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_27_6/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_27_6/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_27_6/_23_  (.A1(\u_multiplier/STAGE1/_0762_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_27_6/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_6/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_27_6/_24_  (.A(\u_multiplier/STAGE1/_0762_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_27_6/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_27_6/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_27_6/_25_  (.A(net125),
    .B(\u_multiplier/STAGE1/E_4_2_pp_27_6/_16_ ),
    .ZN(\u_multiplier/pp1_27 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_27_6/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_27_6/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_27_6/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_27_e42_6_cout ));
 OAI21_X1 \u_multiplier/STAGE1/E_4_2_pp_27_6/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_27_6/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_27_6/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_27_6/_17_ ),
    .ZN(\u_multiplier/pp1_28 [7]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_28_1/_18_  (.A(\u_multiplier/STAGE1/pp1_27_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_28_1/_19_  (.A1(\u_multiplier/STAGE1/_0764_ ),
    .A2(\u_multiplier/STAGE1/_0763_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_28_1/_20_  (.A(\u_multiplier/STAGE1/_0764_ ),
    .B(\u_multiplier/STAGE1/_0763_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_28_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_28_1/_21_  (.A1(\u_multiplier/STAGE1/_0765_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_28_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_28_1/_22_  (.A(\u_multiplier/STAGE1/_0765_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_28_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_28_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_28_1/_23_  (.A1(\u_multiplier/STAGE1/_0766_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_28_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_28_1/_24_  (.A(\u_multiplier/STAGE1/_0766_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_28_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_28_1/_25_  (.A(\u_multiplier/STAGE1/pp1_27_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_28_1/_16_ ),
    .ZN(\u_multiplier/pp1_28 [6]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_28_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_28_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_28_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_28_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_28_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_28_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_28_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_28_1/_17_ ),
    .ZN(\u_multiplier/pp1_29 [13]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_28_2/_18_  (.A(\u_multiplier/STAGE1/pp1_27_e42_2_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_28_2/_19_  (.A1(\u_multiplier/STAGE1/_0768_ ),
    .A2(\u_multiplier/STAGE1/_0767_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_28_2/_20_  (.A(\u_multiplier/STAGE1/_0768_ ),
    .B(\u_multiplier/STAGE1/_0767_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_28_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_28_2/_21_  (.A1(\u_multiplier/STAGE1/_0769_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_28_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_28_2/_22_  (.A(\u_multiplier/STAGE1/_0769_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_28_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_28_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_28_2/_23_  (.A1(\u_multiplier/STAGE1/_0770_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_28_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_28_2/_24_  (.A(\u_multiplier/STAGE1/_0770_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_28_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_28_2/_25_  (.A(\u_multiplier/STAGE1/pp1_27_e42_2_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_28_2/_16_ ),
    .ZN(\u_multiplier/pp1_28 [5]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_28_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_28_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_28_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_28_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_28_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_28_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_28_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_28_2/_17_ ),
    .ZN(\u_multiplier/pp1_29 [12]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_28_3/_18_  (.A(\u_multiplier/STAGE1/pp1_27_e42_3_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_28_3/_19_  (.A1(\u_multiplier/STAGE1/_0772_ ),
    .A2(\u_multiplier/STAGE1/_0771_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_28_3/_20_  (.A(\u_multiplier/STAGE1/_0772_ ),
    .B(\u_multiplier/STAGE1/_0771_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_28_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_28_3/_21_  (.A1(\u_multiplier/STAGE1/_0773_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_28_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_28_3/_22_  (.A(\u_multiplier/STAGE1/_0773_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_28_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_28_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_28_3/_23_  (.A1(\u_multiplier/STAGE1/_0774_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_28_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_28_3/_24_  (.A(\u_multiplier/STAGE1/_0774_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_28_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_28_3/_25_  (.A(\u_multiplier/STAGE1/pp1_27_e42_3_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_28_3/_16_ ),
    .ZN(\u_multiplier/pp1_28 [4]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_28_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_28_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_28_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_28_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_28_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_28_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_28_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_28_3/_17_ ),
    .ZN(\u_multiplier/pp1_29 [11]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_28_4/_18_  (.A(\u_multiplier/STAGE1/pp1_27_e42_4_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_28_4/_19_  (.A1(\u_multiplier/STAGE1/_0776_ ),
    .A2(\u_multiplier/STAGE1/_0775_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_28_4/_20_  (.A(\u_multiplier/STAGE1/_0776_ ),
    .B(\u_multiplier/STAGE1/_0775_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_28_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_28_4/_21_  (.A1(\u_multiplier/STAGE1/_0777_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_28_4/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_28_4/_22_  (.A(\u_multiplier/STAGE1/_0777_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_28_4/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_28_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_28_4/_23_  (.A1(\u_multiplier/STAGE1/_0778_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_28_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_28_4/_24_  (.A(\u_multiplier/STAGE1/_0778_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_28_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_28_4/_25_  (.A(\u_multiplier/STAGE1/pp1_27_e42_4_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_28_4/_16_ ),
    .ZN(\u_multiplier/pp1_28 [3]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_28_4/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_28_4/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_28_4/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_28_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_28_4/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_28_4/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_28_4/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_28_4/_17_ ),
    .ZN(\u_multiplier/pp1_29 [10]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_28_5/_18_  (.A(\u_multiplier/STAGE1/pp1_27_e42_5_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_5/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_28_5/_19_  (.A1(\u_multiplier/STAGE1/_0780_ ),
    .A2(\u_multiplier/STAGE1/_0779_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_5/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_28_5/_20_  (.A(\u_multiplier/STAGE1/_0780_ ),
    .B(\u_multiplier/STAGE1/_0779_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_28_5/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_28_5/_21_  (.A1(\u_multiplier/STAGE1/_0781_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_28_5/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_5/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_28_5/_22_  (.A(\u_multiplier/STAGE1/_0781_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_28_5/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_28_5/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_28_5/_23_  (.A1(\u_multiplier/STAGE1/_0782_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_28_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_5/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_28_5/_24_  (.A(\u_multiplier/STAGE1/_0782_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_28_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_5/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_28_5/_25_  (.A(\u_multiplier/STAGE1/pp1_27_e42_5_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_28_5/_16_ ),
    .ZN(\u_multiplier/pp1_28 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_28_5/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_28_5/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_28_5/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_28_e42_5_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_28_5/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_28_5/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_28_5/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_28_5/_17_ ),
    .ZN(\u_multiplier/pp1_29 [9]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_28_6/_18_  (.A(\u_multiplier/STAGE1/pp1_27_e42_6_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_6/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_28_6/_19_  (.A1(\u_multiplier/STAGE1/_0784_ ),
    .A2(\u_multiplier/STAGE1/_0783_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_6/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_28_6/_20_  (.A(\u_multiplier/STAGE1/_0784_ ),
    .B(\u_multiplier/STAGE1/_0783_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_28_6/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_28_6/_21_  (.A1(\u_multiplier/STAGE1/_0785_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_28_6/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_6/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_28_6/_22_  (.A(\u_multiplier/STAGE1/_0785_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_28_6/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_28_6/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_28_6/_23_  (.A1(\u_multiplier/STAGE1/_0786_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_28_6/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_6/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_28_6/_24_  (.A(\u_multiplier/STAGE1/_0786_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_28_6/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_28_6/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_28_6/_25_  (.A(\u_multiplier/STAGE1/pp1_27_e42_6_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_28_6/_16_ ),
    .ZN(\u_multiplier/pp1_28 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_28_6/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_28_6/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_28_6/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_28_e42_6_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_28_6/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_28_6/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_28_6/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_28_6/_17_ ),
    .ZN(\u_multiplier/pp1_29 [8]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_29_1/_18_  (.A(\u_multiplier/STAGE1/pp1_28_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_29_1/_19_  (.A1(\u_multiplier/STAGE1/_0790_ ),
    .A2(\u_multiplier/STAGE1/_0789_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_1/_20_  (.A(\u_multiplier/STAGE1/_0790_ ),
    .B(\u_multiplier/STAGE1/_0789_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_29_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_29_1/_21_  (.A1(\u_multiplier/STAGE1/_0791_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_29_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_1/_22_  (.A(\u_multiplier/STAGE1/_0791_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_29_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_29_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_29_1/_23_  (.A1(\u_multiplier/STAGE1/_0792_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_29_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_1/_24_  (.A(\u_multiplier/STAGE1/_0792_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_29_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_1/_25_  (.A(\u_multiplier/STAGE1/pp1_28_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_29_1/_16_ ),
    .ZN(\u_multiplier/pp1_29 [6]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_29_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_29_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_29_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_29_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_29_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_29_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_29_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_29_1/_17_ ),
    .ZN(\u_multiplier/pp1_30 [14]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_29_2/_18_  (.A(\u_multiplier/STAGE1/pp1_28_e42_2_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_29_2/_19_  (.A1(\u_multiplier/STAGE1/_0794_ ),
    .A2(\u_multiplier/STAGE1/_0793_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_2/_20_  (.A(\u_multiplier/STAGE1/_0794_ ),
    .B(\u_multiplier/STAGE1/_0793_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_29_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_29_2/_21_  (.A1(\u_multiplier/STAGE1/_0795_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_29_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_2/_22_  (.A(\u_multiplier/STAGE1/_0795_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_29_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_29_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_29_2/_23_  (.A1(\u_multiplier/STAGE1/_0796_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_29_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_2/_24_  (.A(\u_multiplier/STAGE1/_0796_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_29_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_2/_25_  (.A(\u_multiplier/STAGE1/pp1_28_e42_2_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_29_2/_16_ ),
    .ZN(\u_multiplier/pp1_29 [5]));
 NAND2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_29_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_29_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_29_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_29_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_29_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_29_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_29_2/_17_ ),
    .ZN(\u_multiplier/pp1_30 [13]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_29_3/_18_  (.A(\u_multiplier/STAGE1/pp1_28_e42_3_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_29_3/_19_  (.A1(\u_multiplier/STAGE1/_0798_ ),
    .A2(\u_multiplier/STAGE1/_0797_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_3/_20_  (.A(\u_multiplier/STAGE1/_0798_ ),
    .B(\u_multiplier/STAGE1/_0797_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_29_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_29_3/_21_  (.A1(\u_multiplier/STAGE1/_0799_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_29_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_3/_22_  (.A(\u_multiplier/STAGE1/_0799_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_29_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_29_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_29_3/_23_  (.A1(\u_multiplier/STAGE1/_0800_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_29_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_3/_24_  (.A(\u_multiplier/STAGE1/_0800_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_29_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_3/_25_  (.A(\u_multiplier/STAGE1/pp1_28_e42_3_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_29_3/_16_ ),
    .ZN(\u_multiplier/pp1_29 [4]));
 NAND2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_29_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_29_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_29_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_29_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_29_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_29_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_29_3/_17_ ),
    .ZN(\u_multiplier/pp1_30 [12]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_29_4/_18_  (.A(\u_multiplier/STAGE1/pp1_28_e42_4_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_29_4/_19_  (.A1(\u_multiplier/STAGE1/_0802_ ),
    .A2(\u_multiplier/STAGE1/_0801_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_4/_20_  (.A(\u_multiplier/STAGE1/_0802_ ),
    .B(\u_multiplier/STAGE1/_0801_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_29_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_29_4/_21_  (.A1(\u_multiplier/STAGE1/_0803_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_29_4/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_4/_22_  (.A(\u_multiplier/STAGE1/_0803_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_29_4/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_29_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_29_4/_23_  (.A1(\u_multiplier/STAGE1/_0804_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_29_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_4/_24_  (.A(\u_multiplier/STAGE1/_0804_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_29_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_4/_25_  (.A(\u_multiplier/STAGE1/pp1_28_e42_4_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_29_4/_16_ ),
    .ZN(\u_multiplier/pp1_29 [3]));
 NAND2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_4/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_29_4/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_29_4/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_29_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_29_4/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_29_4/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_29_4/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_29_4/_17_ ),
    .ZN(\u_multiplier/pp1_30 [11]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_29_5/_18_  (.A(\u_multiplier/STAGE1/pp1_28_e42_5_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_5/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_29_5/_19_  (.A1(\u_multiplier/STAGE1/_0806_ ),
    .A2(\u_multiplier/STAGE1/_0805_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_5/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_5/_20_  (.A(\u_multiplier/STAGE1/_0806_ ),
    .B(\u_multiplier/STAGE1/_0805_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_29_5/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_29_5/_21_  (.A1(\u_multiplier/STAGE1/_0807_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_29_5/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_5/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_5/_22_  (.A(\u_multiplier/STAGE1/_0807_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_29_5/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_29_5/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_29_5/_23_  (.A1(\u_multiplier/STAGE1/_0808_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_29_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_5/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_5/_24_  (.A(\u_multiplier/STAGE1/_0808_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_29_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_5/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_5/_25_  (.A(\u_multiplier/STAGE1/pp1_28_e42_5_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_29_5/_16_ ),
    .ZN(\u_multiplier/pp1_29 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_29_5/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_29_5/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_29_5/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_29_e42_5_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_29_5/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_29_5/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_29_5/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_29_5/_17_ ),
    .ZN(\u_multiplier/pp1_30 [10]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_29_6/_18_  (.A(\u_multiplier/STAGE1/pp1_28_e42_6_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_6/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_29_6/_19_  (.A1(\u_multiplier/STAGE1/_0810_ ),
    .A2(\u_multiplier/STAGE1/_0809_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_6/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_6/_20_  (.A(\u_multiplier/STAGE1/_0810_ ),
    .B(\u_multiplier/STAGE1/_0809_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_29_6/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_29_6/_21_  (.A1(\u_multiplier/STAGE1/_0811_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_29_6/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_6/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_6/_22_  (.A(\u_multiplier/STAGE1/_0811_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_29_6/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_29_6/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_29_6/_23_  (.A1(\u_multiplier/STAGE1/_0812_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_29_6/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_6/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_6/_24_  (.A(\u_multiplier/STAGE1/_0812_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_29_6/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_6/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_6/_25_  (.A(\u_multiplier/STAGE1/pp1_28_e42_6_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_29_6/_16_ ),
    .ZN(\u_multiplier/pp1_29 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_29_6/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_29_6/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_29_6/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_29_e42_6_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_29_6/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_29_6/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_29_6/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_29_6/_17_ ),
    .ZN(\u_multiplier/pp1_30 [9]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_29_7/_18_  (.A(net126),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_7/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_29_7/_19_  (.A1(\u_multiplier/STAGE1/_0814_ ),
    .A2(\u_multiplier/STAGE1/_0813_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_7/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_7/_20_  (.A(\u_multiplier/STAGE1/_0814_ ),
    .B(\u_multiplier/STAGE1/_0813_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_29_7/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_29_7/_21_  (.A1(\u_multiplier/STAGE1/_0815_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_29_7/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_7/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_7/_22_  (.A(\u_multiplier/STAGE1/_0815_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_29_7/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_29_7/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_29_7/_23_  (.A1(\u_multiplier/STAGE1/_0816_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_29_7/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_7/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_7/_24_  (.A(\u_multiplier/STAGE1/_0816_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_29_7/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_29_7/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_29_7/_25_  (.A(net127),
    .B(\u_multiplier/STAGE1/E_4_2_pp_29_7/_16_ ),
    .ZN(\u_multiplier/pp1_29 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_29_7/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_29_7/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_29_7/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_29_e42_7_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_29_7/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_29_7/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_29_7/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_29_7/_17_ ),
    .ZN(\u_multiplier/pp1_30 [8]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_30_1/_18_  (.A(\u_multiplier/STAGE1/pp1_29_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_30_1/_19_  (.A1(\u_multiplier/STAGE1/_0818_ ),
    .A2(\u_multiplier/STAGE1/_0817_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_1/_20_  (.A(\u_multiplier/STAGE1/_0818_ ),
    .B(\u_multiplier/STAGE1/_0817_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_30_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_30_1/_21_  (.A1(\u_multiplier/STAGE1/_0819_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_30_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_1/_22_  (.A(\u_multiplier/STAGE1/_0819_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_30_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_30_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_30_1/_23_  (.A1(\u_multiplier/STAGE1/_0820_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_30_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_1/_24_  (.A(\u_multiplier/STAGE1/_0820_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_30_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_1/_25_  (.A(\u_multiplier/STAGE1/pp1_29_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_30_1/_16_ ),
    .ZN(\u_multiplier/pp1_30 [7]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_30_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_30_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_30_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_30_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_30_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_30_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_30_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_30_1/_17_ ),
    .ZN(\u_multiplier/pp1_31 [15]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_30_2/_18_  (.A(\u_multiplier/STAGE1/pp1_29_e42_2_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_30_2/_19_  (.A1(\u_multiplier/STAGE1/_0822_ ),
    .A2(\u_multiplier/STAGE1/_0821_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_2/_20_  (.A(\u_multiplier/STAGE1/_0822_ ),
    .B(\u_multiplier/STAGE1/_0821_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_30_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_30_2/_21_  (.A1(\u_multiplier/STAGE1/_0823_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_30_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_2/_22_  (.A(\u_multiplier/STAGE1/_0823_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_30_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_30_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_30_2/_23_  (.A1(\u_multiplier/STAGE1/_0824_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_30_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_2/_24_  (.A(\u_multiplier/STAGE1/_0824_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_30_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_2/_25_  (.A(\u_multiplier/STAGE1/pp1_29_e42_2_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_30_2/_16_ ),
    .ZN(\u_multiplier/pp1_30 [6]));
 NAND2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_30_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_30_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_30_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_30_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_30_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_30_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_30_2/_17_ ),
    .ZN(\u_multiplier/pp1_31 [14]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_30_3/_18_  (.A(\u_multiplier/STAGE1/pp1_29_e42_3_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_30_3/_19_  (.A1(\u_multiplier/STAGE1/_0826_ ),
    .A2(\u_multiplier/STAGE1/_0825_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_3/_20_  (.A(\u_multiplier/STAGE1/_0826_ ),
    .B(\u_multiplier/STAGE1/_0825_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_30_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_30_3/_21_  (.A1(\u_multiplier/STAGE1/_0827_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_30_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_3/_22_  (.A(\u_multiplier/STAGE1/_0827_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_30_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_30_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_30_3/_23_  (.A1(\u_multiplier/STAGE1/_0828_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_30_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_3/_24_  (.A(\u_multiplier/STAGE1/_0828_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_30_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_3/_25_  (.A(\u_multiplier/STAGE1/pp1_29_e42_3_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_30_3/_16_ ),
    .ZN(\u_multiplier/pp1_30 [5]));
 NAND2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_30_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_30_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_30_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_30_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_30_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_30_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_30_3/_17_ ),
    .ZN(\u_multiplier/pp1_31 [13]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_30_4/_18_  (.A(\u_multiplier/STAGE1/pp1_29_e42_4_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_30_4/_19_  (.A1(\u_multiplier/STAGE1/_0830_ ),
    .A2(\u_multiplier/STAGE1/_0829_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_4/_20_  (.A(\u_multiplier/STAGE1/_0830_ ),
    .B(\u_multiplier/STAGE1/_0829_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_30_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_30_4/_21_  (.A1(\u_multiplier/STAGE1/_0831_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_30_4/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_4/_22_  (.A(\u_multiplier/STAGE1/_0831_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_30_4/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_30_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_30_4/_23_  (.A1(\u_multiplier/STAGE1/_0832_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_30_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_4/_24_  (.A(\u_multiplier/STAGE1/_0832_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_30_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_4/_25_  (.A(\u_multiplier/STAGE1/pp1_29_e42_4_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_30_4/_16_ ),
    .ZN(\u_multiplier/pp1_30 [4]));
 NAND2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_4/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_30_4/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_30_4/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_30_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_30_4/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_30_4/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_30_4/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_30_4/_17_ ),
    .ZN(\u_multiplier/pp1_31 [12]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_30_5/_18_  (.A(\u_multiplier/STAGE1/pp1_29_e42_5_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_5/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_30_5/_19_  (.A1(\u_multiplier/STAGE1/_0834_ ),
    .A2(\u_multiplier/STAGE1/_0833_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_5/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_5/_20_  (.A(\u_multiplier/STAGE1/_0834_ ),
    .B(\u_multiplier/STAGE1/_0833_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_30_5/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_30_5/_21_  (.A1(\u_multiplier/STAGE1/_0835_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_30_5/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_5/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_5/_22_  (.A(\u_multiplier/STAGE1/_0835_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_30_5/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_30_5/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_30_5/_23_  (.A1(\u_multiplier/STAGE1/_0836_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_30_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_5/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_5/_24_  (.A(\u_multiplier/STAGE1/_0836_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_30_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_5/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_5/_25_  (.A(\u_multiplier/STAGE1/pp1_29_e42_5_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_30_5/_16_ ),
    .ZN(\u_multiplier/pp1_30 [3]));
 NAND2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_5/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_30_5/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_30_5/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_30_e42_5_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_30_5/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_30_5/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_30_5/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_30_5/_17_ ),
    .ZN(\u_multiplier/pp1_31 [11]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_30_6/_18_  (.A(\u_multiplier/STAGE1/pp1_29_e42_6_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_6/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_30_6/_19_  (.A1(\u_multiplier/STAGE1/_0838_ ),
    .A2(\u_multiplier/STAGE1/_0837_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_6/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_6/_20_  (.A(\u_multiplier/STAGE1/_0838_ ),
    .B(\u_multiplier/STAGE1/_0837_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_30_6/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_30_6/_21_  (.A1(\u_multiplier/STAGE1/_0839_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_30_6/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_6/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_6/_22_  (.A(\u_multiplier/STAGE1/_0839_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_30_6/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_30_6/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_30_6/_23_  (.A1(\u_multiplier/STAGE1/_0840_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_30_6/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_6/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_6/_24_  (.A(\u_multiplier/STAGE1/_0840_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_30_6/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_6/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_6/_25_  (.A(\u_multiplier/STAGE1/pp1_29_e42_6_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_30_6/_16_ ),
    .ZN(\u_multiplier/pp1_30 [2]));
 NAND2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_6/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_30_6/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_30_6/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_30_e42_6_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_30_6/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_30_6/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_30_6/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_30_6/_17_ ),
    .ZN(\u_multiplier/pp1_31 [10]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_30_7/_18_  (.A(\u_multiplier/STAGE1/pp1_29_e42_7_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_7/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_30_7/_19_  (.A1(\u_multiplier/STAGE1/_0842_ ),
    .A2(\u_multiplier/STAGE1/_0841_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_7/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_7/_20_  (.A(\u_multiplier/STAGE1/_0842_ ),
    .B(\u_multiplier/STAGE1/_0841_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_30_7/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_30_7/_21_  (.A1(\u_multiplier/STAGE1/_0843_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_30_7/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_7/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_7/_22_  (.A(\u_multiplier/STAGE1/_0843_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_30_7/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_30_7/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_30_7/_23_  (.A1(\u_multiplier/STAGE1/_0844_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_30_7/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_7/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_7/_24_  (.A(\u_multiplier/STAGE1/_0844_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_30_7/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_30_7/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_7/_25_  (.A(\u_multiplier/STAGE1/pp1_29_e42_7_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_30_7/_16_ ),
    .ZN(\u_multiplier/pp1_30 [1]));
 NAND2_X2 \u_multiplier/STAGE1/E_4_2_pp_30_7/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_30_7/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_30_7/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_30_e42_7_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_30_7/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_30_7/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_30_7/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_30_7/_17_ ),
    .ZN(\u_multiplier/pp1_31 [9]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_31_1/_18_  (.A(\u_multiplier/STAGE1/pp1_30_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_1/_19_  (.A1(\u_multiplier/STAGE1/_0848_ ),
    .A2(\u_multiplier/STAGE1/_0847_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_1/_20_  (.A(\u_multiplier/STAGE1/_0848_ ),
    .B(\u_multiplier/STAGE1/_0847_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_31_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_1/_21_  (.A1(\u_multiplier/STAGE1/_0849_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_31_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_1/_22_  (.A(\u_multiplier/STAGE1/_0849_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_31_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_31_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_1/_23_  (.A1(\u_multiplier/STAGE1/_0850_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_31_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_1/_24_  (.A(\u_multiplier/STAGE1/_0850_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_31_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_1/_25_  (.A(\u_multiplier/STAGE1/pp1_30_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_31_1/_16_ ),
    .ZN(\u_multiplier/pp1_31 [7]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_31_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_31_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_31_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_31_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_31_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_31_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_31_1/_17_ ),
    .ZN(\u_multiplier/pp1_32 [15]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_31_2/_18_  (.A(\u_multiplier/STAGE1/pp1_30_e42_2_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_2/_19_  (.A1(\u_multiplier/STAGE1/_0852_ ),
    .A2(\u_multiplier/STAGE1/_0851_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_2/_20_  (.A(\u_multiplier/STAGE1/_0852_ ),
    .B(\u_multiplier/STAGE1/_0851_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_31_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_2/_21_  (.A1(\u_multiplier/STAGE1/_0853_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_31_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_2/_22_  (.A(\u_multiplier/STAGE1/_0853_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_31_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_31_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_2/_23_  (.A1(\u_multiplier/STAGE1/_0854_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_31_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_2/_24_  (.A(\u_multiplier/STAGE1/_0854_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_31_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_2/_25_  (.A(\u_multiplier/STAGE1/pp1_30_e42_2_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_31_2/_16_ ),
    .ZN(\u_multiplier/pp1_31 [6]));
 NAND2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_31_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_31_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_31_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_31_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_31_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_31_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_31_2/_17_ ),
    .ZN(\u_multiplier/pp1_32 [14]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_31_3/_18_  (.A(\u_multiplier/STAGE1/pp1_30_e42_3_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_3/_19_  (.A1(\u_multiplier/STAGE1/_0856_ ),
    .A2(\u_multiplier/STAGE1/_0855_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_3/_20_  (.A(\u_multiplier/STAGE1/_0856_ ),
    .B(\u_multiplier/STAGE1/_0855_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_31_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_3/_21_  (.A1(\u_multiplier/STAGE1/_0857_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_31_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_3/_22_  (.A(\u_multiplier/STAGE1/_0857_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_31_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_31_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_3/_23_  (.A1(\u_multiplier/STAGE1/_0858_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_31_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_3/_24_  (.A(\u_multiplier/STAGE1/_0858_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_31_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_3/_25_  (.A(\u_multiplier/STAGE1/pp1_30_e42_3_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_31_3/_16_ ),
    .ZN(\u_multiplier/pp1_31 [5]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_31_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_31_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_31_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_31_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_31_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_31_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_31_3/_17_ ),
    .ZN(\u_multiplier/pp1_32 [13]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_31_4/_18_  (.A(\u_multiplier/STAGE1/pp1_30_e42_4_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_4/_19_  (.A1(\u_multiplier/STAGE1/_0860_ ),
    .A2(\u_multiplier/STAGE1/_0859_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_4/_20_  (.A(\u_multiplier/STAGE1/_0860_ ),
    .B(\u_multiplier/STAGE1/_0859_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_31_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_4/_21_  (.A1(\u_multiplier/STAGE1/_0861_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_31_4/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_4/_22_  (.A(\u_multiplier/STAGE1/_0861_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_31_4/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_31_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_4/_23_  (.A1(\u_multiplier/STAGE1/_0862_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_31_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_4/_24_  (.A(\u_multiplier/STAGE1/_0862_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_31_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_4/_25_  (.A(\u_multiplier/STAGE1/pp1_30_e42_4_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_31_4/_16_ ),
    .ZN(\u_multiplier/pp1_31 [4]));
 NAND2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_4/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_31_4/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_31_4/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_31_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_31_4/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_31_4/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_31_4/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_31_4/_17_ ),
    .ZN(\u_multiplier/pp1_32 [12]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_31_5/_18_  (.A(\u_multiplier/STAGE1/pp1_30_e42_5_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_5/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_5/_19_  (.A1(\u_multiplier/STAGE1/_0864_ ),
    .A2(\u_multiplier/STAGE1/_0863_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_5/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_5/_20_  (.A(\u_multiplier/STAGE1/_0864_ ),
    .B(\u_multiplier/STAGE1/_0863_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_31_5/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_5/_21_  (.A1(\u_multiplier/STAGE1/_0865_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_31_5/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_5/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_5/_22_  (.A(\u_multiplier/STAGE1/_0865_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_31_5/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_31_5/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_5/_23_  (.A1(\u_multiplier/STAGE1/_0866_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_31_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_5/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_5/_24_  (.A(\u_multiplier/STAGE1/_0866_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_31_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_5/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_5/_25_  (.A(\u_multiplier/STAGE1/pp1_30_e42_5_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_31_5/_16_ ),
    .ZN(\u_multiplier/pp1_31 [3]));
 NAND2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_5/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_31_5/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_31_5/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_31_e42_5_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_31_5/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_31_5/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_31_5/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_31_5/_17_ ),
    .ZN(\u_multiplier/pp1_32 [11]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_31_6/_18_  (.A(\u_multiplier/STAGE1/pp1_30_e42_6_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_6/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_6/_19_  (.A1(\u_multiplier/STAGE1/_0868_ ),
    .A2(\u_multiplier/STAGE1/_0867_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_6/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_6/_20_  (.A(\u_multiplier/STAGE1/_0868_ ),
    .B(\u_multiplier/STAGE1/_0867_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_31_6/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_6/_21_  (.A1(\u_multiplier/STAGE1/_0869_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_31_6/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_6/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_6/_22_  (.A(\u_multiplier/STAGE1/_0869_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_31_6/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_31_6/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_6/_23_  (.A1(\u_multiplier/STAGE1/_0870_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_31_6/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_6/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_6/_24_  (.A(\u_multiplier/STAGE1/_0870_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_31_6/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_6/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_6/_25_  (.A(\u_multiplier/STAGE1/pp1_30_e42_6_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_31_6/_16_ ),
    .ZN(\u_multiplier/pp1_31 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_6/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_31_6/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_31_6/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_31_e42_6_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_31_6/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_31_6/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_31_6/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_31_6/_17_ ),
    .ZN(\u_multiplier/pp1_32 [10]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_31_7/_18_  (.A(\u_multiplier/STAGE1/pp1_30_e42_7_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_7/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_7/_19_  (.A1(\u_multiplier/STAGE1/_0872_ ),
    .A2(\u_multiplier/STAGE1/_0871_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_7/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_7/_20_  (.A(\u_multiplier/STAGE1/_0872_ ),
    .B(\u_multiplier/STAGE1/_0871_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_31_7/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_7/_21_  (.A1(\u_multiplier/STAGE1/_0873_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_31_7/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_7/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_7/_22_  (.A(\u_multiplier/STAGE1/_0873_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_31_7/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_31_7/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_7/_23_  (.A1(\u_multiplier/STAGE1/_0874_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_31_7/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_7/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_7/_24_  (.A(\u_multiplier/STAGE1/_0874_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_31_7/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_7/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_7/_25_  (.A(\u_multiplier/STAGE1/pp1_30_e42_7_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_31_7/_16_ ),
    .ZN(\u_multiplier/pp1_31 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_7/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_31_7/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_31_7/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_31_e42_7_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_31_7/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_31_7/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_31_7/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_31_7/_17_ ),
    .ZN(\u_multiplier/pp1_32 [9]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_31_8/_18_  (.A(net128),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_8/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_8/_19_  (.A1(\u_multiplier/STAGE1/_0876_ ),
    .A2(\u_multiplier/STAGE1/_0875_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_8/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_8/_20_  (.A(\u_multiplier/STAGE1/_0876_ ),
    .B(\u_multiplier/STAGE1/_0875_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_31_8/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_8/_21_  (.A1(\u_multiplier/STAGE1/_0877_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_31_8/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_8/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_8/_22_  (.A(\u_multiplier/STAGE1/_0877_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_31_8/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_31_8/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_8/_23_  (.A1(\u_multiplier/STAGE1/_0878_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_31_8/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_8/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_8/_24_  (.A(\u_multiplier/STAGE1/_0878_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_31_8/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_31_8/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_31_8/_25_  (.A(net129),
    .B(\u_multiplier/STAGE1/E_4_2_pp_31_8/_16_ ),
    .ZN(\u_multiplier/pp1_31 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_31_8/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_31_8/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_31_8/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_31_e42_8_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_31_8/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_31_8/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_31_8/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_31_8/_17_ ),
    .ZN(\u_multiplier/pp1_32 [8]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_32_1/_18_  (.A(\u_multiplier/STAGE1/pp1_31_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_1/_19_  (.A1(\u_multiplier/STAGE1/_0880_ ),
    .A2(\u_multiplier/STAGE1/_0879_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_1/_20_  (.A(\u_multiplier/STAGE1/_0880_ ),
    .B(\u_multiplier/STAGE1/_0879_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_32_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_1/_21_  (.A1(\u_multiplier/STAGE1/_0881_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_32_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_1/_22_  (.A(\u_multiplier/STAGE1/_0881_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_32_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_32_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_1/_23_  (.A1(\u_multiplier/STAGE1/_0882_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_32_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_1/_24_  (.A(\u_multiplier/STAGE1/_0882_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_32_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_1/_25_  (.A(\u_multiplier/STAGE1/pp1_31_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_32_1/_16_ ),
    .ZN(\u_multiplier/pp1_32 [7]));
 NAND2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_32_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_32_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_32_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_32_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_32_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_32_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_32_1/_17_ ),
    .ZN(\u_multiplier/pp1_33 [15]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_32_2/_18_  (.A(\u_multiplier/STAGE1/pp1_31_e42_2_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_2/_19_  (.A1(\u_multiplier/STAGE1/_0884_ ),
    .A2(\u_multiplier/STAGE1/_0883_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_2/_20_  (.A(\u_multiplier/STAGE1/_0884_ ),
    .B(\u_multiplier/STAGE1/_0883_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_32_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_2/_21_  (.A1(\u_multiplier/STAGE1/_0885_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_32_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_2/_22_  (.A(\u_multiplier/STAGE1/_0885_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_32_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_32_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_2/_23_  (.A1(\u_multiplier/STAGE1/_0886_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_32_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_2/_24_  (.A(\u_multiplier/STAGE1/_0886_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_32_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_2/_25_  (.A(\u_multiplier/STAGE1/pp1_31_e42_2_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_32_2/_16_ ),
    .ZN(\u_multiplier/pp1_32 [6]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_32_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_32_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_32_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_32_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_32_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_32_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_32_2/_17_ ),
    .ZN(\u_multiplier/pp1_33 [14]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_32_3/_18_  (.A(\u_multiplier/STAGE1/pp1_31_e42_3_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_3/_19_  (.A1(\u_multiplier/STAGE1/_0888_ ),
    .A2(\u_multiplier/STAGE1/_0887_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_3/_20_  (.A(\u_multiplier/STAGE1/_0888_ ),
    .B(\u_multiplier/STAGE1/_0887_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_32_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_3/_21_  (.A1(\u_multiplier/STAGE1/_0889_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_32_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_3/_22_  (.A(\u_multiplier/STAGE1/_0889_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_32_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_32_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_3/_23_  (.A1(\u_multiplier/STAGE1/_0890_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_32_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_3/_24_  (.A(\u_multiplier/STAGE1/_0890_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_32_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_3/_25_  (.A(\u_multiplier/STAGE1/pp1_31_e42_3_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_32_3/_16_ ),
    .ZN(\u_multiplier/pp1_32 [5]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_32_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_32_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_32_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_32_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_32_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_32_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_32_3/_17_ ),
    .ZN(\u_multiplier/pp1_33 [13]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_32_4/_18_  (.A(\u_multiplier/STAGE1/pp1_31_e42_4_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_4/_19_  (.A1(\u_multiplier/STAGE1/_0892_ ),
    .A2(\u_multiplier/STAGE1/_0891_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_4/_20_  (.A(\u_multiplier/STAGE1/_0892_ ),
    .B(\u_multiplier/STAGE1/_0891_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_32_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_4/_21_  (.A1(\u_multiplier/STAGE1/_0893_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_32_4/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_4/_22_  (.A(\u_multiplier/STAGE1/_0893_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_32_4/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_32_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_4/_23_  (.A1(\u_multiplier/STAGE1/_0894_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_32_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_4/_24_  (.A(\u_multiplier/STAGE1/_0894_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_32_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_4/_25_  (.A(\u_multiplier/STAGE1/pp1_31_e42_4_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_32_4/_16_ ),
    .ZN(\u_multiplier/pp1_32 [4]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_4/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_32_4/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_32_4/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_32_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_32_4/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_32_4/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_32_4/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_32_4/_17_ ),
    .ZN(\u_multiplier/pp1_33 [12]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_32_5/_18_  (.A(\u_multiplier/STAGE1/pp1_31_e42_5_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_5/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_5/_19_  (.A1(\u_multiplier/STAGE1/_0896_ ),
    .A2(\u_multiplier/STAGE1/_0895_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_5/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_5/_20_  (.A(\u_multiplier/STAGE1/_0896_ ),
    .B(\u_multiplier/STAGE1/_0895_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_32_5/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_5/_21_  (.A1(\u_multiplier/STAGE1/_0897_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_32_5/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_5/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_5/_22_  (.A(\u_multiplier/STAGE1/_0897_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_32_5/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_32_5/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_5/_23_  (.A1(\u_multiplier/STAGE1/_0898_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_32_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_5/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_5/_24_  (.A(\u_multiplier/STAGE1/_0898_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_32_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_5/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_5/_25_  (.A(\u_multiplier/STAGE1/pp1_31_e42_5_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_32_5/_16_ ),
    .ZN(\u_multiplier/pp1_32 [3]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_5/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_32_5/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_32_5/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_32_e42_5_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_32_5/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_32_5/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_32_5/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_32_5/_17_ ),
    .ZN(\u_multiplier/pp1_33 [11]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_32_6/_18_  (.A(\u_multiplier/STAGE1/pp1_31_e42_6_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_6/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_6/_19_  (.A1(\u_multiplier/STAGE1/_0900_ ),
    .A2(\u_multiplier/STAGE1/_0899_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_6/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_6/_20_  (.A(\u_multiplier/STAGE1/_0900_ ),
    .B(\u_multiplier/STAGE1/_0899_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_32_6/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_6/_21_  (.A1(\u_multiplier/STAGE1/_0901_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_32_6/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_6/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_6/_22_  (.A(\u_multiplier/STAGE1/_0901_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_32_6/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_32_6/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_6/_23_  (.A1(\u_multiplier/STAGE1/_0902_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_32_6/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_6/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_6/_24_  (.A(\u_multiplier/STAGE1/_0902_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_32_6/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_6/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_6/_25_  (.A(\u_multiplier/STAGE1/pp1_31_e42_6_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_32_6/_16_ ),
    .ZN(\u_multiplier/pp1_32 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_6/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_32_6/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_32_6/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_32_e42_6_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_32_6/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_32_6/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_32_6/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_32_6/_17_ ),
    .ZN(\u_multiplier/pp1_33 [10]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_32_7/_18_  (.A(\u_multiplier/STAGE1/pp1_31_e42_7_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_7/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_7/_19_  (.A1(\u_multiplier/STAGE1/_0904_ ),
    .A2(\u_multiplier/STAGE1/_0903_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_7/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_7/_20_  (.A(\u_multiplier/STAGE1/_0904_ ),
    .B(\u_multiplier/STAGE1/_0903_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_32_7/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_7/_21_  (.A1(\u_multiplier/STAGE1/_0905_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_32_7/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_7/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_7/_22_  (.A(\u_multiplier/STAGE1/_0905_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_32_7/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_32_7/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_7/_23_  (.A1(\u_multiplier/STAGE1/_0906_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_32_7/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_7/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_7/_24_  (.A(\u_multiplier/STAGE1/_0906_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_32_7/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_7/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_7/_25_  (.A(\u_multiplier/STAGE1/pp1_31_e42_7_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_32_7/_16_ ),
    .ZN(\u_multiplier/pp1_32 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_7/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_32_7/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_32_7/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_32_e42_7_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_32_7/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_32_7/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_32_7/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_32_7/_17_ ),
    .ZN(\u_multiplier/pp1_33 [9]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_32_8/_18_  (.A(\u_multiplier/STAGE1/pp1_31_e42_8_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_8/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_8/_19_  (.A1(\u_multiplier/STAGE1/_0908_ ),
    .A2(\u_multiplier/STAGE1/_0907_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_8/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_8/_20_  (.A(\u_multiplier/STAGE1/_0908_ ),
    .B(\u_multiplier/STAGE1/_0907_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_32_8/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_8/_21_  (.A1(\u_multiplier/STAGE1/_0909_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_32_8/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_8/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_8/_22_  (.A(\u_multiplier/STAGE1/_0909_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_32_8/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_32_8/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_32_8/_23_  (.A1(net130),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_32_8/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_8/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_8/_24_  (.A(net131),
    .B(\u_multiplier/STAGE1/E_4_2_pp_32_8/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_32_8/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_8/_25_  (.A(\u_multiplier/STAGE1/pp1_31_e42_8_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_32_8/_16_ ),
    .ZN(\u_multiplier/pp1_32 [0]));
 NAND2_X2 \u_multiplier/STAGE1/E_4_2_pp_32_8/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_32_8/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_32_8/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_32_e42_8_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_32_8/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_32_8/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_32_8/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_32_8/_17_ ),
    .ZN(\u_multiplier/pp1_33 [8]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_33_1/_18_  (.A(\u_multiplier/STAGE1/pp1_32_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_1/_19_  (.A1(\u_multiplier/STAGE1/_0911_ ),
    .A2(\u_multiplier/STAGE1/_0910_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_1/_20_  (.A(\u_multiplier/STAGE1/_0911_ ),
    .B(\u_multiplier/STAGE1/_0910_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_33_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_1/_21_  (.A1(\u_multiplier/STAGE1/_0912_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_33_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_1/_22_  (.A(\u_multiplier/STAGE1/_0912_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_33_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_33_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_1/_23_  (.A1(\u_multiplier/STAGE1/_0913_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_33_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_1/_24_  (.A(\u_multiplier/STAGE1/_0913_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_33_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_1/_25_  (.A(\u_multiplier/STAGE1/pp1_32_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_33_1/_16_ ),
    .ZN(\u_multiplier/pp1_33 [7]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_33_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_33_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_33_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_33_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_33_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_33_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_33_1/_17_ ),
    .ZN(\u_multiplier/pp1_34 [14]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_33_2/_18_  (.A(\u_multiplier/STAGE1/pp1_32_e42_2_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_2/_19_  (.A1(\u_multiplier/STAGE1/_0915_ ),
    .A2(\u_multiplier/STAGE1/_0914_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_2/_20_  (.A(\u_multiplier/STAGE1/_0915_ ),
    .B(\u_multiplier/STAGE1/_0914_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_33_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_2/_21_  (.A1(\u_multiplier/STAGE1/_0916_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_33_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_2/_22_  (.A(\u_multiplier/STAGE1/_0916_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_33_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_33_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_2/_23_  (.A1(\u_multiplier/STAGE1/_0917_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_33_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_2/_24_  (.A(\u_multiplier/STAGE1/_0917_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_33_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_2/_25_  (.A(\u_multiplier/STAGE1/pp1_32_e42_2_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_33_2/_16_ ),
    .ZN(\u_multiplier/pp1_33 [6]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_33_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_33_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_33_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_33_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_33_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_33_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_33_2/_17_ ),
    .ZN(\u_multiplier/pp1_34 [13]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_33_3/_18_  (.A(\u_multiplier/STAGE1/pp1_32_e42_3_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_3/_19_  (.A1(\u_multiplier/STAGE1/_0919_ ),
    .A2(\u_multiplier/STAGE1/_0918_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_3/_20_  (.A(\u_multiplier/STAGE1/_0919_ ),
    .B(\u_multiplier/STAGE1/_0918_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_33_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_3/_21_  (.A1(\u_multiplier/STAGE1/_0920_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_33_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_3/_22_  (.A(\u_multiplier/STAGE1/_0920_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_33_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_33_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_3/_23_  (.A1(\u_multiplier/STAGE1/_0921_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_33_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_3/_24_  (.A(\u_multiplier/STAGE1/_0921_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_33_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_3/_25_  (.A(\u_multiplier/STAGE1/pp1_32_e42_3_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_33_3/_16_ ),
    .ZN(\u_multiplier/pp1_33 [5]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_33_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_33_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_33_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_33_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_33_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_33_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_33_3/_17_ ),
    .ZN(\u_multiplier/pp1_34 [12]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_33_4/_18_  (.A(\u_multiplier/STAGE1/pp1_32_e42_4_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_4/_19_  (.A1(\u_multiplier/STAGE1/_0923_ ),
    .A2(\u_multiplier/STAGE1/_0922_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_4/_20_  (.A(\u_multiplier/STAGE1/_0923_ ),
    .B(\u_multiplier/STAGE1/_0922_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_33_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_4/_21_  (.A1(\u_multiplier/STAGE1/_0924_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_33_4/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_4/_22_  (.A(\u_multiplier/STAGE1/_0924_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_33_4/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_33_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_4/_23_  (.A1(\u_multiplier/STAGE1/_0925_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_33_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_4/_24_  (.A(\u_multiplier/STAGE1/_0925_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_33_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_4/_25_  (.A(\u_multiplier/STAGE1/pp1_32_e42_4_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_33_4/_16_ ),
    .ZN(\u_multiplier/pp1_33 [4]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_4/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_33_4/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_33_4/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_33_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_33_4/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_33_4/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_33_4/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_33_4/_17_ ),
    .ZN(\u_multiplier/pp1_34 [11]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_33_5/_18_  (.A(\u_multiplier/STAGE1/pp1_32_e42_5_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_5/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_5/_19_  (.A1(\u_multiplier/STAGE1/_0927_ ),
    .A2(\u_multiplier/STAGE1/_0926_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_5/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_5/_20_  (.A(\u_multiplier/STAGE1/_0927_ ),
    .B(\u_multiplier/STAGE1/_0926_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_33_5/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_5/_21_  (.A1(\u_multiplier/STAGE1/_0928_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_33_5/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_5/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_5/_22_  (.A(\u_multiplier/STAGE1/_0928_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_33_5/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_33_5/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_5/_23_  (.A1(\u_multiplier/STAGE1/_0929_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_33_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_5/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_5/_24_  (.A(\u_multiplier/STAGE1/_0929_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_33_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_5/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_5/_25_  (.A(\u_multiplier/STAGE1/pp1_32_e42_5_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_33_5/_16_ ),
    .ZN(\u_multiplier/pp1_33 [3]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_5/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_33_5/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_33_5/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_33_e42_5_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_33_5/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_33_5/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_33_5/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_33_5/_17_ ),
    .ZN(\u_multiplier/pp1_34 [10]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_33_6/_18_  (.A(\u_multiplier/STAGE1/pp1_32_e42_6_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_6/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_6/_19_  (.A1(\u_multiplier/STAGE1/_0931_ ),
    .A2(\u_multiplier/STAGE1/_0930_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_6/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_6/_20_  (.A(\u_multiplier/STAGE1/_0931_ ),
    .B(\u_multiplier/STAGE1/_0930_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_33_6/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_6/_21_  (.A1(\u_multiplier/STAGE1/_0932_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_33_6/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_6/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_6/_22_  (.A(\u_multiplier/STAGE1/_0932_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_33_6/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_33_6/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_6/_23_  (.A1(\u_multiplier/STAGE1/_0933_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_33_6/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_6/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_6/_24_  (.A(\u_multiplier/STAGE1/_0933_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_33_6/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_6/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_6/_25_  (.A(\u_multiplier/STAGE1/pp1_32_e42_6_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_33_6/_16_ ),
    .ZN(\u_multiplier/pp1_33 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_6/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_33_6/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_33_6/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_33_e42_6_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_33_6/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_33_6/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_33_6/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_33_6/_17_ ),
    .ZN(\u_multiplier/pp1_34 [9]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_33_7/_18_  (.A(\u_multiplier/STAGE1/pp1_32_e42_7_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_7/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_7/_19_  (.A1(\u_multiplier/STAGE1/_0935_ ),
    .A2(\u_multiplier/STAGE1/_0934_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_7/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_7/_20_  (.A(\u_multiplier/STAGE1/_0935_ ),
    .B(\u_multiplier/STAGE1/_0934_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_33_7/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_7/_21_  (.A1(\u_multiplier/STAGE1/_0936_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_33_7/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_7/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_7/_22_  (.A(\u_multiplier/STAGE1/_0936_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_33_7/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_33_7/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_7/_23_  (.A1(\u_multiplier/STAGE1/_0937_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_33_7/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_7/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_7/_24_  (.A(\u_multiplier/STAGE1/_0937_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_33_7/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_33_7/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_33_7/_25_  (.A(\u_multiplier/STAGE1/pp1_32_e42_7_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_33_7/_16_ ),
    .ZN(\u_multiplier/pp1_33 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_33_7/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_33_7/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_33_7/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_33_e42_7_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_33_7/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_33_7/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_33_7/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_33_7/_17_ ),
    .ZN(\u_multiplier/pp1_34 [8]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_34_1/_18_  (.A(\u_multiplier/STAGE1/pp1_33_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_1/_19_  (.A1(\u_multiplier/STAGE1/_0941_ ),
    .A2(\u_multiplier/STAGE1/_0940_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_1/_20_  (.A(\u_multiplier/STAGE1/_0941_ ),
    .B(\u_multiplier/STAGE1/_0940_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_34_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_1/_21_  (.A1(\u_multiplier/STAGE1/_0942_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_34_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_1/_22_  (.A(\u_multiplier/STAGE1/_0942_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_34_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_34_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_1/_23_  (.A1(\u_multiplier/STAGE1/_0943_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_34_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_1/_24_  (.A(\u_multiplier/STAGE1/_0943_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_34_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_1/_25_  (.A(\u_multiplier/STAGE1/pp1_33_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_34_1/_16_ ),
    .ZN(\u_multiplier/pp1_34 [6]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_34_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_34_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_34_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_34_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_34_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_34_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_34_1/_17_ ),
    .ZN(\u_multiplier/pp1_35 [13]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_34_2/_18_  (.A(\u_multiplier/STAGE1/pp1_33_e42_2_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_2/_19_  (.A1(\u_multiplier/STAGE1/_0945_ ),
    .A2(\u_multiplier/STAGE1/_0944_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_2/_20_  (.A(\u_multiplier/STAGE1/_0945_ ),
    .B(\u_multiplier/STAGE1/_0944_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_34_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_2/_21_  (.A1(\u_multiplier/STAGE1/_0946_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_34_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_2/_22_  (.A(\u_multiplier/STAGE1/_0946_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_34_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_34_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_2/_23_  (.A1(\u_multiplier/STAGE1/_0947_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_34_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_2/_24_  (.A(\u_multiplier/STAGE1/_0947_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_34_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_2/_25_  (.A(\u_multiplier/STAGE1/pp1_33_e42_2_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_34_2/_16_ ),
    .ZN(\u_multiplier/pp1_34 [5]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_34_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_34_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_34_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_34_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_34_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_34_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_34_2/_17_ ),
    .ZN(\u_multiplier/pp1_35 [12]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_34_3/_18_  (.A(\u_multiplier/STAGE1/pp1_33_e42_3_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_3/_19_  (.A1(\u_multiplier/STAGE1/_0949_ ),
    .A2(\u_multiplier/STAGE1/_0948_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_3/_20_  (.A(\u_multiplier/STAGE1/_0949_ ),
    .B(\u_multiplier/STAGE1/_0948_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_34_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_3/_21_  (.A1(\u_multiplier/STAGE1/_0950_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_34_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_3/_22_  (.A(\u_multiplier/STAGE1/_0950_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_34_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_34_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_3/_23_  (.A1(\u_multiplier/STAGE1/_0951_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_34_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_3/_24_  (.A(\u_multiplier/STAGE1/_0951_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_34_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_3/_25_  (.A(\u_multiplier/STAGE1/pp1_33_e42_3_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_34_3/_16_ ),
    .ZN(\u_multiplier/pp1_34 [4]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_34_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_34_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_34_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_34_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_34_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_34_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_34_3/_17_ ),
    .ZN(\u_multiplier/pp1_35 [11]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_34_4/_18_  (.A(\u_multiplier/STAGE1/pp1_33_e42_4_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_4/_19_  (.A1(\u_multiplier/STAGE1/_0953_ ),
    .A2(\u_multiplier/STAGE1/_0952_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_4/_20_  (.A(\u_multiplier/STAGE1/_0953_ ),
    .B(\u_multiplier/STAGE1/_0952_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_34_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_4/_21_  (.A1(\u_multiplier/STAGE1/_0954_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_34_4/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_4/_22_  (.A(\u_multiplier/STAGE1/_0954_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_34_4/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_34_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_4/_23_  (.A1(\u_multiplier/STAGE1/_0955_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_34_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_4/_24_  (.A(\u_multiplier/STAGE1/_0955_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_34_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_4/_25_  (.A(\u_multiplier/STAGE1/pp1_33_e42_4_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_34_4/_16_ ),
    .ZN(\u_multiplier/pp1_34 [3]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_4/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_34_4/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_34_4/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_34_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_34_4/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_34_4/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_34_4/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_34_4/_17_ ),
    .ZN(\u_multiplier/pp1_35 [10]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_34_5/_18_  (.A(\u_multiplier/STAGE1/pp1_33_e42_5_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_5/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_5/_19_  (.A1(\u_multiplier/STAGE1/_0957_ ),
    .A2(\u_multiplier/STAGE1/_0956_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_5/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_5/_20_  (.A(\u_multiplier/STAGE1/_0957_ ),
    .B(\u_multiplier/STAGE1/_0956_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_34_5/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_5/_21_  (.A1(\u_multiplier/STAGE1/_0958_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_34_5/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_5/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_5/_22_  (.A(\u_multiplier/STAGE1/_0958_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_34_5/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_34_5/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_5/_23_  (.A1(\u_multiplier/STAGE1/_0959_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_34_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_5/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_5/_24_  (.A(\u_multiplier/STAGE1/_0959_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_34_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_5/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_5/_25_  (.A(\u_multiplier/STAGE1/pp1_33_e42_5_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_34_5/_16_ ),
    .ZN(\u_multiplier/pp1_34 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_5/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_34_5/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_34_5/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_34_e42_5_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_34_5/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_34_5/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_34_5/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_34_5/_17_ ),
    .ZN(\u_multiplier/pp1_35 [9]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_34_6/_18_  (.A(\u_multiplier/STAGE1/pp1_33_e42_6_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_6/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_6/_19_  (.A1(\u_multiplier/STAGE1/_0961_ ),
    .A2(\u_multiplier/STAGE1/_0960_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_6/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_6/_20_  (.A(\u_multiplier/STAGE1/_0961_ ),
    .B(\u_multiplier/STAGE1/_0960_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_34_6/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_6/_21_  (.A1(\u_multiplier/STAGE1/_0962_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_34_6/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_6/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_6/_22_  (.A(\u_multiplier/STAGE1/_0962_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_34_6/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_34_6/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_6/_23_  (.A1(\u_multiplier/STAGE1/_0963_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_34_6/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_6/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_6/_24_  (.A(\u_multiplier/STAGE1/_0963_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_34_6/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_6/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_6/_25_  (.A(\u_multiplier/STAGE1/pp1_33_e42_6_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_34_6/_16_ ),
    .ZN(\u_multiplier/pp1_34 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_6/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_34_6/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_34_6/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_34_e42_6_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_34_6/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_34_6/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_34_6/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_34_6/_17_ ),
    .ZN(\u_multiplier/pp1_35 [8]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_34_7/_18_  (.A(\u_multiplier/STAGE1/pp1_33_e42_7_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_7/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_7/_19_  (.A1(\u_multiplier/STAGE1/_0965_ ),
    .A2(\u_multiplier/STAGE1/_0964_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_7/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_7/_20_  (.A(\u_multiplier/STAGE1/_0965_ ),
    .B(\u_multiplier/STAGE1/_0964_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_34_7/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_7/_21_  (.A1(\u_multiplier/STAGE1/_0966_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_34_7/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_7/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_7/_22_  (.A(\u_multiplier/STAGE1/_0966_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_34_7/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_34_7/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_7/_23_  (.A1(\u_multiplier/STAGE1/_0967_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_34_7/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_7/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_7/_24_  (.A(\u_multiplier/STAGE1/_0967_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_34_7/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_34_7/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_34_7/_25_  (.A(\u_multiplier/STAGE1/pp1_33_e42_7_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_34_7/_16_ ),
    .ZN(\u_multiplier/pp1_34 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_34_7/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_34_7/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_34_7/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_34_e42_7_cout ));
 OAI21_X1 \u_multiplier/STAGE1/E_4_2_pp_34_7/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_34_7/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_34_7/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_34_7/_17_ ),
    .ZN(\u_multiplier/pp1_35 [7]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_35_1/_18_  (.A(\u_multiplier/STAGE1/pp1_34_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_35_1/_19_  (.A1(\u_multiplier/STAGE1/_0969_ ),
    .A2(\u_multiplier/STAGE1/_0968_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_35_1/_20_  (.A(\u_multiplier/STAGE1/_0969_ ),
    .B(\u_multiplier/STAGE1/_0968_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_35_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_35_1/_21_  (.A1(\u_multiplier/STAGE1/_0970_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_35_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_35_1/_22_  (.A(\u_multiplier/STAGE1/_0970_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_35_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_35_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_35_1/_23_  (.A1(\u_multiplier/STAGE1/_0971_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_35_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_35_1/_24_  (.A(\u_multiplier/STAGE1/_0971_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_35_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_35_1/_25_  (.A(\u_multiplier/STAGE1/pp1_34_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_35_1/_16_ ),
    .ZN(\u_multiplier/pp1_35 [6]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_35_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_35_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_35_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_35_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_35_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_35_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_35_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_35_1/_17_ ),
    .ZN(\u_multiplier/pp1_36 [12]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_35_2/_18_  (.A(\u_multiplier/STAGE1/pp1_34_e42_2_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_35_2/_19_  (.A1(\u_multiplier/STAGE1/_0973_ ),
    .A2(\u_multiplier/STAGE1/_0972_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_35_2/_20_  (.A(\u_multiplier/STAGE1/_0973_ ),
    .B(\u_multiplier/STAGE1/_0972_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_35_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_35_2/_21_  (.A1(\u_multiplier/STAGE1/_0974_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_35_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_35_2/_22_  (.A(\u_multiplier/STAGE1/_0974_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_35_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_35_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_35_2/_23_  (.A1(\u_multiplier/STAGE1/_0975_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_35_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_35_2/_24_  (.A(\u_multiplier/STAGE1/_0975_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_35_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_35_2/_25_  (.A(\u_multiplier/STAGE1/pp1_34_e42_2_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_35_2/_16_ ),
    .ZN(\u_multiplier/pp1_35 [5]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_35_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_35_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_35_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_35_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_35_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_35_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_35_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_35_2/_17_ ),
    .ZN(\u_multiplier/pp1_36 [11]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_35_3/_18_  (.A(\u_multiplier/STAGE1/pp1_34_e42_3_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_35_3/_19_  (.A1(\u_multiplier/STAGE1/_0977_ ),
    .A2(\u_multiplier/STAGE1/_0976_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_35_3/_20_  (.A(\u_multiplier/STAGE1/_0977_ ),
    .B(\u_multiplier/STAGE1/_0976_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_35_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_35_3/_21_  (.A1(\u_multiplier/STAGE1/_0978_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_35_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_35_3/_22_  (.A(\u_multiplier/STAGE1/_0978_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_35_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_35_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_35_3/_23_  (.A1(\u_multiplier/STAGE1/_0979_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_35_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_35_3/_24_  (.A(\u_multiplier/STAGE1/_0979_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_35_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_35_3/_25_  (.A(\u_multiplier/STAGE1/pp1_34_e42_3_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_35_3/_16_ ),
    .ZN(\u_multiplier/pp1_35 [4]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_35_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_35_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_35_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_35_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_35_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_35_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_35_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_35_3/_17_ ),
    .ZN(\u_multiplier/pp1_36 [10]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_35_4/_18_  (.A(\u_multiplier/STAGE1/pp1_34_e42_4_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_35_4/_19_  (.A1(\u_multiplier/STAGE1/_0981_ ),
    .A2(\u_multiplier/STAGE1/_0980_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_35_4/_20_  (.A(\u_multiplier/STAGE1/_0981_ ),
    .B(\u_multiplier/STAGE1/_0980_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_35_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_35_4/_21_  (.A1(\u_multiplier/STAGE1/_0982_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_35_4/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_35_4/_22_  (.A(\u_multiplier/STAGE1/_0982_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_35_4/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_35_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_35_4/_23_  (.A1(\u_multiplier/STAGE1/_0983_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_35_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_35_4/_24_  (.A(\u_multiplier/STAGE1/_0983_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_35_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_35_4/_25_  (.A(\u_multiplier/STAGE1/pp1_34_e42_4_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_35_4/_16_ ),
    .ZN(\u_multiplier/pp1_35 [3]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_35_4/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_35_4/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_35_4/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_35_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_35_4/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_35_4/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_35_4/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_35_4/_17_ ),
    .ZN(\u_multiplier/pp1_36 [9]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_35_5/_18_  (.A(\u_multiplier/STAGE1/pp1_34_e42_5_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_5/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_35_5/_19_  (.A1(\u_multiplier/STAGE1/_0985_ ),
    .A2(\u_multiplier/STAGE1/_0984_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_5/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_35_5/_20_  (.A(\u_multiplier/STAGE1/_0985_ ),
    .B(\u_multiplier/STAGE1/_0984_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_35_5/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_35_5/_21_  (.A1(\u_multiplier/STAGE1/_0986_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_35_5/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_5/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_35_5/_22_  (.A(\u_multiplier/STAGE1/_0986_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_35_5/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_35_5/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_35_5/_23_  (.A1(\u_multiplier/STAGE1/_0987_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_35_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_5/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_35_5/_24_  (.A(\u_multiplier/STAGE1/_0987_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_35_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_5/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_35_5/_25_  (.A(\u_multiplier/STAGE1/pp1_34_e42_5_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_35_5/_16_ ),
    .ZN(\u_multiplier/pp1_35 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_35_5/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_35_5/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_35_5/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_35_e42_5_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_35_5/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_35_5/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_35_5/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_35_5/_17_ ),
    .ZN(\u_multiplier/pp1_36 [8]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_35_6/_18_  (.A(\u_multiplier/STAGE1/pp1_34_e42_6_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_6/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_35_6/_19_  (.A1(\u_multiplier/STAGE1/_0989_ ),
    .A2(\u_multiplier/STAGE1/_0988_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_6/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_35_6/_20_  (.A(\u_multiplier/STAGE1/_0989_ ),
    .B(\u_multiplier/STAGE1/_0988_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_35_6/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_35_6/_21_  (.A1(\u_multiplier/STAGE1/_0990_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_35_6/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_6/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_35_6/_22_  (.A(\u_multiplier/STAGE1/_0990_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_35_6/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_35_6/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_35_6/_23_  (.A1(\u_multiplier/STAGE1/_0991_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_35_6/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_6/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_35_6/_24_  (.A(\u_multiplier/STAGE1/_0991_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_35_6/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_35_6/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_35_6/_25_  (.A(\u_multiplier/STAGE1/pp1_34_e42_6_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_35_6/_16_ ),
    .ZN(\u_multiplier/pp1_35 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_35_6/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_35_6/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_35_6/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_35_e42_6_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_35_6/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_35_6/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_35_6/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_35_6/_17_ ),
    .ZN(\u_multiplier/pp1_36 [7]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_36_1/_18_  (.A(\u_multiplier/STAGE1/pp1_35_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_36_1/_19_  (.A1(\u_multiplier/STAGE1/_0995_ ),
    .A2(\u_multiplier/STAGE1/_0994_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_36_1/_20_  (.A(\u_multiplier/STAGE1/_0995_ ),
    .B(\u_multiplier/STAGE1/_0994_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_36_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_36_1/_21_  (.A1(\u_multiplier/STAGE1/_0996_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_36_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_36_1/_22_  (.A(\u_multiplier/STAGE1/_0996_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_36_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_36_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_36_1/_23_  (.A1(\u_multiplier/STAGE1/_0997_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_36_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_36_1/_24_  (.A(\u_multiplier/STAGE1/_0997_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_36_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_36_1/_25_  (.A(\u_multiplier/STAGE1/pp1_35_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_36_1/_16_ ),
    .ZN(\u_multiplier/pp1_36 [5]));
 NAND2_X2 \u_multiplier/STAGE1/E_4_2_pp_36_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_36_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_36_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_36_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_36_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_36_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_36_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_36_1/_17_ ),
    .ZN(\u_multiplier/pp1_37 [11]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_36_2/_18_  (.A(\u_multiplier/STAGE1/pp1_35_e42_2_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_36_2/_19_  (.A1(\u_multiplier/STAGE1/_0999_ ),
    .A2(\u_multiplier/STAGE1/_0998_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_36_2/_20_  (.A(\u_multiplier/STAGE1/_0999_ ),
    .B(\u_multiplier/STAGE1/_0998_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_36_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_36_2/_21_  (.A1(\u_multiplier/STAGE1/_1000_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_36_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_36_2/_22_  (.A(\u_multiplier/STAGE1/_1000_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_36_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_36_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_36_2/_23_  (.A1(\u_multiplier/STAGE1/_1001_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_36_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_36_2/_24_  (.A(\u_multiplier/STAGE1/_1001_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_36_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_36_2/_25_  (.A(\u_multiplier/STAGE1/pp1_35_e42_2_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_36_2/_16_ ),
    .ZN(\u_multiplier/pp1_36 [4]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_36_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_36_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_36_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_36_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_36_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_36_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_36_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_36_2/_17_ ),
    .ZN(\u_multiplier/pp1_37 [10]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_36_3/_18_  (.A(\u_multiplier/STAGE1/pp1_35_e42_3_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_36_3/_19_  (.A1(\u_multiplier/STAGE1/_1003_ ),
    .A2(\u_multiplier/STAGE1/_1002_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_36_3/_20_  (.A(\u_multiplier/STAGE1/_1003_ ),
    .B(\u_multiplier/STAGE1/_1002_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_36_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_36_3/_21_  (.A1(\u_multiplier/STAGE1/_1004_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_36_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_36_3/_22_  (.A(\u_multiplier/STAGE1/_1004_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_36_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_36_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_36_3/_23_  (.A1(\u_multiplier/STAGE1/_1005_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_36_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_36_3/_24_  (.A(\u_multiplier/STAGE1/_1005_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_36_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_36_3/_25_  (.A(\u_multiplier/STAGE1/pp1_35_e42_3_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_36_3/_16_ ),
    .ZN(\u_multiplier/pp1_36 [3]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_36_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_36_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_36_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_36_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_36_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_36_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_36_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_36_3/_17_ ),
    .ZN(\u_multiplier/pp1_37 [9]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_36_4/_18_  (.A(\u_multiplier/STAGE1/pp1_35_e42_4_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_36_4/_19_  (.A1(\u_multiplier/STAGE1/_1007_ ),
    .A2(\u_multiplier/STAGE1/_1006_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_36_4/_20_  (.A(\u_multiplier/STAGE1/_1007_ ),
    .B(\u_multiplier/STAGE1/_1006_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_36_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_36_4/_21_  (.A1(\u_multiplier/STAGE1/_1008_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_36_4/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_36_4/_22_  (.A(\u_multiplier/STAGE1/_1008_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_36_4/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_36_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_36_4/_23_  (.A1(\u_multiplier/STAGE1/_1009_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_36_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_36_4/_24_  (.A(\u_multiplier/STAGE1/_1009_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_36_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_36_4/_25_  (.A(\u_multiplier/STAGE1/pp1_35_e42_4_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_36_4/_16_ ),
    .ZN(\u_multiplier/pp1_36 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_36_4/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_36_4/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_36_4/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_36_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_36_4/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_36_4/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_36_4/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_36_4/_17_ ),
    .ZN(\u_multiplier/pp1_37 [8]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_36_5/_18_  (.A(\u_multiplier/STAGE1/pp1_35_e42_5_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_5/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_36_5/_19_  (.A1(\u_multiplier/STAGE1/_1011_ ),
    .A2(\u_multiplier/STAGE1/_1010_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_5/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_36_5/_20_  (.A(\u_multiplier/STAGE1/_1011_ ),
    .B(\u_multiplier/STAGE1/_1010_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_36_5/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_36_5/_21_  (.A1(\u_multiplier/STAGE1/_1012_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_36_5/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_5/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_36_5/_22_  (.A(\u_multiplier/STAGE1/_1012_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_36_5/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_36_5/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_36_5/_23_  (.A1(\u_multiplier/STAGE1/_1013_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_36_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_5/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_36_5/_24_  (.A(\u_multiplier/STAGE1/_1013_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_36_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_5/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_36_5/_25_  (.A(\u_multiplier/STAGE1/pp1_35_e42_5_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_36_5/_16_ ),
    .ZN(\u_multiplier/pp1_36 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_36_5/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_36_5/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_36_5/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_36_e42_5_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_36_5/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_36_5/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_36_5/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_36_5/_17_ ),
    .ZN(\u_multiplier/pp1_37 [7]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_36_6/_18_  (.A(\u_multiplier/STAGE1/pp1_35_e42_6_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_6/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_36_6/_19_  (.A1(\u_multiplier/STAGE1/_1015_ ),
    .A2(\u_multiplier/STAGE1/_1014_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_6/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_36_6/_20_  (.A(\u_multiplier/STAGE1/_1015_ ),
    .B(\u_multiplier/STAGE1/_1014_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_36_6/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_36_6/_21_  (.A1(\u_multiplier/STAGE1/_1016_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_36_6/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_6/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_36_6/_22_  (.A(\u_multiplier/STAGE1/_1016_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_36_6/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_36_6/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_36_6/_23_  (.A1(\u_multiplier/STAGE1/_1017_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_36_6/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_6/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_36_6/_24_  (.A(\u_multiplier/STAGE1/_1017_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_36_6/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_36_6/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_36_6/_25_  (.A(\u_multiplier/STAGE1/pp1_35_e42_6_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_36_6/_16_ ),
    .ZN(\u_multiplier/pp1_36 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_36_6/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_36_6/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_36_6/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_36_e42_6_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_36_6/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_36_6/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_36_6/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_36_6/_17_ ),
    .ZN(\u_multiplier/pp1_37 [6]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_37_1/_18_  (.A(\u_multiplier/STAGE1/pp1_36_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_37_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_37_1/_19_  (.A1(\u_multiplier/STAGE1/_1019_ ),
    .A2(\u_multiplier/STAGE1/_1018_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_37_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_37_1/_20_  (.A(\u_multiplier/STAGE1/_1019_ ),
    .B(\u_multiplier/STAGE1/_1018_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_37_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_37_1/_21_  (.A1(\u_multiplier/STAGE1/_1020_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_37_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_37_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_37_1/_22_  (.A(\u_multiplier/STAGE1/_1020_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_37_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_37_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_37_1/_23_  (.A1(\u_multiplier/STAGE1/_1021_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_37_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_37_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_37_1/_24_  (.A(\u_multiplier/STAGE1/_1021_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_37_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_37_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_37_1/_25_  (.A(\u_multiplier/STAGE1/pp1_36_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_37_1/_16_ ),
    .ZN(\u_multiplier/pp1_37 [5]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_37_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_37_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_37_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_37_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_37_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_37_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_37_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_37_1/_17_ ),
    .ZN(\u_multiplier/pp1_38 [10]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_37_2/_18_  (.A(\u_multiplier/STAGE1/pp1_36_e42_2_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_37_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_37_2/_19_  (.A1(\u_multiplier/STAGE1/_1023_ ),
    .A2(\u_multiplier/STAGE1/_1022_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_37_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_37_2/_20_  (.A(\u_multiplier/STAGE1/_1023_ ),
    .B(\u_multiplier/STAGE1/_1022_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_37_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_37_2/_21_  (.A1(\u_multiplier/STAGE1/_1024_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_37_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_37_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_37_2/_22_  (.A(\u_multiplier/STAGE1/_1024_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_37_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_37_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_37_2/_23_  (.A1(\u_multiplier/STAGE1/_1025_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_37_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_37_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_37_2/_24_  (.A(\u_multiplier/STAGE1/_1025_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_37_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_37_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_37_2/_25_  (.A(\u_multiplier/STAGE1/pp1_36_e42_2_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_37_2/_16_ ),
    .ZN(\u_multiplier/pp1_37 [4]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_37_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_37_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_37_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_37_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_37_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_37_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_37_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_37_2/_17_ ),
    .ZN(\u_multiplier/pp1_38 [9]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_37_3/_18_  (.A(\u_multiplier/STAGE1/pp1_36_e42_3_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_37_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_37_3/_19_  (.A1(\u_multiplier/STAGE1/_1027_ ),
    .A2(\u_multiplier/STAGE1/_1026_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_37_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_37_3/_20_  (.A(\u_multiplier/STAGE1/_1027_ ),
    .B(\u_multiplier/STAGE1/_1026_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_37_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_37_3/_21_  (.A1(\u_multiplier/STAGE1/_1028_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_37_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_37_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_37_3/_22_  (.A(\u_multiplier/STAGE1/_1028_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_37_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_37_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_37_3/_23_  (.A1(\u_multiplier/STAGE1/_1029_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_37_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_37_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_37_3/_24_  (.A(\u_multiplier/STAGE1/_1029_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_37_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_37_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_37_3/_25_  (.A(\u_multiplier/STAGE1/pp1_36_e42_3_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_37_3/_16_ ),
    .ZN(\u_multiplier/pp1_37 [3]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_37_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_37_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_37_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_37_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_37_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_37_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_37_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_37_3/_17_ ),
    .ZN(\u_multiplier/pp1_38 [8]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_37_4/_18_  (.A(\u_multiplier/STAGE1/pp1_36_e42_4_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_37_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_37_4/_19_  (.A1(\u_multiplier/STAGE1/_1031_ ),
    .A2(\u_multiplier/STAGE1/_1030_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_37_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_37_4/_20_  (.A(\u_multiplier/STAGE1/_1031_ ),
    .B(\u_multiplier/STAGE1/_1030_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_37_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_37_4/_21_  (.A1(\u_multiplier/STAGE1/_1032_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_37_4/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_37_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_37_4/_22_  (.A(\u_multiplier/STAGE1/_1032_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_37_4/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_37_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_37_4/_23_  (.A1(\u_multiplier/STAGE1/_1033_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_37_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_37_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_37_4/_24_  (.A(\u_multiplier/STAGE1/_1033_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_37_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_37_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_37_4/_25_  (.A(\u_multiplier/STAGE1/pp1_36_e42_4_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_37_4/_16_ ),
    .ZN(\u_multiplier/pp1_37 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_37_4/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_37_4/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_37_4/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_37_e42_4_cout ));
 OAI21_X1 \u_multiplier/STAGE1/E_4_2_pp_37_4/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_37_4/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_37_4/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_37_4/_17_ ),
    .ZN(\u_multiplier/pp1_38 [7]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_37_5/_18_  (.A(\u_multiplier/STAGE1/pp1_36_e42_5_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_37_5/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_37_5/_19_  (.A1(\u_multiplier/STAGE1/_1035_ ),
    .A2(\u_multiplier/STAGE1/_1034_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_37_5/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_37_5/_20_  (.A(\u_multiplier/STAGE1/_1035_ ),
    .B(\u_multiplier/STAGE1/_1034_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_37_5/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_37_5/_21_  (.A1(\u_multiplier/STAGE1/_1036_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_37_5/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_37_5/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_37_5/_22_  (.A(\u_multiplier/STAGE1/_1036_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_37_5/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_37_5/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_37_5/_23_  (.A1(\u_multiplier/STAGE1/_1037_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_37_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_37_5/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_37_5/_24_  (.A(\u_multiplier/STAGE1/_1037_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_37_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_37_5/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_37_5/_25_  (.A(\u_multiplier/STAGE1/pp1_36_e42_5_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_37_5/_16_ ),
    .ZN(\u_multiplier/pp1_37 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_37_5/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_37_5/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_37_5/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_37_e42_5_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_37_5/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_37_5/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_37_5/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_37_5/_17_ ),
    .ZN(\u_multiplier/pp1_38 [6]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_38_1/_18_  (.A(\u_multiplier/STAGE1/pp1_37_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_38_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_38_1/_19_  (.A1(\u_multiplier/STAGE1/_1041_ ),
    .A2(\u_multiplier/STAGE1/_1040_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_38_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_38_1/_20_  (.A(\u_multiplier/STAGE1/_1041_ ),
    .B(\u_multiplier/STAGE1/_1040_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_38_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_38_1/_21_  (.A1(\u_multiplier/STAGE1/_1042_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_38_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_38_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_38_1/_22_  (.A(\u_multiplier/STAGE1/_1042_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_38_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_38_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_38_1/_23_  (.A1(\u_multiplier/STAGE1/_1043_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_38_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_38_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_38_1/_24_  (.A(\u_multiplier/STAGE1/_1043_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_38_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_38_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_38_1/_25_  (.A(\u_multiplier/STAGE1/pp1_37_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_38_1/_16_ ),
    .ZN(\u_multiplier/pp1_38 [4]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_38_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_38_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_38_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_38_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_38_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_38_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_38_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_38_1/_17_ ),
    .ZN(\u_multiplier/pp1_39 [9]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_38_2/_18_  (.A(\u_multiplier/STAGE1/pp1_37_e42_2_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_38_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_38_2/_19_  (.A1(\u_multiplier/STAGE1/_1045_ ),
    .A2(\u_multiplier/STAGE1/_1044_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_38_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_38_2/_20_  (.A(\u_multiplier/STAGE1/_1045_ ),
    .B(\u_multiplier/STAGE1/_1044_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_38_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_38_2/_21_  (.A1(\u_multiplier/STAGE1/_1046_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_38_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_38_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_38_2/_22_  (.A(\u_multiplier/STAGE1/_1046_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_38_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_38_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_38_2/_23_  (.A1(\u_multiplier/STAGE1/_1047_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_38_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_38_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_38_2/_24_  (.A(\u_multiplier/STAGE1/_1047_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_38_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_38_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_38_2/_25_  (.A(\u_multiplier/STAGE1/pp1_37_e42_2_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_38_2/_16_ ),
    .ZN(\u_multiplier/pp1_38 [3]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_38_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_38_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_38_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_38_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_38_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_38_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_38_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_38_2/_17_ ),
    .ZN(\u_multiplier/pp1_39 [8]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_38_3/_18_  (.A(\u_multiplier/STAGE1/pp1_37_e42_3_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_38_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_38_3/_19_  (.A1(\u_multiplier/STAGE1/_1049_ ),
    .A2(\u_multiplier/STAGE1/_1048_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_38_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_38_3/_20_  (.A(\u_multiplier/STAGE1/_1049_ ),
    .B(\u_multiplier/STAGE1/_1048_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_38_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_38_3/_21_  (.A1(\u_multiplier/STAGE1/_1050_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_38_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_38_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_38_3/_22_  (.A(\u_multiplier/STAGE1/_1050_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_38_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_38_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_38_3/_23_  (.A1(\u_multiplier/STAGE1/_1051_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_38_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_38_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_38_3/_24_  (.A(\u_multiplier/STAGE1/_1051_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_38_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_38_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_38_3/_25_  (.A(\u_multiplier/STAGE1/pp1_37_e42_3_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_38_3/_16_ ),
    .ZN(\u_multiplier/pp1_38 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_38_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_38_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_38_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_38_e42_3_cout ));
 OAI21_X1 \u_multiplier/STAGE1/E_4_2_pp_38_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_38_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_38_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_38_3/_17_ ),
    .ZN(\u_multiplier/pp1_39 [7]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_38_4/_18_  (.A(\u_multiplier/STAGE1/pp1_37_e42_4_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_38_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_38_4/_19_  (.A1(\u_multiplier/STAGE1/_1053_ ),
    .A2(\u_multiplier/STAGE1/_1052_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_38_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_38_4/_20_  (.A(\u_multiplier/STAGE1/_1053_ ),
    .B(\u_multiplier/STAGE1/_1052_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_38_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_38_4/_21_  (.A1(\u_multiplier/STAGE1/_1054_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_38_4/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_38_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_38_4/_22_  (.A(\u_multiplier/STAGE1/_1054_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_38_4/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_38_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_38_4/_23_  (.A1(\u_multiplier/STAGE1/_1055_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_38_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_38_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_38_4/_24_  (.A(\u_multiplier/STAGE1/_1055_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_38_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_38_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_38_4/_25_  (.A(\u_multiplier/STAGE1/pp1_37_e42_4_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_38_4/_16_ ),
    .ZN(\u_multiplier/pp1_38 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_38_4/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_38_4/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_38_4/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_38_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_38_4/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_38_4/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_38_4/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_38_4/_17_ ),
    .ZN(\u_multiplier/pp1_39 [6]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_38_5/_18_  (.A(\u_multiplier/STAGE1/pp1_37_e42_5_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_38_5/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_38_5/_19_  (.A1(\u_multiplier/STAGE1/_1057_ ),
    .A2(\u_multiplier/STAGE1/_1056_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_38_5/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_38_5/_20_  (.A(\u_multiplier/STAGE1/_1057_ ),
    .B(\u_multiplier/STAGE1/_1056_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_38_5/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_38_5/_21_  (.A1(\u_multiplier/STAGE1/_1058_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_38_5/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_38_5/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_38_5/_22_  (.A(\u_multiplier/STAGE1/_1058_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_38_5/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_38_5/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_38_5/_23_  (.A1(\u_multiplier/STAGE1/_1059_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_38_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_38_5/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_38_5/_24_  (.A(\u_multiplier/STAGE1/_1059_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_38_5/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_38_5/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_38_5/_25_  (.A(\u_multiplier/STAGE1/pp1_37_e42_5_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_38_5/_16_ ),
    .ZN(\u_multiplier/pp1_38 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_38_5/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_38_5/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_38_5/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_38_e42_5_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_38_5/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_38_5/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_38_5/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_38_5/_17_ ),
    .ZN(\u_multiplier/pp1_39 [5]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_39_1/_18_  (.A(\u_multiplier/STAGE1/pp1_38_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_39_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_39_1/_19_  (.A1(\u_multiplier/STAGE1/_1061_ ),
    .A2(\u_multiplier/STAGE1/_1060_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_39_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_39_1/_20_  (.A(\u_multiplier/STAGE1/_1061_ ),
    .B(\u_multiplier/STAGE1/_1060_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_39_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_39_1/_21_  (.A1(\u_multiplier/STAGE1/_1062_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_39_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_39_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_39_1/_22_  (.A(\u_multiplier/STAGE1/_1062_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_39_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_39_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_39_1/_23_  (.A1(\u_multiplier/STAGE1/_1063_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_39_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_39_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_39_1/_24_  (.A(\u_multiplier/STAGE1/_1063_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_39_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_39_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_39_1/_25_  (.A(\u_multiplier/STAGE1/pp1_38_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_39_1/_16_ ),
    .ZN(\u_multiplier/pp1_39 [4]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_39_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_39_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_39_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_39_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_39_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_39_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_39_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_39_1/_17_ ),
    .ZN(\u_multiplier/pp1_40 [8]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_39_2/_18_  (.A(\u_multiplier/STAGE1/pp1_38_e42_2_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_39_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_39_2/_19_  (.A1(\u_multiplier/STAGE1/_1065_ ),
    .A2(\u_multiplier/STAGE1/_1064_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_39_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_39_2/_20_  (.A(\u_multiplier/STAGE1/_1065_ ),
    .B(\u_multiplier/STAGE1/_1064_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_39_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_39_2/_21_  (.A1(\u_multiplier/STAGE1/_1066_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_39_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_39_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_39_2/_22_  (.A(\u_multiplier/STAGE1/_1066_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_39_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_39_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_39_2/_23_  (.A1(\u_multiplier/STAGE1/_1067_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_39_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_39_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_39_2/_24_  (.A(\u_multiplier/STAGE1/_1067_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_39_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_39_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_39_2/_25_  (.A(\u_multiplier/STAGE1/pp1_38_e42_2_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_39_2/_16_ ),
    .ZN(\u_multiplier/pp1_39 [3]));
 NAND2_X2 \u_multiplier/STAGE1/E_4_2_pp_39_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_39_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_39_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_39_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_39_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_39_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_39_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_39_2/_17_ ),
    .ZN(\u_multiplier/pp1_40 [7]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_39_3/_18_  (.A(\u_multiplier/STAGE1/pp1_38_e42_3_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_39_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_39_3/_19_  (.A1(\u_multiplier/STAGE1/_1069_ ),
    .A2(\u_multiplier/STAGE1/_1068_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_39_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_39_3/_20_  (.A(\u_multiplier/STAGE1/_1069_ ),
    .B(\u_multiplier/STAGE1/_1068_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_39_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_39_3/_21_  (.A1(\u_multiplier/STAGE1/_1070_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_39_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_39_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_39_3/_22_  (.A(\u_multiplier/STAGE1/_1070_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_39_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_39_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_39_3/_23_  (.A1(\u_multiplier/STAGE1/_1071_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_39_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_39_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_39_3/_24_  (.A(\u_multiplier/STAGE1/_1071_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_39_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_39_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_39_3/_25_  (.A(\u_multiplier/STAGE1/pp1_38_e42_3_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_39_3/_16_ ),
    .ZN(\u_multiplier/pp1_39 [2]));
 NAND2_X2 \u_multiplier/STAGE1/E_4_2_pp_39_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_39_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_39_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_39_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_39_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_39_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_39_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_39_3/_17_ ),
    .ZN(\u_multiplier/pp1_40 [6]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_39_4/_18_  (.A(\u_multiplier/STAGE1/pp1_38_e42_4_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_39_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_39_4/_19_  (.A1(\u_multiplier/STAGE1/_1073_ ),
    .A2(\u_multiplier/STAGE1/_1072_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_39_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_39_4/_20_  (.A(\u_multiplier/STAGE1/_1073_ ),
    .B(\u_multiplier/STAGE1/_1072_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_39_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_39_4/_21_  (.A1(\u_multiplier/STAGE1/_1074_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_39_4/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_39_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_39_4/_22_  (.A(\u_multiplier/STAGE1/_1074_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_39_4/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_39_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_39_4/_23_  (.A1(\u_multiplier/STAGE1/_1075_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_39_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_39_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_39_4/_24_  (.A(\u_multiplier/STAGE1/_1075_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_39_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_39_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_39_4/_25_  (.A(\u_multiplier/STAGE1/pp1_38_e42_4_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_39_4/_16_ ),
    .ZN(\u_multiplier/pp1_39 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_39_4/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_39_4/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_39_4/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_39_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_39_4/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_39_4/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_39_4/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_39_4/_17_ ),
    .ZN(\u_multiplier/pp1_40 [5]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_40_1/_18_  (.A(\u_multiplier/STAGE1/pp1_39_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_40_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_40_1/_19_  (.A1(\u_multiplier/STAGE1/_1079_ ),
    .A2(\u_multiplier/STAGE1/_1078_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_40_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_40_1/_20_  (.A(\u_multiplier/STAGE1/_1079_ ),
    .B(\u_multiplier/STAGE1/_1078_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_40_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_40_1/_21_  (.A1(\u_multiplier/STAGE1/_1080_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_40_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_40_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_40_1/_22_  (.A(\u_multiplier/STAGE1/_1080_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_40_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_40_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_40_1/_23_  (.A1(\u_multiplier/STAGE1/_1081_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_40_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_40_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_40_1/_24_  (.A(\u_multiplier/STAGE1/_1081_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_40_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_40_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_40_1/_25_  (.A(\u_multiplier/STAGE1/pp1_39_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_40_1/_16_ ),
    .ZN(\u_multiplier/pp1_40 [3]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_40_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_40_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_40_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_40_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE1/E_4_2_pp_40_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_40_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_40_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_40_1/_17_ ),
    .ZN(\u_multiplier/pp1_41 [7]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_40_2/_18_  (.A(\u_multiplier/STAGE1/pp1_39_e42_2_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_40_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_40_2/_19_  (.A1(\u_multiplier/STAGE1/_1083_ ),
    .A2(\u_multiplier/STAGE1/_1082_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_40_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_40_2/_20_  (.A(\u_multiplier/STAGE1/_1083_ ),
    .B(\u_multiplier/STAGE1/_1082_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_40_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_40_2/_21_  (.A1(\u_multiplier/STAGE1/_1084_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_40_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_40_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_40_2/_22_  (.A(\u_multiplier/STAGE1/_1084_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_40_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_40_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_40_2/_23_  (.A1(\u_multiplier/STAGE1/_1085_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_40_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_40_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_40_2/_24_  (.A(\u_multiplier/STAGE1/_1085_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_40_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_40_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_40_2/_25_  (.A(\u_multiplier/STAGE1/pp1_39_e42_2_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_40_2/_16_ ),
    .ZN(\u_multiplier/pp1_40 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_40_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_40_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_40_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_40_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_40_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_40_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_40_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_40_2/_17_ ),
    .ZN(\u_multiplier/pp1_41 [6]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_40_3/_18_  (.A(\u_multiplier/STAGE1/pp1_39_e42_3_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_40_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_40_3/_19_  (.A1(\u_multiplier/STAGE1/_1087_ ),
    .A2(\u_multiplier/STAGE1/_1086_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_40_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_40_3/_20_  (.A(\u_multiplier/STAGE1/_1087_ ),
    .B(\u_multiplier/STAGE1/_1086_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_40_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_40_3/_21_  (.A1(\u_multiplier/STAGE1/_1088_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_40_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_40_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_40_3/_22_  (.A(\u_multiplier/STAGE1/_1088_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_40_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_40_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_40_3/_23_  (.A1(\u_multiplier/STAGE1/_1089_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_40_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_40_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_40_3/_24_  (.A(\u_multiplier/STAGE1/_1089_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_40_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_40_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_40_3/_25_  (.A(\u_multiplier/STAGE1/pp1_39_e42_3_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_40_3/_16_ ),
    .ZN(\u_multiplier/pp1_40 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_40_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_40_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_40_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_40_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_40_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_40_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_40_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_40_3/_17_ ),
    .ZN(\u_multiplier/pp1_41 [5]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_40_4/_18_  (.A(\u_multiplier/STAGE1/pp1_39_e42_4_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_40_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_40_4/_19_  (.A1(\u_multiplier/STAGE1/_1091_ ),
    .A2(\u_multiplier/STAGE1/_1090_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_40_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_40_4/_20_  (.A(\u_multiplier/STAGE1/_1091_ ),
    .B(\u_multiplier/STAGE1/_1090_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_40_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_40_4/_21_  (.A1(\u_multiplier/STAGE1/_1092_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_40_4/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_40_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_40_4/_22_  (.A(\u_multiplier/STAGE1/_1092_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_40_4/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_40_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_40_4/_23_  (.A1(\u_multiplier/STAGE1/_1093_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_40_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_40_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_40_4/_24_  (.A(\u_multiplier/STAGE1/_1093_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_40_4/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_40_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_40_4/_25_  (.A(\u_multiplier/STAGE1/pp1_39_e42_4_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_40_4/_16_ ),
    .ZN(\u_multiplier/pp1_40 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_40_4/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_40_4/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_40_4/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_40_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_40_4/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_40_4/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_40_4/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_40_4/_17_ ),
    .ZN(\u_multiplier/pp1_41 [4]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_41_1/_18_  (.A(\u_multiplier/STAGE1/pp1_40_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_41_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_41_1/_19_  (.A1(\u_multiplier/STAGE1/_1095_ ),
    .A2(\u_multiplier/STAGE1/_1094_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_41_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_41_1/_20_  (.A(\u_multiplier/STAGE1/_1095_ ),
    .B(\u_multiplier/STAGE1/_1094_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_41_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_41_1/_21_  (.A1(\u_multiplier/STAGE1/_1096_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_41_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_41_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_41_1/_22_  (.A(\u_multiplier/STAGE1/_1096_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_41_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_41_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_41_1/_23_  (.A1(\u_multiplier/STAGE1/_1097_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_41_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_41_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_41_1/_24_  (.A(\u_multiplier/STAGE1/_1097_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_41_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_41_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_41_1/_25_  (.A(\u_multiplier/STAGE1/pp1_40_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_41_1/_16_ ),
    .ZN(\u_multiplier/pp1_41 [3]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_41_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_41_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_41_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_41_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_41_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_41_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_41_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_41_1/_17_ ),
    .ZN(\u_multiplier/pp1_42 [6]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_41_2/_18_  (.A(\u_multiplier/STAGE1/pp1_40_e42_2_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_41_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_41_2/_19_  (.A1(\u_multiplier/STAGE1/_1099_ ),
    .A2(\u_multiplier/STAGE1/_1098_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_41_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_41_2/_20_  (.A(\u_multiplier/STAGE1/_1099_ ),
    .B(\u_multiplier/STAGE1/_1098_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_41_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_41_2/_21_  (.A1(\u_multiplier/STAGE1/_1100_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_41_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_41_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_41_2/_22_  (.A(\u_multiplier/STAGE1/_1100_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_41_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_41_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_41_2/_23_  (.A1(\u_multiplier/STAGE1/_1101_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_41_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_41_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_41_2/_24_  (.A(\u_multiplier/STAGE1/_1101_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_41_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_41_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_41_2/_25_  (.A(\u_multiplier/STAGE1/pp1_40_e42_2_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_41_2/_16_ ),
    .ZN(\u_multiplier/pp1_41 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_41_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_41_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_41_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_41_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_41_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_41_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_41_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_41_2/_17_ ),
    .ZN(\u_multiplier/pp1_42 [5]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_41_3/_18_  (.A(\u_multiplier/STAGE1/pp1_40_e42_3_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_41_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_41_3/_19_  (.A1(\u_multiplier/STAGE1/_1103_ ),
    .A2(\u_multiplier/STAGE1/_1102_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_41_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_41_3/_20_  (.A(\u_multiplier/STAGE1/_1103_ ),
    .B(\u_multiplier/STAGE1/_1102_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_41_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_41_3/_21_  (.A1(\u_multiplier/STAGE1/_1104_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_41_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_41_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_41_3/_22_  (.A(\u_multiplier/STAGE1/_1104_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_41_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_41_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_41_3/_23_  (.A1(\u_multiplier/STAGE1/_1105_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_41_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_41_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_41_3/_24_  (.A(\u_multiplier/STAGE1/_1105_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_41_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_41_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_41_3/_25_  (.A(\u_multiplier/STAGE1/pp1_40_e42_3_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_41_3/_16_ ),
    .ZN(\u_multiplier/pp1_41 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_41_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_41_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_41_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_41_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_41_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_41_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_41_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_41_3/_17_ ),
    .ZN(\u_multiplier/pp1_42 [4]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_42_1/_18_  (.A(\u_multiplier/STAGE1/pp1_41_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_42_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_42_1/_19_  (.A1(\u_multiplier/STAGE1/_1109_ ),
    .A2(\u_multiplier/STAGE1/_1108_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_42_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_42_1/_20_  (.A(\u_multiplier/STAGE1/_1109_ ),
    .B(\u_multiplier/STAGE1/_1108_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_42_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_42_1/_21_  (.A1(\u_multiplier/STAGE1/_1110_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_42_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_42_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_42_1/_22_  (.A(\u_multiplier/STAGE1/_1110_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_42_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_42_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_42_1/_23_  (.A1(\u_multiplier/STAGE1/_1111_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_42_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_42_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_42_1/_24_  (.A(\u_multiplier/STAGE1/_1111_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_42_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_42_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_42_1/_25_  (.A(\u_multiplier/STAGE1/pp1_41_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_42_1/_16_ ),
    .ZN(\u_multiplier/pp1_42 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_42_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_42_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_42_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_42_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_42_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_42_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_42_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_42_1/_17_ ),
    .ZN(\u_multiplier/pp1_43 [5]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_42_2/_18_  (.A(\u_multiplier/STAGE1/pp1_41_e42_2_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_42_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_42_2/_19_  (.A1(\u_multiplier/STAGE1/_1113_ ),
    .A2(\u_multiplier/STAGE1/_1112_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_42_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_42_2/_20_  (.A(\u_multiplier/STAGE1/_1113_ ),
    .B(\u_multiplier/STAGE1/_1112_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_42_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_42_2/_21_  (.A1(\u_multiplier/STAGE1/_1114_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_42_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_42_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_42_2/_22_  (.A(\u_multiplier/STAGE1/_1114_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_42_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_42_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_42_2/_23_  (.A1(\u_multiplier/STAGE1/_1115_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_42_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_42_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_42_2/_24_  (.A(\u_multiplier/STAGE1/_1115_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_42_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_42_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_42_2/_25_  (.A(\u_multiplier/STAGE1/pp1_41_e42_2_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_42_2/_16_ ),
    .ZN(\u_multiplier/pp1_42 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_42_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_42_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_42_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_42_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_42_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_42_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_42_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_42_2/_17_ ),
    .ZN(\u_multiplier/pp1_43 [4]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_42_3/_18_  (.A(\u_multiplier/STAGE1/pp1_41_e42_3_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_42_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_42_3/_19_  (.A1(\u_multiplier/STAGE1/_1117_ ),
    .A2(\u_multiplier/STAGE1/_1116_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_42_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_42_3/_20_  (.A(\u_multiplier/STAGE1/_1117_ ),
    .B(\u_multiplier/STAGE1/_1116_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_42_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_42_3/_21_  (.A1(\u_multiplier/STAGE1/_1118_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_42_3/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_42_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_42_3/_22_  (.A(\u_multiplier/STAGE1/_1118_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_42_3/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_42_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_42_3/_23_  (.A1(\u_multiplier/STAGE1/_1119_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_42_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_42_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_42_3/_24_  (.A(\u_multiplier/STAGE1/_1119_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_42_3/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_42_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_42_3/_25_  (.A(\u_multiplier/STAGE1/pp1_41_e42_3_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_42_3/_16_ ),
    .ZN(\u_multiplier/pp1_42 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_42_3/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_42_3/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_42_3/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_42_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_42_3/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_42_3/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_42_3/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_42_3/_17_ ),
    .ZN(\u_multiplier/pp1_43 [3]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_43_1/_18_  (.A(\u_multiplier/STAGE1/pp1_42_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_43_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_43_1/_19_  (.A1(\u_multiplier/STAGE1/_1121_ ),
    .A2(\u_multiplier/STAGE1/_1120_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_43_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_43_1/_20_  (.A(\u_multiplier/STAGE1/_1121_ ),
    .B(\u_multiplier/STAGE1/_1120_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_43_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_43_1/_21_  (.A1(\u_multiplier/STAGE1/_1122_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_43_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_43_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_43_1/_22_  (.A(\u_multiplier/STAGE1/_1122_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_43_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_43_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_43_1/_23_  (.A1(\u_multiplier/STAGE1/_1123_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_43_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_43_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_43_1/_24_  (.A(\u_multiplier/STAGE1/_1123_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_43_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_43_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_43_1/_25_  (.A(\u_multiplier/STAGE1/pp1_42_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_43_1/_16_ ),
    .ZN(\u_multiplier/pp1_43 [2]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_43_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_43_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_43_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_43_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_43_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_43_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_43_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_43_1/_17_ ),
    .ZN(\u_multiplier/pp1_44 [4]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_43_2/_18_  (.A(\u_multiplier/STAGE1/pp1_42_e42_2_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_43_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_43_2/_19_  (.A1(\u_multiplier/STAGE1/_1125_ ),
    .A2(\u_multiplier/STAGE1/_1124_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_43_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_43_2/_20_  (.A(\u_multiplier/STAGE1/_1125_ ),
    .B(\u_multiplier/STAGE1/_1124_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_43_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_43_2/_21_  (.A1(\u_multiplier/STAGE1/_1126_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_43_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_43_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_43_2/_22_  (.A(\u_multiplier/STAGE1/_1126_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_43_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_43_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_43_2/_23_  (.A1(\u_multiplier/STAGE1/_1127_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_43_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_43_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_43_2/_24_  (.A(\u_multiplier/STAGE1/_1127_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_43_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_43_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_43_2/_25_  (.A(\u_multiplier/STAGE1/pp1_42_e42_2_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_43_2/_16_ ),
    .ZN(\u_multiplier/pp1_43 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_43_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_43_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_43_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_43_e42_2_cout ));
 OAI21_X1 \u_multiplier/STAGE1/E_4_2_pp_43_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_43_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_43_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_43_2/_17_ ),
    .ZN(\u_multiplier/pp1_44 [3]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_44_1/_18_  (.A(\u_multiplier/STAGE1/pp1_43_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_44_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_44_1/_19_  (.A1(\u_multiplier/STAGE1/_1131_ ),
    .A2(\u_multiplier/STAGE1/_1130_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_44_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_44_1/_20_  (.A(\u_multiplier/STAGE1/_1131_ ),
    .B(\u_multiplier/STAGE1/_1130_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_44_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_44_1/_21_  (.A1(\u_multiplier/STAGE1/_1132_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_44_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_44_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_44_1/_22_  (.A(\u_multiplier/STAGE1/_1132_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_44_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_44_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_44_1/_23_  (.A1(\u_multiplier/STAGE1/_1133_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_44_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_44_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_44_1/_24_  (.A(\u_multiplier/STAGE1/_1133_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_44_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_44_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_44_1/_25_  (.A(\u_multiplier/STAGE1/pp1_43_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_44_1/_16_ ),
    .ZN(\u_multiplier/pp1_44 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_44_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_44_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_44_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_44_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_44_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_44_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_44_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_44_1/_17_ ),
    .ZN(\u_multiplier/pp1_45 [3]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_44_2/_18_  (.A(\u_multiplier/STAGE1/pp1_43_e42_2_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_44_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_44_2/_19_  (.A1(\u_multiplier/STAGE1/_1135_ ),
    .A2(\u_multiplier/STAGE1/_1134_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_44_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_44_2/_20_  (.A(\u_multiplier/STAGE1/_1135_ ),
    .B(\u_multiplier/STAGE1/_1134_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_44_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_44_2/_21_  (.A1(\u_multiplier/STAGE1/_1136_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_44_2/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_44_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_44_2/_22_  (.A(\u_multiplier/STAGE1/_1136_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_44_2/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_44_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_44_2/_23_  (.A1(\u_multiplier/STAGE1/_1137_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_44_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_44_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_44_2/_24_  (.A(\u_multiplier/STAGE1/_1137_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_44_2/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_44_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_44_2/_25_  (.A(\u_multiplier/STAGE1/pp1_43_e42_2_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_44_2/_16_ ),
    .ZN(\u_multiplier/pp1_44 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_44_2/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_44_2/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_44_2/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_44_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_44_2/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_44_2/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_44_2/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_44_2/_17_ ),
    .ZN(\u_multiplier/pp1_45 [2]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_45_1/_18_  (.A(\u_multiplier/STAGE1/pp1_44_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_45_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_45_1/_19_  (.A1(\u_multiplier/STAGE1/_1139_ ),
    .A2(\u_multiplier/STAGE1/_1138_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_45_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_45_1/_20_  (.A(\u_multiplier/STAGE1/_1139_ ),
    .B(\u_multiplier/STAGE1/_1138_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_45_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_45_1/_21_  (.A1(\u_multiplier/STAGE1/_1140_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_45_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_45_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_45_1/_22_  (.A(\u_multiplier/STAGE1/_1140_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_45_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_45_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_45_1/_23_  (.A1(\u_multiplier/STAGE1/_1141_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_45_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_45_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_45_1/_24_  (.A(\u_multiplier/STAGE1/_1141_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_45_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_45_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_45_1/_25_  (.A(\u_multiplier/STAGE1/pp1_44_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_45_1/_16_ ),
    .ZN(\u_multiplier/pp1_45 [1]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_45_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_45_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_45_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_45_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_45_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_45_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_45_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_45_1/_17_ ),
    .ZN(\u_multiplier/pp1_46 [2]));
 INV_X1 \u_multiplier/STAGE1/E_4_2_pp_46_1/_18_  (.A(\u_multiplier/STAGE1/pp1_45_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_46_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_46_1/_19_  (.A1(\u_multiplier/STAGE1/_1145_ ),
    .A2(\u_multiplier/STAGE1/_1144_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_46_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_46_1/_20_  (.A(\u_multiplier/STAGE1/_1145_ ),
    .B(\u_multiplier/STAGE1/_1144_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_46_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_46_1/_21_  (.A1(\u_multiplier/STAGE1/_1146_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_46_1/_12_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_46_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_46_1/_22_  (.A(\u_multiplier/STAGE1/_1146_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_46_1/_12_ ),
    .Z(\u_multiplier/STAGE1/E_4_2_pp_46_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_46_1/_23_  (.A1(\u_multiplier/STAGE1/_1147_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_46_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_46_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_46_1/_24_  (.A(\u_multiplier/STAGE1/_1147_ ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_46_1/_14_ ),
    .ZN(\u_multiplier/STAGE1/E_4_2_pp_46_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE1/E_4_2_pp_46_1/_25_  (.A(\u_multiplier/STAGE1/pp1_45_e42_1_cout ),
    .B(\u_multiplier/STAGE1/E_4_2_pp_46_1/_16_ ),
    .ZN(\u_multiplier/pp1_46 [0]));
 NAND2_X1 \u_multiplier/STAGE1/E_4_2_pp_46_1/_26_  (.A1(\u_multiplier/STAGE1/E_4_2_pp_46_1/_11_ ),
    .A2(\u_multiplier/STAGE1/E_4_2_pp_46_1/_13_ ),
    .ZN(\u_multiplier/STAGE1/pp1_46_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE1/E_4_2_pp_46_1/_27_  (.A(\u_multiplier/STAGE1/E_4_2_pp_46_1/_15_ ),
    .B1(\u_multiplier/STAGE1/E_4_2_pp_46_1/_16_ ),
    .B2(\u_multiplier/STAGE1/E_4_2_pp_46_1/_17_ ),
    .ZN(\u_multiplier/pp1_47 [1]));
 INV_X1 \u_multiplier/STAGE1/Full_adder_pp_33_1/_12_  (.A(\u_multiplier/STAGE1/pp1_32_e42_8_cout ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_33_1/_08_ ));
 NAND3_X2 \u_multiplier/STAGE1/Full_adder_pp_33_1/_13_  (.A1(\u_multiplier/STAGE1/_0939_ ),
    .A2(\u_multiplier/STAGE1/_0938_ ),
    .A3(\u_multiplier/STAGE1/pp1_32_e42_8_cout ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_33_1/_09_ ));
 NOR2_X4 \u_multiplier/STAGE1/Full_adder_pp_33_1/_14_  (.A1(\u_multiplier/STAGE1/_0939_ ),
    .A2(\u_multiplier/STAGE1/_0938_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_33_1/_10_ ));
 AOI21_X2 \u_multiplier/STAGE1/Full_adder_pp_33_1/_15_  (.A(\u_multiplier/STAGE1/pp1_32_e42_8_cout ),
    .B1(\u_multiplier/STAGE1/_0938_ ),
    .B2(\u_multiplier/STAGE1/_0939_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_33_1/_11_ ));
 NOR2_X4 \u_multiplier/STAGE1/Full_adder_pp_33_1/_16_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_33_1/_10_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_33_1/_11_ ),
    .ZN(\u_multiplier/pp1_34 [7]));
 AOI22_X4 \u_multiplier/STAGE1/Full_adder_pp_33_1/_17_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_33_1/_08_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_33_1/_10_ ),
    .B1(\u_multiplier/pp1_34 [7]),
    .B2(\u_multiplier/STAGE1/Full_adder_pp_33_1/_09_ ),
    .ZN(\u_multiplier/pp1_33 [0]));
 INV_X1 \u_multiplier/STAGE1/Full_adder_pp_35_1/_12_  (.A(\u_multiplier/STAGE1/pp1_34_e42_7_cout ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_35_1/_08_ ));
 NAND3_X2 \u_multiplier/STAGE1/Full_adder_pp_35_1/_13_  (.A1(\u_multiplier/STAGE1/_0993_ ),
    .A2(\u_multiplier/STAGE1/_0992_ ),
    .A3(\u_multiplier/STAGE1/pp1_34_e42_7_cout ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_35_1/_09_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_35_1/_14_  (.A1(\u_multiplier/STAGE1/_0993_ ),
    .A2(\u_multiplier/STAGE1/_0992_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_35_1/_10_ ));
 AOI21_X1 \u_multiplier/STAGE1/Full_adder_pp_35_1/_15_  (.A(\u_multiplier/STAGE1/pp1_34_e42_7_cout ),
    .B1(\u_multiplier/STAGE1/_0992_ ),
    .B2(\u_multiplier/STAGE1/_0993_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_35_1/_11_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_35_1/_16_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_35_1/_10_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_35_1/_11_ ),
    .ZN(\u_multiplier/pp1_36 [6]));
 AOI22_X4 \u_multiplier/STAGE1/Full_adder_pp_35_1/_17_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_35_1/_08_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_35_1/_10_ ),
    .B1(\u_multiplier/pp1_36 [6]),
    .B2(\u_multiplier/STAGE1/Full_adder_pp_35_1/_09_ ),
    .ZN(\u_multiplier/pp1_35 [0]));
 INV_X1 \u_multiplier/STAGE1/Full_adder_pp_37_1/_12_  (.A(\u_multiplier/STAGE1/pp1_36_e42_6_cout ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_37_1/_08_ ));
 NAND3_X1 \u_multiplier/STAGE1/Full_adder_pp_37_1/_13_  (.A1(\u_multiplier/STAGE1/_1039_ ),
    .A2(\u_multiplier/STAGE1/_1038_ ),
    .A3(\u_multiplier/STAGE1/pp1_36_e42_6_cout ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_37_1/_09_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_37_1/_14_  (.A1(\u_multiplier/STAGE1/_1039_ ),
    .A2(\u_multiplier/STAGE1/_1038_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_37_1/_10_ ));
 AOI21_X1 \u_multiplier/STAGE1/Full_adder_pp_37_1/_15_  (.A(\u_multiplier/STAGE1/pp1_36_e42_6_cout ),
    .B1(\u_multiplier/STAGE1/_1038_ ),
    .B2(\u_multiplier/STAGE1/_1039_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_37_1/_11_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_37_1/_16_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_37_1/_10_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_37_1/_11_ ),
    .ZN(\u_multiplier/pp1_38 [5]));
 AOI22_X2 \u_multiplier/STAGE1/Full_adder_pp_37_1/_17_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_37_1/_08_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_37_1/_10_ ),
    .B1(\u_multiplier/pp1_38 [5]),
    .B2(\u_multiplier/STAGE1/Full_adder_pp_37_1/_09_ ),
    .ZN(\u_multiplier/pp1_37 [0]));
 INV_X1 \u_multiplier/STAGE1/Full_adder_pp_39_1/_12_  (.A(\u_multiplier/STAGE1/pp1_38_e42_5_cout ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_39_1/_08_ ));
 NAND3_X2 \u_multiplier/STAGE1/Full_adder_pp_39_1/_13_  (.A1(\u_multiplier/STAGE1/_1077_ ),
    .A2(\u_multiplier/STAGE1/_1076_ ),
    .A3(\u_multiplier/STAGE1/pp1_38_e42_5_cout ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_39_1/_09_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_39_1/_14_  (.A1(\u_multiplier/STAGE1/_1077_ ),
    .A2(\u_multiplier/STAGE1/_1076_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_39_1/_10_ ));
 AOI21_X1 \u_multiplier/STAGE1/Full_adder_pp_39_1/_15_  (.A(\u_multiplier/STAGE1/pp1_38_e42_5_cout ),
    .B1(\u_multiplier/STAGE1/_1076_ ),
    .B2(\u_multiplier/STAGE1/_1077_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_39_1/_11_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_39_1/_16_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_39_1/_10_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_39_1/_11_ ),
    .ZN(\u_multiplier/pp1_40 [4]));
 AOI22_X4 \u_multiplier/STAGE1/Full_adder_pp_39_1/_17_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_39_1/_08_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_39_1/_10_ ),
    .B1(\u_multiplier/pp1_40 [4]),
    .B2(\u_multiplier/STAGE1/Full_adder_pp_39_1/_09_ ),
    .ZN(\u_multiplier/pp1_39 [0]));
 INV_X1 \u_multiplier/STAGE1/Full_adder_pp_41_1/_12_  (.A(\u_multiplier/STAGE1/pp1_40_e42_4_cout ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_41_1/_08_ ));
 NAND3_X2 \u_multiplier/STAGE1/Full_adder_pp_41_1/_13_  (.A1(\u_multiplier/STAGE1/_1107_ ),
    .A2(\u_multiplier/STAGE1/_1106_ ),
    .A3(\u_multiplier/STAGE1/pp1_40_e42_4_cout ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_41_1/_09_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_41_1/_14_  (.A1(\u_multiplier/STAGE1/_1107_ ),
    .A2(\u_multiplier/STAGE1/_1106_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_41_1/_10_ ));
 AOI21_X1 \u_multiplier/STAGE1/Full_adder_pp_41_1/_15_  (.A(\u_multiplier/STAGE1/pp1_40_e42_4_cout ),
    .B1(\u_multiplier/STAGE1/_1106_ ),
    .B2(\u_multiplier/STAGE1/_1107_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_41_1/_11_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_41_1/_16_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_41_1/_10_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_41_1/_11_ ),
    .ZN(\u_multiplier/pp1_42 [3]));
 AOI22_X4 \u_multiplier/STAGE1/Full_adder_pp_41_1/_17_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_41_1/_08_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_41_1/_10_ ),
    .B1(\u_multiplier/pp1_42 [3]),
    .B2(\u_multiplier/STAGE1/Full_adder_pp_41_1/_09_ ),
    .ZN(\u_multiplier/pp1_41 [0]));
 INV_X1 \u_multiplier/STAGE1/Full_adder_pp_43_1/_12_  (.A(\u_multiplier/STAGE1/pp1_42_e42_3_cout ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_43_1/_08_ ));
 NAND3_X2 \u_multiplier/STAGE1/Full_adder_pp_43_1/_13_  (.A1(\u_multiplier/STAGE1/_1129_ ),
    .A2(\u_multiplier/STAGE1/_1128_ ),
    .A3(\u_multiplier/STAGE1/pp1_42_e42_3_cout ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_43_1/_09_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_43_1/_14_  (.A1(\u_multiplier/STAGE1/_1129_ ),
    .A2(\u_multiplier/STAGE1/_1128_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_43_1/_10_ ));
 AOI21_X1 \u_multiplier/STAGE1/Full_adder_pp_43_1/_15_  (.A(\u_multiplier/STAGE1/pp1_42_e42_3_cout ),
    .B1(\u_multiplier/STAGE1/_1128_ ),
    .B2(\u_multiplier/STAGE1/_1129_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_43_1/_11_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_43_1/_16_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_43_1/_10_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_43_1/_11_ ),
    .ZN(\u_multiplier/pp1_44 [2]));
 AOI22_X4 \u_multiplier/STAGE1/Full_adder_pp_43_1/_17_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_43_1/_08_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_43_1/_10_ ),
    .B1(\u_multiplier/pp1_44 [2]),
    .B2(\u_multiplier/STAGE1/Full_adder_pp_43_1/_09_ ),
    .ZN(\u_multiplier/pp1_43 [0]));
 INV_X1 \u_multiplier/STAGE1/Full_adder_pp_45_1/_12_  (.A(\u_multiplier/STAGE1/pp1_44_e42_2_cout ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_45_1/_08_ ));
 NAND3_X1 \u_multiplier/STAGE1/Full_adder_pp_45_1/_13_  (.A1(\u_multiplier/STAGE1/_1143_ ),
    .A2(\u_multiplier/STAGE1/_1142_ ),
    .A3(\u_multiplier/STAGE1/pp1_44_e42_2_cout ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_45_1/_09_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_45_1/_14_  (.A1(\u_multiplier/STAGE1/_1143_ ),
    .A2(\u_multiplier/STAGE1/_1142_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_45_1/_10_ ));
 AOI21_X1 \u_multiplier/STAGE1/Full_adder_pp_45_1/_15_  (.A(\u_multiplier/STAGE1/pp1_44_e42_2_cout ),
    .B1(\u_multiplier/STAGE1/_1142_ ),
    .B2(\u_multiplier/STAGE1/_1143_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_45_1/_11_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_45_1/_16_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_45_1/_10_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_45_1/_11_ ),
    .ZN(\u_multiplier/pp1_46 [1]));
 AOI22_X2 \u_multiplier/STAGE1/Full_adder_pp_45_1/_17_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_45_1/_08_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_45_1/_10_ ),
    .B1(\u_multiplier/pp1_46 [1]),
    .B2(\u_multiplier/STAGE1/Full_adder_pp_45_1/_09_ ),
    .ZN(\u_multiplier/pp1_45 [0]));
 INV_X1 \u_multiplier/STAGE1/Full_adder_pp_47_1/_12_  (.A(\u_multiplier/STAGE1/pp1_46_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_47_1/_08_ ));
 NAND3_X2 \u_multiplier/STAGE1/Full_adder_pp_47_1/_13_  (.A1(\u_multiplier/STAGE1/_1149_ ),
    .A2(\u_multiplier/STAGE1/_1148_ ),
    .A3(\u_multiplier/STAGE1/pp1_46_e42_1_cout ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_47_1/_09_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_47_1/_14_  (.A1(\u_multiplier/STAGE1/_1149_ ),
    .A2(\u_multiplier/STAGE1/_1148_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_47_1/_10_ ));
 AOI21_X1 \u_multiplier/STAGE1/Full_adder_pp_47_1/_15_  (.A(\u_multiplier/STAGE1/pp1_46_e42_1_cout ),
    .B1(\u_multiplier/STAGE1/_1148_ ),
    .B2(\u_multiplier/STAGE1/_1149_ ),
    .ZN(\u_multiplier/STAGE1/Full_adder_pp_47_1/_11_ ));
 NOR2_X2 \u_multiplier/STAGE1/Full_adder_pp_47_1/_16_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_47_1/_10_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_47_1/_11_ ),
    .ZN(\u_multiplier/pp1_48 [0]));
 AOI22_X4 \u_multiplier/STAGE1/Full_adder_pp_47_1/_17_  (.A1(\u_multiplier/STAGE1/Full_adder_pp_47_1/_08_ ),
    .A2(\u_multiplier/STAGE1/Full_adder_pp_47_1/_10_ ),
    .B1(\u_multiplier/pp1_48 [0]),
    .B2(\u_multiplier/STAGE1/Full_adder_pp_47_1/_09_ ),
    .ZN(\u_multiplier/pp1_47 [0]));
 AND2_X1 \u_multiplier/STAGE1/Half_adder_pp_16_1/_4_  (.A1(\u_multiplier/STAGE1/_0608_ ),
    .A2(\u_multiplier/STAGE1/_0607_ ),
    .ZN(\u_multiplier/pp1_17 [1]));
 XOR2_X2 \u_multiplier/STAGE1/Half_adder_pp_16_1/_5_  (.A(\u_multiplier/STAGE1/_0608_ ),
    .B(\u_multiplier/STAGE1/_0607_ ),
    .Z(\u_multiplier/pp1_16 [0]));
 AND2_X1 \u_multiplier/STAGE1/Half_adder_pp_18_1/_4_  (.A1(\u_multiplier/STAGE1/_0618_ ),
    .A2(\u_multiplier/STAGE1/_0617_ ),
    .ZN(\u_multiplier/pp1_19 [2]));
 XOR2_X2 \u_multiplier/STAGE1/Half_adder_pp_18_1/_5_  (.A(\u_multiplier/STAGE1/_0618_ ),
    .B(\u_multiplier/STAGE1/_0617_ ),
    .Z(\u_multiplier/pp1_18 [0]));
 AND2_X1 \u_multiplier/STAGE1/Half_adder_pp_20_1/_4_  (.A1(\u_multiplier/STAGE1/_0636_ ),
    .A2(\u_multiplier/STAGE1/_0635_ ),
    .ZN(\u_multiplier/pp1_21 [3]));
 XOR2_X2 \u_multiplier/STAGE1/Half_adder_pp_20_1/_5_  (.A(\u_multiplier/STAGE1/_0636_ ),
    .B(\u_multiplier/STAGE1/_0635_ ),
    .Z(\u_multiplier/pp1_20 [0]));
 AND2_X1 \u_multiplier/STAGE1/Half_adder_pp_22_1/_4_  (.A1(\u_multiplier/STAGE1/_0662_ ),
    .A2(\u_multiplier/STAGE1/_0661_ ),
    .ZN(\u_multiplier/pp1_23 [4]));
 XOR2_X2 \u_multiplier/STAGE1/Half_adder_pp_22_1/_5_  (.A(\u_multiplier/STAGE1/_0662_ ),
    .B(\u_multiplier/STAGE1/_0661_ ),
    .Z(\u_multiplier/pp1_22 [0]));
 AND2_X1 \u_multiplier/STAGE1/Half_adder_pp_24_1/_4_  (.A1(\u_multiplier/STAGE1/_0696_ ),
    .A2(\u_multiplier/STAGE1/_0695_ ),
    .ZN(\u_multiplier/pp1_25 [5]));
 XOR2_X2 \u_multiplier/STAGE1/Half_adder_pp_24_1/_5_  (.A(\u_multiplier/STAGE1/_0696_ ),
    .B(\u_multiplier/STAGE1/_0695_ ),
    .Z(\u_multiplier/pp1_24 [0]));
 AND2_X1 \u_multiplier/STAGE1/Half_adder_pp_26_1/_4_  (.A1(\u_multiplier/STAGE1/_0738_ ),
    .A2(\u_multiplier/STAGE1/_0737_ ),
    .ZN(\u_multiplier/pp1_27 [6]));
 XOR2_X2 \u_multiplier/STAGE1/Half_adder_pp_26_1/_5_  (.A(\u_multiplier/STAGE1/_0738_ ),
    .B(\u_multiplier/STAGE1/_0737_ ),
    .Z(\u_multiplier/pp1_26 [0]));
 AND2_X1 \u_multiplier/STAGE1/Half_adder_pp_28_1/_4_  (.A1(\u_multiplier/STAGE1/_0788_ ),
    .A2(\u_multiplier/STAGE1/_0787_ ),
    .ZN(\u_multiplier/pp1_29 [7]));
 XOR2_X2 \u_multiplier/STAGE1/Half_adder_pp_28_1/_5_  (.A(\u_multiplier/STAGE1/_0788_ ),
    .B(\u_multiplier/STAGE1/_0787_ ),
    .Z(\u_multiplier/pp1_28 [0]));
 AND2_X1 \u_multiplier/STAGE1/Half_adder_pp_30_1/_4_  (.A1(\u_multiplier/STAGE1/_0846_ ),
    .A2(\u_multiplier/STAGE1/_0845_ ),
    .ZN(\u_multiplier/pp1_31 [8]));
 XOR2_X2 \u_multiplier/STAGE1/Half_adder_pp_30_1/_5_  (.A(\u_multiplier/STAGE1/_0846_ ),
    .B(\u_multiplier/STAGE1/_0845_ ),
    .Z(\u_multiplier/pp1_30 [0]));
 AND2_X1 \u_multiplier/STAGE1/_1631_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[0]),
    .ZN(\u_multiplier/pp3_0 ));
 AND2_X1 \u_multiplier/STAGE1/_1632_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[1]),
    .ZN(\u_multiplier/pp3_1 [0]));
 AND2_X1 \u_multiplier/STAGE1/_1633_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[1]),
    .ZN(\u_multiplier/pp3_1 [1]));
 AND2_X1 \u_multiplier/STAGE1/_1634_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[2]),
    .ZN(\u_multiplier/pp3_2 [0]));
 AND2_X1 \u_multiplier/STAGE1/_1635_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[1]),
    .ZN(\u_multiplier/pp3_2 [1]));
 AND2_X1 \u_multiplier/STAGE1/_1636_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[2]),
    .ZN(\u_multiplier/pp3_2 [2]));
 AND2_X1 \u_multiplier/STAGE1/_1637_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[3]),
    .ZN(\u_multiplier/pp3_3 [0]));
 AND2_X1 \u_multiplier/STAGE1/_1638_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[2]),
    .ZN(\u_multiplier/pp3_3 [1]));
 AND2_X1 \u_multiplier/STAGE1/_1639_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[2]),
    .ZN(\u_multiplier/pp3_3 [2]));
 AND2_X1 \u_multiplier/STAGE1/_1640_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[3]),
    .ZN(\u_multiplier/pp3_3 [3]));
 AND2_X1 \u_multiplier/STAGE1/_1641_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[4]),
    .ZN(\u_multiplier/pp3_4 [1]));
 AND2_X1 \u_multiplier/STAGE1/_1642_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[3]),
    .ZN(\u_multiplier/pp3_4 [2]));
 AND2_X1 \u_multiplier/STAGE1/_1643_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[2]),
    .ZN(\u_multiplier/pp3_4 [3]));
 AND2_X1 \u_multiplier/STAGE1/_1644_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[3]),
    .ZN(\u_multiplier/pp2_4 [1]));
 AND2_X1 \u_multiplier/STAGE1/_1645_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[4]),
    .ZN(\u_multiplier/pp2_4 [0]));
 AND2_X1 \u_multiplier/STAGE1/_1646_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[5]),
    .ZN(\u_multiplier/pp3_5 [2]));
 AND2_X1 \u_multiplier/STAGE1/_1647_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[4]),
    .ZN(\u_multiplier/pp3_5 [3]));
 AND2_X1 \u_multiplier/STAGE1/_1648_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[3]),
    .ZN(\u_multiplier/pp2_5 [3]));
 AND2_X1 \u_multiplier/STAGE1/_1649_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[3]),
    .ZN(\u_multiplier/pp2_5 [2]));
 AND2_X1 \u_multiplier/STAGE1/_1650_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[4]),
    .ZN(\u_multiplier/pp2_5 [1]));
 AND2_X1 \u_multiplier/STAGE1/_1651_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[5]),
    .ZN(\u_multiplier/pp2_5 [0]));
 AND2_X1 \u_multiplier/STAGE1/_1652_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[6]),
    .ZN(\u_multiplier/pp3_6 [3]));
 AND2_X1 \u_multiplier/STAGE1/_1653_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[5]),
    .ZN(\u_multiplier/pp2_6 [5]));
 AND2_X1 \u_multiplier/STAGE1/_1654_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[4]),
    .ZN(\u_multiplier/pp2_6 [4]));
 AND2_X1 \u_multiplier/STAGE1/_1655_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[3]),
    .ZN(\u_multiplier/pp2_6 [3]));
 AND2_X1 \u_multiplier/STAGE1/_1656_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[4]),
    .ZN(\u_multiplier/pp2_6 [2]));
 AND2_X1 \u_multiplier/STAGE1/_1657_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[5]),
    .ZN(\u_multiplier/pp2_6 [1]));
 AND2_X1 \u_multiplier/STAGE1/_1658_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[6]),
    .ZN(\u_multiplier/pp2_6 [0]));
 AND2_X1 \u_multiplier/STAGE1/_1659_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[7]),
    .ZN(\u_multiplier/pp2_7 [7]));
 AND2_X1 \u_multiplier/STAGE1/_1660_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[6]),
    .ZN(\u_multiplier/pp2_7 [6]));
 AND2_X1 \u_multiplier/STAGE1/_1661_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[5]),
    .ZN(\u_multiplier/pp2_7 [5]));
 AND2_X1 \u_multiplier/STAGE1/_1662_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[4]),
    .ZN(\u_multiplier/pp2_7 [4]));
 AND2_X1 \u_multiplier/STAGE1/_1663_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[4]),
    .ZN(\u_multiplier/pp2_7 [3]));
 AND2_X1 \u_multiplier/STAGE1/_1664_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[5]),
    .ZN(\u_multiplier/pp2_7 [2]));
 AND2_X1 \u_multiplier/STAGE1/_1665_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[6]),
    .ZN(\u_multiplier/pp2_7 [1]));
 AND2_X1 \u_multiplier/STAGE1/_1666_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[7]),
    .ZN(\u_multiplier/pp2_7 [0]));
 AND2_X1 \u_multiplier/STAGE1/_1667_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/pp1_8 [0]));
 AND2_X1 \u_multiplier/STAGE1/_1668_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[7]),
    .ZN(\u_multiplier/pp1_8 [1]));
 AND2_X1 \u_multiplier/STAGE1/_1669_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[6]),
    .ZN(\u_multiplier/pp2_8 [7]));
 AND2_X1 \u_multiplier/STAGE1/_1670_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[5]),
    .ZN(\u_multiplier/pp2_8 [6]));
 AND2_X1 \u_multiplier/STAGE1/_1671_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[4]),
    .ZN(\u_multiplier/pp2_8 [5]));
 AND2_X1 \u_multiplier/STAGE1/_1672_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[5]),
    .ZN(\u_multiplier/pp2_8 [4]));
 AND2_X1 \u_multiplier/STAGE1/_1673_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[6]),
    .ZN(\u_multiplier/pp2_8 [3]));
 AND2_X1 \u_multiplier/STAGE1/_1674_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[7]),
    .ZN(\u_multiplier/pp2_8 [2]));
 AND2_X1 \u_multiplier/STAGE1/_1675_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/pp2_8 [1]));
 AND2_X1 \u_multiplier/STAGE1/_1676_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/pp1_9 [0]));
 AND2_X1 \u_multiplier/STAGE1/_1677_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/pp1_9 [1]));
 AND2_X1 \u_multiplier/STAGE1/_1678_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[7]),
    .ZN(\u_multiplier/pp1_9 [2]));
 AND2_X1 \u_multiplier/STAGE1/_1679_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[6]),
    .ZN(\u_multiplier/pp1_9 [3]));
 AND2_X1 \u_multiplier/STAGE1/_1680_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[5]),
    .ZN(\u_multiplier/pp2_9 [7]));
 AND2_X1 \u_multiplier/STAGE1/_1681_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[5]),
    .ZN(\u_multiplier/pp2_9 [6]));
 AND2_X1 \u_multiplier/STAGE1/_1682_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[6]),
    .ZN(\u_multiplier/pp2_9 [5]));
 AND2_X1 \u_multiplier/STAGE1/_1683_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[7]),
    .ZN(\u_multiplier/pp2_9 [4]));
 AND2_X1 \u_multiplier/STAGE1/_1684_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/pp2_9 [3]));
 AND2_X1 \u_multiplier/STAGE1/_1685_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/pp2_9 [2]));
 AND2_X1 \u_multiplier/STAGE1/_1686_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/pp1_10 [0]));
 AND2_X1 \u_multiplier/STAGE1/_1687_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/pp1_10 [1]));
 AND2_X1 \u_multiplier/STAGE1/_1688_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/pp1_10 [2]));
 AND2_X1 \u_multiplier/STAGE1/_1689_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[7]),
    .ZN(\u_multiplier/pp1_10 [3]));
 AND2_X1 \u_multiplier/STAGE1/_1690_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[6]),
    .ZN(\u_multiplier/pp1_10 [4]));
 AND2_X1 \u_multiplier/STAGE1/_1691_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[5]),
    .ZN(\u_multiplier/pp1_10 [5]));
 AND2_X1 \u_multiplier/STAGE1/_1692_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[6]),
    .ZN(\u_multiplier/pp2_10 [7]));
 AND2_X1 \u_multiplier/STAGE1/_1693_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[7]),
    .ZN(\u_multiplier/pp2_10 [6]));
 AND2_X1 \u_multiplier/STAGE1/_1694_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/pp2_10 [5]));
 AND2_X1 \u_multiplier/STAGE1/_1695_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/pp2_10 [4]));
 AND2_X1 \u_multiplier/STAGE1/_1696_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/pp2_10 [3]));
 AND2_X1 \u_multiplier/STAGE1/_1697_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/pp1_11 [0]));
 AND2_X1 \u_multiplier/STAGE1/_1698_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/pp1_11 [1]));
 AND2_X1 \u_multiplier/STAGE1/_1699_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/pp1_11 [2]));
 AND2_X1 \u_multiplier/STAGE1/_1700_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/pp1_11 [3]));
 AND2_X1 \u_multiplier/STAGE1/_1701_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[7]),
    .ZN(\u_multiplier/pp1_11 [4]));
 AND2_X1 \u_multiplier/STAGE1/_1702_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[6]),
    .ZN(\u_multiplier/pp1_11 [5]));
 AND2_X1 \u_multiplier/STAGE1/_1703_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[6]),
    .ZN(\u_multiplier/pp1_11 [6]));
 AND2_X1 \u_multiplier/STAGE1/_1704_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[7]),
    .ZN(\u_multiplier/pp1_11 [7]));
 AND2_X1 \u_multiplier/STAGE1/_1705_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/pp2_11 [7]));
 AND2_X1 \u_multiplier/STAGE1/_1706_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/pp2_11 [6]));
 AND2_X1 \u_multiplier/STAGE1/_1707_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/pp2_11 [5]));
 AND2_X1 \u_multiplier/STAGE1/_1708_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/pp2_11 [4]));
 AND2_X1 \u_multiplier/STAGE1/_1709_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/pp1_12 [0]));
 AND2_X1 \u_multiplier/STAGE1/_1710_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/pp1_12 [1]));
 AND2_X1 \u_multiplier/STAGE1/_1711_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/pp1_12 [2]));
 AND2_X1 \u_multiplier/STAGE1/_1712_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/pp1_12 [3]));
 AND2_X1 \u_multiplier/STAGE1/_1713_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/pp1_12 [4]));
 AND2_X1 \u_multiplier/STAGE1/_1714_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[7]),
    .ZN(\u_multiplier/pp1_12 [5]));
 AND2_X1 \u_multiplier/STAGE1/_1715_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[6]),
    .ZN(\u_multiplier/pp1_12 [6]));
 AND2_X1 \u_multiplier/STAGE1/_1716_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[7]),
    .ZN(\u_multiplier/pp1_12 [7]));
 AND2_X1 \u_multiplier/STAGE1/_1717_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/pp1_12 [8]));
 AND2_X1 \u_multiplier/STAGE1/_1718_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/pp1_12 [9]));
 AND2_X1 \u_multiplier/STAGE1/_1719_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/pp2_12 [7]));
 AND2_X1 \u_multiplier/STAGE1/_1720_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/pp2_12 [6]));
 AND2_X1 \u_multiplier/STAGE1/_1721_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/pp2_12 [5]));
 AND2_X1 \u_multiplier/STAGE1/_1722_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/pp1_13 [0]));
 AND2_X1 \u_multiplier/STAGE1/_1723_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/pp1_13 [1]));
 AND2_X1 \u_multiplier/STAGE1/_1724_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/pp1_13 [2]));
 AND2_X1 \u_multiplier/STAGE1/_1725_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/pp1_13 [3]));
 AND2_X1 \u_multiplier/STAGE1/_1726_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/pp1_13 [4]));
 AND2_X1 \u_multiplier/STAGE1/_1727_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/pp1_13 [5]));
 AND2_X1 \u_multiplier/STAGE1/_1728_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[7]),
    .ZN(\u_multiplier/pp1_13 [6]));
 AND2_X1 \u_multiplier/STAGE1/_1729_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[7]),
    .ZN(\u_multiplier/pp1_13 [7]));
 AND2_X1 \u_multiplier/STAGE1/_1730_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/pp1_13 [8]));
 AND2_X1 \u_multiplier/STAGE1/_1731_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/pp1_13 [9]));
 AND2_X1 \u_multiplier/STAGE1/_1732_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/pp1_13 [10]));
 AND2_X1 \u_multiplier/STAGE1/_1733_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/pp1_13 [11]));
 AND2_X1 \u_multiplier/STAGE1/_1734_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/pp2_13 [7]));
 AND2_X1 \u_multiplier/STAGE1/_1735_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/pp2_13 [6]));
 AND2_X1 \u_multiplier/STAGE1/_1736_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/pp1_14 [0]));
 AND2_X1 \u_multiplier/STAGE1/_1737_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/pp1_14 [1]));
 AND2_X1 \u_multiplier/STAGE1/_1738_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/pp1_14 [2]));
 AND2_X1 \u_multiplier/STAGE1/_1739_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/pp1_14 [3]));
 AND2_X1 \u_multiplier/STAGE1/_1740_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/pp1_14 [4]));
 AND2_X1 \u_multiplier/STAGE1/_1741_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/pp1_14 [5]));
 AND2_X1 \u_multiplier/STAGE1/_1742_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/pp1_14 [6]));
 AND2_X1 \u_multiplier/STAGE1/_1743_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[7]),
    .ZN(\u_multiplier/pp1_14 [7]));
 AND2_X1 \u_multiplier/STAGE1/_1744_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/pp1_14 [8]));
 AND2_X1 \u_multiplier/STAGE1/_1745_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/pp1_14 [9]));
 AND2_X1 \u_multiplier/STAGE1/_1746_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/pp1_14 [10]));
 AND2_X1 \u_multiplier/STAGE1/_1747_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/pp1_14 [11]));
 AND2_X1 \u_multiplier/STAGE1/_1748_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/pp1_14 [12]));
 AND2_X1 \u_multiplier/STAGE1/_1749_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/pp1_14 [13]));
 AND2_X1 \u_multiplier/STAGE1/_1750_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/pp2_14 [7]));
 AND2_X1 \u_multiplier/STAGE1/_1751_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/pp1_15 [0]));
 AND2_X1 \u_multiplier/STAGE1/_1752_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/pp1_15 [1]));
 AND2_X1 \u_multiplier/STAGE1/_1753_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/pp1_15 [2]));
 AND2_X1 \u_multiplier/STAGE1/_1754_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/pp1_15 [3]));
 AND2_X1 \u_multiplier/STAGE1/_1755_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/pp1_15 [4]));
 AND2_X1 \u_multiplier/STAGE1/_1756_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/pp1_15 [5]));
 AND2_X1 \u_multiplier/STAGE1/_1757_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/pp1_15 [6]));
 AND2_X1 \u_multiplier/STAGE1/_1758_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[8]),
    .ZN(\u_multiplier/pp1_15 [7]));
 AND2_X1 \u_multiplier/STAGE1/_1759_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/pp1_15 [8]));
 AND2_X1 \u_multiplier/STAGE1/_1760_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/pp1_15 [9]));
 AND2_X1 \u_multiplier/STAGE1/_1761_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/pp1_15 [10]));
 AND2_X1 \u_multiplier/STAGE1/_1762_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/pp1_15 [11]));
 AND2_X1 \u_multiplier/STAGE1/_1763_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/pp1_15 [12]));
 AND2_X1 \u_multiplier/STAGE1/_1764_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/pp1_15 [13]));
 AND2_X1 \u_multiplier/STAGE1/_1765_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/pp1_15 [14]));
 AND2_X1 \u_multiplier/STAGE1/_1766_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/pp1_15 [15]));
 AND2_X1 \u_multiplier/STAGE1/_1767_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[16]),
    .ZN(\u_multiplier/STAGE1/_0607_ ));
 AND2_X1 \u_multiplier/STAGE1/_1768_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/STAGE1/_0608_ ));
 AND2_X1 \u_multiplier/STAGE1/_1769_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[16]),
    .ZN(\u_multiplier/pp1_16 [1]));
 AND2_X1 \u_multiplier/STAGE1/_1770_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/pp1_16 [2]));
 AND2_X1 \u_multiplier/STAGE1/_1771_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/pp1_16 [3]));
 AND2_X1 \u_multiplier/STAGE1/_1772_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/pp1_16 [4]));
 AND2_X1 \u_multiplier/STAGE1/_1773_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/pp1_16 [5]));
 AND2_X1 \u_multiplier/STAGE1/_1774_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/pp1_16 [6]));
 AND2_X1 \u_multiplier/STAGE1/_1775_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/pp1_16 [7]));
 AND2_X1 \u_multiplier/STAGE1/_1776_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/pp1_16 [8]));
 AND2_X1 \u_multiplier/STAGE1/_1777_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[8]),
    .ZN(\u_multiplier/pp1_16 [9]));
 AND2_X1 \u_multiplier/STAGE1/_1778_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/pp1_16 [10]));
 AND2_X1 \u_multiplier/STAGE1/_1779_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/pp1_16 [11]));
 AND2_X1 \u_multiplier/STAGE1/_1780_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/pp1_16 [12]));
 AND2_X1 \u_multiplier/STAGE1/_1781_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/pp1_16 [13]));
 AND2_X1 \u_multiplier/STAGE1/_1782_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/pp1_16 [14]));
 AND2_X1 \u_multiplier/STAGE1/_1783_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/pp1_16 [15]));
 AND2_X1 \u_multiplier/STAGE1/_1784_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0609_ ));
 AND2_X1 \u_multiplier/STAGE1/_1785_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[16]),
    .ZN(\u_multiplier/STAGE1/_0610_ ));
 AND2_X1 \u_multiplier/STAGE1/_1786_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/STAGE1/_0611_ ));
 AND2_X1 \u_multiplier/STAGE1/_1787_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/STAGE1/_0612_ ));
 AND2_X1 \u_multiplier/STAGE1/_1788_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[17]),
    .ZN(\u_multiplier/pp1_17 [2]));
 AND2_X1 \u_multiplier/STAGE1/_1789_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[16]),
    .ZN(\u_multiplier/pp1_17 [3]));
 AND2_X1 \u_multiplier/STAGE1/_1790_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/pp1_17 [4]));
 AND2_X1 \u_multiplier/STAGE1/_1791_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/pp1_17 [5]));
 AND2_X1 \u_multiplier/STAGE1/_1792_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/pp1_17 [6]));
 AND2_X1 \u_multiplier/STAGE1/_1793_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/pp1_17 [7]));
 AND2_X1 \u_multiplier/STAGE1/_1794_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/pp1_17 [8]));
 AND2_X1 \u_multiplier/STAGE1/_1795_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/pp1_17 [9]));
 AND2_X1 \u_multiplier/STAGE1/_1796_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[9]),
    .ZN(\u_multiplier/pp1_17 [10]));
 AND2_X1 \u_multiplier/STAGE1/_1797_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/pp1_17 [11]));
 AND2_X1 \u_multiplier/STAGE1/_1798_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/pp1_17 [12]));
 AND2_X1 \u_multiplier/STAGE1/_1799_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/pp1_17 [13]));
 AND2_X1 \u_multiplier/STAGE1/_1800_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/pp1_17 [14]));
 AND2_X1 \u_multiplier/STAGE1/_1801_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/pp1_17 [15]));
 AND2_X1 \u_multiplier/STAGE1/_1802_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0613_ ));
 AND2_X1 \u_multiplier/STAGE1/_1803_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0614_ ));
 AND2_X1 \u_multiplier/STAGE1/_1804_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[16]),
    .ZN(\u_multiplier/STAGE1/_0615_ ));
 AND2_X1 \u_multiplier/STAGE1/_1805_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/STAGE1/_0616_ ));
 AND2_X1 \u_multiplier/STAGE1/_1806_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/STAGE1/_0617_ ));
 AND2_X1 \u_multiplier/STAGE1/_1807_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/STAGE1/_0618_ ));
 AND2_X1 \u_multiplier/STAGE1/_1808_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[18]),
    .ZN(\u_multiplier/pp1_18 [3]));
 AND2_X1 \u_multiplier/STAGE1/_1809_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[17]),
    .ZN(\u_multiplier/pp1_18 [4]));
 AND2_X1 \u_multiplier/STAGE1/_1810_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[16]),
    .ZN(\u_multiplier/pp1_18 [5]));
 AND2_X1 \u_multiplier/STAGE1/_1811_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/pp1_18 [6]));
 AND2_X1 \u_multiplier/STAGE1/_1812_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/pp1_18 [7]));
 AND2_X1 \u_multiplier/STAGE1/_1813_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/pp1_18 [8]));
 AND2_X1 \u_multiplier/STAGE1/_1814_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/pp1_18 [9]));
 AND2_X1 \u_multiplier/STAGE1/_1815_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/pp1_18 [10]));
 AND2_X1 \u_multiplier/STAGE1/_1816_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/pp1_18 [11]));
 AND2_X1 \u_multiplier/STAGE1/_1817_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[9]),
    .ZN(\u_multiplier/pp1_18 [12]));
 AND2_X1 \u_multiplier/STAGE1/_1818_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/pp1_18 [13]));
 AND2_X1 \u_multiplier/STAGE1/_1819_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/pp1_18 [14]));
 AND2_X1 \u_multiplier/STAGE1/_1820_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/pp1_18 [15]));
 AND2_X1 \u_multiplier/STAGE1/_1821_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0619_ ));
 AND2_X1 \u_multiplier/STAGE1/_1822_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0620_ ));
 AND2_X1 \u_multiplier/STAGE1/_1823_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0621_ ));
 AND2_X1 \u_multiplier/STAGE1/_1824_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[16]),
    .ZN(\u_multiplier/STAGE1/_0622_ ));
 AND2_X1 \u_multiplier/STAGE1/_1825_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/STAGE1/_0623_ ));
 AND2_X1 \u_multiplier/STAGE1/_1826_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/STAGE1/_0624_ ));
 AND2_X1 \u_multiplier/STAGE1/_1827_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/STAGE1/_0625_ ));
 AND2_X1 \u_multiplier/STAGE1/_1828_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/STAGE1/_0626_ ));
 AND2_X1 \u_multiplier/STAGE1/_1829_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[19]),
    .ZN(\u_multiplier/pp1_19 [4]));
 AND2_X1 \u_multiplier/STAGE1/_1830_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[18]),
    .ZN(\u_multiplier/pp1_19 [5]));
 AND2_X1 \u_multiplier/STAGE1/_1831_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[17]),
    .ZN(\u_multiplier/pp1_19 [6]));
 AND2_X1 \u_multiplier/STAGE1/_1832_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[16]),
    .ZN(\u_multiplier/pp1_19 [7]));
 AND2_X1 \u_multiplier/STAGE1/_1833_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/pp1_19 [8]));
 AND2_X1 \u_multiplier/STAGE1/_1834_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/pp1_19 [9]));
 AND2_X1 \u_multiplier/STAGE1/_1835_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/pp1_19 [10]));
 AND2_X1 \u_multiplier/STAGE1/_1836_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/pp1_19 [11]));
 AND2_X1 \u_multiplier/STAGE1/_1837_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/pp1_19 [12]));
 AND2_X1 \u_multiplier/STAGE1/_1838_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[10]),
    .ZN(\u_multiplier/pp1_19 [13]));
 AND2_X1 \u_multiplier/STAGE1/_1839_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/pp1_19 [14]));
 AND2_X1 \u_multiplier/STAGE1/_1840_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/pp1_19 [15]));
 AND2_X1 \u_multiplier/STAGE1/_1841_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[20]),
    .ZN(\u_multiplier/STAGE1/_0627_ ));
 AND2_X1 \u_multiplier/STAGE1/_1842_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0628_ ));
 AND2_X1 \u_multiplier/STAGE1/_1843_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0629_ ));
 AND2_X1 \u_multiplier/STAGE1/_1844_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0630_ ));
 AND2_X1 \u_multiplier/STAGE1/_1845_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[16]),
    .ZN(\u_multiplier/STAGE1/_0631_ ));
 AND2_X1 \u_multiplier/STAGE1/_1846_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/STAGE1/_0632_ ));
 AND2_X1 \u_multiplier/STAGE1/_1847_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/STAGE1/_0633_ ));
 AND2_X1 \u_multiplier/STAGE1/_1848_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/STAGE1/_0634_ ));
 AND2_X1 \u_multiplier/STAGE1/_1849_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/STAGE1/_0635_ ));
 AND2_X1 \u_multiplier/STAGE1/_1850_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/STAGE1/_0636_ ));
 AND2_X1 \u_multiplier/STAGE1/_1851_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[20]),
    .ZN(\u_multiplier/pp1_20 [5]));
 AND2_X1 \u_multiplier/STAGE1/_1852_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[19]),
    .ZN(\u_multiplier/pp1_20 [6]));
 AND2_X1 \u_multiplier/STAGE1/_1853_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[18]),
    .ZN(\u_multiplier/pp1_20 [7]));
 AND2_X1 \u_multiplier/STAGE1/_1854_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[17]),
    .ZN(\u_multiplier/pp1_20 [8]));
 AND2_X1 \u_multiplier/STAGE1/_1855_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[16]),
    .ZN(\u_multiplier/pp1_20 [9]));
 AND2_X1 \u_multiplier/STAGE1/_1856_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/pp1_20 [10]));
 AND2_X1 \u_multiplier/STAGE1/_1857_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/pp1_20 [11]));
 AND2_X1 \u_multiplier/STAGE1/_1858_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/pp1_20 [12]));
 AND2_X1 \u_multiplier/STAGE1/_1859_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/pp1_20 [13]));
 AND2_X1 \u_multiplier/STAGE1/_1860_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/pp1_20 [14]));
 AND2_X1 \u_multiplier/STAGE1/_1861_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[10]),
    .ZN(\u_multiplier/pp1_20 [15]));
 AND2_X1 \u_multiplier/STAGE1/_1862_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[21]),
    .ZN(\u_multiplier/STAGE1/_0637_ ));
 AND2_X1 \u_multiplier/STAGE1/_1863_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[20]),
    .ZN(\u_multiplier/STAGE1/_0638_ ));
 AND2_X1 \u_multiplier/STAGE1/_1864_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0639_ ));
 AND2_X1 \u_multiplier/STAGE1/_1865_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0640_ ));
 AND2_X1 \u_multiplier/STAGE1/_1866_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0641_ ));
 AND2_X1 \u_multiplier/STAGE1/_1867_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[16]),
    .ZN(\u_multiplier/STAGE1/_0642_ ));
 AND2_X1 \u_multiplier/STAGE1/_1868_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/STAGE1/_0643_ ));
 AND2_X1 \u_multiplier/STAGE1/_1869_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/STAGE1/_0644_ ));
 AND2_X1 \u_multiplier/STAGE1/_1870_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/STAGE1/_0645_ ));
 AND2_X1 \u_multiplier/STAGE1/_1871_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/STAGE1/_0646_ ));
 AND2_X1 \u_multiplier/STAGE1/_1872_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/STAGE1/_0647_ ));
 AND2_X1 \u_multiplier/STAGE1/_1873_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[11]),
    .ZN(\u_multiplier/STAGE1/_0648_ ));
 AND2_X1 \u_multiplier/STAGE1/_1874_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[21]),
    .ZN(\u_multiplier/pp1_21 [6]));
 AND2_X1 \u_multiplier/STAGE1/_1875_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[20]),
    .ZN(\u_multiplier/pp1_21 [7]));
 AND2_X1 \u_multiplier/STAGE1/_1876_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[19]),
    .ZN(\u_multiplier/pp1_21 [8]));
 AND2_X1 \u_multiplier/STAGE1/_1877_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[18]),
    .ZN(\u_multiplier/pp1_21 [9]));
 AND2_X1 \u_multiplier/STAGE1/_1878_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[17]),
    .ZN(\u_multiplier/pp1_21 [10]));
 AND2_X1 \u_multiplier/STAGE1/_1879_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[16]),
    .ZN(\u_multiplier/pp1_21 [11]));
 AND2_X1 \u_multiplier/STAGE1/_1880_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/pp1_21 [12]));
 AND2_X1 \u_multiplier/STAGE1/_1881_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/pp1_21 [13]));
 AND2_X1 \u_multiplier/STAGE1/_1882_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/pp1_21 [14]));
 AND2_X1 \u_multiplier/STAGE1/_1883_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/pp1_21 [15]));
 AND2_X1 \u_multiplier/STAGE1/_1884_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[22]),
    .ZN(\u_multiplier/STAGE1/_0649_ ));
 AND2_X1 \u_multiplier/STAGE1/_1885_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[21]),
    .ZN(\u_multiplier/STAGE1/_0650_ ));
 AND2_X1 \u_multiplier/STAGE1/_1886_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[20]),
    .ZN(\u_multiplier/STAGE1/_0651_ ));
 AND2_X1 \u_multiplier/STAGE1/_1887_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0652_ ));
 AND2_X1 \u_multiplier/STAGE1/_1888_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0653_ ));
 AND2_X1 \u_multiplier/STAGE1/_1889_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0654_ ));
 AND2_X1 \u_multiplier/STAGE1/_1890_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[16]),
    .ZN(\u_multiplier/STAGE1/_0655_ ));
 AND2_X1 \u_multiplier/STAGE1/_1891_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/STAGE1/_0656_ ));
 AND2_X1 \u_multiplier/STAGE1/_1892_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/STAGE1/_0657_ ));
 AND2_X1 \u_multiplier/STAGE1/_1893_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/STAGE1/_0658_ ));
 AND2_X1 \u_multiplier/STAGE1/_1894_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/STAGE1/_0659_ ));
 AND2_X1 \u_multiplier/STAGE1/_1895_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[11]),
    .ZN(\u_multiplier/STAGE1/_0660_ ));
 AND2_X1 \u_multiplier/STAGE1/_1896_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/STAGE1/_0661_ ));
 AND2_X1 \u_multiplier/STAGE1/_1897_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/STAGE1/_0662_ ));
 AND2_X1 \u_multiplier/STAGE1/_1898_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[22]),
    .ZN(\u_multiplier/pp1_22 [7]));
 AND2_X1 \u_multiplier/STAGE1/_1899_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[21]),
    .ZN(\u_multiplier/pp1_22 [8]));
 AND2_X1 \u_multiplier/STAGE1/_1900_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[20]),
    .ZN(\u_multiplier/pp1_22 [9]));
 AND2_X1 \u_multiplier/STAGE1/_1901_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[19]),
    .ZN(\u_multiplier/pp1_22 [10]));
 AND2_X1 \u_multiplier/STAGE1/_1902_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[18]),
    .ZN(\u_multiplier/pp1_22 [11]));
 AND2_X1 \u_multiplier/STAGE1/_1903_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[17]),
    .ZN(\u_multiplier/pp1_22 [12]));
 AND2_X1 \u_multiplier/STAGE1/_1904_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[16]),
    .ZN(\u_multiplier/pp1_22 [13]));
 AND2_X1 \u_multiplier/STAGE1/_1905_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/pp1_22 [14]));
 AND2_X1 \u_multiplier/STAGE1/_1906_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/pp1_22 [15]));
 AND2_X1 \u_multiplier/STAGE1/_1907_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[23]),
    .ZN(\u_multiplier/STAGE1/_0663_ ));
 AND2_X1 \u_multiplier/STAGE1/_1908_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[22]),
    .ZN(\u_multiplier/STAGE1/_0664_ ));
 AND2_X1 \u_multiplier/STAGE1/_1909_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[21]),
    .ZN(\u_multiplier/STAGE1/_0665_ ));
 AND2_X1 \u_multiplier/STAGE1/_1910_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[20]),
    .ZN(\u_multiplier/STAGE1/_0666_ ));
 AND2_X1 \u_multiplier/STAGE1/_1911_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0667_ ));
 AND2_X1 \u_multiplier/STAGE1/_1912_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0668_ ));
 AND2_X1 \u_multiplier/STAGE1/_1913_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0669_ ));
 AND2_X1 \u_multiplier/STAGE1/_1914_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[16]),
    .ZN(\u_multiplier/STAGE1/_0670_ ));
 AND2_X1 \u_multiplier/STAGE1/_1915_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/STAGE1/_0671_ ));
 AND2_X1 \u_multiplier/STAGE1/_1916_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/STAGE1/_0672_ ));
 AND2_X1 \u_multiplier/STAGE1/_1917_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/STAGE1/_0673_ ));
 AND2_X1 \u_multiplier/STAGE1/_1918_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/STAGE1/_0674_ ));
 AND2_X1 \u_multiplier/STAGE1/_1919_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[12]),
    .ZN(\u_multiplier/STAGE1/_0675_ ));
 AND2_X1 \u_multiplier/STAGE1/_1920_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/STAGE1/_0676_ ));
 AND2_X1 \u_multiplier/STAGE1/_1921_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/STAGE1/_0677_ ));
 AND2_X1 \u_multiplier/STAGE1/_1922_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/STAGE1/_0678_ ));
 AND2_X1 \u_multiplier/STAGE1/_1923_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[23]),
    .ZN(\u_multiplier/pp1_23 [8]));
 AND2_X1 \u_multiplier/STAGE1/_1924_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[22]),
    .ZN(\u_multiplier/pp1_23 [9]));
 AND2_X1 \u_multiplier/STAGE1/_1925_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[21]),
    .ZN(\u_multiplier/pp1_23 [10]));
 AND2_X1 \u_multiplier/STAGE1/_1926_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[20]),
    .ZN(\u_multiplier/pp1_23 [11]));
 AND2_X1 \u_multiplier/STAGE1/_1927_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[19]),
    .ZN(\u_multiplier/pp1_23 [12]));
 AND2_X1 \u_multiplier/STAGE1/_1928_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[18]),
    .ZN(\u_multiplier/pp1_23 [13]));
 AND2_X1 \u_multiplier/STAGE1/_1929_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[17]),
    .ZN(\u_multiplier/pp1_23 [14]));
 AND2_X1 \u_multiplier/STAGE1/_1930_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[16]),
    .ZN(\u_multiplier/pp1_23 [15]));
 AND2_X1 \u_multiplier/STAGE1/_1931_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[24]),
    .ZN(\u_multiplier/STAGE1/_0679_ ));
 AND2_X1 \u_multiplier/STAGE1/_1932_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[23]),
    .ZN(\u_multiplier/STAGE1/_0680_ ));
 AND2_X1 \u_multiplier/STAGE1/_1933_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[22]),
    .ZN(\u_multiplier/STAGE1/_0681_ ));
 AND2_X1 \u_multiplier/STAGE1/_1934_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[21]),
    .ZN(\u_multiplier/STAGE1/_0682_ ));
 AND2_X1 \u_multiplier/STAGE1/_1935_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[20]),
    .ZN(\u_multiplier/STAGE1/_0683_ ));
 AND2_X1 \u_multiplier/STAGE1/_1936_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0684_ ));
 AND2_X1 \u_multiplier/STAGE1/_1937_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0685_ ));
 AND2_X1 \u_multiplier/STAGE1/_1938_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0686_ ));
 AND2_X1 \u_multiplier/STAGE1/_1939_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[16]),
    .ZN(\u_multiplier/STAGE1/_0687_ ));
 AND2_X1 \u_multiplier/STAGE1/_1940_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/STAGE1/_0688_ ));
 AND2_X1 \u_multiplier/STAGE1/_1941_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/STAGE1/_0689_ ));
 AND2_X1 \u_multiplier/STAGE1/_1942_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/STAGE1/_0690_ ));
 AND2_X1 \u_multiplier/STAGE1/_1943_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[12]),
    .ZN(\u_multiplier/STAGE1/_0691_ ));
 AND2_X1 \u_multiplier/STAGE1/_1944_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/STAGE1/_0692_ ));
 AND2_X1 \u_multiplier/STAGE1/_1945_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/STAGE1/_0693_ ));
 AND2_X1 \u_multiplier/STAGE1/_1946_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/STAGE1/_0694_ ));
 AND2_X1 \u_multiplier/STAGE1/_1947_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[16]),
    .ZN(\u_multiplier/STAGE1/_0695_ ));
 AND2_X1 \u_multiplier/STAGE1/_1948_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0696_ ));
 AND2_X1 \u_multiplier/STAGE1/_1949_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[24]),
    .ZN(\u_multiplier/pp1_24 [9]));
 AND2_X1 \u_multiplier/STAGE1/_1950_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[23]),
    .ZN(\u_multiplier/pp1_24 [10]));
 AND2_X1 \u_multiplier/STAGE1/_1951_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[22]),
    .ZN(\u_multiplier/pp1_24 [11]));
 AND2_X1 \u_multiplier/STAGE1/_1952_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[21]),
    .ZN(\u_multiplier/pp1_24 [12]));
 AND2_X1 \u_multiplier/STAGE1/_1953_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[20]),
    .ZN(\u_multiplier/pp1_24 [13]));
 AND2_X1 \u_multiplier/STAGE1/_1954_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[19]),
    .ZN(\u_multiplier/pp1_24 [14]));
 AND2_X1 \u_multiplier/STAGE1/_1955_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[18]),
    .ZN(\u_multiplier/pp1_24 [15]));
 AND2_X1 \u_multiplier/STAGE1/_1956_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[25]),
    .ZN(\u_multiplier/STAGE1/_0697_ ));
 AND2_X1 \u_multiplier/STAGE1/_1957_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[24]),
    .ZN(\u_multiplier/STAGE1/_0698_ ));
 AND2_X1 \u_multiplier/STAGE1/_1958_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[23]),
    .ZN(\u_multiplier/STAGE1/_0699_ ));
 AND2_X1 \u_multiplier/STAGE1/_1959_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[22]),
    .ZN(\u_multiplier/STAGE1/_0700_ ));
 AND2_X1 \u_multiplier/STAGE1/_1960_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[21]),
    .ZN(\u_multiplier/STAGE1/_0701_ ));
 AND2_X1 \u_multiplier/STAGE1/_1961_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[20]),
    .ZN(\u_multiplier/STAGE1/_0702_ ));
 AND2_X1 \u_multiplier/STAGE1/_1962_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0703_ ));
 AND2_X1 \u_multiplier/STAGE1/_1963_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0704_ ));
 AND2_X1 \u_multiplier/STAGE1/_1964_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0705_ ));
 AND2_X1 \u_multiplier/STAGE1/_1965_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[16]),
    .ZN(\u_multiplier/STAGE1/_0706_ ));
 AND2_X1 \u_multiplier/STAGE1/_1966_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/STAGE1/_0707_ ));
 AND2_X1 \u_multiplier/STAGE1/_1967_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/STAGE1/_0708_ ));
 AND2_X1 \u_multiplier/STAGE1/_1968_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/STAGE1/_0709_ ));
 AND2_X1 \u_multiplier/STAGE1/_1969_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[13]),
    .ZN(\u_multiplier/STAGE1/_0710_ ));
 AND2_X1 \u_multiplier/STAGE1/_1970_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/STAGE1/_0711_ ));
 AND2_X1 \u_multiplier/STAGE1/_1971_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/STAGE1/_0712_ ));
 AND2_X1 \u_multiplier/STAGE1/_1972_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[16]),
    .ZN(\u_multiplier/STAGE1/_0713_ ));
 AND2_X1 \u_multiplier/STAGE1/_1973_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0714_ ));
 AND2_X1 \u_multiplier/STAGE1/_1974_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0715_ ));
 AND2_X1 \u_multiplier/STAGE1/_1975_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0716_ ));
 AND2_X1 \u_multiplier/STAGE1/_1976_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[25]),
    .ZN(\u_multiplier/pp1_25 [10]));
 AND2_X1 \u_multiplier/STAGE1/_1977_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[24]),
    .ZN(\u_multiplier/pp1_25 [11]));
 AND2_X1 \u_multiplier/STAGE1/_1978_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[23]),
    .ZN(\u_multiplier/pp1_25 [12]));
 AND2_X1 \u_multiplier/STAGE1/_1979_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[22]),
    .ZN(\u_multiplier/pp1_25 [13]));
 AND2_X1 \u_multiplier/STAGE1/_1980_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[21]),
    .ZN(\u_multiplier/pp1_25 [14]));
 AND2_X1 \u_multiplier/STAGE1/_1981_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[20]),
    .ZN(\u_multiplier/pp1_25 [15]));
 AND2_X1 \u_multiplier/STAGE1/_1982_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[26]),
    .ZN(\u_multiplier/STAGE1/_0717_ ));
 AND2_X1 \u_multiplier/STAGE1/_1983_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[25]),
    .ZN(\u_multiplier/STAGE1/_0718_ ));
 AND2_X1 \u_multiplier/STAGE1/_1984_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[24]),
    .ZN(\u_multiplier/STAGE1/_0719_ ));
 AND2_X1 \u_multiplier/STAGE1/_1985_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[23]),
    .ZN(\u_multiplier/STAGE1/_0720_ ));
 AND2_X1 \u_multiplier/STAGE1/_1986_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[22]),
    .ZN(\u_multiplier/STAGE1/_0721_ ));
 AND2_X1 \u_multiplier/STAGE1/_1987_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[21]),
    .ZN(\u_multiplier/STAGE1/_0722_ ));
 AND2_X1 \u_multiplier/STAGE1/_1988_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[20]),
    .ZN(\u_multiplier/STAGE1/_0723_ ));
 AND2_X1 \u_multiplier/STAGE1/_1989_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0724_ ));
 AND2_X1 \u_multiplier/STAGE1/_1990_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0725_ ));
 AND2_X1 \u_multiplier/STAGE1/_1991_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0726_ ));
 AND2_X1 \u_multiplier/STAGE1/_1992_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[16]),
    .ZN(\u_multiplier/STAGE1/_0727_ ));
 AND2_X1 \u_multiplier/STAGE1/_1993_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/STAGE1/_0728_ ));
 AND2_X1 \u_multiplier/STAGE1/_1994_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/STAGE1/_0729_ ));
 AND2_X1 \u_multiplier/STAGE1/_1995_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[13]),
    .ZN(\u_multiplier/STAGE1/_0730_ ));
 AND2_X1 \u_multiplier/STAGE1/_1996_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/STAGE1/_0731_ ));
 AND2_X1 \u_multiplier/STAGE1/_1997_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/STAGE1/_0732_ ));
 AND2_X1 \u_multiplier/STAGE1/_1998_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[16]),
    .ZN(\u_multiplier/STAGE1/_0733_ ));
 AND2_X1 \u_multiplier/STAGE1/_1999_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0734_ ));
 AND2_X1 \u_multiplier/STAGE1/_2000_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0735_ ));
 AND2_X1 \u_multiplier/STAGE1/_2001_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0736_ ));
 AND2_X1 \u_multiplier/STAGE1/_2002_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[20]),
    .ZN(\u_multiplier/STAGE1/_0737_ ));
 AND2_X1 \u_multiplier/STAGE1/_2003_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[21]),
    .ZN(\u_multiplier/STAGE1/_0738_ ));
 AND2_X1 \u_multiplier/STAGE1/_2004_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[26]),
    .ZN(\u_multiplier/pp1_26 [11]));
 AND2_X1 \u_multiplier/STAGE1/_2005_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[25]),
    .ZN(\u_multiplier/pp1_26 [12]));
 AND2_X1 \u_multiplier/STAGE1/_2006_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[24]),
    .ZN(\u_multiplier/pp1_26 [13]));
 AND2_X1 \u_multiplier/STAGE1/_2007_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[23]),
    .ZN(\u_multiplier/pp1_26 [14]));
 AND2_X1 \u_multiplier/STAGE1/_2008_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[22]),
    .ZN(\u_multiplier/pp1_26 [15]));
 AND2_X1 \u_multiplier/STAGE1/_2009_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[27]),
    .ZN(\u_multiplier/STAGE1/_0739_ ));
 AND2_X1 \u_multiplier/STAGE1/_2010_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[26]),
    .ZN(\u_multiplier/STAGE1/_0740_ ));
 AND2_X1 \u_multiplier/STAGE1/_2011_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[25]),
    .ZN(\u_multiplier/STAGE1/_0741_ ));
 AND2_X1 \u_multiplier/STAGE1/_2012_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[24]),
    .ZN(\u_multiplier/STAGE1/_0742_ ));
 AND2_X1 \u_multiplier/STAGE1/_2013_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[23]),
    .ZN(\u_multiplier/STAGE1/_0743_ ));
 AND2_X1 \u_multiplier/STAGE1/_2014_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[22]),
    .ZN(\u_multiplier/STAGE1/_0744_ ));
 AND2_X1 \u_multiplier/STAGE1/_2015_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[21]),
    .ZN(\u_multiplier/STAGE1/_0745_ ));
 AND2_X1 \u_multiplier/STAGE1/_2016_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[20]),
    .ZN(\u_multiplier/STAGE1/_0746_ ));
 AND2_X1 \u_multiplier/STAGE1/_2017_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0747_ ));
 AND2_X1 \u_multiplier/STAGE1/_2018_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0748_ ));
 AND2_X1 \u_multiplier/STAGE1/_2019_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0749_ ));
 AND2_X1 \u_multiplier/STAGE1/_2020_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[16]),
    .ZN(\u_multiplier/STAGE1/_0750_ ));
 AND2_X1 \u_multiplier/STAGE1/_2021_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/STAGE1/_0751_ ));
 AND2_X1 \u_multiplier/STAGE1/_2022_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/STAGE1/_0752_ ));
 AND2_X1 \u_multiplier/STAGE1/_2023_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[14]),
    .ZN(\u_multiplier/STAGE1/_0753_ ));
 AND2_X1 \u_multiplier/STAGE1/_2024_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/STAGE1/_0754_ ));
 AND2_X1 \u_multiplier/STAGE1/_2025_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[16]),
    .ZN(\u_multiplier/STAGE1/_0755_ ));
 AND2_X1 \u_multiplier/STAGE1/_2026_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0756_ ));
 AND2_X1 \u_multiplier/STAGE1/_2027_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0757_ ));
 AND2_X1 \u_multiplier/STAGE1/_2028_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0758_ ));
 AND2_X1 \u_multiplier/STAGE1/_2029_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[20]),
    .ZN(\u_multiplier/STAGE1/_0759_ ));
 AND2_X1 \u_multiplier/STAGE1/_2030_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[21]),
    .ZN(\u_multiplier/STAGE1/_0760_ ));
 AND2_X1 \u_multiplier/STAGE1/_2031_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[22]),
    .ZN(\u_multiplier/STAGE1/_0761_ ));
 AND2_X1 \u_multiplier/STAGE1/_2032_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[23]),
    .ZN(\u_multiplier/STAGE1/_0762_ ));
 AND2_X1 \u_multiplier/STAGE1/_2033_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/pp1_27 [12]));
 AND2_X1 \u_multiplier/STAGE1/_2034_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[26]),
    .ZN(\u_multiplier/pp1_27 [13]));
 AND2_X1 \u_multiplier/STAGE1/_2035_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[25]),
    .ZN(\u_multiplier/pp1_27 [14]));
 AND2_X1 \u_multiplier/STAGE1/_2036_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[24]),
    .ZN(\u_multiplier/pp1_27 [15]));
 AND2_X1 \u_multiplier/STAGE1/_2037_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/STAGE1/_0763_ ));
 AND2_X1 \u_multiplier/STAGE1/_2038_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[27]),
    .ZN(\u_multiplier/STAGE1/_0764_ ));
 AND2_X1 \u_multiplier/STAGE1/_2039_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[26]),
    .ZN(\u_multiplier/STAGE1/_0765_ ));
 AND2_X1 \u_multiplier/STAGE1/_2040_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[25]),
    .ZN(\u_multiplier/STAGE1/_0766_ ));
 AND2_X1 \u_multiplier/STAGE1/_2041_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[24]),
    .ZN(\u_multiplier/STAGE1/_0767_ ));
 AND2_X1 \u_multiplier/STAGE1/_2042_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[23]),
    .ZN(\u_multiplier/STAGE1/_0768_ ));
 AND2_X1 \u_multiplier/STAGE1/_2043_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[22]),
    .ZN(\u_multiplier/STAGE1/_0769_ ));
 AND2_X1 \u_multiplier/STAGE1/_2044_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[21]),
    .ZN(\u_multiplier/STAGE1/_0770_ ));
 AND2_X1 \u_multiplier/STAGE1/_2045_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[20]),
    .ZN(\u_multiplier/STAGE1/_0771_ ));
 AND2_X1 \u_multiplier/STAGE1/_2046_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0772_ ));
 AND2_X1 \u_multiplier/STAGE1/_2047_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0773_ ));
 AND2_X1 \u_multiplier/STAGE1/_2048_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0774_ ));
 AND2_X1 \u_multiplier/STAGE1/_2049_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[16]),
    .ZN(\u_multiplier/STAGE1/_0775_ ));
 AND2_X1 \u_multiplier/STAGE1/_2050_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/STAGE1/_0776_ ));
 AND2_X1 \u_multiplier/STAGE1/_2051_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[14]),
    .ZN(\u_multiplier/STAGE1/_0777_ ));
 AND2_X1 \u_multiplier/STAGE1/_2052_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/STAGE1/_0778_ ));
 AND2_X1 \u_multiplier/STAGE1/_2053_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[16]),
    .ZN(\u_multiplier/STAGE1/_0779_ ));
 AND2_X1 \u_multiplier/STAGE1/_2054_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0780_ ));
 AND2_X1 \u_multiplier/STAGE1/_2055_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0781_ ));
 AND2_X1 \u_multiplier/STAGE1/_2056_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0782_ ));
 AND2_X1 \u_multiplier/STAGE1/_2057_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[20]),
    .ZN(\u_multiplier/STAGE1/_0783_ ));
 AND2_X1 \u_multiplier/STAGE1/_2058_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[21]),
    .ZN(\u_multiplier/STAGE1/_0784_ ));
 AND2_X1 \u_multiplier/STAGE1/_2059_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[22]),
    .ZN(\u_multiplier/STAGE1/_0785_ ));
 AND2_X1 \u_multiplier/STAGE1/_2060_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[23]),
    .ZN(\u_multiplier/STAGE1/_0786_ ));
 AND2_X1 \u_multiplier/STAGE1/_2061_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[24]),
    .ZN(\u_multiplier/STAGE1/_0787_ ));
 AND2_X1 \u_multiplier/STAGE1/_2062_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[25]),
    .ZN(\u_multiplier/STAGE1/_0788_ ));
 AND2_X1 \u_multiplier/STAGE1/_2063_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/pp1_28 [13]));
 AND2_X1 \u_multiplier/STAGE1/_2064_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/pp1_28 [14]));
 AND2_X1 \u_multiplier/STAGE1/_2065_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[26]),
    .ZN(\u_multiplier/pp1_28 [15]));
 AND2_X1 \u_multiplier/STAGE1/_2066_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/STAGE1/_0789_ ));
 AND2_X1 \u_multiplier/STAGE1/_2067_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/STAGE1/_0790_ ));
 AND2_X1 \u_multiplier/STAGE1/_2068_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[27]),
    .ZN(\u_multiplier/STAGE1/_0791_ ));
 AND2_X1 \u_multiplier/STAGE1/_2069_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[26]),
    .ZN(\u_multiplier/STAGE1/_0792_ ));
 AND2_X1 \u_multiplier/STAGE1/_2070_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[25]),
    .ZN(\u_multiplier/STAGE1/_0793_ ));
 AND2_X1 \u_multiplier/STAGE1/_2071_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[24]),
    .ZN(\u_multiplier/STAGE1/_0794_ ));
 AND2_X1 \u_multiplier/STAGE1/_2072_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[23]),
    .ZN(\u_multiplier/STAGE1/_0795_ ));
 AND2_X1 \u_multiplier/STAGE1/_2073_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[22]),
    .ZN(\u_multiplier/STAGE1/_0796_ ));
 AND2_X1 \u_multiplier/STAGE1/_2074_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[21]),
    .ZN(\u_multiplier/STAGE1/_0797_ ));
 AND2_X1 \u_multiplier/STAGE1/_2075_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[20]),
    .ZN(\u_multiplier/STAGE1/_0798_ ));
 AND2_X1 \u_multiplier/STAGE1/_2076_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0799_ ));
 AND2_X1 \u_multiplier/STAGE1/_2077_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0800_ ));
 AND2_X1 \u_multiplier/STAGE1/_2078_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0801_ ));
 AND2_X1 \u_multiplier/STAGE1/_2079_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[16]),
    .ZN(\u_multiplier/STAGE1/_0802_ ));
 AND2_X1 \u_multiplier/STAGE1/_2080_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/STAGE1/_0803_ ));
 AND2_X1 \u_multiplier/STAGE1/_2081_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[15]),
    .ZN(\u_multiplier/STAGE1/_0804_ ));
 AND2_X1 \u_multiplier/STAGE1/_2082_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[16]),
    .ZN(\u_multiplier/STAGE1/_0805_ ));
 AND2_X1 \u_multiplier/STAGE1/_2083_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0806_ ));
 AND2_X1 \u_multiplier/STAGE1/_2084_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0807_ ));
 AND2_X1 \u_multiplier/STAGE1/_2085_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0808_ ));
 AND2_X1 \u_multiplier/STAGE1/_2086_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[20]),
    .ZN(\u_multiplier/STAGE1/_0809_ ));
 AND2_X1 \u_multiplier/STAGE1/_2087_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[21]),
    .ZN(\u_multiplier/STAGE1/_0810_ ));
 AND2_X1 \u_multiplier/STAGE1/_2088_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[22]),
    .ZN(\u_multiplier/STAGE1/_0811_ ));
 AND2_X1 \u_multiplier/STAGE1/_2089_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[23]),
    .ZN(\u_multiplier/STAGE1/_0812_ ));
 AND2_X1 \u_multiplier/STAGE1/_2090_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[24]),
    .ZN(\u_multiplier/STAGE1/_0813_ ));
 AND2_X1 \u_multiplier/STAGE1/_2091_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[25]),
    .ZN(\u_multiplier/STAGE1/_0814_ ));
 AND2_X1 \u_multiplier/STAGE1/_2092_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[26]),
    .ZN(\u_multiplier/STAGE1/_0815_ ));
 AND2_X1 \u_multiplier/STAGE1/_2093_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/STAGE1/_0816_ ));
 AND2_X1 \u_multiplier/STAGE1/_2094_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/pp1_29 [14]));
 AND2_X1 \u_multiplier/STAGE1/_2095_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/pp1_29 [15]));
 AND2_X1 \u_multiplier/STAGE1/_2096_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/STAGE1/_0817_ ));
 AND2_X1 \u_multiplier/STAGE1/_2097_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/STAGE1/_0818_ ));
 AND2_X1 \u_multiplier/STAGE1/_2098_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/STAGE1/_0819_ ));
 AND2_X1 \u_multiplier/STAGE1/_2099_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[27]),
    .ZN(\u_multiplier/STAGE1/_0820_ ));
 AND2_X1 \u_multiplier/STAGE1/_2100_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[26]),
    .ZN(\u_multiplier/STAGE1/_0821_ ));
 AND2_X1 \u_multiplier/STAGE1/_2101_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[25]),
    .ZN(\u_multiplier/STAGE1/_0822_ ));
 AND2_X1 \u_multiplier/STAGE1/_2102_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[24]),
    .ZN(\u_multiplier/STAGE1/_0823_ ));
 AND2_X1 \u_multiplier/STAGE1/_2103_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[23]),
    .ZN(\u_multiplier/STAGE1/_0824_ ));
 AND2_X1 \u_multiplier/STAGE1/_2104_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[22]),
    .ZN(\u_multiplier/STAGE1/_0825_ ));
 AND2_X1 \u_multiplier/STAGE1/_2105_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[21]),
    .ZN(\u_multiplier/STAGE1/_0826_ ));
 AND2_X1 \u_multiplier/STAGE1/_2106_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[20]),
    .ZN(\u_multiplier/STAGE1/_0827_ ));
 AND2_X1 \u_multiplier/STAGE1/_2107_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0828_ ));
 AND2_X1 \u_multiplier/STAGE1/_2108_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0829_ ));
 AND2_X1 \u_multiplier/STAGE1/_2109_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0830_ ));
 AND2_X1 \u_multiplier/STAGE1/_2110_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[16]),
    .ZN(\u_multiplier/STAGE1/_0831_ ));
 AND2_X1 \u_multiplier/STAGE1/_2111_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[15]),
    .ZN(\u_multiplier/STAGE1/_0832_ ));
 AND2_X1 \u_multiplier/STAGE1/_2112_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[16]),
    .ZN(\u_multiplier/STAGE1/_0833_ ));
 AND2_X1 \u_multiplier/STAGE1/_2113_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0834_ ));
 AND2_X1 \u_multiplier/STAGE1/_2114_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0835_ ));
 AND2_X1 \u_multiplier/STAGE1/_2115_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0836_ ));
 AND2_X1 \u_multiplier/STAGE1/_2116_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[20]),
    .ZN(\u_multiplier/STAGE1/_0837_ ));
 AND2_X1 \u_multiplier/STAGE1/_2117_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[21]),
    .ZN(\u_multiplier/STAGE1/_0838_ ));
 AND2_X1 \u_multiplier/STAGE1/_2118_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[22]),
    .ZN(\u_multiplier/STAGE1/_0839_ ));
 AND2_X1 \u_multiplier/STAGE1/_2119_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[23]),
    .ZN(\u_multiplier/STAGE1/_0840_ ));
 AND2_X1 \u_multiplier/STAGE1/_2120_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[24]),
    .ZN(\u_multiplier/STAGE1/_0841_ ));
 AND2_X1 \u_multiplier/STAGE1/_2121_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[25]),
    .ZN(\u_multiplier/STAGE1/_0842_ ));
 AND2_X1 \u_multiplier/STAGE1/_2122_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[26]),
    .ZN(\u_multiplier/STAGE1/_0843_ ));
 AND2_X1 \u_multiplier/STAGE1/_2123_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/STAGE1/_0844_ ));
 AND2_X1 \u_multiplier/STAGE1/_2124_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/STAGE1/_0845_ ));
 AND2_X1 \u_multiplier/STAGE1/_2125_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/STAGE1/_0846_ ));
 AND2_X1 \u_multiplier/STAGE1/_2126_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/pp1_30 [15]));
 AND2_X1 \u_multiplier/STAGE1/_2127_  (.A1(data_in_reg[0]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/STAGE1/_0847_ ));
 AND2_X1 \u_multiplier/STAGE1/_2128_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/STAGE1/_0848_ ));
 AND2_X1 \u_multiplier/STAGE1/_2129_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/STAGE1/_0849_ ));
 AND2_X1 \u_multiplier/STAGE1/_2130_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/STAGE1/_0850_ ));
 AND2_X1 \u_multiplier/STAGE1/_2131_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[27]),
    .ZN(\u_multiplier/STAGE1/_0851_ ));
 AND2_X1 \u_multiplier/STAGE1/_2132_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[26]),
    .ZN(\u_multiplier/STAGE1/_0852_ ));
 AND2_X1 \u_multiplier/STAGE1/_2133_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[25]),
    .ZN(\u_multiplier/STAGE1/_0853_ ));
 AND2_X1 \u_multiplier/STAGE1/_2134_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[24]),
    .ZN(\u_multiplier/STAGE1/_0854_ ));
 AND2_X1 \u_multiplier/STAGE1/_2135_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[23]),
    .ZN(\u_multiplier/STAGE1/_0855_ ));
 AND2_X1 \u_multiplier/STAGE1/_2136_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[22]),
    .ZN(\u_multiplier/STAGE1/_0856_ ));
 AND2_X1 \u_multiplier/STAGE1/_2137_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[21]),
    .ZN(\u_multiplier/STAGE1/_0857_ ));
 AND2_X1 \u_multiplier/STAGE1/_2138_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[20]),
    .ZN(\u_multiplier/STAGE1/_0858_ ));
 AND2_X1 \u_multiplier/STAGE1/_2139_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0859_ ));
 AND2_X1 \u_multiplier/STAGE1/_2140_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0860_ ));
 AND2_X1 \u_multiplier/STAGE1/_2141_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0861_ ));
 AND2_X1 \u_multiplier/STAGE1/_2142_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[16]),
    .ZN(\u_multiplier/STAGE1/_0862_ ));
 AND2_X1 \u_multiplier/STAGE1/_2143_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[16]),
    .ZN(\u_multiplier/STAGE1/_0863_ ));
 AND2_X1 \u_multiplier/STAGE1/_2144_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0864_ ));
 AND2_X1 \u_multiplier/STAGE1/_2145_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0865_ ));
 AND2_X1 \u_multiplier/STAGE1/_2146_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0866_ ));
 AND2_X1 \u_multiplier/STAGE1/_2147_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[20]),
    .ZN(\u_multiplier/STAGE1/_0867_ ));
 AND2_X1 \u_multiplier/STAGE1/_2148_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[21]),
    .ZN(\u_multiplier/STAGE1/_0868_ ));
 AND2_X1 \u_multiplier/STAGE1/_2149_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[22]),
    .ZN(\u_multiplier/STAGE1/_0869_ ));
 AND2_X1 \u_multiplier/STAGE1/_2150_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[23]),
    .ZN(\u_multiplier/STAGE1/_0870_ ));
 AND2_X1 \u_multiplier/STAGE1/_2151_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[24]),
    .ZN(\u_multiplier/STAGE1/_0871_ ));
 AND2_X1 \u_multiplier/STAGE1/_2152_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[25]),
    .ZN(\u_multiplier/STAGE1/_0872_ ));
 AND2_X1 \u_multiplier/STAGE1/_2153_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[26]),
    .ZN(\u_multiplier/STAGE1/_0873_ ));
 AND2_X1 \u_multiplier/STAGE1/_2154_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/STAGE1/_0874_ ));
 AND2_X1 \u_multiplier/STAGE1/_2155_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/STAGE1/_0875_ ));
 AND2_X1 \u_multiplier/STAGE1/_2156_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/STAGE1/_0876_ ));
 AND2_X1 \u_multiplier/STAGE1/_2157_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/STAGE1/_0877_ ));
 AND2_X1 \u_multiplier/STAGE1/_2158_  (.A1(sram_rdata_reg[0]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/STAGE1/_0878_ ));
 AND2_X1 \u_multiplier/STAGE1/_2159_  (.A1(data_in_reg[1]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/STAGE1/_0879_ ));
 AND2_X1 \u_multiplier/STAGE1/_2160_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/STAGE1/_0880_ ));
 AND2_X1 \u_multiplier/STAGE1/_2161_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/STAGE1/_0881_ ));
 AND2_X1 \u_multiplier/STAGE1/_2162_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/STAGE1/_0882_ ));
 AND2_X1 \u_multiplier/STAGE1/_2163_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[27]),
    .ZN(\u_multiplier/STAGE1/_0883_ ));
 AND2_X1 \u_multiplier/STAGE1/_2164_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[26]),
    .ZN(\u_multiplier/STAGE1/_0884_ ));
 AND2_X1 \u_multiplier/STAGE1/_2165_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[25]),
    .ZN(\u_multiplier/STAGE1/_0885_ ));
 AND2_X1 \u_multiplier/STAGE1/_2166_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[24]),
    .ZN(\u_multiplier/STAGE1/_0886_ ));
 AND2_X1 \u_multiplier/STAGE1/_2167_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[23]),
    .ZN(\u_multiplier/STAGE1/_0887_ ));
 AND2_X1 \u_multiplier/STAGE1/_2168_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[22]),
    .ZN(\u_multiplier/STAGE1/_0888_ ));
 AND2_X1 \u_multiplier/STAGE1/_2169_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[21]),
    .ZN(\u_multiplier/STAGE1/_0889_ ));
 AND2_X1 \u_multiplier/STAGE1/_2170_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[20]),
    .ZN(\u_multiplier/STAGE1/_0890_ ));
 AND2_X1 \u_multiplier/STAGE1/_2171_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0891_ ));
 AND2_X1 \u_multiplier/STAGE1/_2172_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0892_ ));
 AND2_X1 \u_multiplier/STAGE1/_2173_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0893_ ));
 AND2_X1 \u_multiplier/STAGE1/_2174_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[16]),
    .ZN(\u_multiplier/STAGE1/_0894_ ));
 AND2_X1 \u_multiplier/STAGE1/_2175_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0895_ ));
 AND2_X1 \u_multiplier/STAGE1/_2176_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0896_ ));
 AND2_X1 \u_multiplier/STAGE1/_2177_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0897_ ));
 AND2_X1 \u_multiplier/STAGE1/_2178_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[20]),
    .ZN(\u_multiplier/STAGE1/_0898_ ));
 AND2_X1 \u_multiplier/STAGE1/_2179_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[21]),
    .ZN(\u_multiplier/STAGE1/_0899_ ));
 AND2_X1 \u_multiplier/STAGE1/_2180_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[22]),
    .ZN(\u_multiplier/STAGE1/_0900_ ));
 AND2_X1 \u_multiplier/STAGE1/_2181_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[23]),
    .ZN(\u_multiplier/STAGE1/_0901_ ));
 AND2_X1 \u_multiplier/STAGE1/_2182_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[24]),
    .ZN(\u_multiplier/STAGE1/_0902_ ));
 AND2_X1 \u_multiplier/STAGE1/_2183_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[25]),
    .ZN(\u_multiplier/STAGE1/_0903_ ));
 AND2_X1 \u_multiplier/STAGE1/_2184_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[26]),
    .ZN(\u_multiplier/STAGE1/_0904_ ));
 AND2_X1 \u_multiplier/STAGE1/_2185_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/STAGE1/_0905_ ));
 AND2_X1 \u_multiplier/STAGE1/_2186_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/STAGE1/_0906_ ));
 AND2_X1 \u_multiplier/STAGE1/_2187_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/STAGE1/_0907_ ));
 AND2_X1 \u_multiplier/STAGE1/_2188_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/STAGE1/_0908_ ));
 AND2_X1 \u_multiplier/STAGE1/_2189_  (.A1(sram_rdata_reg[1]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/STAGE1/_0909_ ));
 AND2_X1 \u_multiplier/STAGE1/_2190_  (.A1(data_in_reg[2]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/STAGE1/_0910_ ));
 AND2_X1 \u_multiplier/STAGE1/_2191_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/STAGE1/_0911_ ));
 AND2_X1 \u_multiplier/STAGE1/_2192_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/STAGE1/_0912_ ));
 AND2_X1 \u_multiplier/STAGE1/_2193_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/STAGE1/_0913_ ));
 AND2_X1 \u_multiplier/STAGE1/_2194_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[27]),
    .ZN(\u_multiplier/STAGE1/_0914_ ));
 AND2_X1 \u_multiplier/STAGE1/_2195_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[26]),
    .ZN(\u_multiplier/STAGE1/_0915_ ));
 AND2_X1 \u_multiplier/STAGE1/_2196_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[25]),
    .ZN(\u_multiplier/STAGE1/_0916_ ));
 AND2_X1 \u_multiplier/STAGE1/_2197_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[24]),
    .ZN(\u_multiplier/STAGE1/_0917_ ));
 AND2_X1 \u_multiplier/STAGE1/_2198_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[23]),
    .ZN(\u_multiplier/STAGE1/_0918_ ));
 AND2_X1 \u_multiplier/STAGE1/_2199_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[22]),
    .ZN(\u_multiplier/STAGE1/_0919_ ));
 AND2_X1 \u_multiplier/STAGE1/_2200_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[21]),
    .ZN(\u_multiplier/STAGE1/_0920_ ));
 AND2_X1 \u_multiplier/STAGE1/_2201_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[20]),
    .ZN(\u_multiplier/STAGE1/_0921_ ));
 AND2_X1 \u_multiplier/STAGE1/_2202_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0922_ ));
 AND2_X1 \u_multiplier/STAGE1/_2203_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0923_ ));
 AND2_X1 \u_multiplier/STAGE1/_2204_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0924_ ));
 AND2_X1 \u_multiplier/STAGE1/_2205_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0925_ ));
 AND2_X1 \u_multiplier/STAGE1/_2206_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0926_ ));
 AND2_X1 \u_multiplier/STAGE1/_2207_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0927_ ));
 AND2_X1 \u_multiplier/STAGE1/_2208_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[20]),
    .ZN(\u_multiplier/STAGE1/_0928_ ));
 AND2_X1 \u_multiplier/STAGE1/_2209_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[21]),
    .ZN(\u_multiplier/STAGE1/_0929_ ));
 AND2_X1 \u_multiplier/STAGE1/_2210_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[22]),
    .ZN(\u_multiplier/STAGE1/_0930_ ));
 AND2_X1 \u_multiplier/STAGE1/_2211_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[23]),
    .ZN(\u_multiplier/STAGE1/_0931_ ));
 AND2_X1 \u_multiplier/STAGE1/_2212_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[24]),
    .ZN(\u_multiplier/STAGE1/_0932_ ));
 AND2_X1 \u_multiplier/STAGE1/_2213_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[25]),
    .ZN(\u_multiplier/STAGE1/_0933_ ));
 AND2_X1 \u_multiplier/STAGE1/_2214_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[26]),
    .ZN(\u_multiplier/STAGE1/_0934_ ));
 AND2_X1 \u_multiplier/STAGE1/_2215_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/STAGE1/_0935_ ));
 AND2_X1 \u_multiplier/STAGE1/_2216_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/STAGE1/_0936_ ));
 AND2_X1 \u_multiplier/STAGE1/_2217_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/STAGE1/_0937_ ));
 AND2_X2 \u_multiplier/STAGE1/_2218_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/STAGE1/_0938_ ));
 AND2_X2 \u_multiplier/STAGE1/_2219_  (.A1(sram_rdata_reg[2]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/STAGE1/_0939_ ));
 AND2_X1 \u_multiplier/STAGE1/_2220_  (.A1(data_in_reg[3]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/STAGE1/_0940_ ));
 AND2_X1 \u_multiplier/STAGE1/_2221_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/STAGE1/_0941_ ));
 AND2_X1 \u_multiplier/STAGE1/_2222_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/STAGE1/_0942_ ));
 AND2_X1 \u_multiplier/STAGE1/_2223_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/STAGE1/_0943_ ));
 AND2_X1 \u_multiplier/STAGE1/_2224_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[27]),
    .ZN(\u_multiplier/STAGE1/_0944_ ));
 AND2_X1 \u_multiplier/STAGE1/_2225_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[26]),
    .ZN(\u_multiplier/STAGE1/_0945_ ));
 AND2_X1 \u_multiplier/STAGE1/_2226_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[25]),
    .ZN(\u_multiplier/STAGE1/_0946_ ));
 AND2_X1 \u_multiplier/STAGE1/_2227_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[24]),
    .ZN(\u_multiplier/STAGE1/_0947_ ));
 AND2_X1 \u_multiplier/STAGE1/_2228_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[23]),
    .ZN(\u_multiplier/STAGE1/_0948_ ));
 AND2_X1 \u_multiplier/STAGE1/_2229_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[22]),
    .ZN(\u_multiplier/STAGE1/_0949_ ));
 AND2_X1 \u_multiplier/STAGE1/_2230_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[21]),
    .ZN(\u_multiplier/STAGE1/_0950_ ));
 AND2_X1 \u_multiplier/STAGE1/_2231_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[20]),
    .ZN(\u_multiplier/STAGE1/_0951_ ));
 AND2_X1 \u_multiplier/STAGE1/_2232_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0952_ ));
 AND2_X1 \u_multiplier/STAGE1/_2233_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0953_ ));
 AND2_X1 \u_multiplier/STAGE1/_2234_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[17]),
    .ZN(\u_multiplier/STAGE1/_0954_ ));
 AND2_X1 \u_multiplier/STAGE1/_2235_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0955_ ));
 AND2_X1 \u_multiplier/STAGE1/_2236_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0956_ ));
 AND2_X1 \u_multiplier/STAGE1/_2237_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[20]),
    .ZN(\u_multiplier/STAGE1/_0957_ ));
 AND2_X1 \u_multiplier/STAGE1/_2238_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[21]),
    .ZN(\u_multiplier/STAGE1/_0958_ ));
 AND2_X1 \u_multiplier/STAGE1/_2239_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[22]),
    .ZN(\u_multiplier/STAGE1/_0959_ ));
 AND2_X1 \u_multiplier/STAGE1/_2240_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[23]),
    .ZN(\u_multiplier/STAGE1/_0960_ ));
 AND2_X1 \u_multiplier/STAGE1/_2241_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[24]),
    .ZN(\u_multiplier/STAGE1/_0961_ ));
 AND2_X1 \u_multiplier/STAGE1/_2242_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[25]),
    .ZN(\u_multiplier/STAGE1/_0962_ ));
 AND2_X1 \u_multiplier/STAGE1/_2243_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[26]),
    .ZN(\u_multiplier/STAGE1/_0963_ ));
 AND2_X1 \u_multiplier/STAGE1/_2244_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/STAGE1/_0964_ ));
 AND2_X1 \u_multiplier/STAGE1/_2245_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/STAGE1/_0965_ ));
 AND2_X1 \u_multiplier/STAGE1/_2246_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/STAGE1/_0966_ ));
 AND2_X1 \u_multiplier/STAGE1/_2247_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/STAGE1/_0967_ ));
 AND2_X1 \u_multiplier/STAGE1/_2248_  (.A1(sram_rdata_reg[3]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp1_34 [15]));
 AND2_X1 \u_multiplier/STAGE1/_2249_  (.A1(data_in_reg[4]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/STAGE1/_0968_ ));
 AND2_X1 \u_multiplier/STAGE1/_2250_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/STAGE1/_0969_ ));
 AND2_X1 \u_multiplier/STAGE1/_2251_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/STAGE1/_0970_ ));
 AND2_X1 \u_multiplier/STAGE1/_2252_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/STAGE1/_0971_ ));
 AND2_X1 \u_multiplier/STAGE1/_2253_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[27]),
    .ZN(\u_multiplier/STAGE1/_0972_ ));
 AND2_X1 \u_multiplier/STAGE1/_2254_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[26]),
    .ZN(\u_multiplier/STAGE1/_0973_ ));
 AND2_X1 \u_multiplier/STAGE1/_2255_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[25]),
    .ZN(\u_multiplier/STAGE1/_0974_ ));
 AND2_X1 \u_multiplier/STAGE1/_2256_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[24]),
    .ZN(\u_multiplier/STAGE1/_0975_ ));
 AND2_X1 \u_multiplier/STAGE1/_2257_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[23]),
    .ZN(\u_multiplier/STAGE1/_0976_ ));
 AND2_X1 \u_multiplier/STAGE1/_2258_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[22]),
    .ZN(\u_multiplier/STAGE1/_0977_ ));
 AND2_X1 \u_multiplier/STAGE1/_2259_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[21]),
    .ZN(\u_multiplier/STAGE1/_0978_ ));
 AND2_X1 \u_multiplier/STAGE1/_2260_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[20]),
    .ZN(\u_multiplier/STAGE1/_0979_ ));
 AND2_X1 \u_multiplier/STAGE1/_2261_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0980_ ));
 AND2_X1 \u_multiplier/STAGE1/_2262_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0981_ ));
 AND2_X1 \u_multiplier/STAGE1/_2263_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[18]),
    .ZN(\u_multiplier/STAGE1/_0982_ ));
 AND2_X1 \u_multiplier/STAGE1/_2264_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[19]),
    .ZN(\u_multiplier/STAGE1/_0983_ ));
 AND2_X1 \u_multiplier/STAGE1/_2265_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[20]),
    .ZN(\u_multiplier/STAGE1/_0984_ ));
 AND2_X1 \u_multiplier/STAGE1/_2266_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[21]),
    .ZN(\u_multiplier/STAGE1/_0985_ ));
 AND2_X1 \u_multiplier/STAGE1/_2267_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[22]),
    .ZN(\u_multiplier/STAGE1/_0986_ ));
 AND2_X1 \u_multiplier/STAGE1/_2268_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[23]),
    .ZN(\u_multiplier/STAGE1/_0987_ ));
 AND2_X1 \u_multiplier/STAGE1/_2269_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[24]),
    .ZN(\u_multiplier/STAGE1/_0988_ ));
 AND2_X1 \u_multiplier/STAGE1/_2270_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[25]),
    .ZN(\u_multiplier/STAGE1/_0989_ ));
 AND2_X1 \u_multiplier/STAGE1/_2271_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[26]),
    .ZN(\u_multiplier/STAGE1/_0990_ ));
 AND2_X1 \u_multiplier/STAGE1/_2272_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/STAGE1/_0991_ ));
 AND2_X1 \u_multiplier/STAGE1/_2273_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/STAGE1/_0992_ ));
 AND2_X1 \u_multiplier/STAGE1/_2274_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/STAGE1/_0993_ ));
 AND2_X1 \u_multiplier/STAGE1/_2275_  (.A1(sram_rdata_reg[4]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp1_35 [14]));
 AND2_X1 \u_multiplier/STAGE1/_2276_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/pp1_35 [15]));
 AND2_X1 \u_multiplier/STAGE1/_2277_  (.A1(data_in_reg[5]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/STAGE1/_0994_ ));
 AND2_X1 \u_multiplier/STAGE1/_2278_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/STAGE1/_0995_ ));
 AND2_X1 \u_multiplier/STAGE1/_2279_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/STAGE1/_0996_ ));
 AND2_X1 \u_multiplier/STAGE1/_2280_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/STAGE1/_0997_ ));
 AND2_X1 \u_multiplier/STAGE1/_2281_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[27]),
    .ZN(\u_multiplier/STAGE1/_0998_ ));
 AND2_X1 \u_multiplier/STAGE1/_2282_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[26]),
    .ZN(\u_multiplier/STAGE1/_0999_ ));
 AND2_X1 \u_multiplier/STAGE1/_2283_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[25]),
    .ZN(\u_multiplier/STAGE1/_1000_ ));
 AND2_X1 \u_multiplier/STAGE1/_2284_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[24]),
    .ZN(\u_multiplier/STAGE1/_1001_ ));
 AND2_X1 \u_multiplier/STAGE1/_2285_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[23]),
    .ZN(\u_multiplier/STAGE1/_1002_ ));
 AND2_X1 \u_multiplier/STAGE1/_2286_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[22]),
    .ZN(\u_multiplier/STAGE1/_1003_ ));
 AND2_X1 \u_multiplier/STAGE1/_2287_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[21]),
    .ZN(\u_multiplier/STAGE1/_1004_ ));
 AND2_X1 \u_multiplier/STAGE1/_2288_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[20]),
    .ZN(\u_multiplier/STAGE1/_1005_ ));
 AND2_X1 \u_multiplier/STAGE1/_2289_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[19]),
    .ZN(\u_multiplier/STAGE1/_1006_ ));
 AND2_X1 \u_multiplier/STAGE1/_2290_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[18]),
    .ZN(\u_multiplier/STAGE1/_1007_ ));
 AND2_X1 \u_multiplier/STAGE1/_2291_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[19]),
    .ZN(\u_multiplier/STAGE1/_1008_ ));
 AND2_X1 \u_multiplier/STAGE1/_2292_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[20]),
    .ZN(\u_multiplier/STAGE1/_1009_ ));
 AND2_X1 \u_multiplier/STAGE1/_2293_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[21]),
    .ZN(\u_multiplier/STAGE1/_1010_ ));
 AND2_X1 \u_multiplier/STAGE1/_2294_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[22]),
    .ZN(\u_multiplier/STAGE1/_1011_ ));
 AND2_X1 \u_multiplier/STAGE1/_2295_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[23]),
    .ZN(\u_multiplier/STAGE1/_1012_ ));
 AND2_X1 \u_multiplier/STAGE1/_2296_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[24]),
    .ZN(\u_multiplier/STAGE1/_1013_ ));
 AND2_X1 \u_multiplier/STAGE1/_2297_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[25]),
    .ZN(\u_multiplier/STAGE1/_1014_ ));
 AND2_X1 \u_multiplier/STAGE1/_2298_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[26]),
    .ZN(\u_multiplier/STAGE1/_1015_ ));
 AND2_X1 \u_multiplier/STAGE1/_2299_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/STAGE1/_1016_ ));
 AND2_X1 \u_multiplier/STAGE1/_2300_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/STAGE1/_1017_ ));
 AND2_X1 \u_multiplier/STAGE1/_2301_  (.A1(sram_rdata_reg[5]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp1_36 [13]));
 AND2_X1 \u_multiplier/STAGE1/_2302_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/pp1_36 [14]));
 AND2_X1 \u_multiplier/STAGE1/_2303_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/pp1_36 [15]));
 AND2_X1 \u_multiplier/STAGE1/_2304_  (.A1(data_in_reg[6]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/STAGE1/_1018_ ));
 AND2_X1 \u_multiplier/STAGE1/_2305_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/STAGE1/_1019_ ));
 AND2_X1 \u_multiplier/STAGE1/_2306_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/STAGE1/_1020_ ));
 AND2_X1 \u_multiplier/STAGE1/_2307_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/STAGE1/_1021_ ));
 AND2_X1 \u_multiplier/STAGE1/_2308_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[27]),
    .ZN(\u_multiplier/STAGE1/_1022_ ));
 AND2_X1 \u_multiplier/STAGE1/_2309_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[26]),
    .ZN(\u_multiplier/STAGE1/_1023_ ));
 AND2_X1 \u_multiplier/STAGE1/_2310_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[25]),
    .ZN(\u_multiplier/STAGE1/_1024_ ));
 AND2_X1 \u_multiplier/STAGE1/_2311_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[24]),
    .ZN(\u_multiplier/STAGE1/_1025_ ));
 AND2_X1 \u_multiplier/STAGE1/_2312_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[23]),
    .ZN(\u_multiplier/STAGE1/_1026_ ));
 AND2_X1 \u_multiplier/STAGE1/_2313_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[22]),
    .ZN(\u_multiplier/STAGE1/_1027_ ));
 AND2_X1 \u_multiplier/STAGE1/_2314_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[21]),
    .ZN(\u_multiplier/STAGE1/_1028_ ));
 AND2_X1 \u_multiplier/STAGE1/_2315_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[20]),
    .ZN(\u_multiplier/STAGE1/_1029_ ));
 AND2_X1 \u_multiplier/STAGE1/_2316_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[19]),
    .ZN(\u_multiplier/STAGE1/_1030_ ));
 AND2_X1 \u_multiplier/STAGE1/_2317_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[19]),
    .ZN(\u_multiplier/STAGE1/_1031_ ));
 AND2_X1 \u_multiplier/STAGE1/_2318_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[20]),
    .ZN(\u_multiplier/STAGE1/_1032_ ));
 AND2_X1 \u_multiplier/STAGE1/_2319_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[21]),
    .ZN(\u_multiplier/STAGE1/_1033_ ));
 AND2_X1 \u_multiplier/STAGE1/_2320_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[22]),
    .ZN(\u_multiplier/STAGE1/_1034_ ));
 AND2_X1 \u_multiplier/STAGE1/_2321_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[23]),
    .ZN(\u_multiplier/STAGE1/_1035_ ));
 AND2_X1 \u_multiplier/STAGE1/_2322_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[24]),
    .ZN(\u_multiplier/STAGE1/_1036_ ));
 AND2_X1 \u_multiplier/STAGE1/_2323_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[25]),
    .ZN(\u_multiplier/STAGE1/_1037_ ));
 AND2_X1 \u_multiplier/STAGE1/_2324_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[26]),
    .ZN(\u_multiplier/STAGE1/_1038_ ));
 AND2_X1 \u_multiplier/STAGE1/_2325_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/STAGE1/_1039_ ));
 AND2_X1 \u_multiplier/STAGE1/_2326_  (.A1(sram_rdata_reg[6]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp1_37 [12]));
 AND2_X1 \u_multiplier/STAGE1/_2327_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/pp1_37 [13]));
 AND2_X1 \u_multiplier/STAGE1/_2328_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/pp1_37 [14]));
 AND2_X1 \u_multiplier/STAGE1/_2329_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/pp1_37 [15]));
 AND2_X1 \u_multiplier/STAGE1/_2330_  (.A1(data_in_reg[7]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/STAGE1/_1040_ ));
 AND2_X1 \u_multiplier/STAGE1/_2331_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/STAGE1/_1041_ ));
 AND2_X1 \u_multiplier/STAGE1/_2332_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/STAGE1/_1042_ ));
 AND2_X1 \u_multiplier/STAGE1/_2333_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/STAGE1/_1043_ ));
 AND2_X1 \u_multiplier/STAGE1/_2334_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[27]),
    .ZN(\u_multiplier/STAGE1/_1044_ ));
 AND2_X1 \u_multiplier/STAGE1/_2335_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[26]),
    .ZN(\u_multiplier/STAGE1/_1045_ ));
 AND2_X1 \u_multiplier/STAGE1/_2336_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[25]),
    .ZN(\u_multiplier/STAGE1/_1046_ ));
 AND2_X1 \u_multiplier/STAGE1/_2337_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[24]),
    .ZN(\u_multiplier/STAGE1/_1047_ ));
 AND2_X1 \u_multiplier/STAGE1/_2338_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[23]),
    .ZN(\u_multiplier/STAGE1/_1048_ ));
 AND2_X1 \u_multiplier/STAGE1/_2339_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[22]),
    .ZN(\u_multiplier/STAGE1/_1049_ ));
 AND2_X1 \u_multiplier/STAGE1/_2340_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[21]),
    .ZN(\u_multiplier/STAGE1/_1050_ ));
 AND2_X1 \u_multiplier/STAGE1/_2341_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[20]),
    .ZN(\u_multiplier/STAGE1/_1051_ ));
 AND2_X1 \u_multiplier/STAGE1/_2342_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[19]),
    .ZN(\u_multiplier/STAGE1/_1052_ ));
 AND2_X1 \u_multiplier/STAGE1/_2343_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[20]),
    .ZN(\u_multiplier/STAGE1/_1053_ ));
 AND2_X1 \u_multiplier/STAGE1/_2344_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[21]),
    .ZN(\u_multiplier/STAGE1/_1054_ ));
 AND2_X1 \u_multiplier/STAGE1/_2345_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[22]),
    .ZN(\u_multiplier/STAGE1/_1055_ ));
 AND2_X1 \u_multiplier/STAGE1/_2346_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[23]),
    .ZN(\u_multiplier/STAGE1/_1056_ ));
 AND2_X1 \u_multiplier/STAGE1/_2347_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[24]),
    .ZN(\u_multiplier/STAGE1/_1057_ ));
 AND2_X1 \u_multiplier/STAGE1/_2348_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[25]),
    .ZN(\u_multiplier/STAGE1/_1058_ ));
 AND2_X1 \u_multiplier/STAGE1/_2349_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[26]),
    .ZN(\u_multiplier/STAGE1/_1059_ ));
 AND2_X1 \u_multiplier/STAGE1/_2350_  (.A1(sram_rdata_reg[7]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp1_38 [11]));
 AND2_X1 \u_multiplier/STAGE1/_2351_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/pp1_38 [12]));
 AND2_X1 \u_multiplier/STAGE1/_2352_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/pp1_38 [13]));
 AND2_X1 \u_multiplier/STAGE1/_2353_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/pp1_38 [14]));
 AND2_X1 \u_multiplier/STAGE1/_2354_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/pp1_38 [15]));
 AND2_X1 \u_multiplier/STAGE1/_2355_  (.A1(data_in_reg[8]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/STAGE1/_1060_ ));
 AND2_X1 \u_multiplier/STAGE1/_2356_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/STAGE1/_1061_ ));
 AND2_X1 \u_multiplier/STAGE1/_2357_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/STAGE1/_1062_ ));
 AND2_X1 \u_multiplier/STAGE1/_2358_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/STAGE1/_1063_ ));
 AND2_X1 \u_multiplier/STAGE1/_2359_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[27]),
    .ZN(\u_multiplier/STAGE1/_1064_ ));
 AND2_X1 \u_multiplier/STAGE1/_2360_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[26]),
    .ZN(\u_multiplier/STAGE1/_1065_ ));
 AND2_X1 \u_multiplier/STAGE1/_2361_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[25]),
    .ZN(\u_multiplier/STAGE1/_1066_ ));
 AND2_X1 \u_multiplier/STAGE1/_2362_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[24]),
    .ZN(\u_multiplier/STAGE1/_1067_ ));
 AND2_X1 \u_multiplier/STAGE1/_2363_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[23]),
    .ZN(\u_multiplier/STAGE1/_1068_ ));
 AND2_X1 \u_multiplier/STAGE1/_2364_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[22]),
    .ZN(\u_multiplier/STAGE1/_1069_ ));
 AND2_X1 \u_multiplier/STAGE1/_2365_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[21]),
    .ZN(\u_multiplier/STAGE1/_1070_ ));
 AND2_X1 \u_multiplier/STAGE1/_2366_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[20]),
    .ZN(\u_multiplier/STAGE1/_1071_ ));
 AND2_X1 \u_multiplier/STAGE1/_2367_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[20]),
    .ZN(\u_multiplier/STAGE1/_1072_ ));
 AND2_X1 \u_multiplier/STAGE1/_2368_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[21]),
    .ZN(\u_multiplier/STAGE1/_1073_ ));
 AND2_X1 \u_multiplier/STAGE1/_2369_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[22]),
    .ZN(\u_multiplier/STAGE1/_1074_ ));
 AND2_X1 \u_multiplier/STAGE1/_2370_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[23]),
    .ZN(\u_multiplier/STAGE1/_1075_ ));
 AND2_X1 \u_multiplier/STAGE1/_2371_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[24]),
    .ZN(\u_multiplier/STAGE1/_1076_ ));
 AND2_X1 \u_multiplier/STAGE1/_2372_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[25]),
    .ZN(\u_multiplier/STAGE1/_1077_ ));
 AND2_X1 \u_multiplier/STAGE1/_2373_  (.A1(sram_rdata_reg[8]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp1_39 [10]));
 AND2_X1 \u_multiplier/STAGE1/_2374_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/pp1_39 [11]));
 AND2_X1 \u_multiplier/STAGE1/_2375_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/pp1_39 [12]));
 AND2_X1 \u_multiplier/STAGE1/_2376_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/pp1_39 [13]));
 AND2_X1 \u_multiplier/STAGE1/_2377_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/pp1_39 [14]));
 AND2_X1 \u_multiplier/STAGE1/_2378_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[26]),
    .ZN(\u_multiplier/pp1_39 [15]));
 AND2_X1 \u_multiplier/STAGE1/_2379_  (.A1(data_in_reg[9]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/STAGE1/_1078_ ));
 AND2_X1 \u_multiplier/STAGE1/_2380_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/STAGE1/_1079_ ));
 AND2_X1 \u_multiplier/STAGE1/_2381_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/STAGE1/_1080_ ));
 AND2_X1 \u_multiplier/STAGE1/_2382_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/STAGE1/_1081_ ));
 AND2_X1 \u_multiplier/STAGE1/_2383_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[27]),
    .ZN(\u_multiplier/STAGE1/_1082_ ));
 AND2_X1 \u_multiplier/STAGE1/_2384_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[26]),
    .ZN(\u_multiplier/STAGE1/_1083_ ));
 AND2_X1 \u_multiplier/STAGE1/_2385_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[25]),
    .ZN(\u_multiplier/STAGE1/_1084_ ));
 AND2_X1 \u_multiplier/STAGE1/_2386_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[24]),
    .ZN(\u_multiplier/STAGE1/_1085_ ));
 AND2_X1 \u_multiplier/STAGE1/_2387_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[23]),
    .ZN(\u_multiplier/STAGE1/_1086_ ));
 AND2_X1 \u_multiplier/STAGE1/_2388_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[22]),
    .ZN(\u_multiplier/STAGE1/_1087_ ));
 AND2_X1 \u_multiplier/STAGE1/_2389_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[21]),
    .ZN(\u_multiplier/STAGE1/_1088_ ));
 AND2_X1 \u_multiplier/STAGE1/_2390_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[20]),
    .ZN(\u_multiplier/STAGE1/_1089_ ));
 AND2_X1 \u_multiplier/STAGE1/_2391_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[21]),
    .ZN(\u_multiplier/STAGE1/_1090_ ));
 AND2_X1 \u_multiplier/STAGE1/_2392_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[22]),
    .ZN(\u_multiplier/STAGE1/_1091_ ));
 AND2_X1 \u_multiplier/STAGE1/_2393_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[23]),
    .ZN(\u_multiplier/STAGE1/_1092_ ));
 AND2_X1 \u_multiplier/STAGE1/_2394_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[24]),
    .ZN(\u_multiplier/STAGE1/_1093_ ));
 AND2_X1 \u_multiplier/STAGE1/_2395_  (.A1(sram_rdata_reg[9]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp1_40 [9]));
 AND2_X1 \u_multiplier/STAGE1/_2396_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/pp1_40 [10]));
 AND2_X1 \u_multiplier/STAGE1/_2397_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/pp1_40 [11]));
 AND2_X1 \u_multiplier/STAGE1/_2398_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/pp1_40 [12]));
 AND2_X1 \u_multiplier/STAGE1/_2399_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/pp1_40 [13]));
 AND2_X1 \u_multiplier/STAGE1/_2400_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[26]),
    .ZN(\u_multiplier/pp1_40 [14]));
 AND2_X1 \u_multiplier/STAGE1/_2401_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[25]),
    .ZN(\u_multiplier/pp1_40 [15]));
 AND2_X1 \u_multiplier/STAGE1/_2402_  (.A1(data_in_reg[10]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/STAGE1/_1094_ ));
 AND2_X1 \u_multiplier/STAGE1/_2403_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/STAGE1/_1095_ ));
 AND2_X1 \u_multiplier/STAGE1/_2404_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/STAGE1/_1096_ ));
 AND2_X1 \u_multiplier/STAGE1/_2405_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/STAGE1/_1097_ ));
 AND2_X1 \u_multiplier/STAGE1/_2406_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[27]),
    .ZN(\u_multiplier/STAGE1/_1098_ ));
 AND2_X1 \u_multiplier/STAGE1/_2407_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[26]),
    .ZN(\u_multiplier/STAGE1/_1099_ ));
 AND2_X1 \u_multiplier/STAGE1/_2408_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[25]),
    .ZN(\u_multiplier/STAGE1/_1100_ ));
 AND2_X1 \u_multiplier/STAGE1/_2409_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[24]),
    .ZN(\u_multiplier/STAGE1/_1101_ ));
 AND2_X1 \u_multiplier/STAGE1/_2410_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[23]),
    .ZN(\u_multiplier/STAGE1/_1102_ ));
 AND2_X1 \u_multiplier/STAGE1/_2411_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[22]),
    .ZN(\u_multiplier/STAGE1/_1103_ ));
 AND2_X1 \u_multiplier/STAGE1/_2412_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[21]),
    .ZN(\u_multiplier/STAGE1/_1104_ ));
 AND2_X1 \u_multiplier/STAGE1/_2413_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[21]),
    .ZN(\u_multiplier/STAGE1/_1105_ ));
 AND2_X1 \u_multiplier/STAGE1/_2414_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[22]),
    .ZN(\u_multiplier/STAGE1/_1106_ ));
 AND2_X1 \u_multiplier/STAGE1/_2415_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[23]),
    .ZN(\u_multiplier/STAGE1/_1107_ ));
 AND2_X1 \u_multiplier/STAGE1/_2416_  (.A1(sram_rdata_reg[10]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp1_41 [8]));
 AND2_X1 \u_multiplier/STAGE1/_2417_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/pp1_41 [9]));
 AND2_X1 \u_multiplier/STAGE1/_2418_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/pp1_41 [10]));
 AND2_X1 \u_multiplier/STAGE1/_2419_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/pp1_41 [11]));
 AND2_X1 \u_multiplier/STAGE1/_2420_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/pp1_41 [12]));
 AND2_X1 \u_multiplier/STAGE1/_2421_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[26]),
    .ZN(\u_multiplier/pp1_41 [13]));
 AND2_X1 \u_multiplier/STAGE1/_2422_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[25]),
    .ZN(\u_multiplier/pp1_41 [14]));
 AND2_X1 \u_multiplier/STAGE1/_2423_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[24]),
    .ZN(\u_multiplier/pp1_41 [15]));
 AND2_X1 \u_multiplier/STAGE1/_2424_  (.A1(data_in_reg[11]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/STAGE1/_1108_ ));
 AND2_X1 \u_multiplier/STAGE1/_2425_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/STAGE1/_1109_ ));
 AND2_X1 \u_multiplier/STAGE1/_2426_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/STAGE1/_1110_ ));
 AND2_X1 \u_multiplier/STAGE1/_2427_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/STAGE1/_1111_ ));
 AND2_X1 \u_multiplier/STAGE1/_2428_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[27]),
    .ZN(\u_multiplier/STAGE1/_1112_ ));
 AND2_X1 \u_multiplier/STAGE1/_2429_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[26]),
    .ZN(\u_multiplier/STAGE1/_1113_ ));
 AND2_X1 \u_multiplier/STAGE1/_2430_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[25]),
    .ZN(\u_multiplier/STAGE1/_1114_ ));
 AND2_X1 \u_multiplier/STAGE1/_2431_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[24]),
    .ZN(\u_multiplier/STAGE1/_1115_ ));
 AND2_X1 \u_multiplier/STAGE1/_2432_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[23]),
    .ZN(\u_multiplier/STAGE1/_1116_ ));
 AND2_X1 \u_multiplier/STAGE1/_2433_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[22]),
    .ZN(\u_multiplier/STAGE1/_1117_ ));
 AND2_X1 \u_multiplier/STAGE1/_2434_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[21]),
    .ZN(\u_multiplier/STAGE1/_1118_ ));
 AND2_X1 \u_multiplier/STAGE1/_2435_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[22]),
    .ZN(\u_multiplier/STAGE1/_1119_ ));
 AND2_X1 \u_multiplier/STAGE1/_2436_  (.A1(sram_rdata_reg[11]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp1_42 [7]));
 AND2_X1 \u_multiplier/STAGE1/_2437_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/pp1_42 [8]));
 AND2_X1 \u_multiplier/STAGE1/_2438_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/pp1_42 [9]));
 AND2_X1 \u_multiplier/STAGE1/_2439_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/pp1_42 [10]));
 AND2_X1 \u_multiplier/STAGE1/_2440_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/pp1_42 [11]));
 AND2_X1 \u_multiplier/STAGE1/_2441_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[26]),
    .ZN(\u_multiplier/pp1_42 [12]));
 AND2_X1 \u_multiplier/STAGE1/_2442_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[25]),
    .ZN(\u_multiplier/pp1_42 [13]));
 AND2_X1 \u_multiplier/STAGE1/_2443_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[24]),
    .ZN(\u_multiplier/pp1_42 [14]));
 AND2_X1 \u_multiplier/STAGE1/_2444_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[23]),
    .ZN(\u_multiplier/pp1_42 [15]));
 AND2_X1 \u_multiplier/STAGE1/_2445_  (.A1(data_in_reg[12]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/STAGE1/_1120_ ));
 AND2_X1 \u_multiplier/STAGE1/_2446_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/STAGE1/_1121_ ));
 AND2_X1 \u_multiplier/STAGE1/_2447_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/STAGE1/_1122_ ));
 AND2_X1 \u_multiplier/STAGE1/_2448_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/STAGE1/_1123_ ));
 AND2_X1 \u_multiplier/STAGE1/_2449_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[27]),
    .ZN(\u_multiplier/STAGE1/_1124_ ));
 AND2_X1 \u_multiplier/STAGE1/_2450_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[26]),
    .ZN(\u_multiplier/STAGE1/_1125_ ));
 AND2_X1 \u_multiplier/STAGE1/_2451_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[25]),
    .ZN(\u_multiplier/STAGE1/_1126_ ));
 AND2_X1 \u_multiplier/STAGE1/_2452_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[24]),
    .ZN(\u_multiplier/STAGE1/_1127_ ));
 AND2_X1 \u_multiplier/STAGE1/_2453_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[23]),
    .ZN(\u_multiplier/STAGE1/_1128_ ));
 AND2_X1 \u_multiplier/STAGE1/_2454_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[22]),
    .ZN(\u_multiplier/STAGE1/_1129_ ));
 AND2_X1 \u_multiplier/STAGE1/_2455_  (.A1(sram_rdata_reg[12]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp1_43 [6]));
 AND2_X1 \u_multiplier/STAGE1/_2456_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/pp1_43 [7]));
 AND2_X1 \u_multiplier/STAGE1/_2457_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/pp1_43 [8]));
 AND2_X1 \u_multiplier/STAGE1/_2458_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/pp1_43 [9]));
 AND2_X1 \u_multiplier/STAGE1/_2459_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/pp1_43 [10]));
 AND2_X1 \u_multiplier/STAGE1/_2460_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[26]),
    .ZN(\u_multiplier/pp1_43 [11]));
 AND2_X1 \u_multiplier/STAGE1/_2461_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[25]),
    .ZN(\u_multiplier/pp1_43 [12]));
 AND2_X1 \u_multiplier/STAGE1/_2462_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[24]),
    .ZN(\u_multiplier/pp1_43 [13]));
 AND2_X1 \u_multiplier/STAGE1/_2463_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[23]),
    .ZN(\u_multiplier/pp1_43 [14]));
 AND2_X1 \u_multiplier/STAGE1/_2464_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[22]),
    .ZN(\u_multiplier/pp1_43 [15]));
 AND2_X1 \u_multiplier/STAGE1/_2465_  (.A1(data_in_reg[13]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/STAGE1/_1130_ ));
 AND2_X1 \u_multiplier/STAGE1/_2466_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/STAGE1/_1131_ ));
 AND2_X1 \u_multiplier/STAGE1/_2467_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/STAGE1/_1132_ ));
 AND2_X1 \u_multiplier/STAGE1/_2468_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/STAGE1/_1133_ ));
 AND2_X1 \u_multiplier/STAGE1/_2469_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[27]),
    .ZN(\u_multiplier/STAGE1/_1134_ ));
 AND2_X1 \u_multiplier/STAGE1/_2470_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[26]),
    .ZN(\u_multiplier/STAGE1/_1135_ ));
 AND2_X1 \u_multiplier/STAGE1/_2471_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[25]),
    .ZN(\u_multiplier/STAGE1/_1136_ ));
 AND2_X1 \u_multiplier/STAGE1/_2472_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[24]),
    .ZN(\u_multiplier/STAGE1/_1137_ ));
 AND2_X1 \u_multiplier/STAGE1/_2473_  (.A1(sram_rdata_reg[13]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp1_44 [5]));
 AND2_X1 \u_multiplier/STAGE1/_2474_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/pp1_44 [6]));
 AND2_X1 \u_multiplier/STAGE1/_2475_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/pp1_44 [7]));
 AND2_X1 \u_multiplier/STAGE1/_2476_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/pp1_44 [8]));
 AND2_X1 \u_multiplier/STAGE1/_2477_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/pp1_44 [9]));
 AND2_X1 \u_multiplier/STAGE1/_2478_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[26]),
    .ZN(\u_multiplier/pp1_44 [10]));
 AND2_X1 \u_multiplier/STAGE1/_2479_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[25]),
    .ZN(\u_multiplier/pp1_44 [11]));
 AND2_X1 \u_multiplier/STAGE1/_2480_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[24]),
    .ZN(\u_multiplier/pp1_44 [12]));
 AND2_X1 \u_multiplier/STAGE1/_2481_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[23]),
    .ZN(\u_multiplier/pp1_44 [13]));
 AND2_X1 \u_multiplier/STAGE1/_2482_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[22]),
    .ZN(\u_multiplier/pp1_44 [14]));
 AND2_X1 \u_multiplier/STAGE1/_2483_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[23]),
    .ZN(\u_multiplier/pp1_44 [15]));
 AND2_X1 \u_multiplier/STAGE1/_2484_  (.A1(data_in_reg[14]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/STAGE1/_1138_ ));
 AND2_X1 \u_multiplier/STAGE1/_2485_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/STAGE1/_1139_ ));
 AND2_X1 \u_multiplier/STAGE1/_2486_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/STAGE1/_1140_ ));
 AND2_X1 \u_multiplier/STAGE1/_2487_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/STAGE1/_1141_ ));
 AND2_X1 \u_multiplier/STAGE1/_2488_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[27]),
    .ZN(\u_multiplier/STAGE1/_1142_ ));
 AND2_X1 \u_multiplier/STAGE1/_2489_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[26]),
    .ZN(\u_multiplier/STAGE1/_1143_ ));
 AND2_X1 \u_multiplier/STAGE1/_2490_  (.A1(sram_rdata_reg[14]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp1_45 [4]));
 AND2_X1 \u_multiplier/STAGE1/_2491_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/pp1_45 [5]));
 AND2_X1 \u_multiplier/STAGE1/_2492_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/pp1_45 [6]));
 AND2_X1 \u_multiplier/STAGE1/_2493_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/pp1_45 [7]));
 AND2_X1 \u_multiplier/STAGE1/_2494_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/pp1_45 [8]));
 AND2_X1 \u_multiplier/STAGE1/_2495_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[26]),
    .ZN(\u_multiplier/pp1_45 [9]));
 AND2_X1 \u_multiplier/STAGE1/_2496_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[25]),
    .ZN(\u_multiplier/pp1_45 [10]));
 AND2_X1 \u_multiplier/STAGE1/_2497_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[24]),
    .ZN(\u_multiplier/pp1_45 [11]));
 AND2_X1 \u_multiplier/STAGE1/_2498_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[23]),
    .ZN(\u_multiplier/pp1_45 [12]));
 AND2_X1 \u_multiplier/STAGE1/_2499_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[23]),
    .ZN(\u_multiplier/pp1_45 [13]));
 AND2_X1 \u_multiplier/STAGE1/_2500_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[24]),
    .ZN(\u_multiplier/pp1_45 [14]));
 AND2_X1 \u_multiplier/STAGE1/_2501_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[25]),
    .ZN(\u_multiplier/pp1_45 [15]));
 AND2_X1 \u_multiplier/STAGE1/_2502_  (.A1(data_in_reg[15]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/STAGE1/_1144_ ));
 AND2_X1 \u_multiplier/STAGE1/_2503_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/STAGE1/_1145_ ));
 AND2_X1 \u_multiplier/STAGE1/_2504_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/STAGE1/_1146_ ));
 AND2_X1 \u_multiplier/STAGE1/_2505_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/STAGE1/_1147_ ));
 AND2_X1 \u_multiplier/STAGE1/_2506_  (.A1(sram_rdata_reg[15]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp1_46 [3]));
 AND2_X1 \u_multiplier/STAGE1/_2507_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/pp1_46 [4]));
 AND2_X1 \u_multiplier/STAGE1/_2508_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/pp1_46 [5]));
 AND2_X1 \u_multiplier/STAGE1/_2509_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/pp1_46 [6]));
 AND2_X1 \u_multiplier/STAGE1/_2510_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/pp1_46 [7]));
 AND2_X1 \u_multiplier/STAGE1/_2511_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[26]),
    .ZN(\u_multiplier/pp1_46 [8]));
 AND2_X1 \u_multiplier/STAGE1/_2512_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[25]),
    .ZN(\u_multiplier/pp1_46 [9]));
 AND2_X1 \u_multiplier/STAGE1/_2513_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[24]),
    .ZN(\u_multiplier/pp1_46 [10]));
 AND2_X1 \u_multiplier/STAGE1/_2514_  (.A1(sram_rdata_reg[23]),
    .A2(data_in_reg[23]),
    .ZN(\u_multiplier/pp1_46 [11]));
 AND2_X1 \u_multiplier/STAGE1/_2515_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[24]),
    .ZN(\u_multiplier/pp1_46 [12]));
 AND2_X1 \u_multiplier/STAGE1/_2516_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[25]),
    .ZN(\u_multiplier/pp1_46 [13]));
 AND2_X1 \u_multiplier/STAGE1/_2517_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[26]),
    .ZN(\u_multiplier/pp1_46 [14]));
 AND2_X1 \u_multiplier/STAGE1/_2518_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[27]),
    .ZN(\u_multiplier/pp1_46 [15]));
 AND2_X1 \u_multiplier/STAGE1/_2519_  (.A1(data_in_reg[16]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/STAGE1/_1148_ ));
 AND2_X1 \u_multiplier/STAGE1/_2520_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/STAGE1/_1149_ ));
 AND2_X1 \u_multiplier/STAGE1/_2521_  (.A1(sram_rdata_reg[16]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp1_47 [2]));
 AND2_X1 \u_multiplier/STAGE1/_2522_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/pp1_47 [3]));
 AND2_X1 \u_multiplier/STAGE1/_2523_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/pp1_47 [4]));
 AND2_X1 \u_multiplier/STAGE1/_2524_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/pp1_47 [5]));
 AND2_X1 \u_multiplier/STAGE1/_2525_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/pp1_47 [6]));
 AND2_X1 \u_multiplier/STAGE1/_2526_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[26]),
    .ZN(\u_multiplier/pp1_47 [7]));
 AND2_X1 \u_multiplier/STAGE1/_2527_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[25]),
    .ZN(\u_multiplier/pp1_47 [8]));
 AND2_X1 \u_multiplier/STAGE1/_2528_  (.A1(sram_rdata_reg[23]),
    .A2(data_in_reg[24]),
    .ZN(\u_multiplier/pp1_47 [9]));
 AND2_X1 \u_multiplier/STAGE1/_2529_  (.A1(data_in_reg[23]),
    .A2(sram_rdata_reg[24]),
    .ZN(\u_multiplier/pp1_47 [10]));
 AND2_X1 \u_multiplier/STAGE1/_2530_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[25]),
    .ZN(\u_multiplier/pp1_47 [11]));
 AND2_X1 \u_multiplier/STAGE1/_2531_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[26]),
    .ZN(\u_multiplier/pp1_47 [12]));
 AND2_X1 \u_multiplier/STAGE1/_2532_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[27]),
    .ZN(\u_multiplier/pp1_47 [13]));
 AND2_X1 \u_multiplier/STAGE1/_2533_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/pp1_47 [14]));
 AND2_X1 \u_multiplier/STAGE1/_2534_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/pp1_47 [15]));
 AND2_X1 \u_multiplier/STAGE1/_2535_  (.A1(sram_rdata_reg[17]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp1_48 [1]));
 AND2_X1 \u_multiplier/STAGE1/_2536_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/pp1_48 [2]));
 AND2_X1 \u_multiplier/STAGE1/_2537_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/pp1_48 [3]));
 AND2_X1 \u_multiplier/STAGE1/_2538_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/pp1_48 [4]));
 AND2_X1 \u_multiplier/STAGE1/_2539_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/pp1_48 [5]));
 AND2_X1 \u_multiplier/STAGE1/_2540_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[26]),
    .ZN(\u_multiplier/pp1_48 [6]));
 AND2_X1 \u_multiplier/STAGE1/_2541_  (.A1(sram_rdata_reg[23]),
    .A2(data_in_reg[25]),
    .ZN(\u_multiplier/pp1_48 [7]));
 AND2_X1 \u_multiplier/STAGE1/_2542_  (.A1(sram_rdata_reg[24]),
    .A2(data_in_reg[24]),
    .ZN(\u_multiplier/pp1_48 [8]));
 AND2_X1 \u_multiplier/STAGE1/_2543_  (.A1(data_in_reg[23]),
    .A2(sram_rdata_reg[25]),
    .ZN(\u_multiplier/pp1_48 [9]));
 AND2_X1 \u_multiplier/STAGE1/_2544_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[26]),
    .ZN(\u_multiplier/pp1_48 [10]));
 AND2_X1 \u_multiplier/STAGE1/_2545_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[27]),
    .ZN(\u_multiplier/pp1_48 [11]));
 AND2_X1 \u_multiplier/STAGE1/_2546_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/pp1_48 [12]));
 AND2_X1 \u_multiplier/STAGE1/_2547_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/pp1_48 [13]));
 AND2_X1 \u_multiplier/STAGE1/_2548_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/pp1_48 [14]));
 AND2_X1 \u_multiplier/STAGE1/_2549_  (.A1(data_in_reg[17]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/pp1_48 [15]));
 AND2_X1 \u_multiplier/STAGE1/_2550_  (.A1(sram_rdata_reg[18]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp1_49 [0]));
 AND2_X1 \u_multiplier/STAGE1/_2551_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/pp1_49 [1]));
 AND2_X1 \u_multiplier/STAGE1/_2552_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/pp1_49 [2]));
 AND2_X1 \u_multiplier/STAGE1/_2553_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/pp1_49 [3]));
 AND2_X1 \u_multiplier/STAGE1/_2554_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/pp1_49 [4]));
 AND2_X1 \u_multiplier/STAGE1/_2555_  (.A1(sram_rdata_reg[23]),
    .A2(data_in_reg[26]),
    .ZN(\u_multiplier/pp1_49 [5]));
 AND2_X1 \u_multiplier/STAGE1/_2556_  (.A1(sram_rdata_reg[24]),
    .A2(data_in_reg[25]),
    .ZN(\u_multiplier/pp1_49 [6]));
 AND2_X1 \u_multiplier/STAGE1/_2557_  (.A1(data_in_reg[24]),
    .A2(sram_rdata_reg[25]),
    .ZN(\u_multiplier/pp1_49 [7]));
 AND2_X1 \u_multiplier/STAGE1/_2558_  (.A1(data_in_reg[23]),
    .A2(sram_rdata_reg[26]),
    .ZN(\u_multiplier/pp1_49 [8]));
 AND2_X1 \u_multiplier/STAGE1/_2559_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[27]),
    .ZN(\u_multiplier/pp1_49 [9]));
 AND2_X1 \u_multiplier/STAGE1/_2560_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/pp1_49 [10]));
 AND2_X1 \u_multiplier/STAGE1/_2561_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/pp1_49 [11]));
 AND2_X1 \u_multiplier/STAGE1/_2562_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/pp1_49 [12]));
 AND2_X1 \u_multiplier/STAGE1/_2563_  (.A1(data_in_reg[18]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/pp1_49 [13]));
 AND2_X1 \u_multiplier/STAGE1/_2564_  (.A1(sram_rdata_reg[19]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp1_50 [0]));
 AND2_X1 \u_multiplier/STAGE1/_2565_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/pp1_50 [1]));
 AND2_X1 \u_multiplier/STAGE1/_2566_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/pp1_50 [2]));
 AND2_X1 \u_multiplier/STAGE1/_2567_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/pp1_50 [3]));
 AND2_X1 \u_multiplier/STAGE1/_2568_  (.A1(sram_rdata_reg[23]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/pp1_50 [4]));
 AND2_X1 \u_multiplier/STAGE1/_2569_  (.A1(sram_rdata_reg[24]),
    .A2(data_in_reg[26]),
    .ZN(\u_multiplier/pp1_50 [5]));
 AND2_X1 \u_multiplier/STAGE1/_2570_  (.A1(sram_rdata_reg[25]),
    .A2(data_in_reg[25]),
    .ZN(\u_multiplier/pp1_50 [6]));
 AND2_X1 \u_multiplier/STAGE1/_2571_  (.A1(data_in_reg[24]),
    .A2(sram_rdata_reg[26]),
    .ZN(\u_multiplier/pp1_50 [7]));
 AND2_X1 \u_multiplier/STAGE1/_2572_  (.A1(data_in_reg[23]),
    .A2(sram_rdata_reg[27]),
    .ZN(\u_multiplier/pp1_50 [8]));
 AND2_X1 \u_multiplier/STAGE1/_2573_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/pp1_50 [9]));
 AND2_X1 \u_multiplier/STAGE1/_2574_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/pp1_50 [10]));
 AND2_X1 \u_multiplier/STAGE1/_2575_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/pp1_50 [11]));
 AND2_X1 \u_multiplier/STAGE1/_2576_  (.A1(data_in_reg[19]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/pp2_50 [7]));
 AND2_X1 \u_multiplier/STAGE1/_2577_  (.A1(sram_rdata_reg[20]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp1_51 [0]));
 AND2_X1 \u_multiplier/STAGE1/_2578_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/pp1_51 [1]));
 AND2_X1 \u_multiplier/STAGE1/_2579_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/pp1_51 [2]));
 AND2_X1 \u_multiplier/STAGE1/_2580_  (.A1(sram_rdata_reg[23]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/pp1_51 [3]));
 AND2_X1 \u_multiplier/STAGE1/_2581_  (.A1(sram_rdata_reg[24]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/pp1_51 [4]));
 AND2_X1 \u_multiplier/STAGE1/_2582_  (.A1(sram_rdata_reg[25]),
    .A2(data_in_reg[26]),
    .ZN(\u_multiplier/pp1_51 [5]));
 AND2_X1 \u_multiplier/STAGE1/_2583_  (.A1(data_in_reg[25]),
    .A2(sram_rdata_reg[26]),
    .ZN(\u_multiplier/pp1_51 [6]));
 AND2_X1 \u_multiplier/STAGE1/_2584_  (.A1(data_in_reg[24]),
    .A2(sram_rdata_reg[27]),
    .ZN(\u_multiplier/pp1_51 [7]));
 AND2_X2 \u_multiplier/STAGE1/_2585_  (.A1(data_in_reg[23]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/pp1_51 [8]));
 AND2_X2 \u_multiplier/STAGE1/_2586_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/pp1_51 [9]));
 AND2_X1 \u_multiplier/STAGE1/_2587_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/pp2_51 [7]));
 AND2_X1 \u_multiplier/STAGE1/_2588_  (.A1(data_in_reg[20]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/pp2_51 [6]));
 AND2_X1 \u_multiplier/STAGE1/_2589_  (.A1(sram_rdata_reg[21]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp1_52 [0]));
 AND2_X1 \u_multiplier/STAGE1/_2590_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/pp1_52 [1]));
 AND2_X1 \u_multiplier/STAGE1/_2591_  (.A1(sram_rdata_reg[23]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/pp1_52 [2]));
 AND2_X1 \u_multiplier/STAGE1/_2592_  (.A1(sram_rdata_reg[24]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/pp1_52 [3]));
 AND2_X1 \u_multiplier/STAGE1/_2593_  (.A1(sram_rdata_reg[25]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/pp1_52 [4]));
 AND2_X1 \u_multiplier/STAGE1/_2594_  (.A1(sram_rdata_reg[26]),
    .A2(data_in_reg[26]),
    .ZN(\u_multiplier/pp1_52 [5]));
 AND2_X1 \u_multiplier/STAGE1/_2595_  (.A1(data_in_reg[25]),
    .A2(sram_rdata_reg[27]),
    .ZN(\u_multiplier/pp1_52 [6]));
 AND2_X1 \u_multiplier/STAGE1/_2596_  (.A1(data_in_reg[24]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/pp1_52 [7]));
 AND2_X1 \u_multiplier/STAGE1/_2597_  (.A1(data_in_reg[23]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/pp2_52 [7]));
 AND2_X1 \u_multiplier/STAGE1/_2598_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/pp2_52 [6]));
 AND2_X1 \u_multiplier/STAGE1/_2599_  (.A1(data_in_reg[21]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/pp2_52 [5]));
 AND2_X1 \u_multiplier/STAGE1/_2600_  (.A1(sram_rdata_reg[22]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp1_53 [0]));
 AND2_X1 \u_multiplier/STAGE1/_2601_  (.A1(sram_rdata_reg[23]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/pp1_53 [1]));
 AND2_X1 \u_multiplier/STAGE1/_2602_  (.A1(sram_rdata_reg[24]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/pp1_53 [2]));
 AND2_X1 \u_multiplier/STAGE1/_2603_  (.A1(sram_rdata_reg[25]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/pp1_53 [3]));
 AND2_X1 \u_multiplier/STAGE1/_2604_  (.A1(sram_rdata_reg[26]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/pp1_53 [4]));
 AND2_X1 \u_multiplier/STAGE1/_2605_  (.A1(data_in_reg[26]),
    .A2(sram_rdata_reg[27]),
    .ZN(\u_multiplier/pp1_53 [5]));
 AND2_X1 \u_multiplier/STAGE1/_2606_  (.A1(data_in_reg[25]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/pp2_53 [7]));
 AND2_X1 \u_multiplier/STAGE1/_2607_  (.A1(data_in_reg[24]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/pp2_53 [6]));
 AND2_X1 \u_multiplier/STAGE1/_2608_  (.A1(data_in_reg[23]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/pp2_53 [5]));
 AND2_X1 \u_multiplier/STAGE1/_2609_  (.A1(data_in_reg[22]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/pp2_53 [4]));
 AND2_X1 \u_multiplier/STAGE1/_2610_  (.A1(sram_rdata_reg[23]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp1_54 [0]));
 AND2_X1 \u_multiplier/STAGE1/_2611_  (.A1(sram_rdata_reg[24]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/pp1_54 [1]));
 AND2_X1 \u_multiplier/STAGE1/_2612_  (.A1(sram_rdata_reg[25]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/pp1_54 [2]));
 AND2_X1 \u_multiplier/STAGE1/_2613_  (.A1(sram_rdata_reg[26]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/pp1_54 [3]));
 AND2_X1 \u_multiplier/STAGE1/_2614_  (.A1(sram_rdata_reg[27]),
    .A2(data_in_reg[27]),
    .ZN(\u_multiplier/pp2_54 [7]));
 AND2_X1 \u_multiplier/STAGE1/_2615_  (.A1(data_in_reg[26]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/pp2_54 [6]));
 AND2_X1 \u_multiplier/STAGE1/_2616_  (.A1(data_in_reg[25]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/pp2_54 [5]));
 AND2_X1 \u_multiplier/STAGE1/_2617_  (.A1(data_in_reg[24]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/pp2_54 [4]));
 AND2_X1 \u_multiplier/STAGE1/_2618_  (.A1(data_in_reg[23]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/pp2_54 [3]));
 AND2_X1 \u_multiplier/STAGE1/_2619_  (.A1(sram_rdata_reg[24]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp1_55 [0]));
 AND2_X1 \u_multiplier/STAGE1/_2620_  (.A1(sram_rdata_reg[25]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/pp1_55 [1]));
 AND2_X1 \u_multiplier/STAGE1/_2621_  (.A1(sram_rdata_reg[26]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/pp2_55 [7]));
 AND2_X1 \u_multiplier/STAGE1/_2622_  (.A1(sram_rdata_reg[27]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/pp2_55 [6]));
 AND2_X1 \u_multiplier/STAGE1/_2623_  (.A1(data_in_reg[27]),
    .A2(sram_rdata_reg[28]),
    .ZN(\u_multiplier/pp2_55 [5]));
 AND2_X1 \u_multiplier/STAGE1/_2624_  (.A1(data_in_reg[26]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/pp2_55 [4]));
 AND2_X1 \u_multiplier/STAGE1/_2625_  (.A1(data_in_reg[25]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/pp2_55 [3]));
 AND2_X1 \u_multiplier/STAGE1/_2626_  (.A1(data_in_reg[24]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/pp2_55 [2]));
 AND2_X1 \u_multiplier/STAGE1/_2627_  (.A1(sram_rdata_reg[25]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp2_56 [7]));
 AND2_X1 \u_multiplier/STAGE1/_2628_  (.A1(sram_rdata_reg[26]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/pp2_56 [6]));
 AND2_X1 \u_multiplier/STAGE1/_2629_  (.A1(sram_rdata_reg[27]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/pp2_56 [5]));
 AND2_X1 \u_multiplier/STAGE1/_2630_  (.A1(sram_rdata_reg[28]),
    .A2(data_in_reg[28]),
    .ZN(\u_multiplier/pp2_56 [4]));
 AND2_X1 \u_multiplier/STAGE1/_2631_  (.A1(data_in_reg[27]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/pp2_56 [3]));
 AND2_X1 \u_multiplier/STAGE1/_2632_  (.A1(data_in_reg[26]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/pp2_56 [2]));
 AND2_X1 \u_multiplier/STAGE1/_2633_  (.A1(data_in_reg[25]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/pp2_56 [1]));
 AND2_X1 \u_multiplier/STAGE1/_2634_  (.A1(sram_rdata_reg[26]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp2_57 [5]));
 AND2_X1 \u_multiplier/STAGE1/_2635_  (.A1(sram_rdata_reg[27]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/pp2_57 [4]));
 AND2_X1 \u_multiplier/STAGE1/_2636_  (.A1(sram_rdata_reg[28]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/pp2_57 [3]));
 AND2_X1 \u_multiplier/STAGE1/_2637_  (.A1(data_in_reg[28]),
    .A2(sram_rdata_reg[29]),
    .ZN(\u_multiplier/pp2_57 [2]));
 AND2_X1 \u_multiplier/STAGE1/_2638_  (.A1(data_in_reg[27]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/pp2_57 [1]));
 AND2_X1 \u_multiplier/STAGE1/_2639_  (.A1(data_in_reg[26]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/pp2_57 [0]));
 AND2_X1 \u_multiplier/STAGE1/_2640_  (.A1(sram_rdata_reg[27]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp3_58 [3]));
 AND2_X1 \u_multiplier/STAGE1/_2641_  (.A1(sram_rdata_reg[28]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/pp2_58 [3]));
 AND2_X1 \u_multiplier/STAGE1/_2642_  (.A1(sram_rdata_reg[29]),
    .A2(data_in_reg[29]),
    .ZN(\u_multiplier/pp2_58 [2]));
 AND2_X1 \u_multiplier/STAGE1/_2643_  (.A1(data_in_reg[28]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/pp2_58 [1]));
 AND2_X1 \u_multiplier/STAGE1/_2644_  (.A1(data_in_reg[27]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/pp2_58 [0]));
 AND2_X1 \u_multiplier/STAGE1/_2645_  (.A1(sram_rdata_reg[28]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp3_59 [2]));
 AND2_X1 \u_multiplier/STAGE1/_2646_  (.A1(sram_rdata_reg[29]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/pp3_59 [3]));
 AND2_X1 \u_multiplier/STAGE1/_2647_  (.A1(data_in_reg[29]),
    .A2(sram_rdata_reg[30]),
    .ZN(\u_multiplier/pp2_59 [1]));
 AND2_X1 \u_multiplier/STAGE1/_2648_  (.A1(data_in_reg[28]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/pp2_59 [0]));
 AND2_X1 \u_multiplier/STAGE1/_2649_  (.A1(sram_rdata_reg[29]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp3_60 [1]));
 AND2_X1 \u_multiplier/STAGE1/_2650_  (.A1(sram_rdata_reg[30]),
    .A2(data_in_reg[30]),
    .ZN(\u_multiplier/pp3_60 [2]));
 AND2_X1 \u_multiplier/STAGE1/_2651_  (.A1(data_in_reg[29]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/pp3_60 [3]));
 AND2_X1 \u_multiplier/STAGE1/_2652_  (.A1(sram_rdata_reg[30]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp3_61 [0]));
 AND2_X1 \u_multiplier/STAGE1/_2653_  (.A1(data_in_reg[30]),
    .A2(sram_rdata_reg[31]),
    .ZN(\u_multiplier/pp3_61 [1]));
 AND2_X1 \u_multiplier/STAGE1/_2654_  (.A1(sram_rdata_reg[31]),
    .A2(data_in_reg[31]),
    .ZN(\u_multiplier/pp3_62 ));
 LOGIC0_X1 \u_multiplier/STAGE2/E_4_2_pp2_11_2/_25__133  (.Z(net133));
 LOGIC0_X1 \u_multiplier/STAGE2/E_4_2_pp2_11_2/_18__132  (.Z(net132));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_10_1/_18_  (.A(\u_multiplier/STAGE2/pp2_9_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_10_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_10_1/_19_  (.A1(\u_multiplier/pp1_10 [1]),
    .A2(\u_multiplier/pp1_10 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_10_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_10_1/_20_  (.A(\u_multiplier/pp1_10 [1]),
    .B(\u_multiplier/pp1_10 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_10_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_10_1/_21_  (.A1(\u_multiplier/pp1_10 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_10_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_10_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_10_1/_22_  (.A(\u_multiplier/pp1_10 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_10_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_10_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_10_1/_23_  (.A1(\u_multiplier/pp1_10 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_10_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_10_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_10_1/_24_  (.A(\u_multiplier/pp1_10 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_10_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_10_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_10_1/_25_  (.A(\u_multiplier/STAGE2/pp2_9_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_10_1/_16_ ),
    .ZN(\u_multiplier/pp2_10 [1]));
 NAND2_X2 \u_multiplier/STAGE2/E_4_2_pp2_10_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_10_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_10_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_10_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_10_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_10_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_10_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_10_1/_17_ ),
    .ZN(\u_multiplier/pp2_11 [3]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_11_1/_18_  (.A(\u_multiplier/STAGE2/pp2_10_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_11_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_11_1/_19_  (.A1(\u_multiplier/pp1_11 [1]),
    .A2(\u_multiplier/pp1_11 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_11_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_11_1/_20_  (.A(\u_multiplier/pp1_11 [1]),
    .B(\u_multiplier/pp1_11 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_11_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_11_1/_21_  (.A1(\u_multiplier/pp1_11 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_11_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_11_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_11_1/_22_  (.A(\u_multiplier/pp1_11 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_11_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_11_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_11_1/_23_  (.A1(\u_multiplier/pp1_11 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_11_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_11_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_11_1/_24_  (.A(\u_multiplier/pp1_11 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_11_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_11_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_11_1/_25_  (.A(\u_multiplier/STAGE2/pp2_10_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_11_1/_16_ ),
    .ZN(\u_multiplier/pp2_11 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_11_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_11_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_11_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_11_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_11_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_11_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_11_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_11_1/_17_ ),
    .ZN(\u_multiplier/pp2_12 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_11_2/_18_  (.A(net132),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_11_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_11_2/_19_  (.A1(\u_multiplier/pp1_11 [5]),
    .A2(\u_multiplier/pp1_11 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_11_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_11_2/_20_  (.A(\u_multiplier/pp1_11 [5]),
    .B(\u_multiplier/pp1_11 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_11_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_11_2/_21_  (.A1(\u_multiplier/pp1_11 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_11_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_11_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_11_2/_22_  (.A(\u_multiplier/pp1_11 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_11_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_11_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_11_2/_23_  (.A1(\u_multiplier/pp1_11 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_11_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_11_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_11_2/_24_  (.A(\u_multiplier/pp1_11 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_11_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_11_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_11_2/_25_  (.A(net133),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_11_2/_16_ ),
    .ZN(\u_multiplier/pp2_11 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_11_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_11_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_11_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_11_e42_2_cout ));
 OAI21_X1 \u_multiplier/STAGE2/E_4_2_pp2_11_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_11_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_11_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_11_2/_17_ ),
    .ZN(\u_multiplier/pp2_12 [3]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_12_1/_18_  (.A(\u_multiplier/STAGE2/pp2_11_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_12_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_12_1/_19_  (.A1(\u_multiplier/pp1_12 [1]),
    .A2(\u_multiplier/pp1_12 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_12_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_12_1/_20_  (.A(\u_multiplier/pp1_12 [1]),
    .B(\u_multiplier/pp1_12 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_12_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_12_1/_21_  (.A1(\u_multiplier/pp1_12 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_12_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_12_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_12_1/_22_  (.A(\u_multiplier/pp1_12 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_12_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_12_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_12_1/_23_  (.A1(\u_multiplier/pp1_12 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_12_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_12_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_12_1/_24_  (.A(\u_multiplier/pp1_12 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_12_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_12_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_12_1/_25_  (.A(\u_multiplier/STAGE2/pp2_11_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_12_1/_16_ ),
    .ZN(\u_multiplier/pp2_12 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_12_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_12_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_12_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_12_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_12_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_12_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_12_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_12_1/_17_ ),
    .ZN(\u_multiplier/pp2_13 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_12_2/_18_  (.A(\u_multiplier/STAGE2/pp2_11_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_12_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_12_2/_19_  (.A1(\u_multiplier/pp1_12 [5]),
    .A2(\u_multiplier/pp1_12 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_12_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_12_2/_20_  (.A(\u_multiplier/pp1_12 [5]),
    .B(\u_multiplier/pp1_12 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_12_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_12_2/_21_  (.A1(\u_multiplier/pp1_12 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_12_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_12_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_12_2/_22_  (.A(\u_multiplier/pp1_12 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_12_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_12_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_12_2/_23_  (.A1(\u_multiplier/pp1_12 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_12_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_12_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_12_2/_24_  (.A(\u_multiplier/pp1_12 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_12_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_12_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_12_2/_25_  (.A(\u_multiplier/STAGE2/pp2_11_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_12_2/_16_ ),
    .ZN(\u_multiplier/pp2_12 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_12_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_12_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_12_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_12_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_12_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_12_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_12_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_12_2/_17_ ),
    .ZN(\u_multiplier/pp2_13 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_13_1/_18_  (.A(\u_multiplier/STAGE2/pp2_12_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_13_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_13_1/_19_  (.A1(\u_multiplier/pp1_13 [1]),
    .A2(\u_multiplier/pp1_13 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_13_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_13_1/_20_  (.A(\u_multiplier/pp1_13 [1]),
    .B(\u_multiplier/pp1_13 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_13_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_13_1/_21_  (.A1(\u_multiplier/pp1_13 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_13_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_13_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_13_1/_22_  (.A(\u_multiplier/pp1_13 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_13_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_13_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_13_1/_23_  (.A1(\u_multiplier/pp1_13 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_13_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_13_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_13_1/_24_  (.A(\u_multiplier/pp1_13 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_13_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_13_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_13_1/_25_  (.A(\u_multiplier/STAGE2/pp2_12_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_13_1/_16_ ),
    .ZN(\u_multiplier/pp2_13 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_13_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_13_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_13_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_13_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_13_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_13_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_13_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_13_1/_17_ ),
    .ZN(\u_multiplier/pp2_14 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_13_2/_18_  (.A(\u_multiplier/STAGE2/pp2_12_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_13_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_13_2/_19_  (.A1(\u_multiplier/pp1_13 [5]),
    .A2(\u_multiplier/pp1_13 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_13_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_13_2/_20_  (.A(\u_multiplier/pp1_13 [5]),
    .B(\u_multiplier/pp1_13 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_13_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_13_2/_21_  (.A1(\u_multiplier/pp1_13 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_13_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_13_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_13_2/_22_  (.A(\u_multiplier/pp1_13 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_13_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_13_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_13_2/_23_  (.A1(\u_multiplier/pp1_13 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_13_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_13_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_13_2/_24_  (.A(\u_multiplier/pp1_13 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_13_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_13_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_13_2/_25_  (.A(\u_multiplier/STAGE2/pp2_12_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_13_2/_16_ ),
    .ZN(\u_multiplier/pp2_13 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_13_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_13_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_13_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_13_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_13_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_13_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_13_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_13_2/_17_ ),
    .ZN(\u_multiplier/pp2_14 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_13_3/_18_  (.A(net134),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_13_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_13_3/_19_  (.A1(\u_multiplier/pp1_13 [9]),
    .A2(\u_multiplier/pp1_13 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_13_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_13_3/_20_  (.A(\u_multiplier/pp1_13 [9]),
    .B(\u_multiplier/pp1_13 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_13_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_13_3/_21_  (.A1(\u_multiplier/pp1_13 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_13_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_13_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_13_3/_22_  (.A(\u_multiplier/pp1_13 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_13_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_13_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_13_3/_23_  (.A1(\u_multiplier/pp1_13 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_13_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_13_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_13_3/_24_  (.A(\u_multiplier/pp1_13 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_13_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_13_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_13_3/_25_  (.A(net135),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_13_3/_16_ ),
    .ZN(\u_multiplier/pp2_13 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_13_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_13_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_13_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_13_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_13_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_13_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_13_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_13_3/_17_ ),
    .ZN(\u_multiplier/pp2_14 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_14_1/_18_  (.A(\u_multiplier/STAGE2/pp2_13_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_14_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_14_1/_19_  (.A1(\u_multiplier/pp1_14 [1]),
    .A2(\u_multiplier/pp1_14 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_14_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_14_1/_20_  (.A(\u_multiplier/pp1_14 [1]),
    .B(\u_multiplier/pp1_14 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_14_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_14_1/_21_  (.A1(\u_multiplier/pp1_14 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_14_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_14_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_14_1/_22_  (.A(\u_multiplier/pp1_14 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_14_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_14_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_14_1/_23_  (.A1(\u_multiplier/pp1_14 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_14_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_14_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_14_1/_24_  (.A(\u_multiplier/pp1_14 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_14_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_14_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_14_1/_25_  (.A(\u_multiplier/STAGE2/pp2_13_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_14_1/_16_ ),
    .ZN(\u_multiplier/pp2_14 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_14_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_14_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_14_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_14_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE2/E_4_2_pp2_14_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_14_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_14_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_14_1/_17_ ),
    .ZN(\u_multiplier/pp2_15 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_14_2/_18_  (.A(\u_multiplier/STAGE2/pp2_13_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_14_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_14_2/_19_  (.A1(\u_multiplier/pp1_14 [5]),
    .A2(\u_multiplier/pp1_14 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_14_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_14_2/_20_  (.A(\u_multiplier/pp1_14 [5]),
    .B(\u_multiplier/pp1_14 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_14_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_14_2/_21_  (.A1(\u_multiplier/pp1_14 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_14_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_14_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_14_2/_22_  (.A(\u_multiplier/pp1_14 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_14_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_14_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_14_2/_23_  (.A1(\u_multiplier/pp1_14 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_14_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_14_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_14_2/_24_  (.A(\u_multiplier/pp1_14 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_14_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_14_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_14_2/_25_  (.A(\u_multiplier/STAGE2/pp2_13_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_14_2/_16_ ),
    .ZN(\u_multiplier/pp2_14 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_14_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_14_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_14_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_14_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_14_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_14_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_14_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_14_2/_17_ ),
    .ZN(\u_multiplier/pp2_15 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_14_3/_18_  (.A(\u_multiplier/STAGE2/pp2_13_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_14_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_14_3/_19_  (.A1(\u_multiplier/pp1_14 [9]),
    .A2(\u_multiplier/pp1_14 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_14_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_14_3/_20_  (.A(\u_multiplier/pp1_14 [9]),
    .B(\u_multiplier/pp1_14 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_14_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_14_3/_21_  (.A1(\u_multiplier/pp1_14 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_14_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_14_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_14_3/_22_  (.A(\u_multiplier/pp1_14 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_14_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_14_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_14_3/_23_  (.A1(\u_multiplier/pp1_14 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_14_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_14_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_14_3/_24_  (.A(\u_multiplier/pp1_14 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_14_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_14_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_14_3/_25_  (.A(\u_multiplier/STAGE2/pp2_13_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_14_3/_16_ ),
    .ZN(\u_multiplier/pp2_14 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_14_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_14_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_14_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_14_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_14_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_14_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_14_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_14_3/_17_ ),
    .ZN(\u_multiplier/pp2_15 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_15_1/_18_  (.A(\u_multiplier/STAGE2/pp2_14_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_15_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_15_1/_19_  (.A1(\u_multiplier/pp1_15 [1]),
    .A2(\u_multiplier/pp1_15 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_15_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_15_1/_20_  (.A(\u_multiplier/pp1_15 [1]),
    .B(\u_multiplier/pp1_15 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_15_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_15_1/_21_  (.A1(\u_multiplier/pp1_15 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_15_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_15_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_15_1/_22_  (.A(\u_multiplier/pp1_15 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_15_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_15_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_15_1/_23_  (.A1(\u_multiplier/pp1_15 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_15_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_15_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_15_1/_24_  (.A(\u_multiplier/pp1_15 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_15_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_15_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_15_1/_25_  (.A(\u_multiplier/STAGE2/pp2_14_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_15_1/_16_ ),
    .ZN(\u_multiplier/pp2_15 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_15_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_15_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_15_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_15_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_15_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_15_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_15_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_15_1/_17_ ),
    .ZN(\u_multiplier/pp2_16 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_15_2/_18_  (.A(\u_multiplier/STAGE2/pp2_14_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_15_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_15_2/_19_  (.A1(\u_multiplier/pp1_15 [5]),
    .A2(\u_multiplier/pp1_15 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_15_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_15_2/_20_  (.A(\u_multiplier/pp1_15 [5]),
    .B(\u_multiplier/pp1_15 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_15_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_15_2/_21_  (.A1(\u_multiplier/pp1_15 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_15_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_15_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_15_2/_22_  (.A(\u_multiplier/pp1_15 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_15_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_15_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_15_2/_23_  (.A1(\u_multiplier/pp1_15 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_15_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_15_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_15_2/_24_  (.A(\u_multiplier/pp1_15 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_15_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_15_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_15_2/_25_  (.A(\u_multiplier/STAGE2/pp2_14_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_15_2/_16_ ),
    .ZN(\u_multiplier/pp2_15 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_15_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_15_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_15_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_15_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_15_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_15_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_15_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_15_2/_17_ ),
    .ZN(\u_multiplier/pp2_16 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_15_3/_18_  (.A(\u_multiplier/STAGE2/pp2_14_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_15_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_15_3/_19_  (.A1(\u_multiplier/pp1_15 [9]),
    .A2(\u_multiplier/pp1_15 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_15_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_15_3/_20_  (.A(\u_multiplier/pp1_15 [9]),
    .B(\u_multiplier/pp1_15 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_15_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_15_3/_21_  (.A1(\u_multiplier/pp1_15 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_15_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_15_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_15_3/_22_  (.A(\u_multiplier/pp1_15 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_15_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_15_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_15_3/_23_  (.A1(\u_multiplier/pp1_15 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_15_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_15_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_15_3/_24_  (.A(\u_multiplier/pp1_15 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_15_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_15_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_15_3/_25_  (.A(\u_multiplier/STAGE2/pp2_14_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_15_3/_16_ ),
    .ZN(\u_multiplier/pp2_15 [1]));
 NAND2_X2 \u_multiplier/STAGE2/E_4_2_pp2_15_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_15_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_15_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_15_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_15_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_15_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_15_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_15_3/_17_ ),
    .ZN(\u_multiplier/pp2_16 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_15_4/_18_  (.A(net136),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_15_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_15_4/_19_  (.A1(\u_multiplier/pp1_15 [13]),
    .A2(\u_multiplier/pp1_15 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_15_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_15_4/_20_  (.A(\u_multiplier/pp1_15 [13]),
    .B(\u_multiplier/pp1_15 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_15_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_15_4/_21_  (.A1(\u_multiplier/pp1_15 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_15_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_15_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_15_4/_22_  (.A(\u_multiplier/pp1_15 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_15_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_15_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_15_4/_23_  (.A1(\u_multiplier/pp1_15 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_15_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_15_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_15_4/_24_  (.A(\u_multiplier/pp1_15 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_15_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_15_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_15_4/_25_  (.A(net137),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_15_4/_16_ ),
    .ZN(\u_multiplier/pp2_15 [0]));
 NAND2_X2 \u_multiplier/STAGE2/E_4_2_pp2_15_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_15_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_15_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_15_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_15_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_15_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_15_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_15_4/_17_ ),
    .ZN(\u_multiplier/pp2_16 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_16_1/_18_  (.A(\u_multiplier/STAGE2/pp2_15_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_16_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_16_1/_19_  (.A1(\u_multiplier/pp1_16 [1]),
    .A2(\u_multiplier/pp1_16 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_16_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_16_1/_20_  (.A(\u_multiplier/pp1_16 [1]),
    .B(\u_multiplier/pp1_16 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_16_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_16_1/_21_  (.A1(\u_multiplier/pp1_16 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_16_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_16_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_16_1/_22_  (.A(\u_multiplier/pp1_16 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_16_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_16_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_16_1/_23_  (.A1(\u_multiplier/pp1_16 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_16_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_16_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_16_1/_24_  (.A(\u_multiplier/pp1_16 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_16_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_16_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_16_1/_25_  (.A(\u_multiplier/STAGE2/pp2_15_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_16_1/_16_ ),
    .ZN(\u_multiplier/pp2_16 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_16_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_16_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_16_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_16_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE2/E_4_2_pp2_16_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_16_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_16_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_16_1/_17_ ),
    .ZN(\u_multiplier/pp2_17 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_16_2/_18_  (.A(\u_multiplier/STAGE2/pp2_15_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_16_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_16_2/_19_  (.A1(\u_multiplier/pp1_16 [5]),
    .A2(\u_multiplier/pp1_16 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_16_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_16_2/_20_  (.A(\u_multiplier/pp1_16 [5]),
    .B(\u_multiplier/pp1_16 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_16_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_16_2/_21_  (.A1(\u_multiplier/pp1_16 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_16_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_16_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_16_2/_22_  (.A(\u_multiplier/pp1_16 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_16_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_16_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_16_2/_23_  (.A1(\u_multiplier/pp1_16 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_16_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_16_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_16_2/_24_  (.A(\u_multiplier/pp1_16 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_16_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_16_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_16_2/_25_  (.A(\u_multiplier/STAGE2/pp2_15_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_16_2/_16_ ),
    .ZN(\u_multiplier/pp2_16 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_16_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_16_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_16_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_16_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_16_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_16_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_16_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_16_2/_17_ ),
    .ZN(\u_multiplier/pp2_17 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_16_3/_18_  (.A(\u_multiplier/STAGE2/pp2_15_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_16_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_16_3/_19_  (.A1(\u_multiplier/pp1_16 [9]),
    .A2(\u_multiplier/pp1_16 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_16_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_16_3/_20_  (.A(\u_multiplier/pp1_16 [9]),
    .B(\u_multiplier/pp1_16 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_16_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_16_3/_21_  (.A1(\u_multiplier/pp1_16 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_16_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_16_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_16_3/_22_  (.A(\u_multiplier/pp1_16 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_16_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_16_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_16_3/_23_  (.A1(\u_multiplier/pp1_16 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_16_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_16_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_16_3/_24_  (.A(\u_multiplier/pp1_16 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_16_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_16_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_16_3/_25_  (.A(\u_multiplier/STAGE2/pp2_15_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_16_3/_16_ ),
    .ZN(\u_multiplier/pp2_16 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_16_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_16_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_16_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_16_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_16_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_16_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_16_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_16_3/_17_ ),
    .ZN(\u_multiplier/pp2_17 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_16_4/_18_  (.A(\u_multiplier/STAGE2/pp2_15_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_16_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_16_4/_19_  (.A1(\u_multiplier/pp1_16 [13]),
    .A2(\u_multiplier/pp1_16 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_16_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_16_4/_20_  (.A(\u_multiplier/pp1_16 [13]),
    .B(\u_multiplier/pp1_16 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_16_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_16_4/_21_  (.A1(\u_multiplier/pp1_16 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_16_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_16_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_16_4/_22_  (.A(\u_multiplier/pp1_16 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_16_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_16_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_16_4/_23_  (.A1(\u_multiplier/pp1_16 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_16_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_16_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_16_4/_24_  (.A(\u_multiplier/pp1_16 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_16_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_16_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_16_4/_25_  (.A(\u_multiplier/STAGE2/pp2_15_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_16_4/_16_ ),
    .ZN(\u_multiplier/pp2_16 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_16_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_16_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_16_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_16_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_16_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_16_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_16_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_16_4/_17_ ),
    .ZN(\u_multiplier/pp2_17 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_17_1/_18_  (.A(\u_multiplier/STAGE2/pp2_16_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_17_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_17_1/_19_  (.A1(\u_multiplier/pp1_17 [1]),
    .A2(\u_multiplier/pp1_17 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_17_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_17_1/_20_  (.A(\u_multiplier/pp1_17 [1]),
    .B(\u_multiplier/pp1_17 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_17_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_17_1/_21_  (.A1(\u_multiplier/pp1_17 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_17_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_17_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_17_1/_22_  (.A(\u_multiplier/pp1_17 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_17_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_17_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_17_1/_23_  (.A1(\u_multiplier/pp1_17 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_17_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_17_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_17_1/_24_  (.A(\u_multiplier/pp1_17 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_17_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_17_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_17_1/_25_  (.A(\u_multiplier/STAGE2/pp2_16_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_17_1/_16_ ),
    .ZN(\u_multiplier/pp2_17 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_17_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_17_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_17_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_17_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE2/E_4_2_pp2_17_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_17_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_17_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_17_1/_17_ ),
    .ZN(\u_multiplier/pp2_18 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_17_2/_18_  (.A(\u_multiplier/STAGE2/pp2_16_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_17_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_17_2/_19_  (.A1(\u_multiplier/pp1_17 [5]),
    .A2(\u_multiplier/pp1_17 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_17_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_17_2/_20_  (.A(\u_multiplier/pp1_17 [5]),
    .B(\u_multiplier/pp1_17 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_17_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_17_2/_21_  (.A1(\u_multiplier/pp1_17 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_17_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_17_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_17_2/_22_  (.A(\u_multiplier/pp1_17 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_17_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_17_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_17_2/_23_  (.A1(\u_multiplier/pp1_17 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_17_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_17_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_17_2/_24_  (.A(\u_multiplier/pp1_17 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_17_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_17_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_17_2/_25_  (.A(\u_multiplier/STAGE2/pp2_16_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_17_2/_16_ ),
    .ZN(\u_multiplier/pp2_17 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_17_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_17_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_17_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_17_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_17_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_17_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_17_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_17_2/_17_ ),
    .ZN(\u_multiplier/pp2_18 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_17_3/_18_  (.A(\u_multiplier/STAGE2/pp2_16_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_17_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_17_3/_19_  (.A1(\u_multiplier/pp1_17 [9]),
    .A2(\u_multiplier/pp1_17 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_17_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_17_3/_20_  (.A(\u_multiplier/pp1_17 [9]),
    .B(\u_multiplier/pp1_17 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_17_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_17_3/_21_  (.A1(\u_multiplier/pp1_17 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_17_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_17_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_17_3/_22_  (.A(\u_multiplier/pp1_17 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_17_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_17_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_17_3/_23_  (.A1(\u_multiplier/pp1_17 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_17_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_17_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_17_3/_24_  (.A(\u_multiplier/pp1_17 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_17_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_17_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_17_3/_25_  (.A(\u_multiplier/STAGE2/pp2_16_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_17_3/_16_ ),
    .ZN(\u_multiplier/pp2_17 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_17_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_17_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_17_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_17_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_17_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_17_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_17_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_17_3/_17_ ),
    .ZN(\u_multiplier/pp2_18 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_17_4/_18_  (.A(\u_multiplier/STAGE2/pp2_16_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_17_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_17_4/_19_  (.A1(\u_multiplier/pp1_17 [13]),
    .A2(\u_multiplier/pp1_17 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_17_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_17_4/_20_  (.A(\u_multiplier/pp1_17 [13]),
    .B(\u_multiplier/pp1_17 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_17_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_17_4/_21_  (.A1(\u_multiplier/pp1_17 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_17_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_17_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_17_4/_22_  (.A(\u_multiplier/pp1_17 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_17_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_17_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_17_4/_23_  (.A1(\u_multiplier/pp1_17 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_17_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_17_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_17_4/_24_  (.A(\u_multiplier/pp1_17 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_17_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_17_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_17_4/_25_  (.A(\u_multiplier/STAGE2/pp2_16_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_17_4/_16_ ),
    .ZN(\u_multiplier/pp2_17 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_17_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_17_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_17_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_17_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_17_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_17_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_17_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_17_4/_17_ ),
    .ZN(\u_multiplier/pp2_18 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_18_1/_18_  (.A(\u_multiplier/STAGE2/pp2_17_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_18_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_18_1/_19_  (.A1(\u_multiplier/pp1_18 [1]),
    .A2(\u_multiplier/pp1_18 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_18_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_18_1/_20_  (.A(\u_multiplier/pp1_18 [1]),
    .B(\u_multiplier/pp1_18 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_18_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_18_1/_21_  (.A1(\u_multiplier/pp1_18 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_18_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_18_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_18_1/_22_  (.A(\u_multiplier/pp1_18 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_18_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_18_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_18_1/_23_  (.A1(\u_multiplier/pp1_18 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_18_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_18_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_18_1/_24_  (.A(\u_multiplier/pp1_18 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_18_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_18_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_18_1/_25_  (.A(\u_multiplier/STAGE2/pp2_17_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_18_1/_16_ ),
    .ZN(\u_multiplier/pp2_18 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_18_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_18_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_18_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_18_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE2/E_4_2_pp2_18_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_18_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_18_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_18_1/_17_ ),
    .ZN(\u_multiplier/pp2_19 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_18_2/_18_  (.A(\u_multiplier/STAGE2/pp2_17_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_18_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_18_2/_19_  (.A1(\u_multiplier/pp1_18 [5]),
    .A2(\u_multiplier/pp1_18 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_18_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_18_2/_20_  (.A(\u_multiplier/pp1_18 [5]),
    .B(\u_multiplier/pp1_18 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_18_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_18_2/_21_  (.A1(\u_multiplier/pp1_18 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_18_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_18_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_18_2/_22_  (.A(\u_multiplier/pp1_18 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_18_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_18_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_18_2/_23_  (.A1(\u_multiplier/pp1_18 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_18_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_18_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_18_2/_24_  (.A(\u_multiplier/pp1_18 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_18_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_18_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_18_2/_25_  (.A(\u_multiplier/STAGE2/pp2_17_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_18_2/_16_ ),
    .ZN(\u_multiplier/pp2_18 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_18_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_18_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_18_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_18_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_18_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_18_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_18_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_18_2/_17_ ),
    .ZN(\u_multiplier/pp2_19 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_18_3/_18_  (.A(\u_multiplier/STAGE2/pp2_17_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_18_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_18_3/_19_  (.A1(\u_multiplier/pp1_18 [9]),
    .A2(\u_multiplier/pp1_18 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_18_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_18_3/_20_  (.A(\u_multiplier/pp1_18 [9]),
    .B(\u_multiplier/pp1_18 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_18_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_18_3/_21_  (.A1(\u_multiplier/pp1_18 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_18_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_18_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_18_3/_22_  (.A(\u_multiplier/pp1_18 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_18_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_18_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_18_3/_23_  (.A1(\u_multiplier/pp1_18 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_18_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_18_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_18_3/_24_  (.A(\u_multiplier/pp1_18 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_18_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_18_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_18_3/_25_  (.A(\u_multiplier/STAGE2/pp2_17_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_18_3/_16_ ),
    .ZN(\u_multiplier/pp2_18 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_18_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_18_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_18_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_18_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_18_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_18_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_18_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_18_3/_17_ ),
    .ZN(\u_multiplier/pp2_19 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_18_4/_18_  (.A(\u_multiplier/STAGE2/pp2_17_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_18_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_18_4/_19_  (.A1(\u_multiplier/pp1_18 [13]),
    .A2(\u_multiplier/pp1_18 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_18_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_18_4/_20_  (.A(\u_multiplier/pp1_18 [13]),
    .B(\u_multiplier/pp1_18 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_18_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_18_4/_21_  (.A1(\u_multiplier/pp1_18 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_18_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_18_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_18_4/_22_  (.A(\u_multiplier/pp1_18 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_18_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_18_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_18_4/_23_  (.A1(\u_multiplier/pp1_18 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_18_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_18_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_18_4/_24_  (.A(\u_multiplier/pp1_18 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_18_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_18_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_18_4/_25_  (.A(\u_multiplier/STAGE2/pp2_17_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_18_4/_16_ ),
    .ZN(\u_multiplier/pp2_18 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_18_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_18_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_18_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_18_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_18_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_18_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_18_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_18_4/_17_ ),
    .ZN(\u_multiplier/pp2_19 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_19_1/_18_  (.A(\u_multiplier/STAGE2/pp2_18_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_19_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_19_1/_19_  (.A1(\u_multiplier/pp1_19 [1]),
    .A2(\u_multiplier/pp1_19 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_19_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_19_1/_20_  (.A(\u_multiplier/pp1_19 [1]),
    .B(\u_multiplier/pp1_19 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_19_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_19_1/_21_  (.A1(\u_multiplier/pp1_19 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_19_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_19_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_19_1/_22_  (.A(\u_multiplier/pp1_19 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_19_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_19_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_19_1/_23_  (.A1(\u_multiplier/pp1_19 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_19_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_19_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_19_1/_24_  (.A(\u_multiplier/pp1_19 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_19_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_19_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_19_1/_25_  (.A(\u_multiplier/STAGE2/pp2_18_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_19_1/_16_ ),
    .ZN(\u_multiplier/pp2_19 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_19_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_19_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_19_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_19_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_19_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_19_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_19_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_19_1/_17_ ),
    .ZN(\u_multiplier/pp2_20 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_19_2/_18_  (.A(\u_multiplier/STAGE2/pp2_18_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_19_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_19_2/_19_  (.A1(\u_multiplier/pp1_19 [5]),
    .A2(\u_multiplier/pp1_19 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_19_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_19_2/_20_  (.A(\u_multiplier/pp1_19 [5]),
    .B(\u_multiplier/pp1_19 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_19_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_19_2/_21_  (.A1(\u_multiplier/pp1_19 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_19_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_19_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_19_2/_22_  (.A(\u_multiplier/pp1_19 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_19_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_19_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_19_2/_23_  (.A1(\u_multiplier/pp1_19 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_19_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_19_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_19_2/_24_  (.A(\u_multiplier/pp1_19 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_19_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_19_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_19_2/_25_  (.A(\u_multiplier/STAGE2/pp2_18_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_19_2/_16_ ),
    .ZN(\u_multiplier/pp2_19 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_19_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_19_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_19_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_19_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_19_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_19_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_19_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_19_2/_17_ ),
    .ZN(\u_multiplier/pp2_20 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_19_3/_18_  (.A(\u_multiplier/STAGE2/pp2_18_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_19_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_19_3/_19_  (.A1(\u_multiplier/pp1_19 [9]),
    .A2(\u_multiplier/pp1_19 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_19_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_19_3/_20_  (.A(\u_multiplier/pp1_19 [9]),
    .B(\u_multiplier/pp1_19 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_19_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_19_3/_21_  (.A1(\u_multiplier/pp1_19 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_19_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_19_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_19_3/_22_  (.A(\u_multiplier/pp1_19 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_19_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_19_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_19_3/_23_  (.A1(\u_multiplier/pp1_19 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_19_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_19_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_19_3/_24_  (.A(\u_multiplier/pp1_19 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_19_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_19_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_19_3/_25_  (.A(\u_multiplier/STAGE2/pp2_18_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_19_3/_16_ ),
    .ZN(\u_multiplier/pp2_19 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_19_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_19_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_19_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_19_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_19_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_19_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_19_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_19_3/_17_ ),
    .ZN(\u_multiplier/pp2_20 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_19_4/_18_  (.A(\u_multiplier/STAGE2/pp2_18_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_19_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_19_4/_19_  (.A1(\u_multiplier/pp1_19 [13]),
    .A2(\u_multiplier/pp1_19 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_19_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_19_4/_20_  (.A(\u_multiplier/pp1_19 [13]),
    .B(\u_multiplier/pp1_19 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_19_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_19_4/_21_  (.A1(\u_multiplier/pp1_19 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_19_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_19_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_19_4/_22_  (.A(\u_multiplier/pp1_19 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_19_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_19_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_19_4/_23_  (.A1(\u_multiplier/pp1_19 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_19_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_19_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_19_4/_24_  (.A(\u_multiplier/pp1_19 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_19_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_19_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_19_4/_25_  (.A(\u_multiplier/STAGE2/pp2_18_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_19_4/_16_ ),
    .ZN(\u_multiplier/pp2_19 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_19_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_19_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_19_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_19_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_19_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_19_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_19_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_19_4/_17_ ),
    .ZN(\u_multiplier/pp2_20 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_20_1/_18_  (.A(\u_multiplier/STAGE2/pp2_19_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_20_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_20_1/_19_  (.A1(\u_multiplier/pp1_20 [1]),
    .A2(\u_multiplier/pp1_20 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_20_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_20_1/_20_  (.A(\u_multiplier/pp1_20 [1]),
    .B(\u_multiplier/pp1_20 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_20_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_20_1/_21_  (.A1(\u_multiplier/pp1_20 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_20_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_20_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_20_1/_22_  (.A(\u_multiplier/pp1_20 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_20_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_20_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_20_1/_23_  (.A1(\u_multiplier/pp1_20 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_20_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_20_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_20_1/_24_  (.A(\u_multiplier/pp1_20 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_20_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_20_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_20_1/_25_  (.A(\u_multiplier/STAGE2/pp2_19_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_20_1/_16_ ),
    .ZN(\u_multiplier/pp2_20 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_20_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_20_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_20_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_20_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_20_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_20_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_20_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_20_1/_17_ ),
    .ZN(\u_multiplier/pp2_21 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_20_2/_18_  (.A(\u_multiplier/STAGE2/pp2_19_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_20_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_20_2/_19_  (.A1(\u_multiplier/pp1_20 [5]),
    .A2(\u_multiplier/pp1_20 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_20_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_20_2/_20_  (.A(\u_multiplier/pp1_20 [5]),
    .B(\u_multiplier/pp1_20 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_20_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_20_2/_21_  (.A1(\u_multiplier/pp1_20 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_20_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_20_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_20_2/_22_  (.A(\u_multiplier/pp1_20 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_20_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_20_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_20_2/_23_  (.A1(\u_multiplier/pp1_20 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_20_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_20_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_20_2/_24_  (.A(\u_multiplier/pp1_20 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_20_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_20_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_20_2/_25_  (.A(\u_multiplier/STAGE2/pp2_19_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_20_2/_16_ ),
    .ZN(\u_multiplier/pp2_20 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_20_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_20_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_20_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_20_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_20_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_20_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_20_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_20_2/_17_ ),
    .ZN(\u_multiplier/pp2_21 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_20_3/_18_  (.A(\u_multiplier/STAGE2/pp2_19_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_20_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_20_3/_19_  (.A1(\u_multiplier/pp1_20 [9]),
    .A2(\u_multiplier/pp1_20 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_20_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_20_3/_20_  (.A(\u_multiplier/pp1_20 [9]),
    .B(\u_multiplier/pp1_20 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_20_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_20_3/_21_  (.A1(\u_multiplier/pp1_20 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_20_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_20_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_20_3/_22_  (.A(\u_multiplier/pp1_20 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_20_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_20_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_20_3/_23_  (.A1(\u_multiplier/pp1_20 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_20_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_20_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_20_3/_24_  (.A(\u_multiplier/pp1_20 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_20_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_20_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_20_3/_25_  (.A(\u_multiplier/STAGE2/pp2_19_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_20_3/_16_ ),
    .ZN(\u_multiplier/pp2_20 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_20_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_20_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_20_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_20_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_20_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_20_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_20_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_20_3/_17_ ),
    .ZN(\u_multiplier/pp2_21 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_20_4/_18_  (.A(\u_multiplier/STAGE2/pp2_19_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_20_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_20_4/_19_  (.A1(\u_multiplier/pp1_20 [13]),
    .A2(\u_multiplier/pp1_20 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_20_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_20_4/_20_  (.A(\u_multiplier/pp1_20 [13]),
    .B(\u_multiplier/pp1_20 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_20_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_20_4/_21_  (.A1(\u_multiplier/pp1_20 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_20_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_20_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_20_4/_22_  (.A(\u_multiplier/pp1_20 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_20_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_20_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_20_4/_23_  (.A1(\u_multiplier/pp1_20 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_20_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_20_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_20_4/_24_  (.A(\u_multiplier/pp1_20 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_20_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_20_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_20_4/_25_  (.A(\u_multiplier/STAGE2/pp2_19_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_20_4/_16_ ),
    .ZN(\u_multiplier/pp2_20 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_20_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_20_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_20_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_20_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_20_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_20_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_20_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_20_4/_17_ ),
    .ZN(\u_multiplier/pp2_21 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_21_1/_18_  (.A(\u_multiplier/STAGE2/pp2_20_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_21_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_21_1/_19_  (.A1(\u_multiplier/pp1_21 [1]),
    .A2(\u_multiplier/pp1_21 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_21_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_21_1/_20_  (.A(\u_multiplier/pp1_21 [1]),
    .B(\u_multiplier/pp1_21 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_21_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_21_1/_21_  (.A1(\u_multiplier/pp1_21 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_21_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_21_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_21_1/_22_  (.A(\u_multiplier/pp1_21 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_21_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_21_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_21_1/_23_  (.A1(\u_multiplier/pp1_21 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_21_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_21_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_21_1/_24_  (.A(\u_multiplier/pp1_21 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_21_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_21_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_21_1/_25_  (.A(\u_multiplier/STAGE2/pp2_20_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_21_1/_16_ ),
    .ZN(\u_multiplier/pp2_21 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_21_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_21_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_21_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_21_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_21_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_21_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_21_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_21_1/_17_ ),
    .ZN(\u_multiplier/pp2_22 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_21_2/_18_  (.A(\u_multiplier/STAGE2/pp2_20_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_21_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_21_2/_19_  (.A1(\u_multiplier/pp1_21 [5]),
    .A2(\u_multiplier/pp1_21 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_21_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_21_2/_20_  (.A(\u_multiplier/pp1_21 [5]),
    .B(\u_multiplier/pp1_21 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_21_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_21_2/_21_  (.A1(\u_multiplier/pp1_21 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_21_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_21_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_21_2/_22_  (.A(\u_multiplier/pp1_21 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_21_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_21_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_21_2/_23_  (.A1(\u_multiplier/pp1_21 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_21_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_21_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_21_2/_24_  (.A(\u_multiplier/pp1_21 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_21_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_21_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_21_2/_25_  (.A(\u_multiplier/STAGE2/pp2_20_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_21_2/_16_ ),
    .ZN(\u_multiplier/pp2_21 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_21_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_21_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_21_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_21_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_21_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_21_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_21_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_21_2/_17_ ),
    .ZN(\u_multiplier/pp2_22 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_21_3/_18_  (.A(\u_multiplier/STAGE2/pp2_20_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_21_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_21_3/_19_  (.A1(\u_multiplier/pp1_21 [9]),
    .A2(\u_multiplier/pp1_21 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_21_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_21_3/_20_  (.A(\u_multiplier/pp1_21 [9]),
    .B(\u_multiplier/pp1_21 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_21_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_21_3/_21_  (.A1(\u_multiplier/pp1_21 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_21_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_21_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_21_3/_22_  (.A(\u_multiplier/pp1_21 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_21_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_21_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_21_3/_23_  (.A1(\u_multiplier/pp1_21 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_21_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_21_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_21_3/_24_  (.A(\u_multiplier/pp1_21 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_21_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_21_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_21_3/_25_  (.A(\u_multiplier/STAGE2/pp2_20_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_21_3/_16_ ),
    .ZN(\u_multiplier/pp2_21 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_21_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_21_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_21_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_21_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_21_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_21_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_21_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_21_3/_17_ ),
    .ZN(\u_multiplier/pp2_22 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_21_4/_18_  (.A(\u_multiplier/STAGE2/pp2_20_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_21_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_21_4/_19_  (.A1(\u_multiplier/pp1_21 [13]),
    .A2(\u_multiplier/pp1_21 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_21_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_21_4/_20_  (.A(\u_multiplier/pp1_21 [13]),
    .B(\u_multiplier/pp1_21 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_21_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_21_4/_21_  (.A1(\u_multiplier/pp1_21 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_21_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_21_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_21_4/_22_  (.A(\u_multiplier/pp1_21 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_21_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_21_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_21_4/_23_  (.A1(\u_multiplier/pp1_21 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_21_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_21_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_21_4/_24_  (.A(\u_multiplier/pp1_21 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_21_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_21_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_21_4/_25_  (.A(\u_multiplier/STAGE2/pp2_20_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_21_4/_16_ ),
    .ZN(\u_multiplier/pp2_21 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_21_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_21_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_21_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_21_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_21_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_21_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_21_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_21_4/_17_ ),
    .ZN(\u_multiplier/pp2_22 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_22_1/_18_  (.A(\u_multiplier/STAGE2/pp2_21_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_22_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_22_1/_19_  (.A1(\u_multiplier/pp1_22 [1]),
    .A2(\u_multiplier/pp1_22 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_22_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_22_1/_20_  (.A(\u_multiplier/pp1_22 [1]),
    .B(\u_multiplier/pp1_22 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_22_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_22_1/_21_  (.A1(\u_multiplier/pp1_22 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_22_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_22_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_22_1/_22_  (.A(\u_multiplier/pp1_22 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_22_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_22_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_22_1/_23_  (.A1(\u_multiplier/pp1_22 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_22_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_22_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_22_1/_24_  (.A(\u_multiplier/pp1_22 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_22_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_22_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_22_1/_25_  (.A(\u_multiplier/STAGE2/pp2_21_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_22_1/_16_ ),
    .ZN(\u_multiplier/pp2_22 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_22_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_22_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_22_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_22_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_22_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_22_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_22_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_22_1/_17_ ),
    .ZN(\u_multiplier/pp2_23 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_22_2/_18_  (.A(\u_multiplier/STAGE2/pp2_21_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_22_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_22_2/_19_  (.A1(\u_multiplier/pp1_22 [5]),
    .A2(\u_multiplier/pp1_22 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_22_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_22_2/_20_  (.A(\u_multiplier/pp1_22 [5]),
    .B(\u_multiplier/pp1_22 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_22_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_22_2/_21_  (.A1(\u_multiplier/pp1_22 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_22_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_22_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_22_2/_22_  (.A(\u_multiplier/pp1_22 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_22_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_22_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_22_2/_23_  (.A1(\u_multiplier/pp1_22 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_22_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_22_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_22_2/_24_  (.A(\u_multiplier/pp1_22 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_22_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_22_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_22_2/_25_  (.A(\u_multiplier/STAGE2/pp2_21_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_22_2/_16_ ),
    .ZN(\u_multiplier/pp2_22 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_22_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_22_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_22_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_22_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_22_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_22_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_22_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_22_2/_17_ ),
    .ZN(\u_multiplier/pp2_23 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_22_3/_18_  (.A(\u_multiplier/STAGE2/pp2_21_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_22_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_22_3/_19_  (.A1(\u_multiplier/pp1_22 [9]),
    .A2(\u_multiplier/pp1_22 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_22_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_22_3/_20_  (.A(\u_multiplier/pp1_22 [9]),
    .B(\u_multiplier/pp1_22 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_22_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_22_3/_21_  (.A1(\u_multiplier/pp1_22 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_22_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_22_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_22_3/_22_  (.A(\u_multiplier/pp1_22 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_22_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_22_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_22_3/_23_  (.A1(\u_multiplier/pp1_22 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_22_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_22_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_22_3/_24_  (.A(\u_multiplier/pp1_22 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_22_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_22_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_22_3/_25_  (.A(\u_multiplier/STAGE2/pp2_21_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_22_3/_16_ ),
    .ZN(\u_multiplier/pp2_22 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_22_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_22_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_22_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_22_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_22_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_22_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_22_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_22_3/_17_ ),
    .ZN(\u_multiplier/pp2_23 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_22_4/_18_  (.A(\u_multiplier/STAGE2/pp2_21_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_22_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_22_4/_19_  (.A1(\u_multiplier/pp1_22 [13]),
    .A2(\u_multiplier/pp1_22 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_22_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_22_4/_20_  (.A(\u_multiplier/pp1_22 [13]),
    .B(\u_multiplier/pp1_22 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_22_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_22_4/_21_  (.A1(\u_multiplier/pp1_22 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_22_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_22_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_22_4/_22_  (.A(\u_multiplier/pp1_22 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_22_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_22_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_22_4/_23_  (.A1(\u_multiplier/pp1_22 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_22_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_22_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_22_4/_24_  (.A(\u_multiplier/pp1_22 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_22_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_22_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_22_4/_25_  (.A(\u_multiplier/STAGE2/pp2_21_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_22_4/_16_ ),
    .ZN(\u_multiplier/pp2_22 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_22_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_22_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_22_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_22_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_22_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_22_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_22_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_22_4/_17_ ),
    .ZN(\u_multiplier/pp2_23 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_23_1/_18_  (.A(\u_multiplier/STAGE2/pp2_22_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_23_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_23_1/_19_  (.A1(\u_multiplier/pp1_23 [1]),
    .A2(\u_multiplier/pp1_23 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_23_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_23_1/_20_  (.A(\u_multiplier/pp1_23 [1]),
    .B(\u_multiplier/pp1_23 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_23_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_23_1/_21_  (.A1(\u_multiplier/pp1_23 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_23_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_23_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_23_1/_22_  (.A(\u_multiplier/pp1_23 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_23_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_23_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_23_1/_23_  (.A1(\u_multiplier/pp1_23 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_23_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_23_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_23_1/_24_  (.A(\u_multiplier/pp1_23 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_23_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_23_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_23_1/_25_  (.A(\u_multiplier/STAGE2/pp2_22_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_23_1/_16_ ),
    .ZN(\u_multiplier/pp2_23 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_23_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_23_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_23_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_23_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_23_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_23_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_23_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_23_1/_17_ ),
    .ZN(\u_multiplier/pp2_24 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_23_2/_18_  (.A(\u_multiplier/STAGE2/pp2_22_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_23_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_23_2/_19_  (.A1(\u_multiplier/pp1_23 [5]),
    .A2(\u_multiplier/pp1_23 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_23_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_23_2/_20_  (.A(\u_multiplier/pp1_23 [5]),
    .B(\u_multiplier/pp1_23 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_23_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_23_2/_21_  (.A1(\u_multiplier/pp1_23 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_23_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_23_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_23_2/_22_  (.A(\u_multiplier/pp1_23 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_23_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_23_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_23_2/_23_  (.A1(\u_multiplier/pp1_23 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_23_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_23_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_23_2/_24_  (.A(\u_multiplier/pp1_23 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_23_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_23_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_23_2/_25_  (.A(\u_multiplier/STAGE2/pp2_22_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_23_2/_16_ ),
    .ZN(\u_multiplier/pp2_23 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_23_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_23_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_23_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_23_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_23_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_23_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_23_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_23_2/_17_ ),
    .ZN(\u_multiplier/pp2_24 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_23_3/_18_  (.A(\u_multiplier/STAGE2/pp2_22_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_23_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_23_3/_19_  (.A1(\u_multiplier/pp1_23 [9]),
    .A2(\u_multiplier/pp1_23 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_23_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_23_3/_20_  (.A(\u_multiplier/pp1_23 [9]),
    .B(\u_multiplier/pp1_23 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_23_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_23_3/_21_  (.A1(\u_multiplier/pp1_23 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_23_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_23_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_23_3/_22_  (.A(\u_multiplier/pp1_23 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_23_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_23_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_23_3/_23_  (.A1(\u_multiplier/pp1_23 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_23_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_23_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_23_3/_24_  (.A(\u_multiplier/pp1_23 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_23_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_23_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_23_3/_25_  (.A(\u_multiplier/STAGE2/pp2_22_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_23_3/_16_ ),
    .ZN(\u_multiplier/pp2_23 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_23_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_23_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_23_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_23_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_23_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_23_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_23_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_23_3/_17_ ),
    .ZN(\u_multiplier/pp2_24 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_23_4/_18_  (.A(\u_multiplier/STAGE2/pp2_22_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_23_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_23_4/_19_  (.A1(\u_multiplier/pp1_23 [13]),
    .A2(\u_multiplier/pp1_23 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_23_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_23_4/_20_  (.A(\u_multiplier/pp1_23 [13]),
    .B(\u_multiplier/pp1_23 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_23_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_23_4/_21_  (.A1(\u_multiplier/pp1_23 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_23_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_23_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_23_4/_22_  (.A(\u_multiplier/pp1_23 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_23_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_23_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_23_4/_23_  (.A1(\u_multiplier/pp1_23 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_23_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_23_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_23_4/_24_  (.A(\u_multiplier/pp1_23 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_23_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_23_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_23_4/_25_  (.A(\u_multiplier/STAGE2/pp2_22_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_23_4/_16_ ),
    .ZN(\u_multiplier/pp2_23 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_23_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_23_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_23_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_23_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_23_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_23_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_23_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_23_4/_17_ ),
    .ZN(\u_multiplier/pp2_24 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_24_1/_18_  (.A(\u_multiplier/STAGE2/pp2_23_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_24_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_24_1/_19_  (.A1(\u_multiplier/pp1_24 [1]),
    .A2(\u_multiplier/pp1_24 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_24_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_24_1/_20_  (.A(\u_multiplier/pp1_24 [1]),
    .B(\u_multiplier/pp1_24 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_24_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_24_1/_21_  (.A1(\u_multiplier/pp1_24 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_24_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_24_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_24_1/_22_  (.A(\u_multiplier/pp1_24 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_24_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_24_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_24_1/_23_  (.A1(\u_multiplier/pp1_24 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_24_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_24_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_24_1/_24_  (.A(\u_multiplier/pp1_24 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_24_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_24_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_24_1/_25_  (.A(\u_multiplier/STAGE2/pp2_23_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_24_1/_16_ ),
    .ZN(\u_multiplier/pp2_24 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_24_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_24_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_24_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_24_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_24_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_24_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_24_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_24_1/_17_ ),
    .ZN(\u_multiplier/pp2_25 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_24_2/_18_  (.A(\u_multiplier/STAGE2/pp2_23_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_24_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_24_2/_19_  (.A1(\u_multiplier/pp1_24 [5]),
    .A2(\u_multiplier/pp1_24 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_24_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_24_2/_20_  (.A(\u_multiplier/pp1_24 [5]),
    .B(\u_multiplier/pp1_24 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_24_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_24_2/_21_  (.A1(\u_multiplier/pp1_24 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_24_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_24_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_24_2/_22_  (.A(\u_multiplier/pp1_24 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_24_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_24_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_24_2/_23_  (.A1(\u_multiplier/pp1_24 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_24_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_24_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_24_2/_24_  (.A(\u_multiplier/pp1_24 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_24_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_24_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_24_2/_25_  (.A(\u_multiplier/STAGE2/pp2_23_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_24_2/_16_ ),
    .ZN(\u_multiplier/pp2_24 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_24_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_24_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_24_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_24_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_24_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_24_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_24_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_24_2/_17_ ),
    .ZN(\u_multiplier/pp2_25 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_24_3/_18_  (.A(\u_multiplier/STAGE2/pp2_23_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_24_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_24_3/_19_  (.A1(\u_multiplier/pp1_24 [9]),
    .A2(\u_multiplier/pp1_24 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_24_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_24_3/_20_  (.A(\u_multiplier/pp1_24 [9]),
    .B(\u_multiplier/pp1_24 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_24_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_24_3/_21_  (.A1(\u_multiplier/pp1_24 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_24_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_24_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_24_3/_22_  (.A(\u_multiplier/pp1_24 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_24_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_24_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_24_3/_23_  (.A1(\u_multiplier/pp1_24 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_24_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_24_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_24_3/_24_  (.A(\u_multiplier/pp1_24 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_24_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_24_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_24_3/_25_  (.A(\u_multiplier/STAGE2/pp2_23_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_24_3/_16_ ),
    .ZN(\u_multiplier/pp2_24 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_24_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_24_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_24_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_24_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_24_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_24_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_24_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_24_3/_17_ ),
    .ZN(\u_multiplier/pp2_25 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_24_4/_18_  (.A(\u_multiplier/STAGE2/pp2_23_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_24_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_24_4/_19_  (.A1(\u_multiplier/pp1_24 [13]),
    .A2(\u_multiplier/pp1_24 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_24_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_24_4/_20_  (.A(\u_multiplier/pp1_24 [13]),
    .B(\u_multiplier/pp1_24 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_24_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_24_4/_21_  (.A1(\u_multiplier/pp1_24 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_24_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_24_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_24_4/_22_  (.A(\u_multiplier/pp1_24 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_24_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_24_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_24_4/_23_  (.A1(\u_multiplier/pp1_24 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_24_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_24_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_24_4/_24_  (.A(\u_multiplier/pp1_24 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_24_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_24_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_24_4/_25_  (.A(\u_multiplier/STAGE2/pp2_23_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_24_4/_16_ ),
    .ZN(\u_multiplier/pp2_24 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_24_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_24_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_24_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_24_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_24_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_24_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_24_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_24_4/_17_ ),
    .ZN(\u_multiplier/pp2_25 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_25_1/_18_  (.A(\u_multiplier/STAGE2/pp2_24_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_25_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_25_1/_19_  (.A1(\u_multiplier/pp1_25 [1]),
    .A2(\u_multiplier/pp1_25 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_25_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_25_1/_20_  (.A(\u_multiplier/pp1_25 [1]),
    .B(\u_multiplier/pp1_25 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_25_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_25_1/_21_  (.A1(\u_multiplier/pp1_25 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_25_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_25_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_25_1/_22_  (.A(\u_multiplier/pp1_25 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_25_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_25_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_25_1/_23_  (.A1(\u_multiplier/pp1_25 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_25_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_25_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_25_1/_24_  (.A(\u_multiplier/pp1_25 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_25_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_25_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_25_1/_25_  (.A(\u_multiplier/STAGE2/pp2_24_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_25_1/_16_ ),
    .ZN(\u_multiplier/pp2_25 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_25_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_25_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_25_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_25_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_25_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_25_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_25_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_25_1/_17_ ),
    .ZN(\u_multiplier/pp2_26 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_25_2/_18_  (.A(\u_multiplier/STAGE2/pp2_24_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_25_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_25_2/_19_  (.A1(\u_multiplier/pp1_25 [5]),
    .A2(\u_multiplier/pp1_25 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_25_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_25_2/_20_  (.A(\u_multiplier/pp1_25 [5]),
    .B(\u_multiplier/pp1_25 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_25_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_25_2/_21_  (.A1(\u_multiplier/pp1_25 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_25_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_25_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_25_2/_22_  (.A(\u_multiplier/pp1_25 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_25_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_25_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_25_2/_23_  (.A1(\u_multiplier/pp1_25 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_25_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_25_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_25_2/_24_  (.A(\u_multiplier/pp1_25 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_25_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_25_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_25_2/_25_  (.A(\u_multiplier/STAGE2/pp2_24_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_25_2/_16_ ),
    .ZN(\u_multiplier/pp2_25 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_25_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_25_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_25_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_25_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_25_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_25_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_25_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_25_2/_17_ ),
    .ZN(\u_multiplier/pp2_26 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_25_3/_18_  (.A(\u_multiplier/STAGE2/pp2_24_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_25_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_25_3/_19_  (.A1(\u_multiplier/pp1_25 [9]),
    .A2(\u_multiplier/pp1_25 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_25_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_25_3/_20_  (.A(\u_multiplier/pp1_25 [9]),
    .B(\u_multiplier/pp1_25 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_25_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_25_3/_21_  (.A1(\u_multiplier/pp1_25 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_25_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_25_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_25_3/_22_  (.A(\u_multiplier/pp1_25 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_25_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_25_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_25_3/_23_  (.A1(\u_multiplier/pp1_25 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_25_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_25_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_25_3/_24_  (.A(\u_multiplier/pp1_25 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_25_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_25_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_25_3/_25_  (.A(\u_multiplier/STAGE2/pp2_24_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_25_3/_16_ ),
    .ZN(\u_multiplier/pp2_25 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_25_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_25_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_25_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_25_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_25_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_25_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_25_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_25_3/_17_ ),
    .ZN(\u_multiplier/pp2_26 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_25_4/_18_  (.A(\u_multiplier/STAGE2/pp2_24_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_25_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_25_4/_19_  (.A1(\u_multiplier/pp1_25 [13]),
    .A2(\u_multiplier/pp1_25 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_25_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_25_4/_20_  (.A(\u_multiplier/pp1_25 [13]),
    .B(\u_multiplier/pp1_25 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_25_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_25_4/_21_  (.A1(\u_multiplier/pp1_25 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_25_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_25_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_25_4/_22_  (.A(\u_multiplier/pp1_25 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_25_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_25_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_25_4/_23_  (.A1(\u_multiplier/pp1_25 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_25_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_25_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_25_4/_24_  (.A(\u_multiplier/pp1_25 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_25_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_25_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_25_4/_25_  (.A(\u_multiplier/STAGE2/pp2_24_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_25_4/_16_ ),
    .ZN(\u_multiplier/pp2_25 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_25_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_25_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_25_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_25_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_25_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_25_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_25_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_25_4/_17_ ),
    .ZN(\u_multiplier/pp2_26 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_26_1/_18_  (.A(\u_multiplier/STAGE2/pp2_25_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_26_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_26_1/_19_  (.A1(\u_multiplier/pp1_26 [1]),
    .A2(\u_multiplier/pp1_26 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_26_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_26_1/_20_  (.A(\u_multiplier/pp1_26 [1]),
    .B(\u_multiplier/pp1_26 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_26_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_26_1/_21_  (.A1(\u_multiplier/pp1_26 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_26_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_26_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_26_1/_22_  (.A(\u_multiplier/pp1_26 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_26_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_26_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_26_1/_23_  (.A1(\u_multiplier/pp1_26 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_26_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_26_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_26_1/_24_  (.A(\u_multiplier/pp1_26 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_26_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_26_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_26_1/_25_  (.A(\u_multiplier/STAGE2/pp2_25_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_26_1/_16_ ),
    .ZN(\u_multiplier/pp2_26 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_26_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_26_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_26_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_26_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_26_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_26_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_26_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_26_1/_17_ ),
    .ZN(\u_multiplier/pp2_27 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_26_2/_18_  (.A(\u_multiplier/STAGE2/pp2_25_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_26_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_26_2/_19_  (.A1(\u_multiplier/pp1_26 [5]),
    .A2(\u_multiplier/pp1_26 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_26_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_26_2/_20_  (.A(\u_multiplier/pp1_26 [5]),
    .B(\u_multiplier/pp1_26 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_26_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_26_2/_21_  (.A1(\u_multiplier/pp1_26 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_26_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_26_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_26_2/_22_  (.A(\u_multiplier/pp1_26 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_26_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_26_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_26_2/_23_  (.A1(\u_multiplier/pp1_26 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_26_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_26_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_26_2/_24_  (.A(\u_multiplier/pp1_26 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_26_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_26_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_26_2/_25_  (.A(\u_multiplier/STAGE2/pp2_25_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_26_2/_16_ ),
    .ZN(\u_multiplier/pp2_26 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_26_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_26_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_26_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_26_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_26_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_26_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_26_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_26_2/_17_ ),
    .ZN(\u_multiplier/pp2_27 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_26_3/_18_  (.A(\u_multiplier/STAGE2/pp2_25_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_26_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_26_3/_19_  (.A1(\u_multiplier/pp1_26 [9]),
    .A2(\u_multiplier/pp1_26 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_26_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_26_3/_20_  (.A(\u_multiplier/pp1_26 [9]),
    .B(\u_multiplier/pp1_26 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_26_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_26_3/_21_  (.A1(\u_multiplier/pp1_26 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_26_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_26_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_26_3/_22_  (.A(\u_multiplier/pp1_26 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_26_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_26_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_26_3/_23_  (.A1(\u_multiplier/pp1_26 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_26_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_26_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_26_3/_24_  (.A(\u_multiplier/pp1_26 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_26_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_26_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_26_3/_25_  (.A(\u_multiplier/STAGE2/pp2_25_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_26_3/_16_ ),
    .ZN(\u_multiplier/pp2_26 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_26_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_26_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_26_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_26_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_26_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_26_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_26_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_26_3/_17_ ),
    .ZN(\u_multiplier/pp2_27 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_26_4/_18_  (.A(\u_multiplier/STAGE2/pp2_25_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_26_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_26_4/_19_  (.A1(\u_multiplier/pp1_26 [13]),
    .A2(\u_multiplier/pp1_26 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_26_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_26_4/_20_  (.A(\u_multiplier/pp1_26 [13]),
    .B(\u_multiplier/pp1_26 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_26_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_26_4/_21_  (.A1(\u_multiplier/pp1_26 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_26_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_26_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_26_4/_22_  (.A(\u_multiplier/pp1_26 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_26_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_26_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_26_4/_23_  (.A1(\u_multiplier/pp1_26 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_26_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_26_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_26_4/_24_  (.A(\u_multiplier/pp1_26 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_26_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_26_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_26_4/_25_  (.A(\u_multiplier/STAGE2/pp2_25_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_26_4/_16_ ),
    .ZN(\u_multiplier/pp2_26 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_26_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_26_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_26_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_26_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_26_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_26_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_26_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_26_4/_17_ ),
    .ZN(\u_multiplier/pp2_27 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_27_1/_18_  (.A(\u_multiplier/STAGE2/pp2_26_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_27_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_27_1/_19_  (.A1(\u_multiplier/pp1_27 [1]),
    .A2(\u_multiplier/pp1_27 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_27_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_27_1/_20_  (.A(\u_multiplier/pp1_27 [1]),
    .B(\u_multiplier/pp1_27 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_27_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_27_1/_21_  (.A1(\u_multiplier/pp1_27 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_27_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_27_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_27_1/_22_  (.A(\u_multiplier/pp1_27 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_27_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_27_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_27_1/_23_  (.A1(\u_multiplier/pp1_27 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_27_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_27_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_27_1/_24_  (.A(\u_multiplier/pp1_27 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_27_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_27_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_27_1/_25_  (.A(\u_multiplier/STAGE2/pp2_26_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_27_1/_16_ ),
    .ZN(\u_multiplier/pp2_27 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_27_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_27_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_27_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_27_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_27_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_27_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_27_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_27_1/_17_ ),
    .ZN(\u_multiplier/pp2_28 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_27_2/_18_  (.A(\u_multiplier/STAGE2/pp2_26_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_27_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_27_2/_19_  (.A1(\u_multiplier/pp1_27 [5]),
    .A2(\u_multiplier/pp1_27 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_27_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_27_2/_20_  (.A(\u_multiplier/pp1_27 [5]),
    .B(\u_multiplier/pp1_27 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_27_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_27_2/_21_  (.A1(\u_multiplier/pp1_27 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_27_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_27_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_27_2/_22_  (.A(\u_multiplier/pp1_27 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_27_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_27_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_27_2/_23_  (.A1(\u_multiplier/pp1_27 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_27_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_27_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_27_2/_24_  (.A(\u_multiplier/pp1_27 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_27_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_27_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_27_2/_25_  (.A(\u_multiplier/STAGE2/pp2_26_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_27_2/_16_ ),
    .ZN(\u_multiplier/pp2_27 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_27_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_27_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_27_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_27_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_27_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_27_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_27_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_27_2/_17_ ),
    .ZN(\u_multiplier/pp2_28 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_27_3/_18_  (.A(\u_multiplier/STAGE2/pp2_26_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_27_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_27_3/_19_  (.A1(\u_multiplier/pp1_27 [9]),
    .A2(\u_multiplier/pp1_27 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_27_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_27_3/_20_  (.A(\u_multiplier/pp1_27 [9]),
    .B(\u_multiplier/pp1_27 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_27_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_27_3/_21_  (.A1(\u_multiplier/pp1_27 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_27_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_27_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_27_3/_22_  (.A(\u_multiplier/pp1_27 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_27_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_27_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_27_3/_23_  (.A1(\u_multiplier/pp1_27 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_27_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_27_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_27_3/_24_  (.A(\u_multiplier/pp1_27 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_27_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_27_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_27_3/_25_  (.A(\u_multiplier/STAGE2/pp2_26_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_27_3/_16_ ),
    .ZN(\u_multiplier/pp2_27 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_27_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_27_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_27_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_27_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_27_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_27_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_27_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_27_3/_17_ ),
    .ZN(\u_multiplier/pp2_28 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_27_4/_18_  (.A(\u_multiplier/STAGE2/pp2_26_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_27_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_27_4/_19_  (.A1(\u_multiplier/pp1_27 [13]),
    .A2(\u_multiplier/pp1_27 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_27_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_27_4/_20_  (.A(\u_multiplier/pp1_27 [13]),
    .B(\u_multiplier/pp1_27 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_27_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_27_4/_21_  (.A1(\u_multiplier/pp1_27 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_27_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_27_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_27_4/_22_  (.A(\u_multiplier/pp1_27 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_27_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_27_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_27_4/_23_  (.A1(\u_multiplier/pp1_27 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_27_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_27_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_27_4/_24_  (.A(\u_multiplier/pp1_27 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_27_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_27_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_27_4/_25_  (.A(\u_multiplier/STAGE2/pp2_26_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_27_4/_16_ ),
    .ZN(\u_multiplier/pp2_27 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_27_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_27_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_27_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_27_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_27_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_27_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_27_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_27_4/_17_ ),
    .ZN(\u_multiplier/pp2_28 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_28_1/_18_  (.A(\u_multiplier/STAGE2/pp2_27_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_28_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_28_1/_19_  (.A1(\u_multiplier/pp1_28 [1]),
    .A2(\u_multiplier/pp1_28 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_28_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_28_1/_20_  (.A(\u_multiplier/pp1_28 [1]),
    .B(\u_multiplier/pp1_28 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_28_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_28_1/_21_  (.A1(\u_multiplier/pp1_28 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_28_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_28_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_28_1/_22_  (.A(\u_multiplier/pp1_28 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_28_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_28_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_28_1/_23_  (.A1(\u_multiplier/pp1_28 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_28_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_28_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_28_1/_24_  (.A(\u_multiplier/pp1_28 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_28_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_28_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_28_1/_25_  (.A(\u_multiplier/STAGE2/pp2_27_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_28_1/_16_ ),
    .ZN(\u_multiplier/pp2_28 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_28_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_28_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_28_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_28_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_28_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_28_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_28_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_28_1/_17_ ),
    .ZN(\u_multiplier/pp2_29 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_28_2/_18_  (.A(\u_multiplier/STAGE2/pp2_27_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_28_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_28_2/_19_  (.A1(\u_multiplier/pp1_28 [5]),
    .A2(\u_multiplier/pp1_28 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_28_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_28_2/_20_  (.A(\u_multiplier/pp1_28 [5]),
    .B(\u_multiplier/pp1_28 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_28_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_28_2/_21_  (.A1(\u_multiplier/pp1_28 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_28_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_28_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_28_2/_22_  (.A(\u_multiplier/pp1_28 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_28_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_28_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_28_2/_23_  (.A1(\u_multiplier/pp1_28 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_28_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_28_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_28_2/_24_  (.A(\u_multiplier/pp1_28 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_28_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_28_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_28_2/_25_  (.A(\u_multiplier/STAGE2/pp2_27_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_28_2/_16_ ),
    .ZN(\u_multiplier/pp2_28 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_28_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_28_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_28_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_28_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_28_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_28_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_28_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_28_2/_17_ ),
    .ZN(\u_multiplier/pp2_29 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_28_3/_18_  (.A(\u_multiplier/STAGE2/pp2_27_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_28_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_28_3/_19_  (.A1(\u_multiplier/pp1_28 [9]),
    .A2(\u_multiplier/pp1_28 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_28_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_28_3/_20_  (.A(\u_multiplier/pp1_28 [9]),
    .B(\u_multiplier/pp1_28 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_28_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_28_3/_21_  (.A1(\u_multiplier/pp1_28 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_28_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_28_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_28_3/_22_  (.A(\u_multiplier/pp1_28 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_28_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_28_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_28_3/_23_  (.A1(\u_multiplier/pp1_28 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_28_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_28_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_28_3/_24_  (.A(\u_multiplier/pp1_28 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_28_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_28_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_28_3/_25_  (.A(\u_multiplier/STAGE2/pp2_27_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_28_3/_16_ ),
    .ZN(\u_multiplier/pp2_28 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_28_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_28_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_28_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_28_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_28_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_28_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_28_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_28_3/_17_ ),
    .ZN(\u_multiplier/pp2_29 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_28_4/_18_  (.A(\u_multiplier/STAGE2/pp2_27_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_28_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_28_4/_19_  (.A1(\u_multiplier/pp1_28 [13]),
    .A2(\u_multiplier/pp1_28 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_28_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_28_4/_20_  (.A(\u_multiplier/pp1_28 [13]),
    .B(\u_multiplier/pp1_28 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_28_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_28_4/_21_  (.A1(\u_multiplier/pp1_28 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_28_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_28_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_28_4/_22_  (.A(\u_multiplier/pp1_28 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_28_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_28_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_28_4/_23_  (.A1(\u_multiplier/pp1_28 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_28_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_28_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_28_4/_24_  (.A(\u_multiplier/pp1_28 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_28_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_28_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_28_4/_25_  (.A(\u_multiplier/STAGE2/pp2_27_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_28_4/_16_ ),
    .ZN(\u_multiplier/pp2_28 [0]));
 NAND2_X2 \u_multiplier/STAGE2/E_4_2_pp2_28_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_28_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_28_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_28_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_28_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_28_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_28_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_28_4/_17_ ),
    .ZN(\u_multiplier/pp2_29 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_29_1/_18_  (.A(\u_multiplier/STAGE2/pp2_28_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_29_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_29_1/_19_  (.A1(\u_multiplier/pp1_29 [1]),
    .A2(\u_multiplier/pp1_29 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_29_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_29_1/_20_  (.A(\u_multiplier/pp1_29 [1]),
    .B(\u_multiplier/pp1_29 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_29_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_29_1/_21_  (.A1(\u_multiplier/pp1_29 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_29_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_29_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_29_1/_22_  (.A(\u_multiplier/pp1_29 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_29_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_29_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_29_1/_23_  (.A1(\u_multiplier/pp1_29 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_29_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_29_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_29_1/_24_  (.A(\u_multiplier/pp1_29 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_29_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_29_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_29_1/_25_  (.A(\u_multiplier/STAGE2/pp2_28_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_29_1/_16_ ),
    .ZN(\u_multiplier/pp2_29 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_29_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_29_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_29_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_29_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_29_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_29_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_29_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_29_1/_17_ ),
    .ZN(\u_multiplier/pp2_30 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_29_2/_18_  (.A(\u_multiplier/STAGE2/pp2_28_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_29_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_29_2/_19_  (.A1(\u_multiplier/pp1_29 [5]),
    .A2(\u_multiplier/pp1_29 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_29_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_29_2/_20_  (.A(\u_multiplier/pp1_29 [5]),
    .B(\u_multiplier/pp1_29 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_29_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_29_2/_21_  (.A1(\u_multiplier/pp1_29 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_29_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_29_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_29_2/_22_  (.A(\u_multiplier/pp1_29 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_29_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_29_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_29_2/_23_  (.A1(\u_multiplier/pp1_29 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_29_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_29_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_29_2/_24_  (.A(\u_multiplier/pp1_29 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_29_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_29_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_29_2/_25_  (.A(\u_multiplier/STAGE2/pp2_28_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_29_2/_16_ ),
    .ZN(\u_multiplier/pp2_29 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_29_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_29_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_29_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_29_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_29_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_29_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_29_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_29_2/_17_ ),
    .ZN(\u_multiplier/pp2_30 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_29_3/_18_  (.A(\u_multiplier/STAGE2/pp2_28_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_29_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_29_3/_19_  (.A1(\u_multiplier/pp1_29 [9]),
    .A2(\u_multiplier/pp1_29 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_29_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_29_3/_20_  (.A(\u_multiplier/pp1_29 [9]),
    .B(\u_multiplier/pp1_29 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_29_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_29_3/_21_  (.A1(\u_multiplier/pp1_29 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_29_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_29_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_29_3/_22_  (.A(\u_multiplier/pp1_29 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_29_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_29_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_29_3/_23_  (.A1(\u_multiplier/pp1_29 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_29_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_29_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_29_3/_24_  (.A(\u_multiplier/pp1_29 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_29_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_29_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_29_3/_25_  (.A(\u_multiplier/STAGE2/pp2_28_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_29_3/_16_ ),
    .ZN(\u_multiplier/pp2_29 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_29_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_29_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_29_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_29_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_29_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_29_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_29_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_29_3/_17_ ),
    .ZN(\u_multiplier/pp2_30 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_29_4/_18_  (.A(\u_multiplier/STAGE2/pp2_28_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_29_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_29_4/_19_  (.A1(\u_multiplier/pp1_29 [13]),
    .A2(\u_multiplier/pp1_29 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_29_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_29_4/_20_  (.A(\u_multiplier/pp1_29 [13]),
    .B(\u_multiplier/pp1_29 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_29_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_29_4/_21_  (.A1(\u_multiplier/pp1_29 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_29_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_29_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_29_4/_22_  (.A(\u_multiplier/pp1_29 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_29_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_29_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_29_4/_23_  (.A1(\u_multiplier/pp1_29 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_29_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_29_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_29_4/_24_  (.A(\u_multiplier/pp1_29 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_29_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_29_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_29_4/_25_  (.A(\u_multiplier/STAGE2/pp2_28_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_29_4/_16_ ),
    .ZN(\u_multiplier/pp2_29 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_29_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_29_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_29_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_29_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_29_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_29_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_29_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_29_4/_17_ ),
    .ZN(\u_multiplier/pp2_30 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_30_1/_18_  (.A(\u_multiplier/STAGE2/pp2_29_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_30_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_30_1/_19_  (.A1(\u_multiplier/pp1_30 [1]),
    .A2(\u_multiplier/pp1_30 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_30_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_30_1/_20_  (.A(\u_multiplier/pp1_30 [1]),
    .B(\u_multiplier/pp1_30 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_30_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_30_1/_21_  (.A1(\u_multiplier/pp1_30 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_30_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_30_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_30_1/_22_  (.A(\u_multiplier/pp1_30 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_30_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_30_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_30_1/_23_  (.A1(\u_multiplier/pp1_30 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_30_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_30_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_30_1/_24_  (.A(\u_multiplier/pp1_30 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_30_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_30_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_30_1/_25_  (.A(\u_multiplier/STAGE2/pp2_29_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_30_1/_16_ ),
    .ZN(\u_multiplier/pp2_30 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_30_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_30_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_30_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_30_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE2/E_4_2_pp2_30_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_30_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_30_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_30_1/_17_ ),
    .ZN(\u_multiplier/pp2_31 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_30_2/_18_  (.A(\u_multiplier/STAGE2/pp2_29_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_30_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_30_2/_19_  (.A1(\u_multiplier/pp1_30 [5]),
    .A2(\u_multiplier/pp1_30 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_30_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_30_2/_20_  (.A(\u_multiplier/pp1_30 [5]),
    .B(\u_multiplier/pp1_30 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_30_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_30_2/_21_  (.A1(\u_multiplier/pp1_30 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_30_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_30_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_30_2/_22_  (.A(\u_multiplier/pp1_30 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_30_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_30_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_30_2/_23_  (.A1(\u_multiplier/pp1_30 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_30_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_30_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_30_2/_24_  (.A(\u_multiplier/pp1_30 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_30_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_30_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_30_2/_25_  (.A(\u_multiplier/STAGE2/pp2_29_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_30_2/_16_ ),
    .ZN(\u_multiplier/pp2_30 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_30_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_30_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_30_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_30_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_30_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_30_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_30_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_30_2/_17_ ),
    .ZN(\u_multiplier/pp2_31 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_30_3/_18_  (.A(\u_multiplier/STAGE2/pp2_29_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_30_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_30_3/_19_  (.A1(\u_multiplier/pp1_30 [9]),
    .A2(\u_multiplier/pp1_30 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_30_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_30_3/_20_  (.A(\u_multiplier/pp1_30 [9]),
    .B(\u_multiplier/pp1_30 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_30_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_30_3/_21_  (.A1(\u_multiplier/pp1_30 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_30_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_30_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_30_3/_22_  (.A(\u_multiplier/pp1_30 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_30_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_30_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_30_3/_23_  (.A1(\u_multiplier/pp1_30 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_30_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_30_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_30_3/_24_  (.A(\u_multiplier/pp1_30 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_30_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_30_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_30_3/_25_  (.A(\u_multiplier/STAGE2/pp2_29_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_30_3/_16_ ),
    .ZN(\u_multiplier/pp2_30 [1]));
 NAND2_X2 \u_multiplier/STAGE2/E_4_2_pp2_30_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_30_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_30_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_30_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_30_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_30_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_30_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_30_3/_17_ ),
    .ZN(\u_multiplier/pp2_31 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_30_4/_18_  (.A(\u_multiplier/STAGE2/pp2_29_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_30_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_30_4/_19_  (.A1(\u_multiplier/pp1_30 [13]),
    .A2(\u_multiplier/pp1_30 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_30_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_30_4/_20_  (.A(\u_multiplier/pp1_30 [13]),
    .B(\u_multiplier/pp1_30 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_30_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_30_4/_21_  (.A1(\u_multiplier/pp1_30 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_30_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_30_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_30_4/_22_  (.A(\u_multiplier/pp1_30 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_30_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_30_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_30_4/_23_  (.A1(\u_multiplier/pp1_30 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_30_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_30_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_30_4/_24_  (.A(\u_multiplier/pp1_30 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_30_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_30_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_30_4/_25_  (.A(\u_multiplier/STAGE2/pp2_29_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_30_4/_16_ ),
    .ZN(\u_multiplier/pp2_30 [0]));
 NAND2_X2 \u_multiplier/STAGE2/E_4_2_pp2_30_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_30_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_30_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_30_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_30_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_30_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_30_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_30_4/_17_ ),
    .ZN(\u_multiplier/pp2_31 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_31_1/_18_  (.A(\u_multiplier/STAGE2/pp2_30_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_31_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_31_1/_19_  (.A1(\u_multiplier/pp1_31 [1]),
    .A2(\u_multiplier/pp1_31 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_31_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_31_1/_20_  (.A(\u_multiplier/pp1_31 [1]),
    .B(\u_multiplier/pp1_31 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_31_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_31_1/_21_  (.A1(\u_multiplier/pp1_31 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_31_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_31_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_31_1/_22_  (.A(\u_multiplier/pp1_31 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_31_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_31_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_31_1/_23_  (.A1(\u_multiplier/pp1_31 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_31_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_31_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_31_1/_24_  (.A(\u_multiplier/pp1_31 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_31_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_31_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_31_1/_25_  (.A(\u_multiplier/STAGE2/pp2_30_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_31_1/_16_ ),
    .ZN(\u_multiplier/pp2_31 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_31_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_31_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_31_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_31_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE2/E_4_2_pp2_31_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_31_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_31_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_31_1/_17_ ),
    .ZN(\u_multiplier/pp2_32 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_31_2/_18_  (.A(\u_multiplier/STAGE2/pp2_30_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_31_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_31_2/_19_  (.A1(\u_multiplier/pp1_31 [5]),
    .A2(\u_multiplier/pp1_31 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_31_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_31_2/_20_  (.A(\u_multiplier/pp1_31 [5]),
    .B(\u_multiplier/pp1_31 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_31_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_31_2/_21_  (.A1(\u_multiplier/pp1_31 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_31_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_31_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_31_2/_22_  (.A(\u_multiplier/pp1_31 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_31_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_31_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_31_2/_23_  (.A1(\u_multiplier/pp1_31 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_31_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_31_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_31_2/_24_  (.A(\u_multiplier/pp1_31 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_31_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_31_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_31_2/_25_  (.A(\u_multiplier/STAGE2/pp2_30_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_31_2/_16_ ),
    .ZN(\u_multiplier/pp2_31 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_31_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_31_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_31_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_31_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_31_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_31_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_31_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_31_2/_17_ ),
    .ZN(\u_multiplier/pp2_32 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_31_3/_18_  (.A(\u_multiplier/STAGE2/pp2_30_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_31_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_31_3/_19_  (.A1(\u_multiplier/pp1_31 [9]),
    .A2(\u_multiplier/pp1_31 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_31_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_31_3/_20_  (.A(\u_multiplier/pp1_31 [9]),
    .B(\u_multiplier/pp1_31 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_31_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_31_3/_21_  (.A1(\u_multiplier/pp1_31 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_31_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_31_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_31_3/_22_  (.A(\u_multiplier/pp1_31 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_31_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_31_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_31_3/_23_  (.A1(\u_multiplier/pp1_31 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_31_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_31_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_31_3/_24_  (.A(\u_multiplier/pp1_31 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_31_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_31_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_31_3/_25_  (.A(\u_multiplier/STAGE2/pp2_30_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_31_3/_16_ ),
    .ZN(\u_multiplier/pp2_31 [1]));
 NAND2_X2 \u_multiplier/STAGE2/E_4_2_pp2_31_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_31_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_31_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_31_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_31_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_31_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_31_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_31_3/_17_ ),
    .ZN(\u_multiplier/pp2_32 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_31_4/_18_  (.A(\u_multiplier/STAGE2/pp2_30_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_31_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_31_4/_19_  (.A1(\u_multiplier/pp1_31 [13]),
    .A2(\u_multiplier/pp1_31 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_31_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_31_4/_20_  (.A(\u_multiplier/pp1_31 [13]),
    .B(\u_multiplier/pp1_31 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_31_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_31_4/_21_  (.A1(\u_multiplier/pp1_31 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_31_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_31_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_31_4/_22_  (.A(\u_multiplier/pp1_31 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_31_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_31_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_31_4/_23_  (.A1(\u_multiplier/pp1_31 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_31_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_31_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_31_4/_24_  (.A(\u_multiplier/pp1_31 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_31_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_31_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_31_4/_25_  (.A(\u_multiplier/STAGE2/pp2_30_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_31_4/_16_ ),
    .ZN(\u_multiplier/pp2_31 [0]));
 NAND2_X2 \u_multiplier/STAGE2/E_4_2_pp2_31_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_31_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_31_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_31_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_31_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_31_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_31_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_31_4/_17_ ),
    .ZN(\u_multiplier/pp2_32 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_32_1/_18_  (.A(\u_multiplier/STAGE2/pp2_31_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_32_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_32_1/_19_  (.A1(\u_multiplier/pp1_32 [1]),
    .A2(\u_multiplier/pp1_32 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_32_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_32_1/_20_  (.A(\u_multiplier/pp1_32 [1]),
    .B(\u_multiplier/pp1_32 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_32_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_32_1/_21_  (.A1(\u_multiplier/pp1_32 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_32_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_32_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_32_1/_22_  (.A(\u_multiplier/pp1_32 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_32_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_32_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_32_1/_23_  (.A1(\u_multiplier/pp1_32 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_32_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_32_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_32_1/_24_  (.A(\u_multiplier/pp1_32 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_32_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_32_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_32_1/_25_  (.A(\u_multiplier/STAGE2/pp2_31_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_32_1/_16_ ),
    .ZN(\u_multiplier/pp2_32 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_32_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_32_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_32_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_32_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_32_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_32_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_32_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_32_1/_17_ ),
    .ZN(\u_multiplier/pp2_33 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_32_2/_18_  (.A(\u_multiplier/STAGE2/pp2_31_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_32_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_32_2/_19_  (.A1(\u_multiplier/pp1_32 [5]),
    .A2(\u_multiplier/pp1_32 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_32_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_32_2/_20_  (.A(\u_multiplier/pp1_32 [5]),
    .B(\u_multiplier/pp1_32 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_32_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_32_2/_21_  (.A1(\u_multiplier/pp1_32 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_32_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_32_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_32_2/_22_  (.A(\u_multiplier/pp1_32 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_32_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_32_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_32_2/_23_  (.A1(\u_multiplier/pp1_32 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_32_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_32_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_32_2/_24_  (.A(\u_multiplier/pp1_32 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_32_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_32_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_32_2/_25_  (.A(\u_multiplier/STAGE2/pp2_31_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_32_2/_16_ ),
    .ZN(\u_multiplier/pp2_32 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_32_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_32_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_32_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_32_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_32_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_32_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_32_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_32_2/_17_ ),
    .ZN(\u_multiplier/pp2_33 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_32_3/_18_  (.A(\u_multiplier/STAGE2/pp2_31_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_32_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_32_3/_19_  (.A1(\u_multiplier/pp1_32 [9]),
    .A2(\u_multiplier/pp1_32 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_32_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_32_3/_20_  (.A(\u_multiplier/pp1_32 [9]),
    .B(\u_multiplier/pp1_32 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_32_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_32_3/_21_  (.A1(\u_multiplier/pp1_32 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_32_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_32_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_32_3/_22_  (.A(\u_multiplier/pp1_32 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_32_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_32_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_32_3/_23_  (.A1(\u_multiplier/pp1_32 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_32_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_32_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_32_3/_24_  (.A(\u_multiplier/pp1_32 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_32_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_32_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_32_3/_25_  (.A(\u_multiplier/STAGE2/pp2_31_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_32_3/_16_ ),
    .ZN(\u_multiplier/pp2_32 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_32_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_32_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_32_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_32_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_32_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_32_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_32_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_32_3/_17_ ),
    .ZN(\u_multiplier/pp2_33 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_32_4/_18_  (.A(\u_multiplier/STAGE2/pp2_31_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_32_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_32_4/_19_  (.A1(\u_multiplier/pp1_32 [13]),
    .A2(\u_multiplier/pp1_32 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_32_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_32_4/_20_  (.A(\u_multiplier/pp1_32 [13]),
    .B(\u_multiplier/pp1_32 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_32_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_32_4/_21_  (.A1(\u_multiplier/pp1_32 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_32_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_32_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_32_4/_22_  (.A(\u_multiplier/pp1_32 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_32_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_32_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_32_4/_23_  (.A1(\u_multiplier/pp1_32 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_32_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_32_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_32_4/_24_  (.A(\u_multiplier/pp1_32 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_32_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_32_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_32_4/_25_  (.A(\u_multiplier/STAGE2/pp2_31_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_32_4/_16_ ),
    .ZN(\u_multiplier/pp2_32 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_32_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_32_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_32_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_32_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_32_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_32_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_32_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_32_4/_17_ ),
    .ZN(\u_multiplier/pp2_33 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_33_1/_18_  (.A(\u_multiplier/STAGE2/pp2_32_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_33_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_33_1/_19_  (.A1(\u_multiplier/pp1_33 [1]),
    .A2(\u_multiplier/pp1_33 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_33_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_33_1/_20_  (.A(\u_multiplier/pp1_33 [1]),
    .B(\u_multiplier/pp1_33 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_33_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_33_1/_21_  (.A1(\u_multiplier/pp1_33 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_33_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_33_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_33_1/_22_  (.A(\u_multiplier/pp1_33 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_33_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_33_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_33_1/_23_  (.A1(\u_multiplier/pp1_33 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_33_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_33_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_33_1/_24_  (.A(\u_multiplier/pp1_33 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_33_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_33_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_33_1/_25_  (.A(\u_multiplier/STAGE2/pp2_32_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_33_1/_16_ ),
    .ZN(\u_multiplier/pp2_33 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_33_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_33_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_33_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_33_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_33_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_33_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_33_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_33_1/_17_ ),
    .ZN(\u_multiplier/pp2_34 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_33_2/_18_  (.A(\u_multiplier/STAGE2/pp2_32_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_33_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_33_2/_19_  (.A1(\u_multiplier/pp1_33 [5]),
    .A2(\u_multiplier/pp1_33 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_33_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_33_2/_20_  (.A(\u_multiplier/pp1_33 [5]),
    .B(\u_multiplier/pp1_33 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_33_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_33_2/_21_  (.A1(\u_multiplier/pp1_33 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_33_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_33_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_33_2/_22_  (.A(\u_multiplier/pp1_33 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_33_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_33_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_33_2/_23_  (.A1(\u_multiplier/pp1_33 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_33_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_33_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_33_2/_24_  (.A(\u_multiplier/pp1_33 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_33_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_33_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_33_2/_25_  (.A(\u_multiplier/STAGE2/pp2_32_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_33_2/_16_ ),
    .ZN(\u_multiplier/pp2_33 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_33_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_33_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_33_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_33_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_33_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_33_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_33_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_33_2/_17_ ),
    .ZN(\u_multiplier/pp2_34 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_33_3/_18_  (.A(\u_multiplier/STAGE2/pp2_32_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_33_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_33_3/_19_  (.A1(\u_multiplier/pp1_33 [9]),
    .A2(\u_multiplier/pp1_33 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_33_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_33_3/_20_  (.A(\u_multiplier/pp1_33 [9]),
    .B(\u_multiplier/pp1_33 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_33_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_33_3/_21_  (.A1(\u_multiplier/pp1_33 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_33_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_33_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_33_3/_22_  (.A(\u_multiplier/pp1_33 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_33_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_33_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_33_3/_23_  (.A1(\u_multiplier/pp1_33 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_33_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_33_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_33_3/_24_  (.A(\u_multiplier/pp1_33 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_33_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_33_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_33_3/_25_  (.A(\u_multiplier/STAGE2/pp2_32_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_33_3/_16_ ),
    .ZN(\u_multiplier/pp2_33 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_33_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_33_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_33_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_33_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_33_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_33_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_33_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_33_3/_17_ ),
    .ZN(\u_multiplier/pp2_34 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_33_4/_18_  (.A(\u_multiplier/STAGE2/pp2_32_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_33_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_33_4/_19_  (.A1(\u_multiplier/pp1_33 [13]),
    .A2(\u_multiplier/pp1_33 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_33_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_33_4/_20_  (.A(\u_multiplier/pp1_33 [13]),
    .B(\u_multiplier/pp1_33 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_33_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_33_4/_21_  (.A1(\u_multiplier/pp1_33 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_33_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_33_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_33_4/_22_  (.A(\u_multiplier/pp1_33 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_33_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_33_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_33_4/_23_  (.A1(\u_multiplier/pp1_33 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_33_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_33_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_33_4/_24_  (.A(\u_multiplier/pp1_33 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_33_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_33_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_33_4/_25_  (.A(\u_multiplier/STAGE2/pp2_32_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_33_4/_16_ ),
    .ZN(\u_multiplier/pp2_33 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_33_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_33_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_33_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_33_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_33_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_33_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_33_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_33_4/_17_ ),
    .ZN(\u_multiplier/pp2_34 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_34_1/_18_  (.A(\u_multiplier/STAGE2/pp2_33_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_34_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_34_1/_19_  (.A1(\u_multiplier/pp1_34 [1]),
    .A2(\u_multiplier/pp1_34 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_34_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_34_1/_20_  (.A(\u_multiplier/pp1_34 [1]),
    .B(\u_multiplier/pp1_34 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_34_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_34_1/_21_  (.A1(\u_multiplier/pp1_34 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_34_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_34_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_34_1/_22_  (.A(\u_multiplier/pp1_34 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_34_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_34_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_34_1/_23_  (.A1(\u_multiplier/pp1_34 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_34_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_34_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_34_1/_24_  (.A(\u_multiplier/pp1_34 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_34_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_34_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_34_1/_25_  (.A(\u_multiplier/STAGE2/pp2_33_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_34_1/_16_ ),
    .ZN(\u_multiplier/pp2_34 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_34_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_34_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_34_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_34_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_34_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_34_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_34_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_34_1/_17_ ),
    .ZN(\u_multiplier/pp2_35 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_34_2/_18_  (.A(\u_multiplier/STAGE2/pp2_33_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_34_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_34_2/_19_  (.A1(\u_multiplier/pp1_34 [5]),
    .A2(\u_multiplier/pp1_34 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_34_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_34_2/_20_  (.A(\u_multiplier/pp1_34 [5]),
    .B(\u_multiplier/pp1_34 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_34_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_34_2/_21_  (.A1(\u_multiplier/pp1_34 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_34_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_34_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_34_2/_22_  (.A(\u_multiplier/pp1_34 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_34_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_34_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_34_2/_23_  (.A1(\u_multiplier/pp1_34 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_34_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_34_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_34_2/_24_  (.A(\u_multiplier/pp1_34 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_34_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_34_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_34_2/_25_  (.A(\u_multiplier/STAGE2/pp2_33_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_34_2/_16_ ),
    .ZN(\u_multiplier/pp2_34 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_34_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_34_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_34_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_34_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_34_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_34_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_34_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_34_2/_17_ ),
    .ZN(\u_multiplier/pp2_35 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_34_3/_18_  (.A(\u_multiplier/STAGE2/pp2_33_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_34_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_34_3/_19_  (.A1(\u_multiplier/pp1_34 [9]),
    .A2(\u_multiplier/pp1_34 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_34_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_34_3/_20_  (.A(\u_multiplier/pp1_34 [9]),
    .B(\u_multiplier/pp1_34 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_34_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_34_3/_21_  (.A1(\u_multiplier/pp1_34 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_34_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_34_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_34_3/_22_  (.A(\u_multiplier/pp1_34 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_34_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_34_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_34_3/_23_  (.A1(\u_multiplier/pp1_34 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_34_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_34_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_34_3/_24_  (.A(\u_multiplier/pp1_34 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_34_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_34_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_34_3/_25_  (.A(\u_multiplier/STAGE2/pp2_33_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_34_3/_16_ ),
    .ZN(\u_multiplier/pp2_34 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_34_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_34_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_34_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_34_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_34_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_34_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_34_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_34_3/_17_ ),
    .ZN(\u_multiplier/pp2_35 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_34_4/_18_  (.A(\u_multiplier/STAGE2/pp2_33_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_34_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_34_4/_19_  (.A1(\u_multiplier/pp1_34 [13]),
    .A2(\u_multiplier/pp1_34 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_34_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_34_4/_20_  (.A(\u_multiplier/pp1_34 [13]),
    .B(\u_multiplier/pp1_34 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_34_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_34_4/_21_  (.A1(\u_multiplier/pp1_34 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_34_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_34_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_34_4/_22_  (.A(\u_multiplier/pp1_34 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_34_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_34_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_34_4/_23_  (.A1(\u_multiplier/pp1_34 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_34_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_34_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_34_4/_24_  (.A(\u_multiplier/pp1_34 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_34_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_34_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_34_4/_25_  (.A(\u_multiplier/STAGE2/pp2_33_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_34_4/_16_ ),
    .ZN(\u_multiplier/pp2_34 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_34_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_34_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_34_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_34_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_34_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_34_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_34_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_34_4/_17_ ),
    .ZN(\u_multiplier/pp2_35 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_35_1/_18_  (.A(\u_multiplier/STAGE2/pp2_34_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_35_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_35_1/_19_  (.A1(\u_multiplier/pp1_35 [1]),
    .A2(\u_multiplier/pp1_35 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_35_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_35_1/_20_  (.A(\u_multiplier/pp1_35 [1]),
    .B(\u_multiplier/pp1_35 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_35_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_35_1/_21_  (.A1(\u_multiplier/pp1_35 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_35_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_35_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_35_1/_22_  (.A(\u_multiplier/pp1_35 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_35_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_35_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_35_1/_23_  (.A1(\u_multiplier/pp1_35 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_35_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_35_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_35_1/_24_  (.A(\u_multiplier/pp1_35 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_35_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_35_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_35_1/_25_  (.A(\u_multiplier/STAGE2/pp2_34_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_35_1/_16_ ),
    .ZN(\u_multiplier/pp2_35 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_35_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_35_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_35_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_35_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_35_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_35_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_35_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_35_1/_17_ ),
    .ZN(\u_multiplier/pp2_36 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_35_2/_18_  (.A(\u_multiplier/STAGE2/pp2_34_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_35_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_35_2/_19_  (.A1(\u_multiplier/pp1_35 [5]),
    .A2(\u_multiplier/pp1_35 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_35_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_35_2/_20_  (.A(\u_multiplier/pp1_35 [5]),
    .B(\u_multiplier/pp1_35 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_35_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_35_2/_21_  (.A1(\u_multiplier/pp1_35 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_35_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_35_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_35_2/_22_  (.A(\u_multiplier/pp1_35 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_35_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_35_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_35_2/_23_  (.A1(\u_multiplier/pp1_35 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_35_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_35_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_35_2/_24_  (.A(\u_multiplier/pp1_35 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_35_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_35_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_35_2/_25_  (.A(\u_multiplier/STAGE2/pp2_34_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_35_2/_16_ ),
    .ZN(\u_multiplier/pp2_35 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_35_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_35_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_35_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_35_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_35_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_35_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_35_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_35_2/_17_ ),
    .ZN(\u_multiplier/pp2_36 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_35_3/_18_  (.A(\u_multiplier/STAGE2/pp2_34_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_35_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_35_3/_19_  (.A1(\u_multiplier/pp1_35 [9]),
    .A2(\u_multiplier/pp1_35 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_35_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_35_3/_20_  (.A(\u_multiplier/pp1_35 [9]),
    .B(\u_multiplier/pp1_35 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_35_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_35_3/_21_  (.A1(\u_multiplier/pp1_35 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_35_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_35_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_35_3/_22_  (.A(\u_multiplier/pp1_35 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_35_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_35_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_35_3/_23_  (.A1(\u_multiplier/pp1_35 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_35_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_35_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_35_3/_24_  (.A(\u_multiplier/pp1_35 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_35_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_35_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_35_3/_25_  (.A(\u_multiplier/STAGE2/pp2_34_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_35_3/_16_ ),
    .ZN(\u_multiplier/pp2_35 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_35_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_35_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_35_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_35_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_35_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_35_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_35_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_35_3/_17_ ),
    .ZN(\u_multiplier/pp2_36 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_35_4/_18_  (.A(\u_multiplier/STAGE2/pp2_34_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_35_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_35_4/_19_  (.A1(\u_multiplier/pp1_35 [13]),
    .A2(\u_multiplier/pp1_35 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_35_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_35_4/_20_  (.A(\u_multiplier/pp1_35 [13]),
    .B(\u_multiplier/pp1_35 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_35_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_35_4/_21_  (.A1(\u_multiplier/pp1_35 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_35_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_35_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_35_4/_22_  (.A(\u_multiplier/pp1_35 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_35_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_35_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_35_4/_23_  (.A1(\u_multiplier/pp1_35 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_35_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_35_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_35_4/_24_  (.A(\u_multiplier/pp1_35 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_35_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_35_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_35_4/_25_  (.A(\u_multiplier/STAGE2/pp2_34_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_35_4/_16_ ),
    .ZN(\u_multiplier/pp2_35 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_35_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_35_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_35_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_35_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_35_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_35_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_35_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_35_4/_17_ ),
    .ZN(\u_multiplier/pp2_36 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_36_1/_18_  (.A(\u_multiplier/STAGE2/pp2_35_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_36_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_36_1/_19_  (.A1(\u_multiplier/pp1_36 [1]),
    .A2(\u_multiplier/pp1_36 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_36_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_36_1/_20_  (.A(\u_multiplier/pp1_36 [1]),
    .B(\u_multiplier/pp1_36 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_36_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_36_1/_21_  (.A1(\u_multiplier/pp1_36 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_36_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_36_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_36_1/_22_  (.A(\u_multiplier/pp1_36 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_36_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_36_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_36_1/_23_  (.A1(\u_multiplier/pp1_36 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_36_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_36_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_36_1/_24_  (.A(\u_multiplier/pp1_36 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_36_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_36_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_36_1/_25_  (.A(\u_multiplier/STAGE2/pp2_35_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_36_1/_16_ ),
    .ZN(\u_multiplier/pp2_36 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_36_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_36_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_36_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_36_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_36_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_36_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_36_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_36_1/_17_ ),
    .ZN(\u_multiplier/pp2_37 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_36_2/_18_  (.A(\u_multiplier/STAGE2/pp2_35_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_36_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_36_2/_19_  (.A1(\u_multiplier/pp1_36 [5]),
    .A2(\u_multiplier/pp1_36 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_36_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_36_2/_20_  (.A(\u_multiplier/pp1_36 [5]),
    .B(\u_multiplier/pp1_36 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_36_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_36_2/_21_  (.A1(\u_multiplier/pp1_36 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_36_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_36_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_36_2/_22_  (.A(\u_multiplier/pp1_36 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_36_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_36_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_36_2/_23_  (.A1(\u_multiplier/pp1_36 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_36_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_36_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_36_2/_24_  (.A(\u_multiplier/pp1_36 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_36_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_36_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_36_2/_25_  (.A(\u_multiplier/STAGE2/pp2_35_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_36_2/_16_ ),
    .ZN(\u_multiplier/pp2_36 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_36_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_36_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_36_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_36_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_36_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_36_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_36_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_36_2/_17_ ),
    .ZN(\u_multiplier/pp2_37 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_36_3/_18_  (.A(\u_multiplier/STAGE2/pp2_35_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_36_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_36_3/_19_  (.A1(\u_multiplier/pp1_36 [9]),
    .A2(\u_multiplier/pp1_36 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_36_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_36_3/_20_  (.A(\u_multiplier/pp1_36 [9]),
    .B(\u_multiplier/pp1_36 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_36_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_36_3/_21_  (.A1(\u_multiplier/pp1_36 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_36_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_36_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_36_3/_22_  (.A(\u_multiplier/pp1_36 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_36_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_36_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_36_3/_23_  (.A1(\u_multiplier/pp1_36 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_36_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_36_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_36_3/_24_  (.A(\u_multiplier/pp1_36 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_36_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_36_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_36_3/_25_  (.A(\u_multiplier/STAGE2/pp2_35_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_36_3/_16_ ),
    .ZN(\u_multiplier/pp2_36 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_36_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_36_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_36_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_36_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_36_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_36_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_36_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_36_3/_17_ ),
    .ZN(\u_multiplier/pp2_37 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_36_4/_18_  (.A(\u_multiplier/STAGE2/pp2_35_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_36_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_36_4/_19_  (.A1(\u_multiplier/pp1_36 [13]),
    .A2(\u_multiplier/pp1_36 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_36_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_36_4/_20_  (.A(\u_multiplier/pp1_36 [13]),
    .B(\u_multiplier/pp1_36 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_36_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_36_4/_21_  (.A1(\u_multiplier/pp1_36 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_36_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_36_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_36_4/_22_  (.A(\u_multiplier/pp1_36 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_36_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_36_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_36_4/_23_  (.A1(\u_multiplier/pp1_36 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_36_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_36_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_36_4/_24_  (.A(\u_multiplier/pp1_36 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_36_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_36_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_36_4/_25_  (.A(\u_multiplier/STAGE2/pp2_35_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_36_4/_16_ ),
    .ZN(\u_multiplier/pp2_36 [0]));
 NAND2_X2 \u_multiplier/STAGE2/E_4_2_pp2_36_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_36_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_36_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_36_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_36_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_36_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_36_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_36_4/_17_ ),
    .ZN(\u_multiplier/pp2_37 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_37_1/_18_  (.A(\u_multiplier/STAGE2/pp2_36_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_37_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_37_1/_19_  (.A1(\u_multiplier/pp1_37 [1]),
    .A2(\u_multiplier/pp1_37 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_37_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_37_1/_20_  (.A(\u_multiplier/pp1_37 [1]),
    .B(\u_multiplier/pp1_37 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_37_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_37_1/_21_  (.A1(\u_multiplier/pp1_37 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_37_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_37_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_37_1/_22_  (.A(\u_multiplier/pp1_37 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_37_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_37_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_37_1/_23_  (.A1(\u_multiplier/pp1_37 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_37_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_37_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_37_1/_24_  (.A(\u_multiplier/pp1_37 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_37_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_37_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_37_1/_25_  (.A(\u_multiplier/STAGE2/pp2_36_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_37_1/_16_ ),
    .ZN(\u_multiplier/pp2_37 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_37_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_37_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_37_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_37_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_37_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_37_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_37_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_37_1/_17_ ),
    .ZN(\u_multiplier/pp2_38 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_37_2/_18_  (.A(\u_multiplier/STAGE2/pp2_36_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_37_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_37_2/_19_  (.A1(\u_multiplier/pp1_37 [5]),
    .A2(\u_multiplier/pp1_37 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_37_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_37_2/_20_  (.A(\u_multiplier/pp1_37 [5]),
    .B(\u_multiplier/pp1_37 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_37_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_37_2/_21_  (.A1(\u_multiplier/pp1_37 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_37_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_37_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_37_2/_22_  (.A(\u_multiplier/pp1_37 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_37_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_37_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_37_2/_23_  (.A1(\u_multiplier/pp1_37 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_37_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_37_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_37_2/_24_  (.A(\u_multiplier/pp1_37 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_37_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_37_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_37_2/_25_  (.A(\u_multiplier/STAGE2/pp2_36_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_37_2/_16_ ),
    .ZN(\u_multiplier/pp2_37 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_37_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_37_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_37_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_37_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_37_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_37_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_37_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_37_2/_17_ ),
    .ZN(\u_multiplier/pp2_38 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_37_3/_18_  (.A(\u_multiplier/STAGE2/pp2_36_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_37_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_37_3/_19_  (.A1(\u_multiplier/pp1_37 [9]),
    .A2(\u_multiplier/pp1_37 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_37_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_37_3/_20_  (.A(\u_multiplier/pp1_37 [9]),
    .B(\u_multiplier/pp1_37 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_37_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_37_3/_21_  (.A1(\u_multiplier/pp1_37 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_37_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_37_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_37_3/_22_  (.A(\u_multiplier/pp1_37 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_37_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_37_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_37_3/_23_  (.A1(\u_multiplier/pp1_37 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_37_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_37_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_37_3/_24_  (.A(\u_multiplier/pp1_37 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_37_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_37_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_37_3/_25_  (.A(\u_multiplier/STAGE2/pp2_36_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_37_3/_16_ ),
    .ZN(\u_multiplier/pp2_37 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_37_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_37_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_37_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_37_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_37_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_37_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_37_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_37_3/_17_ ),
    .ZN(\u_multiplier/pp2_38 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_37_4/_18_  (.A(\u_multiplier/STAGE2/pp2_36_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_37_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_37_4/_19_  (.A1(\u_multiplier/pp1_37 [13]),
    .A2(\u_multiplier/pp1_37 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_37_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_37_4/_20_  (.A(\u_multiplier/pp1_37 [13]),
    .B(\u_multiplier/pp1_37 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_37_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_37_4/_21_  (.A1(\u_multiplier/pp1_37 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_37_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_37_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_37_4/_22_  (.A(\u_multiplier/pp1_37 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_37_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_37_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_37_4/_23_  (.A1(\u_multiplier/pp1_37 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_37_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_37_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_37_4/_24_  (.A(\u_multiplier/pp1_37 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_37_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_37_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_37_4/_25_  (.A(\u_multiplier/STAGE2/pp2_36_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_37_4/_16_ ),
    .ZN(\u_multiplier/pp2_37 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_37_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_37_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_37_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_37_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_37_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_37_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_37_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_37_4/_17_ ),
    .ZN(\u_multiplier/pp2_38 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_38_1/_18_  (.A(\u_multiplier/STAGE2/pp2_37_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_38_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_38_1/_19_  (.A1(\u_multiplier/pp1_38 [1]),
    .A2(\u_multiplier/pp1_38 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_38_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_38_1/_20_  (.A(\u_multiplier/pp1_38 [1]),
    .B(\u_multiplier/pp1_38 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_38_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_38_1/_21_  (.A1(\u_multiplier/pp1_38 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_38_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_38_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_38_1/_22_  (.A(\u_multiplier/pp1_38 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_38_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_38_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_38_1/_23_  (.A1(\u_multiplier/pp1_38 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_38_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_38_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_38_1/_24_  (.A(\u_multiplier/pp1_38 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_38_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_38_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_38_1/_25_  (.A(\u_multiplier/STAGE2/pp2_37_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_38_1/_16_ ),
    .ZN(\u_multiplier/pp2_38 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_38_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_38_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_38_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_38_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE2/E_4_2_pp2_38_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_38_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_38_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_38_1/_17_ ),
    .ZN(\u_multiplier/pp2_39 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_38_2/_18_  (.A(\u_multiplier/STAGE2/pp2_37_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_38_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_38_2/_19_  (.A1(\u_multiplier/pp1_38 [5]),
    .A2(\u_multiplier/pp1_38 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_38_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_38_2/_20_  (.A(\u_multiplier/pp1_38 [5]),
    .B(\u_multiplier/pp1_38 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_38_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_38_2/_21_  (.A1(\u_multiplier/pp1_38 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_38_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_38_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_38_2/_22_  (.A(\u_multiplier/pp1_38 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_38_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_38_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_38_2/_23_  (.A1(\u_multiplier/pp1_38 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_38_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_38_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_38_2/_24_  (.A(\u_multiplier/pp1_38 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_38_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_38_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_38_2/_25_  (.A(\u_multiplier/STAGE2/pp2_37_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_38_2/_16_ ),
    .ZN(\u_multiplier/pp2_38 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_38_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_38_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_38_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_38_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_38_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_38_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_38_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_38_2/_17_ ),
    .ZN(\u_multiplier/pp2_39 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_38_3/_18_  (.A(\u_multiplier/STAGE2/pp2_37_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_38_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_38_3/_19_  (.A1(\u_multiplier/pp1_38 [9]),
    .A2(\u_multiplier/pp1_38 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_38_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_38_3/_20_  (.A(\u_multiplier/pp1_38 [9]),
    .B(\u_multiplier/pp1_38 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_38_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_38_3/_21_  (.A1(\u_multiplier/pp1_38 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_38_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_38_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_38_3/_22_  (.A(\u_multiplier/pp1_38 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_38_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_38_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_38_3/_23_  (.A1(\u_multiplier/pp1_38 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_38_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_38_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_38_3/_24_  (.A(\u_multiplier/pp1_38 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_38_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_38_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_38_3/_25_  (.A(\u_multiplier/STAGE2/pp2_37_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_38_3/_16_ ),
    .ZN(\u_multiplier/pp2_38 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_38_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_38_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_38_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_38_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_38_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_38_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_38_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_38_3/_17_ ),
    .ZN(\u_multiplier/pp2_39 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_38_4/_18_  (.A(\u_multiplier/STAGE2/pp2_37_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_38_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_38_4/_19_  (.A1(\u_multiplier/pp1_38 [13]),
    .A2(\u_multiplier/pp1_38 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_38_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_38_4/_20_  (.A(\u_multiplier/pp1_38 [13]),
    .B(\u_multiplier/pp1_38 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_38_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_38_4/_21_  (.A1(\u_multiplier/pp1_38 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_38_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_38_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_38_4/_22_  (.A(\u_multiplier/pp1_38 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_38_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_38_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_38_4/_23_  (.A1(\u_multiplier/pp1_38 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_38_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_38_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_38_4/_24_  (.A(\u_multiplier/pp1_38 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_38_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_38_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_38_4/_25_  (.A(\u_multiplier/STAGE2/pp2_37_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_38_4/_16_ ),
    .ZN(\u_multiplier/pp2_38 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_38_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_38_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_38_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_38_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_38_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_38_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_38_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_38_4/_17_ ),
    .ZN(\u_multiplier/pp2_39 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_39_1/_18_  (.A(\u_multiplier/STAGE2/pp2_38_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_39_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_39_1/_19_  (.A1(\u_multiplier/pp1_39 [1]),
    .A2(\u_multiplier/pp1_39 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_39_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_39_1/_20_  (.A(\u_multiplier/pp1_39 [1]),
    .B(\u_multiplier/pp1_39 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_39_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_39_1/_21_  (.A1(\u_multiplier/pp1_39 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_39_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_39_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_39_1/_22_  (.A(\u_multiplier/pp1_39 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_39_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_39_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_39_1/_23_  (.A1(\u_multiplier/pp1_39 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_39_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_39_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_39_1/_24_  (.A(\u_multiplier/pp1_39 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_39_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_39_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_39_1/_25_  (.A(\u_multiplier/STAGE2/pp2_38_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_39_1/_16_ ),
    .ZN(\u_multiplier/pp2_39 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_39_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_39_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_39_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_39_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_39_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_39_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_39_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_39_1/_17_ ),
    .ZN(\u_multiplier/pp2_40 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_39_2/_18_  (.A(\u_multiplier/STAGE2/pp2_38_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_39_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_39_2/_19_  (.A1(\u_multiplier/pp1_39 [5]),
    .A2(\u_multiplier/pp1_39 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_39_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_39_2/_20_  (.A(\u_multiplier/pp1_39 [5]),
    .B(\u_multiplier/pp1_39 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_39_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_39_2/_21_  (.A1(\u_multiplier/pp1_39 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_39_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_39_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_39_2/_22_  (.A(\u_multiplier/pp1_39 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_39_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_39_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_39_2/_23_  (.A1(\u_multiplier/pp1_39 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_39_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_39_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_39_2/_24_  (.A(\u_multiplier/pp1_39 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_39_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_39_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_39_2/_25_  (.A(\u_multiplier/STAGE2/pp2_38_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_39_2/_16_ ),
    .ZN(\u_multiplier/pp2_39 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_39_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_39_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_39_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_39_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_39_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_39_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_39_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_39_2/_17_ ),
    .ZN(\u_multiplier/pp2_40 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_39_3/_18_  (.A(\u_multiplier/STAGE2/pp2_38_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_39_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_39_3/_19_  (.A1(\u_multiplier/pp1_39 [9]),
    .A2(\u_multiplier/pp1_39 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_39_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_39_3/_20_  (.A(\u_multiplier/pp1_39 [9]),
    .B(\u_multiplier/pp1_39 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_39_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_39_3/_21_  (.A1(\u_multiplier/pp1_39 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_39_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_39_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_39_3/_22_  (.A(\u_multiplier/pp1_39 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_39_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_39_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_39_3/_23_  (.A1(\u_multiplier/pp1_39 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_39_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_39_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_39_3/_24_  (.A(\u_multiplier/pp1_39 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_39_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_39_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_39_3/_25_  (.A(\u_multiplier/STAGE2/pp2_38_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_39_3/_16_ ),
    .ZN(\u_multiplier/pp2_39 [1]));
 NAND2_X2 \u_multiplier/STAGE2/E_4_2_pp2_39_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_39_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_39_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_39_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_39_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_39_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_39_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_39_3/_17_ ),
    .ZN(\u_multiplier/pp2_40 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_39_4/_18_  (.A(\u_multiplier/STAGE2/pp2_38_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_39_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_39_4/_19_  (.A1(\u_multiplier/pp1_39 [13]),
    .A2(\u_multiplier/pp1_39 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_39_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_39_4/_20_  (.A(\u_multiplier/pp1_39 [13]),
    .B(\u_multiplier/pp1_39 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_39_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_39_4/_21_  (.A1(\u_multiplier/pp1_39 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_39_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_39_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_39_4/_22_  (.A(\u_multiplier/pp1_39 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_39_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_39_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_39_4/_23_  (.A1(\u_multiplier/pp1_39 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_39_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_39_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_39_4/_24_  (.A(\u_multiplier/pp1_39 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_39_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_39_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_39_4/_25_  (.A(\u_multiplier/STAGE2/pp2_38_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_39_4/_16_ ),
    .ZN(\u_multiplier/pp2_39 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_39_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_39_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_39_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_39_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_39_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_39_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_39_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_39_4/_17_ ),
    .ZN(\u_multiplier/pp2_40 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_40_1/_18_  (.A(\u_multiplier/STAGE2/pp2_39_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_40_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_40_1/_19_  (.A1(\u_multiplier/pp1_40 [1]),
    .A2(\u_multiplier/pp1_40 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_40_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_40_1/_20_  (.A(\u_multiplier/pp1_40 [1]),
    .B(\u_multiplier/pp1_40 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_40_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_40_1/_21_  (.A1(\u_multiplier/pp1_40 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_40_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_40_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_40_1/_22_  (.A(\u_multiplier/pp1_40 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_40_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_40_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_40_1/_23_  (.A1(\u_multiplier/pp1_40 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_40_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_40_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_40_1/_24_  (.A(\u_multiplier/pp1_40 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_40_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_40_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_40_1/_25_  (.A(\u_multiplier/STAGE2/pp2_39_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_40_1/_16_ ),
    .ZN(\u_multiplier/pp2_40 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_40_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_40_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_40_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_40_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE2/E_4_2_pp2_40_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_40_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_40_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_40_1/_17_ ),
    .ZN(\u_multiplier/pp2_41 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_40_2/_18_  (.A(\u_multiplier/STAGE2/pp2_39_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_40_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_40_2/_19_  (.A1(\u_multiplier/pp1_40 [5]),
    .A2(\u_multiplier/pp1_40 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_40_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_40_2/_20_  (.A(\u_multiplier/pp1_40 [5]),
    .B(\u_multiplier/pp1_40 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_40_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_40_2/_21_  (.A1(\u_multiplier/pp1_40 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_40_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_40_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_40_2/_22_  (.A(\u_multiplier/pp1_40 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_40_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_40_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_40_2/_23_  (.A1(\u_multiplier/pp1_40 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_40_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_40_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_40_2/_24_  (.A(\u_multiplier/pp1_40 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_40_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_40_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_40_2/_25_  (.A(\u_multiplier/STAGE2/pp2_39_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_40_2/_16_ ),
    .ZN(\u_multiplier/pp2_40 [2]));
 NAND2_X2 \u_multiplier/STAGE2/E_4_2_pp2_40_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_40_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_40_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_40_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_40_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_40_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_40_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_40_2/_17_ ),
    .ZN(\u_multiplier/pp2_41 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_40_3/_18_  (.A(\u_multiplier/STAGE2/pp2_39_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_40_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_40_3/_19_  (.A1(\u_multiplier/pp1_40 [9]),
    .A2(\u_multiplier/pp1_40 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_40_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_40_3/_20_  (.A(\u_multiplier/pp1_40 [9]),
    .B(\u_multiplier/pp1_40 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_40_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_40_3/_21_  (.A1(\u_multiplier/pp1_40 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_40_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_40_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_40_3/_22_  (.A(\u_multiplier/pp1_40 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_40_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_40_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_40_3/_23_  (.A1(\u_multiplier/pp1_40 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_40_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_40_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_40_3/_24_  (.A(\u_multiplier/pp1_40 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_40_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_40_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_40_3/_25_  (.A(\u_multiplier/STAGE2/pp2_39_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_40_3/_16_ ),
    .ZN(\u_multiplier/pp2_40 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_40_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_40_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_40_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_40_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_40_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_40_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_40_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_40_3/_17_ ),
    .ZN(\u_multiplier/pp2_41 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_40_4/_18_  (.A(\u_multiplier/STAGE2/pp2_39_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_40_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_40_4/_19_  (.A1(\u_multiplier/pp1_40 [13]),
    .A2(\u_multiplier/pp1_40 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_40_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_40_4/_20_  (.A(\u_multiplier/pp1_40 [13]),
    .B(\u_multiplier/pp1_40 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_40_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_40_4/_21_  (.A1(\u_multiplier/pp1_40 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_40_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_40_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_40_4/_22_  (.A(\u_multiplier/pp1_40 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_40_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_40_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_40_4/_23_  (.A1(\u_multiplier/pp1_40 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_40_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_40_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_40_4/_24_  (.A(\u_multiplier/pp1_40 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_40_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_40_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_40_4/_25_  (.A(\u_multiplier/STAGE2/pp2_39_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_40_4/_16_ ),
    .ZN(\u_multiplier/pp2_40 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_40_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_40_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_40_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_40_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_40_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_40_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_40_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_40_4/_17_ ),
    .ZN(\u_multiplier/pp2_41 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_41_1/_18_  (.A(\u_multiplier/STAGE2/pp2_40_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_41_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_41_1/_19_  (.A1(\u_multiplier/pp1_41 [1]),
    .A2(\u_multiplier/pp1_41 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_41_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_41_1/_20_  (.A(\u_multiplier/pp1_41 [1]),
    .B(\u_multiplier/pp1_41 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_41_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_41_1/_21_  (.A1(\u_multiplier/pp1_41 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_41_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_41_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_41_1/_22_  (.A(\u_multiplier/pp1_41 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_41_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_41_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_41_1/_23_  (.A1(\u_multiplier/pp1_41 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_41_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_41_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_41_1/_24_  (.A(\u_multiplier/pp1_41 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_41_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_41_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_41_1/_25_  (.A(\u_multiplier/STAGE2/pp2_40_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_41_1/_16_ ),
    .ZN(\u_multiplier/pp2_41 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_41_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_41_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_41_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_41_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_41_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_41_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_41_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_41_1/_17_ ),
    .ZN(\u_multiplier/pp2_42 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_41_2/_18_  (.A(\u_multiplier/STAGE2/pp2_40_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_41_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_41_2/_19_  (.A1(\u_multiplier/pp1_41 [5]),
    .A2(\u_multiplier/pp1_41 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_41_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_41_2/_20_  (.A(\u_multiplier/pp1_41 [5]),
    .B(\u_multiplier/pp1_41 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_41_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_41_2/_21_  (.A1(\u_multiplier/pp1_41 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_41_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_41_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_41_2/_22_  (.A(\u_multiplier/pp1_41 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_41_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_41_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_41_2/_23_  (.A1(\u_multiplier/pp1_41 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_41_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_41_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_41_2/_24_  (.A(\u_multiplier/pp1_41 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_41_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_41_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_41_2/_25_  (.A(\u_multiplier/STAGE2/pp2_40_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_41_2/_16_ ),
    .ZN(\u_multiplier/pp2_41 [2]));
 NAND2_X2 \u_multiplier/STAGE2/E_4_2_pp2_41_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_41_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_41_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_41_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_41_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_41_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_41_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_41_2/_17_ ),
    .ZN(\u_multiplier/pp2_42 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_41_3/_18_  (.A(\u_multiplier/STAGE2/pp2_40_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_41_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_41_3/_19_  (.A1(\u_multiplier/pp1_41 [9]),
    .A2(\u_multiplier/pp1_41 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_41_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_41_3/_20_  (.A(\u_multiplier/pp1_41 [9]),
    .B(\u_multiplier/pp1_41 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_41_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_41_3/_21_  (.A1(\u_multiplier/pp1_41 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_41_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_41_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_41_3/_22_  (.A(\u_multiplier/pp1_41 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_41_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_41_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_41_3/_23_  (.A1(\u_multiplier/pp1_41 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_41_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_41_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_41_3/_24_  (.A(\u_multiplier/pp1_41 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_41_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_41_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_41_3/_25_  (.A(\u_multiplier/STAGE2/pp2_40_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_41_3/_16_ ),
    .ZN(\u_multiplier/pp2_41 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_41_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_41_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_41_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_41_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_41_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_41_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_41_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_41_3/_17_ ),
    .ZN(\u_multiplier/pp2_42 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_41_4/_18_  (.A(\u_multiplier/STAGE2/pp2_40_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_41_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_41_4/_19_  (.A1(\u_multiplier/pp1_41 [13]),
    .A2(\u_multiplier/pp1_41 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_41_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_41_4/_20_  (.A(\u_multiplier/pp1_41 [13]),
    .B(\u_multiplier/pp1_41 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_41_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_41_4/_21_  (.A1(\u_multiplier/pp1_41 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_41_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_41_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_41_4/_22_  (.A(\u_multiplier/pp1_41 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_41_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_41_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_41_4/_23_  (.A1(\u_multiplier/pp1_41 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_41_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_41_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_41_4/_24_  (.A(\u_multiplier/pp1_41 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_41_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_41_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_41_4/_25_  (.A(\u_multiplier/STAGE2/pp2_40_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_41_4/_16_ ),
    .ZN(\u_multiplier/pp2_41 [0]));
 NAND2_X2 \u_multiplier/STAGE2/E_4_2_pp2_41_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_41_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_41_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_41_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_41_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_41_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_41_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_41_4/_17_ ),
    .ZN(\u_multiplier/pp2_42 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_42_1/_18_  (.A(\u_multiplier/STAGE2/pp2_41_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_42_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_42_1/_19_  (.A1(\u_multiplier/pp1_42 [1]),
    .A2(\u_multiplier/pp1_42 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_42_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_42_1/_20_  (.A(\u_multiplier/pp1_42 [1]),
    .B(\u_multiplier/pp1_42 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_42_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_42_1/_21_  (.A1(\u_multiplier/pp1_42 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_42_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_42_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_42_1/_22_  (.A(\u_multiplier/pp1_42 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_42_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_42_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_42_1/_23_  (.A1(\u_multiplier/pp1_42 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_42_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_42_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_42_1/_24_  (.A(\u_multiplier/pp1_42 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_42_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_42_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_42_1/_25_  (.A(\u_multiplier/STAGE2/pp2_41_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_42_1/_16_ ),
    .ZN(\u_multiplier/pp2_42 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_42_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_42_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_42_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_42_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE2/E_4_2_pp2_42_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_42_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_42_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_42_1/_17_ ),
    .ZN(\u_multiplier/pp2_43 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_42_2/_18_  (.A(\u_multiplier/STAGE2/pp2_41_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_42_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_42_2/_19_  (.A1(\u_multiplier/pp1_42 [5]),
    .A2(\u_multiplier/pp1_42 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_42_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_42_2/_20_  (.A(\u_multiplier/pp1_42 [5]),
    .B(\u_multiplier/pp1_42 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_42_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_42_2/_21_  (.A1(\u_multiplier/pp1_42 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_42_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_42_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_42_2/_22_  (.A(\u_multiplier/pp1_42 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_42_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_42_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_42_2/_23_  (.A1(\u_multiplier/pp1_42 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_42_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_42_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_42_2/_24_  (.A(\u_multiplier/pp1_42 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_42_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_42_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_42_2/_25_  (.A(\u_multiplier/STAGE2/pp2_41_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_42_2/_16_ ),
    .ZN(\u_multiplier/pp2_42 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_42_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_42_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_42_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_42_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_42_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_42_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_42_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_42_2/_17_ ),
    .ZN(\u_multiplier/pp2_43 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_42_3/_18_  (.A(\u_multiplier/STAGE2/pp2_41_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_42_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_42_3/_19_  (.A1(\u_multiplier/pp1_42 [9]),
    .A2(\u_multiplier/pp1_42 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_42_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_42_3/_20_  (.A(\u_multiplier/pp1_42 [9]),
    .B(\u_multiplier/pp1_42 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_42_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_42_3/_21_  (.A1(\u_multiplier/pp1_42 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_42_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_42_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_42_3/_22_  (.A(\u_multiplier/pp1_42 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_42_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_42_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_42_3/_23_  (.A1(\u_multiplier/pp1_42 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_42_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_42_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_42_3/_24_  (.A(\u_multiplier/pp1_42 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_42_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_42_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_42_3/_25_  (.A(\u_multiplier/STAGE2/pp2_41_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_42_3/_16_ ),
    .ZN(\u_multiplier/pp2_42 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_42_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_42_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_42_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_42_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_42_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_42_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_42_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_42_3/_17_ ),
    .ZN(\u_multiplier/pp2_43 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_42_4/_18_  (.A(\u_multiplier/STAGE2/pp2_41_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_42_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_42_4/_19_  (.A1(\u_multiplier/pp1_42 [13]),
    .A2(\u_multiplier/pp1_42 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_42_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_42_4/_20_  (.A(\u_multiplier/pp1_42 [13]),
    .B(\u_multiplier/pp1_42 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_42_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_42_4/_21_  (.A1(\u_multiplier/pp1_42 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_42_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_42_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_42_4/_22_  (.A(\u_multiplier/pp1_42 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_42_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_42_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_42_4/_23_  (.A1(\u_multiplier/pp1_42 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_42_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_42_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_42_4/_24_  (.A(\u_multiplier/pp1_42 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_42_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_42_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_42_4/_25_  (.A(\u_multiplier/STAGE2/pp2_41_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_42_4/_16_ ),
    .ZN(\u_multiplier/pp2_42 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_42_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_42_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_42_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_42_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_42_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_42_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_42_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_42_4/_17_ ),
    .ZN(\u_multiplier/pp2_43 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_43_1/_18_  (.A(\u_multiplier/STAGE2/pp2_42_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_43_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_43_1/_19_  (.A1(\u_multiplier/pp1_43 [1]),
    .A2(\u_multiplier/pp1_43 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_43_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_43_1/_20_  (.A(\u_multiplier/pp1_43 [1]),
    .B(\u_multiplier/pp1_43 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_43_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_43_1/_21_  (.A1(\u_multiplier/pp1_43 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_43_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_43_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_43_1/_22_  (.A(\u_multiplier/pp1_43 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_43_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_43_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_43_1/_23_  (.A1(\u_multiplier/pp1_43 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_43_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_43_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_43_1/_24_  (.A(\u_multiplier/pp1_43 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_43_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_43_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_43_1/_25_  (.A(\u_multiplier/STAGE2/pp2_42_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_43_1/_16_ ),
    .ZN(\u_multiplier/pp2_43 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_43_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_43_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_43_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_43_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE2/E_4_2_pp2_43_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_43_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_43_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_43_1/_17_ ),
    .ZN(\u_multiplier/pp2_44 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_43_2/_18_  (.A(\u_multiplier/STAGE2/pp2_42_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_43_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_43_2/_19_  (.A1(\u_multiplier/pp1_43 [5]),
    .A2(\u_multiplier/pp1_43 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_43_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_43_2/_20_  (.A(\u_multiplier/pp1_43 [5]),
    .B(\u_multiplier/pp1_43 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_43_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_43_2/_21_  (.A1(\u_multiplier/pp1_43 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_43_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_43_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_43_2/_22_  (.A(\u_multiplier/pp1_43 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_43_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_43_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_43_2/_23_  (.A1(\u_multiplier/pp1_43 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_43_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_43_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_43_2/_24_  (.A(\u_multiplier/pp1_43 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_43_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_43_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_43_2/_25_  (.A(\u_multiplier/STAGE2/pp2_42_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_43_2/_16_ ),
    .ZN(\u_multiplier/pp2_43 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_43_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_43_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_43_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_43_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_43_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_43_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_43_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_43_2/_17_ ),
    .ZN(\u_multiplier/pp2_44 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_43_3/_18_  (.A(\u_multiplier/STAGE2/pp2_42_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_43_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_43_3/_19_  (.A1(\u_multiplier/pp1_43 [9]),
    .A2(\u_multiplier/pp1_43 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_43_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_43_3/_20_  (.A(\u_multiplier/pp1_43 [9]),
    .B(\u_multiplier/pp1_43 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_43_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_43_3/_21_  (.A1(\u_multiplier/pp1_43 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_43_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_43_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_43_3/_22_  (.A(\u_multiplier/pp1_43 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_43_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_43_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_43_3/_23_  (.A1(\u_multiplier/pp1_43 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_43_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_43_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_43_3/_24_  (.A(\u_multiplier/pp1_43 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_43_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_43_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_43_3/_25_  (.A(\u_multiplier/STAGE2/pp2_42_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_43_3/_16_ ),
    .ZN(\u_multiplier/pp2_43 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_43_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_43_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_43_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_43_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_43_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_43_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_43_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_43_3/_17_ ),
    .ZN(\u_multiplier/pp2_44 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_43_4/_18_  (.A(\u_multiplier/STAGE2/pp2_42_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_43_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_43_4/_19_  (.A1(\u_multiplier/pp1_43 [13]),
    .A2(\u_multiplier/pp1_43 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_43_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_43_4/_20_  (.A(\u_multiplier/pp1_43 [13]),
    .B(\u_multiplier/pp1_43 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_43_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_43_4/_21_  (.A1(\u_multiplier/pp1_43 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_43_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_43_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_43_4/_22_  (.A(\u_multiplier/pp1_43 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_43_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_43_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_43_4/_23_  (.A1(\u_multiplier/pp1_43 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_43_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_43_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_43_4/_24_  (.A(\u_multiplier/pp1_43 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_43_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_43_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_43_4/_25_  (.A(\u_multiplier/STAGE2/pp2_42_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_43_4/_16_ ),
    .ZN(\u_multiplier/pp2_43 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_43_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_43_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_43_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_43_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_43_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_43_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_43_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_43_4/_17_ ),
    .ZN(\u_multiplier/pp2_44 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_44_1/_18_  (.A(\u_multiplier/STAGE2/pp2_43_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_44_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_44_1/_19_  (.A1(\u_multiplier/pp1_44 [1]),
    .A2(\u_multiplier/pp1_44 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_44_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_44_1/_20_  (.A(\u_multiplier/pp1_44 [1]),
    .B(\u_multiplier/pp1_44 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_44_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_44_1/_21_  (.A1(\u_multiplier/pp1_44 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_44_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_44_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_44_1/_22_  (.A(\u_multiplier/pp1_44 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_44_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_44_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_44_1/_23_  (.A1(\u_multiplier/pp1_44 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_44_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_44_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_44_1/_24_  (.A(\u_multiplier/pp1_44 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_44_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_44_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_44_1/_25_  (.A(\u_multiplier/STAGE2/pp2_43_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_44_1/_16_ ),
    .ZN(\u_multiplier/pp2_44 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_44_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_44_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_44_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_44_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE2/E_4_2_pp2_44_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_44_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_44_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_44_1/_17_ ),
    .ZN(\u_multiplier/pp2_45 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_44_2/_18_  (.A(\u_multiplier/STAGE2/pp2_43_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_44_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_44_2/_19_  (.A1(\u_multiplier/pp1_44 [5]),
    .A2(\u_multiplier/pp1_44 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_44_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_44_2/_20_  (.A(\u_multiplier/pp1_44 [5]),
    .B(\u_multiplier/pp1_44 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_44_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_44_2/_21_  (.A1(\u_multiplier/pp1_44 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_44_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_44_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_44_2/_22_  (.A(\u_multiplier/pp1_44 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_44_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_44_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_44_2/_23_  (.A1(\u_multiplier/pp1_44 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_44_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_44_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_44_2/_24_  (.A(\u_multiplier/pp1_44 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_44_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_44_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_44_2/_25_  (.A(\u_multiplier/STAGE2/pp2_43_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_44_2/_16_ ),
    .ZN(\u_multiplier/pp2_44 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_44_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_44_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_44_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_44_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_44_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_44_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_44_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_44_2/_17_ ),
    .ZN(\u_multiplier/pp2_45 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_44_3/_18_  (.A(\u_multiplier/STAGE2/pp2_43_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_44_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_44_3/_19_  (.A1(\u_multiplier/pp1_44 [9]),
    .A2(\u_multiplier/pp1_44 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_44_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_44_3/_20_  (.A(\u_multiplier/pp1_44 [9]),
    .B(\u_multiplier/pp1_44 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_44_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_44_3/_21_  (.A1(\u_multiplier/pp1_44 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_44_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_44_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_44_3/_22_  (.A(\u_multiplier/pp1_44 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_44_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_44_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_44_3/_23_  (.A1(\u_multiplier/pp1_44 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_44_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_44_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_44_3/_24_  (.A(\u_multiplier/pp1_44 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_44_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_44_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_44_3/_25_  (.A(\u_multiplier/STAGE2/pp2_43_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_44_3/_16_ ),
    .ZN(\u_multiplier/pp2_44 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_44_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_44_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_44_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_44_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_44_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_44_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_44_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_44_3/_17_ ),
    .ZN(\u_multiplier/pp2_45 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_44_4/_18_  (.A(\u_multiplier/STAGE2/pp2_43_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_44_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_44_4/_19_  (.A1(\u_multiplier/pp1_44 [13]),
    .A2(\u_multiplier/pp1_44 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_44_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_44_4/_20_  (.A(\u_multiplier/pp1_44 [13]),
    .B(\u_multiplier/pp1_44 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_44_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_44_4/_21_  (.A1(\u_multiplier/pp1_44 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_44_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_44_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_44_4/_22_  (.A(\u_multiplier/pp1_44 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_44_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_44_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_44_4/_23_  (.A1(\u_multiplier/pp1_44 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_44_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_44_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_44_4/_24_  (.A(\u_multiplier/pp1_44 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_44_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_44_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_44_4/_25_  (.A(\u_multiplier/STAGE2/pp2_43_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_44_4/_16_ ),
    .ZN(\u_multiplier/pp2_44 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_44_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_44_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_44_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_44_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_44_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_44_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_44_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_44_4/_17_ ),
    .ZN(\u_multiplier/pp2_45 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_45_1/_18_  (.A(\u_multiplier/STAGE2/pp2_44_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_45_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_45_1/_19_  (.A1(\u_multiplier/pp1_45 [1]),
    .A2(\u_multiplier/pp1_45 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_45_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_45_1/_20_  (.A(\u_multiplier/pp1_45 [1]),
    .B(\u_multiplier/pp1_45 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_45_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_45_1/_21_  (.A1(\u_multiplier/pp1_45 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_45_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_45_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_45_1/_22_  (.A(\u_multiplier/pp1_45 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_45_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_45_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_45_1/_23_  (.A1(\u_multiplier/pp1_45 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_45_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_45_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_45_1/_24_  (.A(\u_multiplier/pp1_45 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_45_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_45_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_45_1/_25_  (.A(\u_multiplier/STAGE2/pp2_44_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_45_1/_16_ ),
    .ZN(\u_multiplier/pp2_45 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_45_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_45_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_45_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_45_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_45_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_45_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_45_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_45_1/_17_ ),
    .ZN(\u_multiplier/pp2_46 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_45_2/_18_  (.A(\u_multiplier/STAGE2/pp2_44_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_45_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_45_2/_19_  (.A1(\u_multiplier/pp1_45 [5]),
    .A2(\u_multiplier/pp1_45 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_45_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_45_2/_20_  (.A(\u_multiplier/pp1_45 [5]),
    .B(\u_multiplier/pp1_45 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_45_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_45_2/_21_  (.A1(\u_multiplier/pp1_45 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_45_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_45_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_45_2/_22_  (.A(\u_multiplier/pp1_45 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_45_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_45_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_45_2/_23_  (.A1(\u_multiplier/pp1_45 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_45_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_45_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_45_2/_24_  (.A(\u_multiplier/pp1_45 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_45_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_45_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_45_2/_25_  (.A(\u_multiplier/STAGE2/pp2_44_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_45_2/_16_ ),
    .ZN(\u_multiplier/pp2_45 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_45_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_45_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_45_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_45_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_45_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_45_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_45_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_45_2/_17_ ),
    .ZN(\u_multiplier/pp2_46 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_45_3/_18_  (.A(\u_multiplier/STAGE2/pp2_44_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_45_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_45_3/_19_  (.A1(\u_multiplier/pp1_45 [9]),
    .A2(\u_multiplier/pp1_45 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_45_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_45_3/_20_  (.A(\u_multiplier/pp1_45 [9]),
    .B(\u_multiplier/pp1_45 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_45_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_45_3/_21_  (.A1(\u_multiplier/pp1_45 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_45_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_45_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_45_3/_22_  (.A(\u_multiplier/pp1_45 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_45_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_45_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_45_3/_23_  (.A1(\u_multiplier/pp1_45 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_45_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_45_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_45_3/_24_  (.A(\u_multiplier/pp1_45 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_45_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_45_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_45_3/_25_  (.A(\u_multiplier/STAGE2/pp2_44_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_45_3/_16_ ),
    .ZN(\u_multiplier/pp2_45 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_45_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_45_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_45_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_45_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_45_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_45_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_45_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_45_3/_17_ ),
    .ZN(\u_multiplier/pp2_46 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_45_4/_18_  (.A(\u_multiplier/STAGE2/pp2_44_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_45_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_45_4/_19_  (.A1(\u_multiplier/pp1_45 [13]),
    .A2(\u_multiplier/pp1_45 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_45_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_45_4/_20_  (.A(\u_multiplier/pp1_45 [13]),
    .B(\u_multiplier/pp1_45 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_45_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_45_4/_21_  (.A1(\u_multiplier/pp1_45 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_45_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_45_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_45_4/_22_  (.A(\u_multiplier/pp1_45 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_45_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_45_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_45_4/_23_  (.A1(\u_multiplier/pp1_45 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_45_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_45_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_45_4/_24_  (.A(\u_multiplier/pp1_45 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_45_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_45_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_45_4/_25_  (.A(\u_multiplier/STAGE2/pp2_44_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_45_4/_16_ ),
    .ZN(\u_multiplier/pp2_45 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_45_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_45_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_45_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_45_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_45_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_45_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_45_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_45_4/_17_ ),
    .ZN(\u_multiplier/pp2_46 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_46_1/_18_  (.A(\u_multiplier/STAGE2/pp2_45_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_46_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_46_1/_19_  (.A1(\u_multiplier/pp1_46 [1]),
    .A2(\u_multiplier/pp1_46 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_46_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_46_1/_20_  (.A(\u_multiplier/pp1_46 [1]),
    .B(\u_multiplier/pp1_46 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_46_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_46_1/_21_  (.A1(\u_multiplier/pp1_46 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_46_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_46_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_46_1/_22_  (.A(\u_multiplier/pp1_46 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_46_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_46_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_46_1/_23_  (.A1(\u_multiplier/pp1_46 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_46_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_46_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_46_1/_24_  (.A(\u_multiplier/pp1_46 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_46_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_46_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_46_1/_25_  (.A(\u_multiplier/STAGE2/pp2_45_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_46_1/_16_ ),
    .ZN(\u_multiplier/pp2_46 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_46_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_46_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_46_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_46_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_46_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_46_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_46_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_46_1/_17_ ),
    .ZN(\u_multiplier/pp2_47 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_46_2/_18_  (.A(\u_multiplier/STAGE2/pp2_45_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_46_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_46_2/_19_  (.A1(\u_multiplier/pp1_46 [5]),
    .A2(\u_multiplier/pp1_46 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_46_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_46_2/_20_  (.A(\u_multiplier/pp1_46 [5]),
    .B(\u_multiplier/pp1_46 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_46_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_46_2/_21_  (.A1(\u_multiplier/pp1_46 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_46_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_46_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_46_2/_22_  (.A(\u_multiplier/pp1_46 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_46_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_46_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_46_2/_23_  (.A1(\u_multiplier/pp1_46 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_46_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_46_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_46_2/_24_  (.A(\u_multiplier/pp1_46 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_46_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_46_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_46_2/_25_  (.A(\u_multiplier/STAGE2/pp2_45_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_46_2/_16_ ),
    .ZN(\u_multiplier/pp2_46 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_46_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_46_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_46_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_46_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_46_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_46_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_46_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_46_2/_17_ ),
    .ZN(\u_multiplier/pp2_47 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_46_3/_18_  (.A(\u_multiplier/STAGE2/pp2_45_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_46_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_46_3/_19_  (.A1(\u_multiplier/pp1_46 [9]),
    .A2(\u_multiplier/pp1_46 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_46_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_46_3/_20_  (.A(\u_multiplier/pp1_46 [9]),
    .B(\u_multiplier/pp1_46 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_46_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_46_3/_21_  (.A1(\u_multiplier/pp1_46 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_46_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_46_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_46_3/_22_  (.A(\u_multiplier/pp1_46 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_46_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_46_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_46_3/_23_  (.A1(\u_multiplier/pp1_46 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_46_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_46_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_46_3/_24_  (.A(\u_multiplier/pp1_46 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_46_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_46_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_46_3/_25_  (.A(\u_multiplier/STAGE2/pp2_45_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_46_3/_16_ ),
    .ZN(\u_multiplier/pp2_46 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_46_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_46_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_46_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_46_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_46_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_46_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_46_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_46_3/_17_ ),
    .ZN(\u_multiplier/pp2_47 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_46_4/_18_  (.A(\u_multiplier/STAGE2/pp2_45_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_46_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_46_4/_19_  (.A1(\u_multiplier/pp1_46 [13]),
    .A2(\u_multiplier/pp1_46 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_46_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_46_4/_20_  (.A(\u_multiplier/pp1_46 [13]),
    .B(\u_multiplier/pp1_46 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_46_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_46_4/_21_  (.A1(\u_multiplier/pp1_46 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_46_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_46_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_46_4/_22_  (.A(\u_multiplier/pp1_46 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_46_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_46_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_46_4/_23_  (.A1(\u_multiplier/pp1_46 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_46_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_46_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_46_4/_24_  (.A(\u_multiplier/pp1_46 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_46_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_46_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_46_4/_25_  (.A(\u_multiplier/STAGE2/pp2_45_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_46_4/_16_ ),
    .ZN(\u_multiplier/pp2_46 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_46_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_46_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_46_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_46_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_46_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_46_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_46_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_46_4/_17_ ),
    .ZN(\u_multiplier/pp2_47 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_47_1/_18_  (.A(\u_multiplier/STAGE2/pp2_46_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_47_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_47_1/_19_  (.A1(\u_multiplier/pp1_47 [1]),
    .A2(\u_multiplier/pp1_47 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_47_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_47_1/_20_  (.A(\u_multiplier/pp1_47 [1]),
    .B(\u_multiplier/pp1_47 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_47_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_47_1/_21_  (.A1(\u_multiplier/pp1_47 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_47_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_47_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_47_1/_22_  (.A(\u_multiplier/pp1_47 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_47_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_47_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_47_1/_23_  (.A1(\u_multiplier/pp1_47 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_47_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_47_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_47_1/_24_  (.A(\u_multiplier/pp1_47 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_47_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_47_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_47_1/_25_  (.A(\u_multiplier/STAGE2/pp2_46_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_47_1/_16_ ),
    .ZN(\u_multiplier/pp2_47 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_47_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_47_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_47_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_47_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_47_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_47_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_47_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_47_1/_17_ ),
    .ZN(\u_multiplier/pp2_48 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_47_2/_18_  (.A(\u_multiplier/STAGE2/pp2_46_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_47_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_47_2/_19_  (.A1(\u_multiplier/pp1_47 [5]),
    .A2(\u_multiplier/pp1_47 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_47_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_47_2/_20_  (.A(\u_multiplier/pp1_47 [5]),
    .B(\u_multiplier/pp1_47 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_47_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_47_2/_21_  (.A1(\u_multiplier/pp1_47 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_47_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_47_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_47_2/_22_  (.A(\u_multiplier/pp1_47 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_47_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_47_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_47_2/_23_  (.A1(\u_multiplier/pp1_47 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_47_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_47_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_47_2/_24_  (.A(\u_multiplier/pp1_47 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_47_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_47_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_47_2/_25_  (.A(\u_multiplier/STAGE2/pp2_46_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_47_2/_16_ ),
    .ZN(\u_multiplier/pp2_47 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_47_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_47_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_47_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_47_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_47_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_47_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_47_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_47_2/_17_ ),
    .ZN(\u_multiplier/pp2_48 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_47_3/_18_  (.A(\u_multiplier/STAGE2/pp2_46_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_47_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_47_3/_19_  (.A1(\u_multiplier/pp1_47 [9]),
    .A2(\u_multiplier/pp1_47 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_47_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_47_3/_20_  (.A(\u_multiplier/pp1_47 [9]),
    .B(\u_multiplier/pp1_47 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_47_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_47_3/_21_  (.A1(\u_multiplier/pp1_47 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_47_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_47_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_47_3/_22_  (.A(\u_multiplier/pp1_47 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_47_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_47_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_47_3/_23_  (.A1(\u_multiplier/pp1_47 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_47_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_47_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_47_3/_24_  (.A(\u_multiplier/pp1_47 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_47_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_47_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_47_3/_25_  (.A(\u_multiplier/STAGE2/pp2_46_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_47_3/_16_ ),
    .ZN(\u_multiplier/pp2_47 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_47_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_47_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_47_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_47_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_47_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_47_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_47_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_47_3/_17_ ),
    .ZN(\u_multiplier/pp2_48 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_47_4/_18_  (.A(\u_multiplier/STAGE2/pp2_46_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_47_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_47_4/_19_  (.A1(\u_multiplier/pp1_47 [13]),
    .A2(\u_multiplier/pp1_47 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_47_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_47_4/_20_  (.A(\u_multiplier/pp1_47 [13]),
    .B(\u_multiplier/pp1_47 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_47_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_47_4/_21_  (.A1(\u_multiplier/pp1_47 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_47_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_47_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_47_4/_22_  (.A(\u_multiplier/pp1_47 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_47_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_47_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_47_4/_23_  (.A1(\u_multiplier/pp1_47 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_47_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_47_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_47_4/_24_  (.A(\u_multiplier/pp1_47 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_47_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_47_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_47_4/_25_  (.A(\u_multiplier/STAGE2/pp2_46_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_47_4/_16_ ),
    .ZN(\u_multiplier/pp2_47 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_47_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_47_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_47_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_47_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_47_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_47_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_47_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_47_4/_17_ ),
    .ZN(\u_multiplier/pp2_48 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_48_1/_18_  (.A(\u_multiplier/STAGE2/pp2_47_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_48_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_48_1/_19_  (.A1(\u_multiplier/pp1_48 [1]),
    .A2(\u_multiplier/pp1_48 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_48_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_48_1/_20_  (.A(\u_multiplier/pp1_48 [1]),
    .B(\u_multiplier/pp1_48 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_48_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_48_1/_21_  (.A1(\u_multiplier/pp1_48 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_48_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_48_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_48_1/_22_  (.A(\u_multiplier/pp1_48 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_48_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_48_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_48_1/_23_  (.A1(\u_multiplier/pp1_48 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_48_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_48_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_48_1/_24_  (.A(\u_multiplier/pp1_48 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_48_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_48_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_48_1/_25_  (.A(\u_multiplier/STAGE2/pp2_47_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_48_1/_16_ ),
    .ZN(\u_multiplier/pp2_48 [3]));
 NAND2_X2 \u_multiplier/STAGE2/E_4_2_pp2_48_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_48_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_48_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_48_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_48_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_48_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_48_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_48_1/_17_ ),
    .ZN(\u_multiplier/pp2_49 [7]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_48_2/_18_  (.A(\u_multiplier/STAGE2/pp2_47_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_48_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_48_2/_19_  (.A1(\u_multiplier/pp1_48 [5]),
    .A2(\u_multiplier/pp1_48 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_48_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_48_2/_20_  (.A(\u_multiplier/pp1_48 [5]),
    .B(\u_multiplier/pp1_48 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_48_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_48_2/_21_  (.A1(\u_multiplier/pp1_48 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_48_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_48_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_48_2/_22_  (.A(\u_multiplier/pp1_48 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_48_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_48_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_48_2/_23_  (.A1(\u_multiplier/pp1_48 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_48_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_48_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_48_2/_24_  (.A(\u_multiplier/pp1_48 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_48_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_48_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_48_2/_25_  (.A(\u_multiplier/STAGE2/pp2_47_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_48_2/_16_ ),
    .ZN(\u_multiplier/pp2_48 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_48_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_48_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_48_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_48_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_48_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_48_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_48_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_48_2/_17_ ),
    .ZN(\u_multiplier/pp2_49 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_48_3/_18_  (.A(\u_multiplier/STAGE2/pp2_47_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_48_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_48_3/_19_  (.A1(\u_multiplier/pp1_48 [9]),
    .A2(\u_multiplier/pp1_48 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_48_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_48_3/_20_  (.A(\u_multiplier/pp1_48 [9]),
    .B(\u_multiplier/pp1_48 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_48_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_48_3/_21_  (.A1(\u_multiplier/pp1_48 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_48_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_48_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_48_3/_22_  (.A(\u_multiplier/pp1_48 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_48_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_48_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_48_3/_23_  (.A1(\u_multiplier/pp1_48 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_48_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_48_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_48_3/_24_  (.A(\u_multiplier/pp1_48 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_48_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_48_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_48_3/_25_  (.A(\u_multiplier/STAGE2/pp2_47_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_48_3/_16_ ),
    .ZN(\u_multiplier/pp2_48 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_48_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_48_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_48_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_48_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_48_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_48_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_48_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_48_3/_17_ ),
    .ZN(\u_multiplier/pp2_49 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_48_4/_18_  (.A(\u_multiplier/STAGE2/pp2_47_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_48_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_48_4/_19_  (.A1(\u_multiplier/pp1_48 [13]),
    .A2(\u_multiplier/pp1_48 [12]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_48_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_48_4/_20_  (.A(\u_multiplier/pp1_48 [13]),
    .B(\u_multiplier/pp1_48 [12]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_48_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_48_4/_21_  (.A1(\u_multiplier/pp1_48 [14]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_48_4/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_48_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_48_4/_22_  (.A(\u_multiplier/pp1_48 [14]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_48_4/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_48_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_48_4/_23_  (.A1(\u_multiplier/pp1_48 [15]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_48_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_48_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_48_4/_24_  (.A(\u_multiplier/pp1_48 [15]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_48_4/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_48_4/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_48_4/_25_  (.A(\u_multiplier/STAGE2/pp2_47_e42_4_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_48_4/_16_ ),
    .ZN(\u_multiplier/pp2_48 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_48_4/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_48_4/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_48_4/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_48_e42_4_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_48_4/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_48_4/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_48_4/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_48_4/_17_ ),
    .ZN(\u_multiplier/pp2_49 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_49_1/_18_  (.A(\u_multiplier/STAGE2/pp2_48_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_49_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_49_1/_19_  (.A1(\u_multiplier/pp1_49 [1]),
    .A2(\u_multiplier/pp1_49 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_49_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_49_1/_20_  (.A(\u_multiplier/pp1_49 [1]),
    .B(\u_multiplier/pp1_49 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_49_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_49_1/_21_  (.A1(\u_multiplier/pp1_49 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_49_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_49_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_49_1/_22_  (.A(\u_multiplier/pp1_49 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_49_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_49_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_49_1/_23_  (.A1(\u_multiplier/pp1_49 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_49_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_49_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_49_1/_24_  (.A(\u_multiplier/pp1_49 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_49_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_49_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_49_1/_25_  (.A(\u_multiplier/STAGE2/pp2_48_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_49_1/_16_ ),
    .ZN(\u_multiplier/pp2_49 [3]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_49_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_49_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_49_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_49_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_49_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_49_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_49_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_49_1/_17_ ),
    .ZN(\u_multiplier/pp2_50 [6]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_49_2/_18_  (.A(\u_multiplier/STAGE2/pp2_48_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_49_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_49_2/_19_  (.A1(\u_multiplier/pp1_49 [5]),
    .A2(\u_multiplier/pp1_49 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_49_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_49_2/_20_  (.A(\u_multiplier/pp1_49 [5]),
    .B(\u_multiplier/pp1_49 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_49_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_49_2/_21_  (.A1(\u_multiplier/pp1_49 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_49_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_49_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_49_2/_22_  (.A(\u_multiplier/pp1_49 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_49_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_49_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_49_2/_23_  (.A1(\u_multiplier/pp1_49 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_49_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_49_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_49_2/_24_  (.A(\u_multiplier/pp1_49 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_49_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_49_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_49_2/_25_  (.A(\u_multiplier/STAGE2/pp2_48_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_49_2/_16_ ),
    .ZN(\u_multiplier/pp2_49 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_49_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_49_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_49_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_49_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_49_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_49_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_49_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_49_2/_17_ ),
    .ZN(\u_multiplier/pp2_50 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_49_3/_18_  (.A(\u_multiplier/STAGE2/pp2_48_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_49_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_49_3/_19_  (.A1(\u_multiplier/pp1_49 [9]),
    .A2(\u_multiplier/pp1_49 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_49_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_49_3/_20_  (.A(\u_multiplier/pp1_49 [9]),
    .B(\u_multiplier/pp1_49 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_49_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_49_3/_21_  (.A1(\u_multiplier/pp1_49 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_49_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_49_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_49_3/_22_  (.A(\u_multiplier/pp1_49 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_49_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_49_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_49_3/_23_  (.A1(\u_multiplier/pp1_49 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_49_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_49_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_49_3/_24_  (.A(\u_multiplier/pp1_49 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_49_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_49_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_49_3/_25_  (.A(\u_multiplier/STAGE2/pp2_48_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_49_3/_16_ ),
    .ZN(\u_multiplier/pp2_49 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_49_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_49_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_49_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_49_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_49_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_49_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_49_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_49_3/_17_ ),
    .ZN(\u_multiplier/pp2_50 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_50_1/_18_  (.A(\u_multiplier/STAGE2/pp2_49_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_50_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_50_1/_19_  (.A1(\u_multiplier/pp1_50 [1]),
    .A2(\u_multiplier/pp1_50 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_50_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_50_1/_20_  (.A(\u_multiplier/pp1_50 [1]),
    .B(\u_multiplier/pp1_50 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_50_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_50_1/_21_  (.A1(\u_multiplier/pp1_50 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_50_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_50_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_50_1/_22_  (.A(\u_multiplier/pp1_50 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_50_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_50_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_50_1/_23_  (.A1(\u_multiplier/pp1_50 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_50_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_50_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_50_1/_24_  (.A(\u_multiplier/pp1_50 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_50_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_50_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_50_1/_25_  (.A(\u_multiplier/STAGE2/pp2_49_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_50_1/_16_ ),
    .ZN(\u_multiplier/pp2_50 [2]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_50_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_50_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_50_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_50_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_50_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_50_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_50_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_50_1/_17_ ),
    .ZN(\u_multiplier/pp2_51 [5]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_50_2/_18_  (.A(\u_multiplier/STAGE2/pp2_49_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_50_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_50_2/_19_  (.A1(\u_multiplier/pp1_50 [5]),
    .A2(\u_multiplier/pp1_50 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_50_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_50_2/_20_  (.A(\u_multiplier/pp1_50 [5]),
    .B(\u_multiplier/pp1_50 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_50_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_50_2/_21_  (.A1(\u_multiplier/pp1_50 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_50_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_50_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_50_2/_22_  (.A(\u_multiplier/pp1_50 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_50_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_50_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_50_2/_23_  (.A1(\u_multiplier/pp1_50 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_50_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_50_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_50_2/_24_  (.A(\u_multiplier/pp1_50 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_50_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_50_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_50_2/_25_  (.A(\u_multiplier/STAGE2/pp2_49_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_50_2/_16_ ),
    .ZN(\u_multiplier/pp2_50 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_50_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_50_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_50_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_50_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_50_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_50_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_50_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_50_2/_17_ ),
    .ZN(\u_multiplier/pp2_51 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_50_3/_18_  (.A(\u_multiplier/STAGE2/pp2_49_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_50_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_50_3/_19_  (.A1(\u_multiplier/pp1_50 [9]),
    .A2(\u_multiplier/pp1_50 [8]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_50_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_50_3/_20_  (.A(\u_multiplier/pp1_50 [9]),
    .B(\u_multiplier/pp1_50 [8]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_50_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_50_3/_21_  (.A1(\u_multiplier/pp1_50 [10]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_50_3/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_50_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_50_3/_22_  (.A(\u_multiplier/pp1_50 [10]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_50_3/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_50_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_50_3/_23_  (.A1(\u_multiplier/pp1_50 [11]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_50_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_50_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_50_3/_24_  (.A(\u_multiplier/pp1_50 [11]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_50_3/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_50_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_50_3/_25_  (.A(\u_multiplier/STAGE2/pp2_49_e42_3_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_50_3/_16_ ),
    .ZN(\u_multiplier/pp2_50 [0]));
 NAND2_X2 \u_multiplier/STAGE2/E_4_2_pp2_50_3/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_50_3/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_50_3/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_50_e42_3_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_50_3/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_50_3/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_50_3/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_50_3/_17_ ),
    .ZN(\u_multiplier/pp2_51 [3]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_51_1/_18_  (.A(\u_multiplier/STAGE2/pp2_50_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_51_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_51_1/_19_  (.A1(\u_multiplier/pp1_51 [1]),
    .A2(\u_multiplier/pp1_51 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_51_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_51_1/_20_  (.A(\u_multiplier/pp1_51 [1]),
    .B(\u_multiplier/pp1_51 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_51_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_51_1/_21_  (.A1(\u_multiplier/pp1_51 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_51_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_51_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_51_1/_22_  (.A(\u_multiplier/pp1_51 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_51_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_51_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_51_1/_23_  (.A1(\u_multiplier/pp1_51 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_51_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_51_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_51_1/_24_  (.A(\u_multiplier/pp1_51 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_51_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_51_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_51_1/_25_  (.A(\u_multiplier/STAGE2/pp2_50_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_51_1/_16_ ),
    .ZN(\u_multiplier/pp2_51 [2]));
 NAND2_X2 \u_multiplier/STAGE2/E_4_2_pp2_51_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_51_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_51_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_51_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_51_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_51_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_51_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_51_1/_17_ ),
    .ZN(\u_multiplier/pp2_52 [4]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_51_2/_18_  (.A(\u_multiplier/STAGE2/pp2_50_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_51_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_51_2/_19_  (.A1(\u_multiplier/pp1_51 [5]),
    .A2(\u_multiplier/pp1_51 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_51_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_51_2/_20_  (.A(\u_multiplier/pp1_51 [5]),
    .B(\u_multiplier/pp1_51 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_51_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_51_2/_21_  (.A1(\u_multiplier/pp1_51 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_51_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_51_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_51_2/_22_  (.A(\u_multiplier/pp1_51 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_51_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_51_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_51_2/_23_  (.A1(\u_multiplier/pp1_51 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_51_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_51_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_51_2/_24_  (.A(\u_multiplier/pp1_51 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_51_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_51_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_51_2/_25_  (.A(\u_multiplier/STAGE2/pp2_50_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_51_2/_16_ ),
    .ZN(\u_multiplier/pp2_51 [1]));
 NAND2_X2 \u_multiplier/STAGE2/E_4_2_pp2_51_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_51_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_51_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_51_e42_2_cout ));
 OAI21_X1 \u_multiplier/STAGE2/E_4_2_pp2_51_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_51_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_51_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_51_2/_17_ ),
    .ZN(\u_multiplier/pp2_52 [3]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_52_1/_18_  (.A(\u_multiplier/STAGE2/pp2_51_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_52_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_52_1/_19_  (.A1(\u_multiplier/pp1_52 [1]),
    .A2(\u_multiplier/pp1_52 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_52_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_52_1/_20_  (.A(\u_multiplier/pp1_52 [1]),
    .B(\u_multiplier/pp1_52 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_52_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_52_1/_21_  (.A1(\u_multiplier/pp1_52 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_52_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_52_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_52_1/_22_  (.A(\u_multiplier/pp1_52 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_52_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_52_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_52_1/_23_  (.A1(\u_multiplier/pp1_52 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_52_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_52_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_52_1/_24_  (.A(\u_multiplier/pp1_52 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_52_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_52_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_52_1/_25_  (.A(\u_multiplier/STAGE2/pp2_51_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_52_1/_16_ ),
    .ZN(\u_multiplier/pp2_52 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_52_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_52_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_52_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_52_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE2/E_4_2_pp2_52_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_52_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_52_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_52_1/_17_ ),
    .ZN(\u_multiplier/pp2_53 [3]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_52_2/_18_  (.A(\u_multiplier/STAGE2/pp2_51_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_52_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_52_2/_19_  (.A1(\u_multiplier/pp1_52 [5]),
    .A2(\u_multiplier/pp1_52 [4]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_52_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_52_2/_20_  (.A(\u_multiplier/pp1_52 [5]),
    .B(\u_multiplier/pp1_52 [4]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_52_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_52_2/_21_  (.A1(\u_multiplier/pp1_52 [6]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_52_2/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_52_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_52_2/_22_  (.A(\u_multiplier/pp1_52 [6]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_52_2/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_52_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_52_2/_23_  (.A1(\u_multiplier/pp1_52 [7]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_52_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_52_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_52_2/_24_  (.A(\u_multiplier/pp1_52 [7]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_52_2/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_52_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_52_2/_25_  (.A(\u_multiplier/STAGE2/pp2_51_e42_2_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_52_2/_16_ ),
    .ZN(\u_multiplier/pp2_52 [0]));
 NAND2_X2 \u_multiplier/STAGE2/E_4_2_pp2_52_2/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_52_2/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_52_2/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_52_e42_2_cout ));
 OAI21_X4 \u_multiplier/STAGE2/E_4_2_pp2_52_2/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_52_2/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_52_2/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_52_2/_17_ ),
    .ZN(\u_multiplier/pp2_53 [2]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_53_1/_18_  (.A(\u_multiplier/STAGE2/pp2_52_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_53_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_53_1/_19_  (.A1(\u_multiplier/pp1_53 [1]),
    .A2(\u_multiplier/pp1_53 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_53_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_53_1/_20_  (.A(\u_multiplier/pp1_53 [1]),
    .B(\u_multiplier/pp1_53 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_53_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_53_1/_21_  (.A1(\u_multiplier/pp1_53 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_53_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_53_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_53_1/_22_  (.A(\u_multiplier/pp1_53 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_53_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_53_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_53_1/_23_  (.A1(\u_multiplier/pp1_53 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_53_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_53_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_53_1/_24_  (.A(\u_multiplier/pp1_53 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_53_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_53_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_53_1/_25_  (.A(\u_multiplier/STAGE2/pp2_52_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_53_1/_16_ ),
    .ZN(\u_multiplier/pp2_53 [1]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_53_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_53_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_53_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_53_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_53_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_53_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_53_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_53_1/_17_ ),
    .ZN(\u_multiplier/pp2_54 [2]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_54_1/_18_  (.A(\u_multiplier/STAGE2/pp2_53_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_54_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_54_1/_19_  (.A1(\u_multiplier/pp1_54 [1]),
    .A2(\u_multiplier/pp1_54 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_54_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_54_1/_20_  (.A(\u_multiplier/pp1_54 [1]),
    .B(\u_multiplier/pp1_54 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_54_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_54_1/_21_  (.A1(\u_multiplier/pp1_54 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_54_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_54_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_54_1/_22_  (.A(\u_multiplier/pp1_54 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_54_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_54_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_54_1/_23_  (.A1(\u_multiplier/pp1_54 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_54_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_54_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_54_1/_24_  (.A(\u_multiplier/pp1_54 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_54_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_54_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_54_1/_25_  (.A(\u_multiplier/STAGE2/pp2_53_e42_1_cout ),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_54_1/_16_ ),
    .ZN(\u_multiplier/pp2_54 [0]));
 NAND2_X2 \u_multiplier/STAGE2/E_4_2_pp2_54_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_54_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_54_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_54_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_54_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_54_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_54_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_54_1/_17_ ),
    .ZN(\u_multiplier/pp2_55 [1]));
 INV_X1 \u_multiplier/STAGE2/E_4_2_pp2_9_1/_18_  (.A(net138),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_9_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_9_1/_19_  (.A1(\u_multiplier/pp1_9 [1]),
    .A2(\u_multiplier/pp1_9 [0]),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_9_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_9_1/_20_  (.A(\u_multiplier/pp1_9 [1]),
    .B(\u_multiplier/pp1_9 [0]),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_9_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_9_1/_21_  (.A1(\u_multiplier/pp1_9 [2]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_9_1/_12_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_9_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_9_1/_22_  (.A(\u_multiplier/pp1_9 [2]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_9_1/_12_ ),
    .Z(\u_multiplier/STAGE2/E_4_2_pp2_9_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_9_1/_23_  (.A1(\u_multiplier/pp1_9 [3]),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_9_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_9_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_9_1/_24_  (.A(\u_multiplier/pp1_9 [3]),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_9_1/_14_ ),
    .ZN(\u_multiplier/STAGE2/E_4_2_pp2_9_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE2/E_4_2_pp2_9_1/_25_  (.A(net139),
    .B(\u_multiplier/STAGE2/E_4_2_pp2_9_1/_16_ ),
    .ZN(\u_multiplier/pp2_9 [0]));
 NAND2_X1 \u_multiplier/STAGE2/E_4_2_pp2_9_1/_26_  (.A1(\u_multiplier/STAGE2/E_4_2_pp2_9_1/_11_ ),
    .A2(\u_multiplier/STAGE2/E_4_2_pp2_9_1/_13_ ),
    .ZN(\u_multiplier/STAGE2/pp2_9_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE2/E_4_2_pp2_9_1/_27_  (.A(\u_multiplier/STAGE2/E_4_2_pp2_9_1/_15_ ),
    .B1(\u_multiplier/STAGE2/E_4_2_pp2_9_1/_16_ ),
    .B2(\u_multiplier/STAGE2/E_4_2_pp2_9_1/_17_ ),
    .ZN(\u_multiplier/pp2_10 [2]));
 INV_X1 \u_multiplier/STAGE2/Full_adder_pp2_49_1/_12_  (.A(\u_multiplier/STAGE2/pp2_48_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp2_49_1/_08_ ));
 NAND3_X2 \u_multiplier/STAGE2/Full_adder_pp2_49_1/_13_  (.A1(\u_multiplier/pp1_49 [13]),
    .A2(\u_multiplier/pp1_49 [12]),
    .A3(\u_multiplier/STAGE2/pp2_48_e42_4_cout ),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp2_49_1/_09_ ));
 NOR2_X2 \u_multiplier/STAGE2/Full_adder_pp2_49_1/_14_  (.A1(\u_multiplier/pp1_49 [13]),
    .A2(\u_multiplier/pp1_49 [12]),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp2_49_1/_10_ ));
 AOI21_X1 \u_multiplier/STAGE2/Full_adder_pp2_49_1/_15_  (.A(\u_multiplier/STAGE2/pp2_48_e42_4_cout ),
    .B1(\u_multiplier/pp1_49 [12]),
    .B2(\u_multiplier/pp1_49 [13]),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp2_49_1/_11_ ));
 NOR2_X2 \u_multiplier/STAGE2/Full_adder_pp2_49_1/_16_  (.A1(\u_multiplier/STAGE2/Full_adder_pp2_49_1/_10_ ),
    .A2(\u_multiplier/STAGE2/Full_adder_pp2_49_1/_11_ ),
    .ZN(\u_multiplier/pp2_50 [3]));
 AOI22_X4 \u_multiplier/STAGE2/Full_adder_pp2_49_1/_17_  (.A1(\u_multiplier/STAGE2/Full_adder_pp2_49_1/_08_ ),
    .A2(\u_multiplier/STAGE2/Full_adder_pp2_49_1/_10_ ),
    .B1(\u_multiplier/pp2_50 [3]),
    .B2(\u_multiplier/STAGE2/Full_adder_pp2_49_1/_09_ ),
    .ZN(\u_multiplier/pp2_49 [0]));
 INV_X1 \u_multiplier/STAGE2/Full_adder_pp2_51_1/_12_  (.A(\u_multiplier/STAGE2/pp2_50_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp2_51_1/_08_ ));
 NAND3_X2 \u_multiplier/STAGE2/Full_adder_pp2_51_1/_13_  (.A1(\u_multiplier/pp1_51 [9]),
    .A2(\u_multiplier/pp1_51 [8]),
    .A3(\u_multiplier/STAGE2/pp2_50_e42_3_cout ),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp2_51_1/_09_ ));
 NOR2_X4 \u_multiplier/STAGE2/Full_adder_pp2_51_1/_14_  (.A1(\u_multiplier/pp1_51 [9]),
    .A2(\u_multiplier/pp1_51 [8]),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp2_51_1/_10_ ));
 AOI21_X2 \u_multiplier/STAGE2/Full_adder_pp2_51_1/_15_  (.A(\u_multiplier/STAGE2/pp2_50_e42_3_cout ),
    .B1(\u_multiplier/pp1_51 [8]),
    .B2(\u_multiplier/pp1_51 [9]),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp2_51_1/_11_ ));
 NOR2_X4 \u_multiplier/STAGE2/Full_adder_pp2_51_1/_16_  (.A1(\u_multiplier/STAGE2/Full_adder_pp2_51_1/_10_ ),
    .A2(\u_multiplier/STAGE2/Full_adder_pp2_51_1/_11_ ),
    .ZN(\u_multiplier/pp2_52 [2]));
 AOI22_X4 \u_multiplier/STAGE2/Full_adder_pp2_51_1/_17_  (.A1(\u_multiplier/STAGE2/Full_adder_pp2_51_1/_08_ ),
    .A2(\u_multiplier/STAGE2/Full_adder_pp2_51_1/_10_ ),
    .B1(\u_multiplier/pp2_52 [2]),
    .B2(\u_multiplier/STAGE2/Full_adder_pp2_51_1/_09_ ),
    .ZN(\u_multiplier/pp2_51 [0]));
 INV_X1 \u_multiplier/STAGE2/Full_adder_pp2_53_1/_12_  (.A(\u_multiplier/STAGE2/pp2_52_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp2_53_1/_08_ ));
 NAND3_X2 \u_multiplier/STAGE2/Full_adder_pp2_53_1/_13_  (.A1(\u_multiplier/pp1_53 [5]),
    .A2(\u_multiplier/pp1_53 [4]),
    .A3(\u_multiplier/STAGE2/pp2_52_e42_2_cout ),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp2_53_1/_09_ ));
 NOR2_X2 \u_multiplier/STAGE2/Full_adder_pp2_53_1/_14_  (.A1(\u_multiplier/pp1_53 [5]),
    .A2(\u_multiplier/pp1_53 [4]),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp2_53_1/_10_ ));
 AOI21_X1 \u_multiplier/STAGE2/Full_adder_pp2_53_1/_15_  (.A(\u_multiplier/STAGE2/pp2_52_e42_2_cout ),
    .B1(\u_multiplier/pp1_53 [4]),
    .B2(\u_multiplier/pp1_53 [5]),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp2_53_1/_11_ ));
 NOR2_X2 \u_multiplier/STAGE2/Full_adder_pp2_53_1/_16_  (.A1(\u_multiplier/STAGE2/Full_adder_pp2_53_1/_10_ ),
    .A2(\u_multiplier/STAGE2/Full_adder_pp2_53_1/_11_ ),
    .ZN(\u_multiplier/pp2_54 [1]));
 AOI22_X4 \u_multiplier/STAGE2/Full_adder_pp2_53_1/_17_  (.A1(\u_multiplier/STAGE2/Full_adder_pp2_53_1/_08_ ),
    .A2(\u_multiplier/STAGE2/Full_adder_pp2_53_1/_10_ ),
    .B1(\u_multiplier/pp2_54 [1]),
    .B2(\u_multiplier/STAGE2/Full_adder_pp2_53_1/_09_ ),
    .ZN(\u_multiplier/pp2_53 [0]));
 INV_X1 \u_multiplier/STAGE2/Full_adder_pp2_55_1/_12_  (.A(\u_multiplier/STAGE2/pp2_54_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp2_55_1/_08_ ));
 NAND3_X2 \u_multiplier/STAGE2/Full_adder_pp2_55_1/_13_  (.A1(\u_multiplier/pp1_55 [1]),
    .A2(\u_multiplier/pp1_55 [0]),
    .A3(\u_multiplier/STAGE2/pp2_54_e42_1_cout ),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp2_55_1/_09_ ));
 NOR2_X2 \u_multiplier/STAGE2/Full_adder_pp2_55_1/_14_  (.A1(\u_multiplier/pp1_55 [1]),
    .A2(\u_multiplier/pp1_55 [0]),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp2_55_1/_10_ ));
 AOI21_X1 \u_multiplier/STAGE2/Full_adder_pp2_55_1/_15_  (.A(\u_multiplier/STAGE2/pp2_54_e42_1_cout ),
    .B1(\u_multiplier/pp1_55 [0]),
    .B2(\u_multiplier/pp1_55 [1]),
    .ZN(\u_multiplier/STAGE2/Full_adder_pp2_55_1/_11_ ));
 NOR2_X2 \u_multiplier/STAGE2/Full_adder_pp2_55_1/_16_  (.A1(\u_multiplier/STAGE2/Full_adder_pp2_55_1/_10_ ),
    .A2(\u_multiplier/STAGE2/Full_adder_pp2_55_1/_11_ ),
    .ZN(\u_multiplier/pp2_56 [0]));
 AOI22_X4 \u_multiplier/STAGE2/Full_adder_pp2_55_1/_17_  (.A1(\u_multiplier/STAGE2/Full_adder_pp2_55_1/_08_ ),
    .A2(\u_multiplier/STAGE2/Full_adder_pp2_55_1/_10_ ),
    .B1(\u_multiplier/pp2_56 [0]),
    .B2(\u_multiplier/STAGE2/Full_adder_pp2_55_1/_09_ ),
    .ZN(\u_multiplier/pp2_55 [0]));
 AND2_X1 \u_multiplier/STAGE2/Half_adder_pp2_10_1/_4_  (.A1(\u_multiplier/pp1_10 [5]),
    .A2(\u_multiplier/pp1_10 [4]),
    .ZN(\u_multiplier/pp2_11 [2]));
 XOR2_X2 \u_multiplier/STAGE2/Half_adder_pp2_10_1/_5_  (.A(\u_multiplier/pp1_10 [5]),
    .B(\u_multiplier/pp1_10 [4]),
    .Z(\u_multiplier/pp2_10 [0]));
 AND2_X1 \u_multiplier/STAGE2/Half_adder_pp2_12_1/_4_  (.A1(\u_multiplier/pp1_12 [9]),
    .A2(\u_multiplier/pp1_12 [8]),
    .ZN(\u_multiplier/pp2_13 [3]));
 XOR2_X2 \u_multiplier/STAGE2/Half_adder_pp2_12_1/_5_  (.A(\u_multiplier/pp1_12 [9]),
    .B(\u_multiplier/pp1_12 [8]),
    .Z(\u_multiplier/pp2_12 [0]));
 AND2_X1 \u_multiplier/STAGE2/Half_adder_pp2_14_1/_4_  (.A1(\u_multiplier/pp1_14 [13]),
    .A2(\u_multiplier/pp1_14 [12]),
    .ZN(\u_multiplier/pp2_15 [4]));
 XOR2_X2 \u_multiplier/STAGE2/Half_adder_pp2_14_1/_5_  (.A(\u_multiplier/pp1_14 [13]),
    .B(\u_multiplier/pp1_14 [12]),
    .Z(\u_multiplier/pp2_14 [0]));
 AND2_X1 \u_multiplier/STAGE2/Half_adder_pp2_8_1/_4_  (.A1(\u_multiplier/pp1_8 [1]),
    .A2(\u_multiplier/pp1_8 [0]),
    .ZN(\u_multiplier/pp2_9 [1]));
 XOR2_X2 \u_multiplier/STAGE2/Half_adder_pp2_8_1/_5_  (.A(\u_multiplier/pp1_8 [1]),
    .B(\u_multiplier/pp1_8 [0]),
    .Z(\u_multiplier/pp2_8 [0]));
 LOGIC0_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_55__140  (.Z(net140));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_10_1/_18_  (.A(\u_multiplier/STAGE3/pp3_9_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_10_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_10_1/_19_  (.A1(\u_multiplier/pp2_10 [1]),
    .A2(\u_multiplier/pp2_10 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_10_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_10_1/_20_  (.A(\u_multiplier/pp2_10 [1]),
    .B(\u_multiplier/pp2_10 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_10_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_10_1/_21_  (.A1(\u_multiplier/pp2_10 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_10_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_10_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_10_1/_22_  (.A(\u_multiplier/pp2_10 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_10_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_10_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_10_1/_23_  (.A1(\u_multiplier/pp2_10 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_10_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_10_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_10_1/_24_  (.A(\u_multiplier/pp2_10 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_10_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_10_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_10_1/_25_  (.A(\u_multiplier/STAGE3/pp3_9_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_10_1/_16_ ),
    .ZN(\u_multiplier/pp3_10 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_10_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_10_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_10_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_10_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_10_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_10_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_10_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_10_1/_17_ ),
    .ZN(\u_multiplier/pp3_11 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_10_2/_18_  (.A(\u_multiplier/STAGE3/pp3_9_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_10_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_10_2/_19_  (.A1(\u_multiplier/pp2_10 [5]),
    .A2(\u_multiplier/pp2_10 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_10_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_10_2/_20_  (.A(\u_multiplier/pp2_10 [5]),
    .B(\u_multiplier/pp2_10 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_10_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_10_2/_21_  (.A1(\u_multiplier/pp2_10 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_10_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_10_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_10_2/_22_  (.A(\u_multiplier/pp2_10 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_10_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_10_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_10_2/_23_  (.A1(\u_multiplier/pp2_10 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_10_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_10_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_10_2/_24_  (.A(\u_multiplier/pp2_10 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_10_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_10_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_10_2/_25_  (.A(\u_multiplier/STAGE3/pp3_9_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_10_2/_16_ ),
    .ZN(\u_multiplier/pp3_10 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_10_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_10_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_10_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_10_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_10_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_10_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_10_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_10_2/_17_ ),
    .ZN(\u_multiplier/pp3_11 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_11_1/_18_  (.A(\u_multiplier/STAGE3/pp3_10_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_11_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_11_1/_19_  (.A1(\u_multiplier/pp2_11 [1]),
    .A2(\u_multiplier/pp2_11 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_11_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_11_1/_20_  (.A(\u_multiplier/pp2_11 [1]),
    .B(\u_multiplier/pp2_11 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_11_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_11_1/_21_  (.A1(\u_multiplier/pp2_11 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_11_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_11_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_11_1/_22_  (.A(\u_multiplier/pp2_11 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_11_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_11_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_11_1/_23_  (.A1(\u_multiplier/pp2_11 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_11_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_11_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_11_1/_24_  (.A(\u_multiplier/pp2_11 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_11_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_11_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_11_1/_25_  (.A(\u_multiplier/STAGE3/pp3_10_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_11_1/_16_ ),
    .ZN(\u_multiplier/pp3_11 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_11_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_11_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_11_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_11_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_11_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_11_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_11_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_11_1/_17_ ),
    .ZN(\u_multiplier/pp3_12 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_11_2/_18_  (.A(\u_multiplier/STAGE3/pp3_10_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_11_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_11_2/_19_  (.A1(\u_multiplier/pp2_11 [5]),
    .A2(\u_multiplier/pp2_11 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_11_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_11_2/_20_  (.A(\u_multiplier/pp2_11 [5]),
    .B(\u_multiplier/pp2_11 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_11_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_11_2/_21_  (.A1(\u_multiplier/pp2_11 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_11_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_11_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_11_2/_22_  (.A(\u_multiplier/pp2_11 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_11_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_11_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_11_2/_23_  (.A1(\u_multiplier/pp2_11 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_11_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_11_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_11_2/_24_  (.A(\u_multiplier/pp2_11 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_11_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_11_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_11_2/_25_  (.A(\u_multiplier/STAGE3/pp3_10_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_11_2/_16_ ),
    .ZN(\u_multiplier/pp3_11 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_11_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_11_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_11_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_11_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_11_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_11_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_11_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_11_2/_17_ ),
    .ZN(\u_multiplier/pp3_12 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_12_1/_18_  (.A(\u_multiplier/STAGE3/pp3_11_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_12_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_12_1/_19_  (.A1(\u_multiplier/pp2_12 [1]),
    .A2(\u_multiplier/pp2_12 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_12_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_12_1/_20_  (.A(\u_multiplier/pp2_12 [1]),
    .B(\u_multiplier/pp2_12 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_12_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_12_1/_21_  (.A1(\u_multiplier/pp2_12 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_12_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_12_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_12_1/_22_  (.A(\u_multiplier/pp2_12 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_12_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_12_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_12_1/_23_  (.A1(\u_multiplier/pp2_12 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_12_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_12_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_12_1/_24_  (.A(\u_multiplier/pp2_12 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_12_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_12_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_12_1/_25_  (.A(\u_multiplier/STAGE3/pp3_11_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_12_1/_16_ ),
    .ZN(\u_multiplier/pp3_12 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_12_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_12_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_12_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_12_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_12_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_12_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_12_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_12_1/_17_ ),
    .ZN(\u_multiplier/pp3_13 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_12_2/_18_  (.A(\u_multiplier/STAGE3/pp3_11_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_12_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_12_2/_19_  (.A1(\u_multiplier/pp2_12 [5]),
    .A2(\u_multiplier/pp2_12 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_12_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_12_2/_20_  (.A(\u_multiplier/pp2_12 [5]),
    .B(\u_multiplier/pp2_12 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_12_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_12_2/_21_  (.A1(\u_multiplier/pp2_12 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_12_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_12_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_12_2/_22_  (.A(\u_multiplier/pp2_12 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_12_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_12_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_12_2/_23_  (.A1(\u_multiplier/pp2_12 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_12_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_12_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_12_2/_24_  (.A(\u_multiplier/pp2_12 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_12_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_12_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_12_2/_25_  (.A(\u_multiplier/STAGE3/pp3_11_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_12_2/_16_ ),
    .ZN(\u_multiplier/pp3_12 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_12_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_12_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_12_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_12_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_12_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_12_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_12_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_12_2/_17_ ),
    .ZN(\u_multiplier/pp3_13 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_13_1/_18_  (.A(\u_multiplier/STAGE3/pp3_12_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_13_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_13_1/_19_  (.A1(\u_multiplier/pp2_13 [1]),
    .A2(\u_multiplier/pp2_13 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_13_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_13_1/_20_  (.A(\u_multiplier/pp2_13 [1]),
    .B(\u_multiplier/pp2_13 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_13_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_13_1/_21_  (.A1(\u_multiplier/pp2_13 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_13_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_13_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_13_1/_22_  (.A(\u_multiplier/pp2_13 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_13_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_13_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_13_1/_23_  (.A1(\u_multiplier/pp2_13 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_13_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_13_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_13_1/_24_  (.A(\u_multiplier/pp2_13 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_13_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_13_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_13_1/_25_  (.A(\u_multiplier/STAGE3/pp3_12_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_13_1/_16_ ),
    .ZN(\u_multiplier/pp3_13 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_13_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_13_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_13_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_13_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_13_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_13_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_13_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_13_1/_17_ ),
    .ZN(\u_multiplier/pp3_14 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_13_2/_18_  (.A(\u_multiplier/STAGE3/pp3_12_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_13_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_13_2/_19_  (.A1(\u_multiplier/pp2_13 [5]),
    .A2(\u_multiplier/pp2_13 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_13_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_13_2/_20_  (.A(\u_multiplier/pp2_13 [5]),
    .B(\u_multiplier/pp2_13 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_13_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_13_2/_21_  (.A1(\u_multiplier/pp2_13 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_13_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_13_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_13_2/_22_  (.A(\u_multiplier/pp2_13 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_13_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_13_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_13_2/_23_  (.A1(\u_multiplier/pp2_13 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_13_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_13_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_13_2/_24_  (.A(\u_multiplier/pp2_13 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_13_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_13_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_13_2/_25_  (.A(\u_multiplier/STAGE3/pp3_12_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_13_2/_16_ ),
    .ZN(\u_multiplier/pp3_13 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_13_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_13_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_13_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_13_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_13_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_13_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_13_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_13_2/_17_ ),
    .ZN(\u_multiplier/pp3_14 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_14_1/_18_  (.A(\u_multiplier/STAGE3/pp3_13_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_14_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_14_1/_19_  (.A1(\u_multiplier/pp2_14 [1]),
    .A2(\u_multiplier/pp2_14 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_14_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_14_1/_20_  (.A(\u_multiplier/pp2_14 [1]),
    .B(\u_multiplier/pp2_14 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_14_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_14_1/_21_  (.A1(\u_multiplier/pp2_14 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_14_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_14_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_14_1/_22_  (.A(\u_multiplier/pp2_14 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_14_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_14_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_14_1/_23_  (.A1(\u_multiplier/pp2_14 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_14_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_14_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_14_1/_24_  (.A(\u_multiplier/pp2_14 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_14_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_14_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_14_1/_25_  (.A(\u_multiplier/STAGE3/pp3_13_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_14_1/_16_ ),
    .ZN(\u_multiplier/pp3_14 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_14_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_14_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_14_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_14_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_14_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_14_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_14_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_14_1/_17_ ),
    .ZN(\u_multiplier/pp3_15 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_14_2/_18_  (.A(\u_multiplier/STAGE3/pp3_13_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_14_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_14_2/_19_  (.A1(\u_multiplier/pp2_14 [5]),
    .A2(\u_multiplier/pp2_14 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_14_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_14_2/_20_  (.A(\u_multiplier/pp2_14 [5]),
    .B(\u_multiplier/pp2_14 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_14_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_14_2/_21_  (.A1(\u_multiplier/pp2_14 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_14_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_14_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_14_2/_22_  (.A(\u_multiplier/pp2_14 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_14_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_14_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_14_2/_23_  (.A1(\u_multiplier/pp2_14 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_14_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_14_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_14_2/_24_  (.A(\u_multiplier/pp2_14 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_14_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_14_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_14_2/_25_  (.A(\u_multiplier/STAGE3/pp3_13_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_14_2/_16_ ),
    .ZN(\u_multiplier/pp3_14 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_14_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_14_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_14_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_14_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_14_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_14_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_14_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_14_2/_17_ ),
    .ZN(\u_multiplier/pp3_15 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_15_1/_18_  (.A(\u_multiplier/STAGE3/pp3_14_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_15_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_15_1/_19_  (.A1(\u_multiplier/pp2_15 [1]),
    .A2(\u_multiplier/pp2_15 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_15_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_15_1/_20_  (.A(\u_multiplier/pp2_15 [1]),
    .B(\u_multiplier/pp2_15 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_15_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_15_1/_21_  (.A1(\u_multiplier/pp2_15 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_15_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_15_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_15_1/_22_  (.A(\u_multiplier/pp2_15 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_15_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_15_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_15_1/_23_  (.A1(\u_multiplier/pp2_15 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_15_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_15_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_15_1/_24_  (.A(\u_multiplier/pp2_15 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_15_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_15_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_15_1/_25_  (.A(\u_multiplier/STAGE3/pp3_14_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_15_1/_16_ ),
    .ZN(\u_multiplier/pp3_15 [1]));
 NAND2_X2 \u_multiplier/STAGE3/E_4_2_pp3_15_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_15_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_15_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_15_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_15_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_15_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_15_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_15_1/_17_ ),
    .ZN(\u_multiplier/pp3_16 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_15_2/_18_  (.A(\u_multiplier/STAGE3/pp3_14_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_15_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_15_2/_19_  (.A1(\u_multiplier/pp2_15 [5]),
    .A2(\u_multiplier/pp2_15 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_15_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_15_2/_20_  (.A(\u_multiplier/pp2_15 [5]),
    .B(\u_multiplier/pp2_15 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_15_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_15_2/_21_  (.A1(\u_multiplier/pp2_15 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_15_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_15_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_15_2/_22_  (.A(\u_multiplier/pp2_15 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_15_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_15_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_15_2/_23_  (.A1(\u_multiplier/pp2_15 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_15_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_15_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_15_2/_24_  (.A(\u_multiplier/pp2_15 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_15_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_15_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_15_2/_25_  (.A(\u_multiplier/STAGE3/pp3_14_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_15_2/_16_ ),
    .ZN(\u_multiplier/pp3_15 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_15_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_15_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_15_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_15_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_15_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_15_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_15_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_15_2/_17_ ),
    .ZN(\u_multiplier/pp3_16 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_16_1/_18_  (.A(\u_multiplier/STAGE3/pp3_15_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_16_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_16_1/_19_  (.A1(\u_multiplier/pp2_16 [1]),
    .A2(\u_multiplier/pp2_16 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_16_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_16_1/_20_  (.A(\u_multiplier/pp2_16 [1]),
    .B(\u_multiplier/pp2_16 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_16_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_16_1/_21_  (.A1(\u_multiplier/pp2_16 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_16_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_16_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_16_1/_22_  (.A(\u_multiplier/pp2_16 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_16_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_16_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_16_1/_23_  (.A1(\u_multiplier/pp2_16 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_16_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_16_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_16_1/_24_  (.A(\u_multiplier/pp2_16 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_16_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_16_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_16_1/_25_  (.A(\u_multiplier/STAGE3/pp3_15_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_16_1/_16_ ),
    .ZN(\u_multiplier/pp3_16 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_16_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_16_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_16_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_16_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_16_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_16_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_16_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_16_1/_17_ ),
    .ZN(\u_multiplier/pp3_17 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_16_2/_18_  (.A(\u_multiplier/STAGE3/pp3_15_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_16_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_16_2/_19_  (.A1(\u_multiplier/pp2_16 [5]),
    .A2(\u_multiplier/pp2_16 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_16_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_16_2/_20_  (.A(\u_multiplier/pp2_16 [5]),
    .B(\u_multiplier/pp2_16 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_16_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_16_2/_21_  (.A1(\u_multiplier/pp2_16 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_16_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_16_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_16_2/_22_  (.A(\u_multiplier/pp2_16 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_16_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_16_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_16_2/_23_  (.A1(\u_multiplier/pp2_16 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_16_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_16_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_16_2/_24_  (.A(\u_multiplier/pp2_16 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_16_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_16_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_16_2/_25_  (.A(\u_multiplier/STAGE3/pp3_15_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_16_2/_16_ ),
    .ZN(\u_multiplier/pp3_16 [0]));
 NAND2_X2 \u_multiplier/STAGE3/E_4_2_pp3_16_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_16_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_16_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_16_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_16_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_16_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_16_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_16_2/_17_ ),
    .ZN(\u_multiplier/pp3_17 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_17_1/_18_  (.A(\u_multiplier/STAGE3/pp3_16_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_17_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_17_1/_19_  (.A1(\u_multiplier/pp2_17 [1]),
    .A2(\u_multiplier/pp2_17 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_17_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_17_1/_20_  (.A(\u_multiplier/pp2_17 [1]),
    .B(\u_multiplier/pp2_17 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_17_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_17_1/_21_  (.A1(\u_multiplier/pp2_17 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_17_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_17_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_17_1/_22_  (.A(\u_multiplier/pp2_17 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_17_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_17_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_17_1/_23_  (.A1(\u_multiplier/pp2_17 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_17_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_17_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_17_1/_24_  (.A(\u_multiplier/pp2_17 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_17_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_17_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_17_1/_25_  (.A(\u_multiplier/STAGE3/pp3_16_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_17_1/_16_ ),
    .ZN(\u_multiplier/pp3_17 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_17_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_17_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_17_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_17_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_17_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_17_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_17_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_17_1/_17_ ),
    .ZN(\u_multiplier/pp3_18 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_17_2/_18_  (.A(\u_multiplier/STAGE3/pp3_16_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_17_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_17_2/_19_  (.A1(\u_multiplier/pp2_17 [5]),
    .A2(\u_multiplier/pp2_17 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_17_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_17_2/_20_  (.A(\u_multiplier/pp2_17 [5]),
    .B(\u_multiplier/pp2_17 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_17_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_17_2/_21_  (.A1(\u_multiplier/pp2_17 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_17_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_17_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_17_2/_22_  (.A(\u_multiplier/pp2_17 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_17_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_17_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_17_2/_23_  (.A1(\u_multiplier/pp2_17 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_17_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_17_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_17_2/_24_  (.A(\u_multiplier/pp2_17 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_17_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_17_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_17_2/_25_  (.A(\u_multiplier/STAGE3/pp3_16_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_17_2/_16_ ),
    .ZN(\u_multiplier/pp3_17 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_17_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_17_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_17_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_17_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_17_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_17_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_17_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_17_2/_17_ ),
    .ZN(\u_multiplier/pp3_18 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_18_1/_18_  (.A(\u_multiplier/STAGE3/pp3_17_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_18_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_18_1/_19_  (.A1(\u_multiplier/pp2_18 [1]),
    .A2(\u_multiplier/pp2_18 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_18_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_18_1/_20_  (.A(\u_multiplier/pp2_18 [1]),
    .B(\u_multiplier/pp2_18 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_18_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_18_1/_21_  (.A1(\u_multiplier/pp2_18 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_18_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_18_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_18_1/_22_  (.A(\u_multiplier/pp2_18 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_18_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_18_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_18_1/_23_  (.A1(\u_multiplier/pp2_18 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_18_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_18_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_18_1/_24_  (.A(\u_multiplier/pp2_18 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_18_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_18_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_18_1/_25_  (.A(\u_multiplier/STAGE3/pp3_17_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_18_1/_16_ ),
    .ZN(\u_multiplier/pp3_18 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_18_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_18_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_18_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_18_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_18_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_18_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_18_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_18_1/_17_ ),
    .ZN(\u_multiplier/pp3_19 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_18_2/_18_  (.A(\u_multiplier/STAGE3/pp3_17_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_18_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_18_2/_19_  (.A1(\u_multiplier/pp2_18 [5]),
    .A2(\u_multiplier/pp2_18 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_18_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_18_2/_20_  (.A(\u_multiplier/pp2_18 [5]),
    .B(\u_multiplier/pp2_18 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_18_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_18_2/_21_  (.A1(\u_multiplier/pp2_18 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_18_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_18_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_18_2/_22_  (.A(\u_multiplier/pp2_18 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_18_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_18_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_18_2/_23_  (.A1(\u_multiplier/pp2_18 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_18_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_18_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_18_2/_24_  (.A(\u_multiplier/pp2_18 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_18_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_18_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_18_2/_25_  (.A(\u_multiplier/STAGE3/pp3_17_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_18_2/_16_ ),
    .ZN(\u_multiplier/pp3_18 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_18_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_18_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_18_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_18_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_18_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_18_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_18_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_18_2/_17_ ),
    .ZN(\u_multiplier/pp3_19 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_19_1/_18_  (.A(\u_multiplier/STAGE3/pp3_18_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_19_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_19_1/_19_  (.A1(\u_multiplier/pp2_19 [1]),
    .A2(\u_multiplier/pp2_19 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_19_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_19_1/_20_  (.A(\u_multiplier/pp2_19 [1]),
    .B(\u_multiplier/pp2_19 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_19_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_19_1/_21_  (.A1(\u_multiplier/pp2_19 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_19_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_19_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_19_1/_22_  (.A(\u_multiplier/pp2_19 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_19_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_19_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_19_1/_23_  (.A1(\u_multiplier/pp2_19 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_19_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_19_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_19_1/_24_  (.A(\u_multiplier/pp2_19 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_19_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_19_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_19_1/_25_  (.A(\u_multiplier/STAGE3/pp3_18_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_19_1/_16_ ),
    .ZN(\u_multiplier/pp3_19 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_19_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_19_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_19_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_19_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_19_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_19_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_19_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_19_1/_17_ ),
    .ZN(\u_multiplier/pp3_20 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_19_2/_18_  (.A(\u_multiplier/STAGE3/pp3_18_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_19_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_19_2/_19_  (.A1(\u_multiplier/pp2_19 [5]),
    .A2(\u_multiplier/pp2_19 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_19_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_19_2/_20_  (.A(\u_multiplier/pp2_19 [5]),
    .B(\u_multiplier/pp2_19 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_19_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_19_2/_21_  (.A1(\u_multiplier/pp2_19 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_19_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_19_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_19_2/_22_  (.A(\u_multiplier/pp2_19 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_19_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_19_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_19_2/_23_  (.A1(\u_multiplier/pp2_19 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_19_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_19_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_19_2/_24_  (.A(\u_multiplier/pp2_19 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_19_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_19_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_19_2/_25_  (.A(\u_multiplier/STAGE3/pp3_18_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_19_2/_16_ ),
    .ZN(\u_multiplier/pp3_19 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_19_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_19_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_19_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_19_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_19_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_19_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_19_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_19_2/_17_ ),
    .ZN(\u_multiplier/pp3_20 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_20_1/_18_  (.A(\u_multiplier/STAGE3/pp3_19_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_20_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_20_1/_19_  (.A1(\u_multiplier/pp2_20 [1]),
    .A2(\u_multiplier/pp2_20 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_20_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_20_1/_20_  (.A(\u_multiplier/pp2_20 [1]),
    .B(\u_multiplier/pp2_20 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_20_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_20_1/_21_  (.A1(\u_multiplier/pp2_20 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_20_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_20_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_20_1/_22_  (.A(\u_multiplier/pp2_20 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_20_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_20_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_20_1/_23_  (.A1(\u_multiplier/pp2_20 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_20_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_20_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_20_1/_24_  (.A(\u_multiplier/pp2_20 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_20_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_20_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_20_1/_25_  (.A(\u_multiplier/STAGE3/pp3_19_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_20_1/_16_ ),
    .ZN(\u_multiplier/pp3_20 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_20_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_20_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_20_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_20_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_20_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_20_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_20_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_20_1/_17_ ),
    .ZN(\u_multiplier/pp3_21 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_20_2/_18_  (.A(\u_multiplier/STAGE3/pp3_19_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_20_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_20_2/_19_  (.A1(\u_multiplier/pp2_20 [5]),
    .A2(\u_multiplier/pp2_20 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_20_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_20_2/_20_  (.A(\u_multiplier/pp2_20 [5]),
    .B(\u_multiplier/pp2_20 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_20_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_20_2/_21_  (.A1(\u_multiplier/pp2_20 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_20_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_20_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_20_2/_22_  (.A(\u_multiplier/pp2_20 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_20_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_20_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_20_2/_23_  (.A1(\u_multiplier/pp2_20 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_20_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_20_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_20_2/_24_  (.A(\u_multiplier/pp2_20 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_20_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_20_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_20_2/_25_  (.A(\u_multiplier/STAGE3/pp3_19_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_20_2/_16_ ),
    .ZN(\u_multiplier/pp3_20 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_20_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_20_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_20_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_20_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_20_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_20_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_20_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_20_2/_17_ ),
    .ZN(\u_multiplier/pp3_21 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_21_1/_18_  (.A(\u_multiplier/STAGE3/pp3_20_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_21_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_21_1/_19_  (.A1(\u_multiplier/pp2_21 [1]),
    .A2(\u_multiplier/pp2_21 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_21_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_21_1/_20_  (.A(\u_multiplier/pp2_21 [1]),
    .B(\u_multiplier/pp2_21 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_21_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_21_1/_21_  (.A1(\u_multiplier/pp2_21 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_21_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_21_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_21_1/_22_  (.A(\u_multiplier/pp2_21 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_21_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_21_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_21_1/_23_  (.A1(\u_multiplier/pp2_21 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_21_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_21_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_21_1/_24_  (.A(\u_multiplier/pp2_21 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_21_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_21_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_21_1/_25_  (.A(\u_multiplier/STAGE3/pp3_20_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_21_1/_16_ ),
    .ZN(\u_multiplier/pp3_21 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_21_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_21_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_21_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_21_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_21_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_21_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_21_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_21_1/_17_ ),
    .ZN(\u_multiplier/pp3_22 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_21_2/_18_  (.A(\u_multiplier/STAGE3/pp3_20_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_21_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_21_2/_19_  (.A1(\u_multiplier/pp2_21 [5]),
    .A2(\u_multiplier/pp2_21 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_21_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_21_2/_20_  (.A(\u_multiplier/pp2_21 [5]),
    .B(\u_multiplier/pp2_21 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_21_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_21_2/_21_  (.A1(\u_multiplier/pp2_21 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_21_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_21_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_21_2/_22_  (.A(\u_multiplier/pp2_21 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_21_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_21_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_21_2/_23_  (.A1(\u_multiplier/pp2_21 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_21_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_21_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_21_2/_24_  (.A(\u_multiplier/pp2_21 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_21_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_21_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_21_2/_25_  (.A(\u_multiplier/STAGE3/pp3_20_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_21_2/_16_ ),
    .ZN(\u_multiplier/pp3_21 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_21_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_21_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_21_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_21_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_21_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_21_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_21_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_21_2/_17_ ),
    .ZN(\u_multiplier/pp3_22 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_22_1/_18_  (.A(\u_multiplier/STAGE3/pp3_21_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_22_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_22_1/_19_  (.A1(\u_multiplier/pp2_22 [1]),
    .A2(\u_multiplier/pp2_22 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_22_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_22_1/_20_  (.A(\u_multiplier/pp2_22 [1]),
    .B(\u_multiplier/pp2_22 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_22_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_22_1/_21_  (.A1(\u_multiplier/pp2_22 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_22_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_22_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_22_1/_22_  (.A(\u_multiplier/pp2_22 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_22_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_22_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_22_1/_23_  (.A1(\u_multiplier/pp2_22 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_22_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_22_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_22_1/_24_  (.A(\u_multiplier/pp2_22 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_22_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_22_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_22_1/_25_  (.A(\u_multiplier/STAGE3/pp3_21_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_22_1/_16_ ),
    .ZN(\u_multiplier/pp3_22 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_22_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_22_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_22_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_22_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_22_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_22_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_22_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_22_1/_17_ ),
    .ZN(\u_multiplier/pp3_23 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_22_2/_18_  (.A(\u_multiplier/STAGE3/pp3_21_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_22_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_22_2/_19_  (.A1(\u_multiplier/pp2_22 [5]),
    .A2(\u_multiplier/pp2_22 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_22_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_22_2/_20_  (.A(\u_multiplier/pp2_22 [5]),
    .B(\u_multiplier/pp2_22 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_22_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_22_2/_21_  (.A1(\u_multiplier/pp2_22 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_22_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_22_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_22_2/_22_  (.A(\u_multiplier/pp2_22 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_22_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_22_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_22_2/_23_  (.A1(\u_multiplier/pp2_22 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_22_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_22_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_22_2/_24_  (.A(\u_multiplier/pp2_22 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_22_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_22_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_22_2/_25_  (.A(\u_multiplier/STAGE3/pp3_21_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_22_2/_16_ ),
    .ZN(\u_multiplier/pp3_22 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_22_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_22_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_22_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_22_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_22_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_22_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_22_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_22_2/_17_ ),
    .ZN(\u_multiplier/pp3_23 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_23_1/_18_  (.A(\u_multiplier/STAGE3/pp3_22_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_23_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_23_1/_19_  (.A1(\u_multiplier/pp2_23 [1]),
    .A2(\u_multiplier/pp2_23 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_23_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_23_1/_20_  (.A(\u_multiplier/pp2_23 [1]),
    .B(\u_multiplier/pp2_23 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_23_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_23_1/_21_  (.A1(\u_multiplier/pp2_23 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_23_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_23_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_23_1/_22_  (.A(\u_multiplier/pp2_23 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_23_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_23_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_23_1/_23_  (.A1(\u_multiplier/pp2_23 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_23_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_23_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_23_1/_24_  (.A(\u_multiplier/pp2_23 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_23_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_23_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_23_1/_25_  (.A(\u_multiplier/STAGE3/pp3_22_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_23_1/_16_ ),
    .ZN(\u_multiplier/pp3_23 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_23_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_23_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_23_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_23_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_23_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_23_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_23_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_23_1/_17_ ),
    .ZN(\u_multiplier/pp3_24 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_23_2/_18_  (.A(\u_multiplier/STAGE3/pp3_22_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_23_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_23_2/_19_  (.A1(\u_multiplier/pp2_23 [5]),
    .A2(\u_multiplier/pp2_23 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_23_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_23_2/_20_  (.A(\u_multiplier/pp2_23 [5]),
    .B(\u_multiplier/pp2_23 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_23_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_23_2/_21_  (.A1(\u_multiplier/pp2_23 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_23_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_23_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_23_2/_22_  (.A(\u_multiplier/pp2_23 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_23_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_23_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_23_2/_23_  (.A1(\u_multiplier/pp2_23 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_23_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_23_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_23_2/_24_  (.A(\u_multiplier/pp2_23 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_23_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_23_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_23_2/_25_  (.A(\u_multiplier/STAGE3/pp3_22_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_23_2/_16_ ),
    .ZN(\u_multiplier/pp3_23 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_23_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_23_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_23_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_23_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_23_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_23_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_23_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_23_2/_17_ ),
    .ZN(\u_multiplier/pp3_24 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_24_1/_18_  (.A(\u_multiplier/STAGE3/pp3_23_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_24_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_24_1/_19_  (.A1(\u_multiplier/pp2_24 [1]),
    .A2(\u_multiplier/pp2_24 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_24_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_24_1/_20_  (.A(\u_multiplier/pp2_24 [1]),
    .B(\u_multiplier/pp2_24 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_24_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_24_1/_21_  (.A1(\u_multiplier/pp2_24 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_24_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_24_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_24_1/_22_  (.A(\u_multiplier/pp2_24 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_24_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_24_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_24_1/_23_  (.A1(\u_multiplier/pp2_24 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_24_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_24_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_24_1/_24_  (.A(\u_multiplier/pp2_24 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_24_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_24_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_24_1/_25_  (.A(\u_multiplier/STAGE3/pp3_23_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_24_1/_16_ ),
    .ZN(\u_multiplier/pp3_24 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_24_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_24_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_24_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_24_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_24_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_24_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_24_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_24_1/_17_ ),
    .ZN(\u_multiplier/pp3_25 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_24_2/_18_  (.A(\u_multiplier/STAGE3/pp3_23_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_24_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_24_2/_19_  (.A1(\u_multiplier/pp2_24 [5]),
    .A2(\u_multiplier/pp2_24 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_24_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_24_2/_20_  (.A(\u_multiplier/pp2_24 [5]),
    .B(\u_multiplier/pp2_24 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_24_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_24_2/_21_  (.A1(\u_multiplier/pp2_24 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_24_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_24_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_24_2/_22_  (.A(\u_multiplier/pp2_24 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_24_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_24_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_24_2/_23_  (.A1(\u_multiplier/pp2_24 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_24_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_24_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_24_2/_24_  (.A(\u_multiplier/pp2_24 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_24_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_24_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_24_2/_25_  (.A(\u_multiplier/STAGE3/pp3_23_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_24_2/_16_ ),
    .ZN(\u_multiplier/pp3_24 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_24_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_24_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_24_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_24_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_24_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_24_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_24_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_24_2/_17_ ),
    .ZN(\u_multiplier/pp3_25 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_25_1/_18_  (.A(\u_multiplier/STAGE3/pp3_24_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_25_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_25_1/_19_  (.A1(\u_multiplier/pp2_25 [1]),
    .A2(\u_multiplier/pp2_25 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_25_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_25_1/_20_  (.A(\u_multiplier/pp2_25 [1]),
    .B(\u_multiplier/pp2_25 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_25_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_25_1/_21_  (.A1(\u_multiplier/pp2_25 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_25_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_25_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_25_1/_22_  (.A(\u_multiplier/pp2_25 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_25_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_25_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_25_1/_23_  (.A1(\u_multiplier/pp2_25 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_25_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_25_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_25_1/_24_  (.A(\u_multiplier/pp2_25 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_25_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_25_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_25_1/_25_  (.A(\u_multiplier/STAGE3/pp3_24_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_25_1/_16_ ),
    .ZN(\u_multiplier/pp3_25 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_25_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_25_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_25_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_25_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_25_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_25_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_25_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_25_1/_17_ ),
    .ZN(\u_multiplier/pp3_26 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_25_2/_18_  (.A(\u_multiplier/STAGE3/pp3_24_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_25_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_25_2/_19_  (.A1(\u_multiplier/pp2_25 [5]),
    .A2(\u_multiplier/pp2_25 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_25_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_25_2/_20_  (.A(\u_multiplier/pp2_25 [5]),
    .B(\u_multiplier/pp2_25 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_25_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_25_2/_21_  (.A1(\u_multiplier/pp2_25 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_25_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_25_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_25_2/_22_  (.A(\u_multiplier/pp2_25 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_25_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_25_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_25_2/_23_  (.A1(\u_multiplier/pp2_25 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_25_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_25_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_25_2/_24_  (.A(\u_multiplier/pp2_25 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_25_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_25_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_25_2/_25_  (.A(\u_multiplier/STAGE3/pp3_24_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_25_2/_16_ ),
    .ZN(\u_multiplier/pp3_25 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_25_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_25_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_25_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_25_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_25_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_25_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_25_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_25_2/_17_ ),
    .ZN(\u_multiplier/pp3_26 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_26_1/_18_  (.A(\u_multiplier/STAGE3/pp3_25_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_26_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_26_1/_19_  (.A1(\u_multiplier/pp2_26 [1]),
    .A2(\u_multiplier/pp2_26 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_26_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_26_1/_20_  (.A(\u_multiplier/pp2_26 [1]),
    .B(\u_multiplier/pp2_26 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_26_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_26_1/_21_  (.A1(\u_multiplier/pp2_26 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_26_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_26_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_26_1/_22_  (.A(\u_multiplier/pp2_26 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_26_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_26_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_26_1/_23_  (.A1(\u_multiplier/pp2_26 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_26_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_26_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_26_1/_24_  (.A(\u_multiplier/pp2_26 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_26_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_26_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_26_1/_25_  (.A(\u_multiplier/STAGE3/pp3_25_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_26_1/_16_ ),
    .ZN(\u_multiplier/pp3_26 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_26_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_26_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_26_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_26_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_26_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_26_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_26_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_26_1/_17_ ),
    .ZN(\u_multiplier/pp3_27 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_26_2/_18_  (.A(\u_multiplier/STAGE3/pp3_25_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_26_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_26_2/_19_  (.A1(\u_multiplier/pp2_26 [5]),
    .A2(\u_multiplier/pp2_26 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_26_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_26_2/_20_  (.A(\u_multiplier/pp2_26 [5]),
    .B(\u_multiplier/pp2_26 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_26_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_26_2/_21_  (.A1(\u_multiplier/pp2_26 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_26_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_26_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_26_2/_22_  (.A(\u_multiplier/pp2_26 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_26_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_26_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_26_2/_23_  (.A1(\u_multiplier/pp2_26 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_26_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_26_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_26_2/_24_  (.A(\u_multiplier/pp2_26 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_26_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_26_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_26_2/_25_  (.A(\u_multiplier/STAGE3/pp3_25_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_26_2/_16_ ),
    .ZN(\u_multiplier/pp3_26 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_26_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_26_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_26_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_26_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_26_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_26_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_26_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_26_2/_17_ ),
    .ZN(\u_multiplier/pp3_27 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_27_1/_18_  (.A(\u_multiplier/STAGE3/pp3_26_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_27_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_27_1/_19_  (.A1(\u_multiplier/pp2_27 [1]),
    .A2(\u_multiplier/pp2_27 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_27_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_27_1/_20_  (.A(\u_multiplier/pp2_27 [1]),
    .B(\u_multiplier/pp2_27 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_27_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_27_1/_21_  (.A1(\u_multiplier/pp2_27 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_27_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_27_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_27_1/_22_  (.A(\u_multiplier/pp2_27 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_27_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_27_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_27_1/_23_  (.A1(\u_multiplier/pp2_27 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_27_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_27_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_27_1/_24_  (.A(\u_multiplier/pp2_27 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_27_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_27_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_27_1/_25_  (.A(\u_multiplier/STAGE3/pp3_26_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_27_1/_16_ ),
    .ZN(\u_multiplier/pp3_27 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_27_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_27_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_27_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_27_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_27_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_27_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_27_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_27_1/_17_ ),
    .ZN(\u_multiplier/pp3_28 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_27_2/_18_  (.A(\u_multiplier/STAGE3/pp3_26_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_27_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_27_2/_19_  (.A1(\u_multiplier/pp2_27 [5]),
    .A2(\u_multiplier/pp2_27 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_27_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_27_2/_20_  (.A(\u_multiplier/pp2_27 [5]),
    .B(\u_multiplier/pp2_27 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_27_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_27_2/_21_  (.A1(\u_multiplier/pp2_27 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_27_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_27_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_27_2/_22_  (.A(\u_multiplier/pp2_27 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_27_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_27_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_27_2/_23_  (.A1(\u_multiplier/pp2_27 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_27_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_27_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_27_2/_24_  (.A(\u_multiplier/pp2_27 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_27_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_27_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_27_2/_25_  (.A(\u_multiplier/STAGE3/pp3_26_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_27_2/_16_ ),
    .ZN(\u_multiplier/pp3_27 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_27_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_27_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_27_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_27_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_27_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_27_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_27_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_27_2/_17_ ),
    .ZN(\u_multiplier/pp3_28 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_28_1/_18_  (.A(\u_multiplier/STAGE3/pp3_27_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_28_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_28_1/_19_  (.A1(\u_multiplier/pp2_28 [1]),
    .A2(\u_multiplier/pp2_28 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_28_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_28_1/_20_  (.A(\u_multiplier/pp2_28 [1]),
    .B(\u_multiplier/pp2_28 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_28_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_28_1/_21_  (.A1(\u_multiplier/pp2_28 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_28_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_28_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_28_1/_22_  (.A(\u_multiplier/pp2_28 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_28_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_28_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_28_1/_23_  (.A1(\u_multiplier/pp2_28 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_28_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_28_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_28_1/_24_  (.A(\u_multiplier/pp2_28 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_28_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_28_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_28_1/_25_  (.A(\u_multiplier/STAGE3/pp3_27_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_28_1/_16_ ),
    .ZN(\u_multiplier/pp3_28 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_28_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_28_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_28_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_28_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_28_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_28_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_28_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_28_1/_17_ ),
    .ZN(\u_multiplier/pp3_29 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_28_2/_18_  (.A(\u_multiplier/STAGE3/pp3_27_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_28_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_28_2/_19_  (.A1(\u_multiplier/pp2_28 [5]),
    .A2(\u_multiplier/pp2_28 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_28_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_28_2/_20_  (.A(\u_multiplier/pp2_28 [5]),
    .B(\u_multiplier/pp2_28 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_28_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_28_2/_21_  (.A1(\u_multiplier/pp2_28 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_28_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_28_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_28_2/_22_  (.A(\u_multiplier/pp2_28 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_28_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_28_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_28_2/_23_  (.A1(\u_multiplier/pp2_28 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_28_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_28_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_28_2/_24_  (.A(\u_multiplier/pp2_28 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_28_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_28_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_28_2/_25_  (.A(\u_multiplier/STAGE3/pp3_27_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_28_2/_16_ ),
    .ZN(\u_multiplier/pp3_28 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_28_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_28_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_28_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_28_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_28_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_28_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_28_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_28_2/_17_ ),
    .ZN(\u_multiplier/pp3_29 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_29_1/_18_  (.A(\u_multiplier/STAGE3/pp3_28_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_29_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_29_1/_19_  (.A1(\u_multiplier/pp2_29 [1]),
    .A2(\u_multiplier/pp2_29 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_29_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_29_1/_20_  (.A(\u_multiplier/pp2_29 [1]),
    .B(\u_multiplier/pp2_29 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_29_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_29_1/_21_  (.A1(\u_multiplier/pp2_29 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_29_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_29_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_29_1/_22_  (.A(\u_multiplier/pp2_29 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_29_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_29_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_29_1/_23_  (.A1(\u_multiplier/pp2_29 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_29_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_29_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_29_1/_24_  (.A(\u_multiplier/pp2_29 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_29_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_29_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_29_1/_25_  (.A(\u_multiplier/STAGE3/pp3_28_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_29_1/_16_ ),
    .ZN(\u_multiplier/pp3_29 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_29_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_29_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_29_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_29_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_29_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_29_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_29_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_29_1/_17_ ),
    .ZN(\u_multiplier/pp3_30 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_29_2/_18_  (.A(\u_multiplier/STAGE3/pp3_28_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_29_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_29_2/_19_  (.A1(\u_multiplier/pp2_29 [5]),
    .A2(\u_multiplier/pp2_29 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_29_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_29_2/_20_  (.A(\u_multiplier/pp2_29 [5]),
    .B(\u_multiplier/pp2_29 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_29_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_29_2/_21_  (.A1(\u_multiplier/pp2_29 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_29_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_29_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_29_2/_22_  (.A(\u_multiplier/pp2_29 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_29_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_29_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_29_2/_23_  (.A1(\u_multiplier/pp2_29 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_29_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_29_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_29_2/_24_  (.A(\u_multiplier/pp2_29 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_29_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_29_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_29_2/_25_  (.A(\u_multiplier/STAGE3/pp3_28_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_29_2/_16_ ),
    .ZN(\u_multiplier/pp3_29 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_29_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_29_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_29_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_29_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_29_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_29_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_29_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_29_2/_17_ ),
    .ZN(\u_multiplier/pp3_30 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_30_1/_18_  (.A(\u_multiplier/STAGE3/pp3_29_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_30_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_30_1/_19_  (.A1(\u_multiplier/pp2_30 [1]),
    .A2(\u_multiplier/pp2_30 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_30_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_30_1/_20_  (.A(\u_multiplier/pp2_30 [1]),
    .B(\u_multiplier/pp2_30 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_30_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_30_1/_21_  (.A1(\u_multiplier/pp2_30 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_30_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_30_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_30_1/_22_  (.A(\u_multiplier/pp2_30 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_30_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_30_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_30_1/_23_  (.A1(\u_multiplier/pp2_30 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_30_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_30_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_30_1/_24_  (.A(\u_multiplier/pp2_30 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_30_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_30_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_30_1/_25_  (.A(\u_multiplier/STAGE3/pp3_29_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_30_1/_16_ ),
    .ZN(\u_multiplier/pp3_30 [1]));
 NAND2_X2 \u_multiplier/STAGE3/E_4_2_pp3_30_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_30_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_30_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_30_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_30_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_30_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_30_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_30_1/_17_ ),
    .ZN(\u_multiplier/pp3_31 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_30_2/_18_  (.A(\u_multiplier/STAGE3/pp3_29_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_30_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_30_2/_19_  (.A1(\u_multiplier/pp2_30 [5]),
    .A2(\u_multiplier/pp2_30 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_30_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_30_2/_20_  (.A(\u_multiplier/pp2_30 [5]),
    .B(\u_multiplier/pp2_30 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_30_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_30_2/_21_  (.A1(\u_multiplier/pp2_30 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_30_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_30_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_30_2/_22_  (.A(\u_multiplier/pp2_30 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_30_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_30_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_30_2/_23_  (.A1(\u_multiplier/pp2_30 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_30_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_30_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_30_2/_24_  (.A(\u_multiplier/pp2_30 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_30_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_30_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_30_2/_25_  (.A(\u_multiplier/STAGE3/pp3_29_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_30_2/_16_ ),
    .ZN(\u_multiplier/pp3_30 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_30_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_30_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_30_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_30_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_30_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_30_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_30_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_30_2/_17_ ),
    .ZN(\u_multiplier/pp3_31 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_31_1/_18_  (.A(\u_multiplier/STAGE3/pp3_30_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_31_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_31_1/_19_  (.A1(\u_multiplier/pp2_31 [1]),
    .A2(\u_multiplier/pp2_31 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_31_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_31_1/_20_  (.A(\u_multiplier/pp2_31 [1]),
    .B(\u_multiplier/pp2_31 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_31_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_31_1/_21_  (.A1(\u_multiplier/pp2_31 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_31_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_31_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_31_1/_22_  (.A(\u_multiplier/pp2_31 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_31_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_31_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_31_1/_23_  (.A1(\u_multiplier/pp2_31 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_31_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_31_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_31_1/_24_  (.A(\u_multiplier/pp2_31 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_31_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_31_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_31_1/_25_  (.A(\u_multiplier/STAGE3/pp3_30_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_31_1/_16_ ),
    .ZN(\u_multiplier/pp3_31 [1]));
 NAND2_X2 \u_multiplier/STAGE3/E_4_2_pp3_31_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_31_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_31_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_31_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_31_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_31_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_31_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_31_1/_17_ ),
    .ZN(\u_multiplier/pp3_32 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_31_2/_18_  (.A(\u_multiplier/STAGE3/pp3_30_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_31_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_31_2/_19_  (.A1(\u_multiplier/pp2_31 [5]),
    .A2(\u_multiplier/pp2_31 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_31_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_31_2/_20_  (.A(\u_multiplier/pp2_31 [5]),
    .B(\u_multiplier/pp2_31 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_31_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_31_2/_21_  (.A1(\u_multiplier/pp2_31 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_31_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_31_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_31_2/_22_  (.A(\u_multiplier/pp2_31 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_31_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_31_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_31_2/_23_  (.A1(\u_multiplier/pp2_31 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_31_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_31_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_31_2/_24_  (.A(\u_multiplier/pp2_31 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_31_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_31_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_31_2/_25_  (.A(\u_multiplier/STAGE3/pp3_30_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_31_2/_16_ ),
    .ZN(\u_multiplier/pp3_31 [0]));
 NAND2_X2 \u_multiplier/STAGE3/E_4_2_pp3_31_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_31_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_31_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_31_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_31_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_31_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_31_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_31_2/_17_ ),
    .ZN(\u_multiplier/pp3_32 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_32_1/_18_  (.A(\u_multiplier/STAGE3/pp3_31_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_32_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_32_1/_19_  (.A1(\u_multiplier/pp2_32 [1]),
    .A2(\u_multiplier/pp2_32 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_32_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_32_1/_20_  (.A(\u_multiplier/pp2_32 [1]),
    .B(\u_multiplier/pp2_32 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_32_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_32_1/_21_  (.A1(\u_multiplier/pp2_32 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_32_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_32_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_32_1/_22_  (.A(\u_multiplier/pp2_32 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_32_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_32_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_32_1/_23_  (.A1(\u_multiplier/pp2_32 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_32_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_32_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_32_1/_24_  (.A(\u_multiplier/pp2_32 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_32_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_32_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_32_1/_25_  (.A(\u_multiplier/STAGE3/pp3_31_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_32_1/_16_ ),
    .ZN(\u_multiplier/pp3_32 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_32_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_32_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_32_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_32_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_32_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_32_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_32_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_32_1/_17_ ),
    .ZN(\u_multiplier/pp3_33 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_32_2/_18_  (.A(\u_multiplier/STAGE3/pp3_31_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_32_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_32_2/_19_  (.A1(\u_multiplier/pp2_32 [5]),
    .A2(\u_multiplier/pp2_32 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_32_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_32_2/_20_  (.A(\u_multiplier/pp2_32 [5]),
    .B(\u_multiplier/pp2_32 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_32_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_32_2/_21_  (.A1(\u_multiplier/pp2_32 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_32_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_32_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_32_2/_22_  (.A(\u_multiplier/pp2_32 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_32_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_32_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_32_2/_23_  (.A1(\u_multiplier/pp2_32 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_32_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_32_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_32_2/_24_  (.A(\u_multiplier/pp2_32 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_32_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_32_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_32_2/_25_  (.A(\u_multiplier/STAGE3/pp3_31_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_32_2/_16_ ),
    .ZN(\u_multiplier/pp3_32 [0]));
 NAND2_X2 \u_multiplier/STAGE3/E_4_2_pp3_32_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_32_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_32_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_32_e42_2_cout ));
 OAI21_X4 \u_multiplier/STAGE3/E_4_2_pp3_32_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_32_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_32_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_32_2/_17_ ),
    .ZN(\u_multiplier/pp3_33 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_33_1/_18_  (.A(\u_multiplier/STAGE3/pp3_32_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_33_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_33_1/_19_  (.A1(\u_multiplier/pp2_33 [1]),
    .A2(\u_multiplier/pp2_33 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_33_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_33_1/_20_  (.A(\u_multiplier/pp2_33 [1]),
    .B(\u_multiplier/pp2_33 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_33_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_33_1/_21_  (.A1(\u_multiplier/pp2_33 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_33_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_33_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_33_1/_22_  (.A(\u_multiplier/pp2_33 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_33_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_33_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_33_1/_23_  (.A1(\u_multiplier/pp2_33 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_33_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_33_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_33_1/_24_  (.A(\u_multiplier/pp2_33 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_33_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_33_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_33_1/_25_  (.A(\u_multiplier/STAGE3/pp3_32_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_33_1/_16_ ),
    .ZN(\u_multiplier/pp3_33 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_33_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_33_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_33_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_33_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_33_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_33_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_33_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_33_1/_17_ ),
    .ZN(\u_multiplier/pp3_34 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_33_2/_18_  (.A(\u_multiplier/STAGE3/pp3_32_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_33_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_33_2/_19_  (.A1(\u_multiplier/pp2_33 [5]),
    .A2(\u_multiplier/pp2_33 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_33_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_33_2/_20_  (.A(\u_multiplier/pp2_33 [5]),
    .B(\u_multiplier/pp2_33 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_33_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_33_2/_21_  (.A1(\u_multiplier/pp2_33 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_33_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_33_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_33_2/_22_  (.A(\u_multiplier/pp2_33 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_33_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_33_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_33_2/_23_  (.A1(\u_multiplier/pp2_33 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_33_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_33_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_33_2/_24_  (.A(\u_multiplier/pp2_33 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_33_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_33_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_33_2/_25_  (.A(\u_multiplier/STAGE3/pp3_32_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_33_2/_16_ ),
    .ZN(\u_multiplier/pp3_33 [0]));
 NAND2_X2 \u_multiplier/STAGE3/E_4_2_pp3_33_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_33_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_33_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_33_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_33_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_33_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_33_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_33_2/_17_ ),
    .ZN(\u_multiplier/pp3_34 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_34_1/_18_  (.A(\u_multiplier/STAGE3/pp3_33_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_34_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_34_1/_19_  (.A1(\u_multiplier/pp2_34 [1]),
    .A2(\u_multiplier/pp2_34 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_34_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_34_1/_20_  (.A(\u_multiplier/pp2_34 [1]),
    .B(\u_multiplier/pp2_34 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_34_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_34_1/_21_  (.A1(\u_multiplier/pp2_34 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_34_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_34_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_34_1/_22_  (.A(\u_multiplier/pp2_34 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_34_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_34_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_34_1/_23_  (.A1(\u_multiplier/pp2_34 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_34_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_34_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_34_1/_24_  (.A(\u_multiplier/pp2_34 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_34_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_34_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_34_1/_25_  (.A(\u_multiplier/STAGE3/pp3_33_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_34_1/_16_ ),
    .ZN(\u_multiplier/pp3_34 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_34_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_34_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_34_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_34_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_34_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_34_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_34_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_34_1/_17_ ),
    .ZN(\u_multiplier/pp3_35 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_34_2/_18_  (.A(\u_multiplier/STAGE3/pp3_33_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_34_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_34_2/_19_  (.A1(\u_multiplier/pp2_34 [5]),
    .A2(\u_multiplier/pp2_34 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_34_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_34_2/_20_  (.A(\u_multiplier/pp2_34 [5]),
    .B(\u_multiplier/pp2_34 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_34_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_34_2/_21_  (.A1(\u_multiplier/pp2_34 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_34_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_34_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_34_2/_22_  (.A(\u_multiplier/pp2_34 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_34_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_34_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_34_2/_23_  (.A1(\u_multiplier/pp2_34 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_34_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_34_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_34_2/_24_  (.A(\u_multiplier/pp2_34 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_34_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_34_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_34_2/_25_  (.A(\u_multiplier/STAGE3/pp3_33_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_34_2/_16_ ),
    .ZN(\u_multiplier/pp3_34 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_34_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_34_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_34_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_34_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_34_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_34_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_34_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_34_2/_17_ ),
    .ZN(\u_multiplier/pp3_35 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_35_1/_18_  (.A(\u_multiplier/STAGE3/pp3_34_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_35_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_35_1/_19_  (.A1(\u_multiplier/pp2_35 [1]),
    .A2(\u_multiplier/pp2_35 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_35_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_35_1/_20_  (.A(\u_multiplier/pp2_35 [1]),
    .B(\u_multiplier/pp2_35 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_35_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_35_1/_21_  (.A1(\u_multiplier/pp2_35 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_35_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_35_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_35_1/_22_  (.A(\u_multiplier/pp2_35 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_35_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_35_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_35_1/_23_  (.A1(\u_multiplier/pp2_35 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_35_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_35_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_35_1/_24_  (.A(\u_multiplier/pp2_35 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_35_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_35_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_35_1/_25_  (.A(\u_multiplier/STAGE3/pp3_34_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_35_1/_16_ ),
    .ZN(\u_multiplier/pp3_35 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_35_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_35_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_35_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_35_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_35_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_35_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_35_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_35_1/_17_ ),
    .ZN(\u_multiplier/pp3_36 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_35_2/_18_  (.A(\u_multiplier/STAGE3/pp3_34_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_35_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_35_2/_19_  (.A1(\u_multiplier/pp2_35 [5]),
    .A2(\u_multiplier/pp2_35 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_35_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_35_2/_20_  (.A(\u_multiplier/pp2_35 [5]),
    .B(\u_multiplier/pp2_35 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_35_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_35_2/_21_  (.A1(\u_multiplier/pp2_35 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_35_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_35_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_35_2/_22_  (.A(\u_multiplier/pp2_35 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_35_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_35_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_35_2/_23_  (.A1(\u_multiplier/pp2_35 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_35_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_35_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_35_2/_24_  (.A(\u_multiplier/pp2_35 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_35_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_35_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_35_2/_25_  (.A(\u_multiplier/STAGE3/pp3_34_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_35_2/_16_ ),
    .ZN(\u_multiplier/pp3_35 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_35_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_35_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_35_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_35_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_35_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_35_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_35_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_35_2/_17_ ),
    .ZN(\u_multiplier/pp3_36 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_36_1/_18_  (.A(\u_multiplier/STAGE3/pp3_35_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_36_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_36_1/_19_  (.A1(\u_multiplier/pp2_36 [1]),
    .A2(\u_multiplier/pp2_36 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_36_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_36_1/_20_  (.A(\u_multiplier/pp2_36 [1]),
    .B(\u_multiplier/pp2_36 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_36_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_36_1/_21_  (.A1(\u_multiplier/pp2_36 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_36_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_36_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_36_1/_22_  (.A(\u_multiplier/pp2_36 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_36_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_36_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_36_1/_23_  (.A1(\u_multiplier/pp2_36 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_36_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_36_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_36_1/_24_  (.A(\u_multiplier/pp2_36 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_36_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_36_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_36_1/_25_  (.A(\u_multiplier/STAGE3/pp3_35_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_36_1/_16_ ),
    .ZN(\u_multiplier/pp3_36 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_36_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_36_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_36_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_36_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_36_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_36_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_36_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_36_1/_17_ ),
    .ZN(\u_multiplier/pp3_37 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_36_2/_18_  (.A(\u_multiplier/STAGE3/pp3_35_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_36_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_36_2/_19_  (.A1(\u_multiplier/pp2_36 [5]),
    .A2(\u_multiplier/pp2_36 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_36_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_36_2/_20_  (.A(\u_multiplier/pp2_36 [5]),
    .B(\u_multiplier/pp2_36 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_36_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_36_2/_21_  (.A1(\u_multiplier/pp2_36 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_36_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_36_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_36_2/_22_  (.A(\u_multiplier/pp2_36 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_36_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_36_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_36_2/_23_  (.A1(\u_multiplier/pp2_36 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_36_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_36_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_36_2/_24_  (.A(\u_multiplier/pp2_36 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_36_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_36_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_36_2/_25_  (.A(\u_multiplier/STAGE3/pp3_35_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_36_2/_16_ ),
    .ZN(\u_multiplier/pp3_36 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_36_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_36_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_36_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_36_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_36_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_36_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_36_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_36_2/_17_ ),
    .ZN(\u_multiplier/pp3_37 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_37_1/_18_  (.A(\u_multiplier/STAGE3/pp3_36_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_37_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_37_1/_19_  (.A1(\u_multiplier/pp2_37 [1]),
    .A2(\u_multiplier/pp2_37 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_37_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_37_1/_20_  (.A(\u_multiplier/pp2_37 [1]),
    .B(\u_multiplier/pp2_37 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_37_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_37_1/_21_  (.A1(\u_multiplier/pp2_37 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_37_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_37_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_37_1/_22_  (.A(\u_multiplier/pp2_37 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_37_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_37_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_37_1/_23_  (.A1(\u_multiplier/pp2_37 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_37_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_37_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_37_1/_24_  (.A(\u_multiplier/pp2_37 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_37_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_37_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_37_1/_25_  (.A(\u_multiplier/STAGE3/pp3_36_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_37_1/_16_ ),
    .ZN(\u_multiplier/pp3_37 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_37_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_37_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_37_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_37_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_37_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_37_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_37_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_37_1/_17_ ),
    .ZN(\u_multiplier/pp3_38 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_37_2/_18_  (.A(\u_multiplier/STAGE3/pp3_36_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_37_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_37_2/_19_  (.A1(\u_multiplier/pp2_37 [5]),
    .A2(\u_multiplier/pp2_37 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_37_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_37_2/_20_  (.A(\u_multiplier/pp2_37 [5]),
    .B(\u_multiplier/pp2_37 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_37_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_37_2/_21_  (.A1(\u_multiplier/pp2_37 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_37_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_37_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_37_2/_22_  (.A(\u_multiplier/pp2_37 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_37_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_37_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_37_2/_23_  (.A1(\u_multiplier/pp2_37 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_37_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_37_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_37_2/_24_  (.A(\u_multiplier/pp2_37 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_37_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_37_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_37_2/_25_  (.A(\u_multiplier/STAGE3/pp3_36_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_37_2/_16_ ),
    .ZN(\u_multiplier/pp3_37 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_37_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_37_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_37_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_37_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_37_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_37_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_37_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_37_2/_17_ ),
    .ZN(\u_multiplier/pp3_38 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_38_1/_18_  (.A(\u_multiplier/STAGE3/pp3_37_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_38_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_38_1/_19_  (.A1(\u_multiplier/pp2_38 [1]),
    .A2(\u_multiplier/pp2_38 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_38_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_38_1/_20_  (.A(\u_multiplier/pp2_38 [1]),
    .B(\u_multiplier/pp2_38 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_38_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_38_1/_21_  (.A1(\u_multiplier/pp2_38 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_38_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_38_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_38_1/_22_  (.A(\u_multiplier/pp2_38 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_38_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_38_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_38_1/_23_  (.A1(\u_multiplier/pp2_38 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_38_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_38_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_38_1/_24_  (.A(\u_multiplier/pp2_38 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_38_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_38_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_38_1/_25_  (.A(\u_multiplier/STAGE3/pp3_37_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_38_1/_16_ ),
    .ZN(\u_multiplier/pp3_38 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_38_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_38_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_38_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_38_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_38_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_38_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_38_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_38_1/_17_ ),
    .ZN(\u_multiplier/pp3_39 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_38_2/_18_  (.A(\u_multiplier/STAGE3/pp3_37_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_38_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_38_2/_19_  (.A1(\u_multiplier/pp2_38 [5]),
    .A2(\u_multiplier/pp2_38 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_38_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_38_2/_20_  (.A(\u_multiplier/pp2_38 [5]),
    .B(\u_multiplier/pp2_38 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_38_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_38_2/_21_  (.A1(\u_multiplier/pp2_38 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_38_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_38_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_38_2/_22_  (.A(\u_multiplier/pp2_38 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_38_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_38_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_38_2/_23_  (.A1(\u_multiplier/pp2_38 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_38_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_38_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_38_2/_24_  (.A(\u_multiplier/pp2_38 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_38_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_38_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_38_2/_25_  (.A(\u_multiplier/STAGE3/pp3_37_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_38_2/_16_ ),
    .ZN(\u_multiplier/pp3_38 [0]));
 NAND2_X2 \u_multiplier/STAGE3/E_4_2_pp3_38_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_38_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_38_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_38_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_38_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_38_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_38_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_38_2/_17_ ),
    .ZN(\u_multiplier/pp3_39 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_39_1/_18_  (.A(\u_multiplier/STAGE3/pp3_38_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_39_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_39_1/_19_  (.A1(\u_multiplier/pp2_39 [1]),
    .A2(\u_multiplier/pp2_39 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_39_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_39_1/_20_  (.A(\u_multiplier/pp2_39 [1]),
    .B(\u_multiplier/pp2_39 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_39_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_39_1/_21_  (.A1(\u_multiplier/pp2_39 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_39_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_39_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_39_1/_22_  (.A(\u_multiplier/pp2_39 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_39_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_39_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_39_1/_23_  (.A1(\u_multiplier/pp2_39 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_39_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_39_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_39_1/_24_  (.A(\u_multiplier/pp2_39 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_39_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_39_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_39_1/_25_  (.A(\u_multiplier/STAGE3/pp3_38_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_39_1/_16_ ),
    .ZN(\u_multiplier/pp3_39 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_39_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_39_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_39_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_39_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_39_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_39_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_39_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_39_1/_17_ ),
    .ZN(\u_multiplier/pp3_40 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_39_2/_18_  (.A(\u_multiplier/STAGE3/pp3_38_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_39_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_39_2/_19_  (.A1(\u_multiplier/pp2_39 [5]),
    .A2(\u_multiplier/pp2_39 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_39_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_39_2/_20_  (.A(\u_multiplier/pp2_39 [5]),
    .B(\u_multiplier/pp2_39 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_39_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_39_2/_21_  (.A1(\u_multiplier/pp2_39 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_39_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_39_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_39_2/_22_  (.A(\u_multiplier/pp2_39 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_39_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_39_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_39_2/_23_  (.A1(\u_multiplier/pp2_39 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_39_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_39_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_39_2/_24_  (.A(\u_multiplier/pp2_39 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_39_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_39_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_39_2/_25_  (.A(\u_multiplier/STAGE3/pp3_38_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_39_2/_16_ ),
    .ZN(\u_multiplier/pp3_39 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_39_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_39_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_39_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_39_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_39_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_39_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_39_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_39_2/_17_ ),
    .ZN(\u_multiplier/pp3_40 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_40_1/_18_  (.A(\u_multiplier/STAGE3/pp3_39_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_40_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_40_1/_19_  (.A1(\u_multiplier/pp2_40 [1]),
    .A2(\u_multiplier/pp2_40 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_40_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_40_1/_20_  (.A(\u_multiplier/pp2_40 [1]),
    .B(\u_multiplier/pp2_40 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_40_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_40_1/_21_  (.A1(\u_multiplier/pp2_40 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_40_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_40_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_40_1/_22_  (.A(\u_multiplier/pp2_40 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_40_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_40_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_40_1/_23_  (.A1(\u_multiplier/pp2_40 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_40_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_40_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_40_1/_24_  (.A(\u_multiplier/pp2_40 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_40_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_40_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_40_1/_25_  (.A(\u_multiplier/STAGE3/pp3_39_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_40_1/_16_ ),
    .ZN(\u_multiplier/pp3_40 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_40_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_40_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_40_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_40_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_40_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_40_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_40_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_40_1/_17_ ),
    .ZN(\u_multiplier/pp3_41 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_40_2/_18_  (.A(\u_multiplier/STAGE3/pp3_39_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_40_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_40_2/_19_  (.A1(\u_multiplier/pp2_40 [5]),
    .A2(\u_multiplier/pp2_40 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_40_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_40_2/_20_  (.A(\u_multiplier/pp2_40 [5]),
    .B(\u_multiplier/pp2_40 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_40_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_40_2/_21_  (.A1(\u_multiplier/pp2_40 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_40_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_40_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_40_2/_22_  (.A(\u_multiplier/pp2_40 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_40_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_40_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_40_2/_23_  (.A1(\u_multiplier/pp2_40 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_40_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_40_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_40_2/_24_  (.A(\u_multiplier/pp2_40 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_40_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_40_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_40_2/_25_  (.A(\u_multiplier/STAGE3/pp3_39_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_40_2/_16_ ),
    .ZN(\u_multiplier/pp3_40 [0]));
 NAND2_X2 \u_multiplier/STAGE3/E_4_2_pp3_40_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_40_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_40_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_40_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_40_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_40_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_40_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_40_2/_17_ ),
    .ZN(\u_multiplier/pp3_41 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_41_1/_18_  (.A(\u_multiplier/STAGE3/pp3_40_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_41_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_41_1/_19_  (.A1(\u_multiplier/pp2_41 [1]),
    .A2(\u_multiplier/pp2_41 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_41_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_41_1/_20_  (.A(\u_multiplier/pp2_41 [1]),
    .B(\u_multiplier/pp2_41 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_41_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_41_1/_21_  (.A1(\u_multiplier/pp2_41 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_41_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_41_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_41_1/_22_  (.A(\u_multiplier/pp2_41 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_41_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_41_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_41_1/_23_  (.A1(\u_multiplier/pp2_41 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_41_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_41_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_41_1/_24_  (.A(\u_multiplier/pp2_41 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_41_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_41_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_41_1/_25_  (.A(\u_multiplier/STAGE3/pp3_40_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_41_1/_16_ ),
    .ZN(\u_multiplier/pp3_41 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_41_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_41_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_41_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_41_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_41_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_41_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_41_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_41_1/_17_ ),
    .ZN(\u_multiplier/pp3_42 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_41_2/_18_  (.A(\u_multiplier/STAGE3/pp3_40_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_41_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_41_2/_19_  (.A1(\u_multiplier/pp2_41 [5]),
    .A2(\u_multiplier/pp2_41 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_41_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_41_2/_20_  (.A(\u_multiplier/pp2_41 [5]),
    .B(\u_multiplier/pp2_41 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_41_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_41_2/_21_  (.A1(\u_multiplier/pp2_41 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_41_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_41_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_41_2/_22_  (.A(\u_multiplier/pp2_41 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_41_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_41_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_41_2/_23_  (.A1(\u_multiplier/pp2_41 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_41_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_41_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_41_2/_24_  (.A(\u_multiplier/pp2_41 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_41_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_41_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_41_2/_25_  (.A(\u_multiplier/STAGE3/pp3_40_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_41_2/_16_ ),
    .ZN(\u_multiplier/pp3_41 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_41_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_41_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_41_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_41_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_41_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_41_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_41_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_41_2/_17_ ),
    .ZN(\u_multiplier/pp3_42 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_42_1/_18_  (.A(\u_multiplier/STAGE3/pp3_41_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_42_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_42_1/_19_  (.A1(\u_multiplier/pp2_42 [1]),
    .A2(\u_multiplier/pp2_42 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_42_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_42_1/_20_  (.A(\u_multiplier/pp2_42 [1]),
    .B(\u_multiplier/pp2_42 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_42_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_42_1/_21_  (.A1(\u_multiplier/pp2_42 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_42_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_42_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_42_1/_22_  (.A(\u_multiplier/pp2_42 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_42_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_42_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_42_1/_23_  (.A1(\u_multiplier/pp2_42 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_42_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_42_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_42_1/_24_  (.A(\u_multiplier/pp2_42 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_42_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_42_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_42_1/_25_  (.A(\u_multiplier/STAGE3/pp3_41_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_42_1/_16_ ),
    .ZN(\u_multiplier/pp3_42 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_42_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_42_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_42_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_42_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_42_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_42_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_42_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_42_1/_17_ ),
    .ZN(\u_multiplier/pp3_43 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_42_2/_18_  (.A(\u_multiplier/STAGE3/pp3_41_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_42_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_42_2/_19_  (.A1(\u_multiplier/pp2_42 [5]),
    .A2(\u_multiplier/pp2_42 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_42_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_42_2/_20_  (.A(\u_multiplier/pp2_42 [5]),
    .B(\u_multiplier/pp2_42 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_42_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_42_2/_21_  (.A1(\u_multiplier/pp2_42 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_42_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_42_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_42_2/_22_  (.A(\u_multiplier/pp2_42 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_42_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_42_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_42_2/_23_  (.A1(\u_multiplier/pp2_42 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_42_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_42_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_42_2/_24_  (.A(\u_multiplier/pp2_42 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_42_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_42_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_42_2/_25_  (.A(\u_multiplier/STAGE3/pp3_41_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_42_2/_16_ ),
    .ZN(\u_multiplier/pp3_42 [0]));
 NAND2_X2 \u_multiplier/STAGE3/E_4_2_pp3_42_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_42_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_42_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_42_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_42_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_42_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_42_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_42_2/_17_ ),
    .ZN(\u_multiplier/pp3_43 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_43_1/_18_  (.A(\u_multiplier/STAGE3/pp3_42_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_43_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_43_1/_19_  (.A1(\u_multiplier/pp2_43 [1]),
    .A2(\u_multiplier/pp2_43 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_43_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_43_1/_20_  (.A(\u_multiplier/pp2_43 [1]),
    .B(\u_multiplier/pp2_43 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_43_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_43_1/_21_  (.A1(\u_multiplier/pp2_43 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_43_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_43_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_43_1/_22_  (.A(\u_multiplier/pp2_43 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_43_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_43_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_43_1/_23_  (.A1(\u_multiplier/pp2_43 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_43_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_43_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_43_1/_24_  (.A(\u_multiplier/pp2_43 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_43_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_43_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_43_1/_25_  (.A(\u_multiplier/STAGE3/pp3_42_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_43_1/_16_ ),
    .ZN(\u_multiplier/pp3_43 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_43_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_43_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_43_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_43_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_43_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_43_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_43_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_43_1/_17_ ),
    .ZN(\u_multiplier/pp3_44 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_43_2/_18_  (.A(\u_multiplier/STAGE3/pp3_42_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_43_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_43_2/_19_  (.A1(\u_multiplier/pp2_43 [5]),
    .A2(\u_multiplier/pp2_43 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_43_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_43_2/_20_  (.A(\u_multiplier/pp2_43 [5]),
    .B(\u_multiplier/pp2_43 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_43_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_43_2/_21_  (.A1(\u_multiplier/pp2_43 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_43_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_43_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_43_2/_22_  (.A(\u_multiplier/pp2_43 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_43_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_43_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_43_2/_23_  (.A1(\u_multiplier/pp2_43 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_43_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_43_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_43_2/_24_  (.A(\u_multiplier/pp2_43 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_43_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_43_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_43_2/_25_  (.A(\u_multiplier/STAGE3/pp3_42_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_43_2/_16_ ),
    .ZN(\u_multiplier/pp3_43 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_43_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_43_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_43_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_43_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_43_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_43_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_43_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_43_2/_17_ ),
    .ZN(\u_multiplier/pp3_44 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_44_1/_18_  (.A(\u_multiplier/STAGE3/pp3_43_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_44_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_44_1/_19_  (.A1(\u_multiplier/pp2_44 [1]),
    .A2(\u_multiplier/pp2_44 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_44_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_44_1/_20_  (.A(\u_multiplier/pp2_44 [1]),
    .B(\u_multiplier/pp2_44 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_44_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_44_1/_21_  (.A1(\u_multiplier/pp2_44 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_44_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_44_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_44_1/_22_  (.A(\u_multiplier/pp2_44 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_44_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_44_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_44_1/_23_  (.A1(\u_multiplier/pp2_44 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_44_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_44_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_44_1/_24_  (.A(\u_multiplier/pp2_44 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_44_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_44_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_44_1/_25_  (.A(\u_multiplier/STAGE3/pp3_43_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_44_1/_16_ ),
    .ZN(\u_multiplier/pp3_44 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_44_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_44_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_44_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_44_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_44_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_44_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_44_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_44_1/_17_ ),
    .ZN(\u_multiplier/pp3_45 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_44_2/_18_  (.A(\u_multiplier/STAGE3/pp3_43_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_44_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_44_2/_19_  (.A1(\u_multiplier/pp2_44 [5]),
    .A2(\u_multiplier/pp2_44 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_44_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_44_2/_20_  (.A(\u_multiplier/pp2_44 [5]),
    .B(\u_multiplier/pp2_44 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_44_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_44_2/_21_  (.A1(\u_multiplier/pp2_44 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_44_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_44_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_44_2/_22_  (.A(\u_multiplier/pp2_44 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_44_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_44_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_44_2/_23_  (.A1(\u_multiplier/pp2_44 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_44_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_44_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_44_2/_24_  (.A(\u_multiplier/pp2_44 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_44_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_44_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_44_2/_25_  (.A(\u_multiplier/STAGE3/pp3_43_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_44_2/_16_ ),
    .ZN(\u_multiplier/pp3_44 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_44_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_44_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_44_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_44_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_44_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_44_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_44_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_44_2/_17_ ),
    .ZN(\u_multiplier/pp3_45 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_45_1/_18_  (.A(\u_multiplier/STAGE3/pp3_44_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_45_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_45_1/_19_  (.A1(\u_multiplier/pp2_45 [1]),
    .A2(\u_multiplier/pp2_45 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_45_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_45_1/_20_  (.A(\u_multiplier/pp2_45 [1]),
    .B(\u_multiplier/pp2_45 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_45_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_45_1/_21_  (.A1(\u_multiplier/pp2_45 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_45_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_45_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_45_1/_22_  (.A(\u_multiplier/pp2_45 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_45_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_45_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_45_1/_23_  (.A1(\u_multiplier/pp2_45 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_45_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_45_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_45_1/_24_  (.A(\u_multiplier/pp2_45 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_45_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_45_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_45_1/_25_  (.A(\u_multiplier/STAGE3/pp3_44_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_45_1/_16_ ),
    .ZN(\u_multiplier/pp3_45 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_45_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_45_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_45_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_45_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_45_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_45_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_45_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_45_1/_17_ ),
    .ZN(\u_multiplier/pp3_46 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_45_2/_18_  (.A(\u_multiplier/STAGE3/pp3_44_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_45_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_45_2/_19_  (.A1(\u_multiplier/pp2_45 [5]),
    .A2(\u_multiplier/pp2_45 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_45_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_45_2/_20_  (.A(\u_multiplier/pp2_45 [5]),
    .B(\u_multiplier/pp2_45 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_45_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_45_2/_21_  (.A1(\u_multiplier/pp2_45 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_45_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_45_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_45_2/_22_  (.A(\u_multiplier/pp2_45 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_45_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_45_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_45_2/_23_  (.A1(\u_multiplier/pp2_45 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_45_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_45_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_45_2/_24_  (.A(\u_multiplier/pp2_45 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_45_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_45_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_45_2/_25_  (.A(\u_multiplier/STAGE3/pp3_44_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_45_2/_16_ ),
    .ZN(\u_multiplier/pp3_45 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_45_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_45_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_45_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_45_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_45_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_45_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_45_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_45_2/_17_ ),
    .ZN(\u_multiplier/pp3_46 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_46_1/_18_  (.A(\u_multiplier/STAGE3/pp3_45_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_46_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_46_1/_19_  (.A1(\u_multiplier/pp2_46 [1]),
    .A2(\u_multiplier/pp2_46 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_46_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_46_1/_20_  (.A(\u_multiplier/pp2_46 [1]),
    .B(\u_multiplier/pp2_46 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_46_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_46_1/_21_  (.A1(\u_multiplier/pp2_46 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_46_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_46_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_46_1/_22_  (.A(\u_multiplier/pp2_46 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_46_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_46_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_46_1/_23_  (.A1(\u_multiplier/pp2_46 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_46_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_46_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_46_1/_24_  (.A(\u_multiplier/pp2_46 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_46_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_46_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_46_1/_25_  (.A(\u_multiplier/STAGE3/pp3_45_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_46_1/_16_ ),
    .ZN(\u_multiplier/pp3_46 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_46_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_46_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_46_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_46_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_46_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_46_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_46_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_46_1/_17_ ),
    .ZN(\u_multiplier/pp3_47 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_46_2/_18_  (.A(\u_multiplier/STAGE3/pp3_45_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_46_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_46_2/_19_  (.A1(\u_multiplier/pp2_46 [5]),
    .A2(\u_multiplier/pp2_46 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_46_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_46_2/_20_  (.A(\u_multiplier/pp2_46 [5]),
    .B(\u_multiplier/pp2_46 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_46_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_46_2/_21_  (.A1(\u_multiplier/pp2_46 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_46_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_46_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_46_2/_22_  (.A(\u_multiplier/pp2_46 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_46_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_46_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_46_2/_23_  (.A1(\u_multiplier/pp2_46 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_46_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_46_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_46_2/_24_  (.A(\u_multiplier/pp2_46 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_46_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_46_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_46_2/_25_  (.A(\u_multiplier/STAGE3/pp3_45_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_46_2/_16_ ),
    .ZN(\u_multiplier/pp3_46 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_46_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_46_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_46_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_46_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_46_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_46_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_46_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_46_2/_17_ ),
    .ZN(\u_multiplier/pp3_47 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_47_1/_18_  (.A(\u_multiplier/STAGE3/pp3_46_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_47_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_47_1/_19_  (.A1(\u_multiplier/pp2_47 [1]),
    .A2(\u_multiplier/pp2_47 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_47_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_47_1/_20_  (.A(\u_multiplier/pp2_47 [1]),
    .B(\u_multiplier/pp2_47 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_47_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_47_1/_21_  (.A1(\u_multiplier/pp2_47 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_47_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_47_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_47_1/_22_  (.A(\u_multiplier/pp2_47 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_47_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_47_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_47_1/_23_  (.A1(\u_multiplier/pp2_47 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_47_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_47_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_47_1/_24_  (.A(\u_multiplier/pp2_47 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_47_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_47_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_47_1/_25_  (.A(\u_multiplier/STAGE3/pp3_46_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_47_1/_16_ ),
    .ZN(\u_multiplier/pp3_47 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_47_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_47_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_47_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_47_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_47_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_47_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_47_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_47_1/_17_ ),
    .ZN(\u_multiplier/pp3_48 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_47_2/_18_  (.A(\u_multiplier/STAGE3/pp3_46_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_47_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_47_2/_19_  (.A1(\u_multiplier/pp2_47 [5]),
    .A2(\u_multiplier/pp2_47 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_47_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_47_2/_20_  (.A(\u_multiplier/pp2_47 [5]),
    .B(\u_multiplier/pp2_47 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_47_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_47_2/_21_  (.A1(\u_multiplier/pp2_47 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_47_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_47_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_47_2/_22_  (.A(\u_multiplier/pp2_47 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_47_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_47_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_47_2/_23_  (.A1(\u_multiplier/pp2_47 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_47_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_47_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_47_2/_24_  (.A(\u_multiplier/pp2_47 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_47_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_47_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_47_2/_25_  (.A(\u_multiplier/STAGE3/pp3_46_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_47_2/_16_ ),
    .ZN(\u_multiplier/pp3_47 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_47_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_47_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_47_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_47_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_47_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_47_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_47_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_47_2/_17_ ),
    .ZN(\u_multiplier/pp3_48 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_48_1/_18_  (.A(\u_multiplier/STAGE3/pp3_47_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_48_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_48_1/_19_  (.A1(\u_multiplier/pp2_48 [1]),
    .A2(\u_multiplier/pp2_48 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_48_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_48_1/_20_  (.A(\u_multiplier/pp2_48 [1]),
    .B(\u_multiplier/pp2_48 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_48_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_48_1/_21_  (.A1(\u_multiplier/pp2_48 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_48_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_48_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_48_1/_22_  (.A(\u_multiplier/pp2_48 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_48_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_48_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_48_1/_23_  (.A1(\u_multiplier/pp2_48 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_48_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_48_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_48_1/_24_  (.A(\u_multiplier/pp2_48 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_48_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_48_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_48_1/_25_  (.A(\u_multiplier/STAGE3/pp3_47_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_48_1/_16_ ),
    .ZN(\u_multiplier/pp3_48 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_48_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_48_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_48_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_48_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_48_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_48_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_48_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_48_1/_17_ ),
    .ZN(\u_multiplier/pp3_49 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_48_2/_18_  (.A(\u_multiplier/STAGE3/pp3_47_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_48_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_48_2/_19_  (.A1(\u_multiplier/pp2_48 [5]),
    .A2(\u_multiplier/pp2_48 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_48_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_48_2/_20_  (.A(\u_multiplier/pp2_48 [5]),
    .B(\u_multiplier/pp2_48 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_48_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_48_2/_21_  (.A1(\u_multiplier/pp2_48 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_48_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_48_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_48_2/_22_  (.A(\u_multiplier/pp2_48 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_48_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_48_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_48_2/_23_  (.A1(\u_multiplier/pp2_48 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_48_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_48_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_48_2/_24_  (.A(\u_multiplier/pp2_48 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_48_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_48_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_48_2/_25_  (.A(\u_multiplier/STAGE3/pp3_47_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_48_2/_16_ ),
    .ZN(\u_multiplier/pp3_48 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_48_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_48_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_48_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_48_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_48_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_48_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_48_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_48_2/_17_ ),
    .ZN(\u_multiplier/pp3_49 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_49_1/_18_  (.A(\u_multiplier/STAGE3/pp3_48_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_49_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_49_1/_19_  (.A1(\u_multiplier/pp2_49 [1]),
    .A2(\u_multiplier/pp2_49 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_49_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_49_1/_20_  (.A(\u_multiplier/pp2_49 [1]),
    .B(\u_multiplier/pp2_49 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_49_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_49_1/_21_  (.A1(\u_multiplier/pp2_49 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_49_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_49_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_49_1/_22_  (.A(\u_multiplier/pp2_49 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_49_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_49_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_49_1/_23_  (.A1(\u_multiplier/pp2_49 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_49_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_49_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_49_1/_24_  (.A(\u_multiplier/pp2_49 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_49_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_49_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_49_1/_25_  (.A(\u_multiplier/STAGE3/pp3_48_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_49_1/_16_ ),
    .ZN(\u_multiplier/pp3_49 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_49_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_49_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_49_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_49_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_49_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_49_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_49_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_49_1/_17_ ),
    .ZN(\u_multiplier/pp3_50 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_49_2/_18_  (.A(\u_multiplier/STAGE3/pp3_48_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_49_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_49_2/_19_  (.A1(\u_multiplier/pp2_49 [5]),
    .A2(\u_multiplier/pp2_49 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_49_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_49_2/_20_  (.A(\u_multiplier/pp2_49 [5]),
    .B(\u_multiplier/pp2_49 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_49_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_49_2/_21_  (.A1(\u_multiplier/pp2_49 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_49_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_49_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_49_2/_22_  (.A(\u_multiplier/pp2_49 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_49_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_49_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_49_2/_23_  (.A1(\u_multiplier/pp2_49 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_49_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_49_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_49_2/_24_  (.A(\u_multiplier/pp2_49 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_49_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_49_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_49_2/_25_  (.A(\u_multiplier/STAGE3/pp3_48_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_49_2/_16_ ),
    .ZN(\u_multiplier/pp3_49 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_49_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_49_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_49_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_49_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_49_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_49_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_49_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_49_2/_17_ ),
    .ZN(\u_multiplier/pp3_50 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_50_1/_18_  (.A(\u_multiplier/STAGE3/pp3_49_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_50_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_50_1/_19_  (.A1(\u_multiplier/pp2_50 [1]),
    .A2(\u_multiplier/pp2_50 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_50_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_50_1/_20_  (.A(\u_multiplier/pp2_50 [1]),
    .B(\u_multiplier/pp2_50 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_50_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_50_1/_21_  (.A1(\u_multiplier/pp2_50 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_50_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_50_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_50_1/_22_  (.A(\u_multiplier/pp2_50 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_50_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_50_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_50_1/_23_  (.A1(\u_multiplier/pp2_50 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_50_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_50_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_50_1/_24_  (.A(\u_multiplier/pp2_50 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_50_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_50_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_50_1/_25_  (.A(\u_multiplier/STAGE3/pp3_49_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_50_1/_16_ ),
    .ZN(\u_multiplier/pp3_50 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_50_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_50_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_50_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_50_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_50_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_50_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_50_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_50_1/_17_ ),
    .ZN(\u_multiplier/pp3_51 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_50_2/_18_  (.A(\u_multiplier/STAGE3/pp3_49_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_50_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_50_2/_19_  (.A1(\u_multiplier/pp2_50 [5]),
    .A2(\u_multiplier/pp2_50 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_50_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_50_2/_20_  (.A(\u_multiplier/pp2_50 [5]),
    .B(\u_multiplier/pp2_50 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_50_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_50_2/_21_  (.A1(\u_multiplier/pp2_50 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_50_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_50_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_50_2/_22_  (.A(\u_multiplier/pp2_50 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_50_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_50_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_50_2/_23_  (.A1(\u_multiplier/pp2_50 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_50_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_50_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_50_2/_24_  (.A(\u_multiplier/pp2_50 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_50_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_50_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_50_2/_25_  (.A(\u_multiplier/STAGE3/pp3_49_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_50_2/_16_ ),
    .ZN(\u_multiplier/pp3_50 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_50_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_50_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_50_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_50_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_50_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_50_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_50_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_50_2/_17_ ),
    .ZN(\u_multiplier/pp3_51 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_51_1/_18_  (.A(\u_multiplier/STAGE3/pp3_50_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_51_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_51_1/_19_  (.A1(\u_multiplier/pp2_51 [1]),
    .A2(\u_multiplier/pp2_51 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_51_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_51_1/_20_  (.A(\u_multiplier/pp2_51 [1]),
    .B(\u_multiplier/pp2_51 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_51_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_51_1/_21_  (.A1(\u_multiplier/pp2_51 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_51_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_51_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_51_1/_22_  (.A(\u_multiplier/pp2_51 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_51_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_51_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_51_1/_23_  (.A1(\u_multiplier/pp2_51 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_51_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_51_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_51_1/_24_  (.A(\u_multiplier/pp2_51 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_51_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_51_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_51_1/_25_  (.A(\u_multiplier/STAGE3/pp3_50_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_51_1/_16_ ),
    .ZN(\u_multiplier/pp3_51 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_51_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_51_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_51_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_51_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_51_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_51_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_51_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_51_1/_17_ ),
    .ZN(\u_multiplier/pp3_52 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_51_2/_18_  (.A(\u_multiplier/STAGE3/pp3_50_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_51_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_51_2/_19_  (.A1(\u_multiplier/pp2_51 [5]),
    .A2(\u_multiplier/pp2_51 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_51_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_51_2/_20_  (.A(\u_multiplier/pp2_51 [5]),
    .B(\u_multiplier/pp2_51 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_51_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_51_2/_21_  (.A1(\u_multiplier/pp2_51 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_51_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_51_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_51_2/_22_  (.A(\u_multiplier/pp2_51 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_51_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_51_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_51_2/_23_  (.A1(\u_multiplier/pp2_51 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_51_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_51_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_51_2/_24_  (.A(\u_multiplier/pp2_51 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_51_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_51_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_51_2/_25_  (.A(\u_multiplier/STAGE3/pp3_50_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_51_2/_16_ ),
    .ZN(\u_multiplier/pp3_51 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_51_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_51_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_51_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_51_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_51_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_51_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_51_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_51_2/_17_ ),
    .ZN(\u_multiplier/pp3_52 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_52_1/_18_  (.A(\u_multiplier/STAGE3/pp3_51_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_52_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_52_1/_19_  (.A1(\u_multiplier/pp2_52 [1]),
    .A2(\u_multiplier/pp2_52 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_52_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_52_1/_20_  (.A(\u_multiplier/pp2_52 [1]),
    .B(\u_multiplier/pp2_52 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_52_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_52_1/_21_  (.A1(\u_multiplier/pp2_52 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_52_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_52_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_52_1/_22_  (.A(\u_multiplier/pp2_52 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_52_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_52_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_52_1/_23_  (.A1(\u_multiplier/pp2_52 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_52_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_52_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_52_1/_24_  (.A(\u_multiplier/pp2_52 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_52_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_52_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_52_1/_25_  (.A(\u_multiplier/STAGE3/pp3_51_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_52_1/_16_ ),
    .ZN(\u_multiplier/pp3_52 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_52_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_52_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_52_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_52_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_52_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_52_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_52_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_52_1/_17_ ),
    .ZN(\u_multiplier/pp3_53 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_52_2/_18_  (.A(\u_multiplier/STAGE3/pp3_51_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_52_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_52_2/_19_  (.A1(\u_multiplier/pp2_52 [5]),
    .A2(\u_multiplier/pp2_52 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_52_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_52_2/_20_  (.A(\u_multiplier/pp2_52 [5]),
    .B(\u_multiplier/pp2_52 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_52_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_52_2/_21_  (.A1(\u_multiplier/pp2_52 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_52_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_52_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_52_2/_22_  (.A(\u_multiplier/pp2_52 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_52_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_52_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_52_2/_23_  (.A1(\u_multiplier/pp2_52 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_52_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_52_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_52_2/_24_  (.A(\u_multiplier/pp2_52 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_52_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_52_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_52_2/_25_  (.A(\u_multiplier/STAGE3/pp3_51_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_52_2/_16_ ),
    .ZN(\u_multiplier/pp3_52 [0]));
 NAND2_X2 \u_multiplier/STAGE3/E_4_2_pp3_52_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_52_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_52_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_52_e42_2_cout ));
 OAI21_X4 \u_multiplier/STAGE3/E_4_2_pp3_52_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_52_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_52_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_52_2/_17_ ),
    .ZN(\u_multiplier/pp3_53 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_53_1/_18_  (.A(\u_multiplier/STAGE3/pp3_52_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_53_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_53_1/_19_  (.A1(\u_multiplier/pp2_53 [1]),
    .A2(\u_multiplier/pp2_53 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_53_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_53_1/_20_  (.A(\u_multiplier/pp2_53 [1]),
    .B(\u_multiplier/pp2_53 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_53_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_53_1/_21_  (.A1(\u_multiplier/pp2_53 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_53_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_53_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_53_1/_22_  (.A(\u_multiplier/pp2_53 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_53_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_53_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_53_1/_23_  (.A1(\u_multiplier/pp2_53 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_53_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_53_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_53_1/_24_  (.A(\u_multiplier/pp2_53 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_53_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_53_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_53_1/_25_  (.A(\u_multiplier/STAGE3/pp3_52_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_53_1/_16_ ),
    .ZN(\u_multiplier/pp3_53 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_53_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_53_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_53_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_53_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_53_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_53_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_53_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_53_1/_17_ ),
    .ZN(\u_multiplier/pp3_54 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_53_2/_18_  (.A(\u_multiplier/STAGE3/pp3_52_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_53_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_53_2/_19_  (.A1(\u_multiplier/pp2_53 [5]),
    .A2(\u_multiplier/pp2_53 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_53_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_53_2/_20_  (.A(\u_multiplier/pp2_53 [5]),
    .B(\u_multiplier/pp2_53 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_53_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_53_2/_21_  (.A1(\u_multiplier/pp2_53 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_53_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_53_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_53_2/_22_  (.A(\u_multiplier/pp2_53 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_53_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_53_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_53_2/_23_  (.A1(\u_multiplier/pp2_53 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_53_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_53_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_53_2/_24_  (.A(\u_multiplier/pp2_53 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_53_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_53_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_53_2/_25_  (.A(\u_multiplier/STAGE3/pp3_52_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_53_2/_16_ ),
    .ZN(\u_multiplier/pp3_53 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_53_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_53_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_53_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_53_e42_2_cout ));
 OAI21_X4 \u_multiplier/STAGE3/E_4_2_pp3_53_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_53_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_53_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_53_2/_17_ ),
    .ZN(\u_multiplier/pp3_54 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_54_1/_18_  (.A(\u_multiplier/STAGE3/pp3_53_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_54_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_54_1/_19_  (.A1(\u_multiplier/pp2_54 [1]),
    .A2(\u_multiplier/pp2_54 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_54_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_54_1/_20_  (.A(\u_multiplier/pp2_54 [1]),
    .B(\u_multiplier/pp2_54 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_54_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_54_1/_21_  (.A1(\u_multiplier/pp2_54 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_54_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_54_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_54_1/_22_  (.A(\u_multiplier/pp2_54 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_54_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_54_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_54_1/_23_  (.A1(\u_multiplier/pp2_54 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_54_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_54_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_54_1/_24_  (.A(\u_multiplier/pp2_54 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_54_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_54_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_54_1/_25_  (.A(\u_multiplier/STAGE3/pp3_53_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_54_1/_16_ ),
    .ZN(\u_multiplier/pp3_54 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_54_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_54_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_54_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_54_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_54_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_54_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_54_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_54_1/_17_ ),
    .ZN(\u_multiplier/pp3_55 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_54_2/_18_  (.A(\u_multiplier/STAGE3/pp3_53_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_54_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_54_2/_19_  (.A1(\u_multiplier/pp2_54 [5]),
    .A2(\u_multiplier/pp2_54 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_54_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_54_2/_20_  (.A(\u_multiplier/pp2_54 [5]),
    .B(\u_multiplier/pp2_54 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_54_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_54_2/_21_  (.A1(\u_multiplier/pp2_54 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_54_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_54_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_54_2/_22_  (.A(\u_multiplier/pp2_54 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_54_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_54_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_54_2/_23_  (.A1(\u_multiplier/pp2_54 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_54_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_54_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_54_2/_24_  (.A(\u_multiplier/pp2_54 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_54_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_54_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_54_2/_25_  (.A(\u_multiplier/STAGE3/pp3_53_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_54_2/_16_ ),
    .ZN(\u_multiplier/pp3_54 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_54_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_54_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_54_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_54_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_54_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_54_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_54_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_54_2/_17_ ),
    .ZN(\u_multiplier/pp3_55 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_55_1/_18_  (.A(\u_multiplier/STAGE3/pp3_54_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_55_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_55_1/_19_  (.A1(\u_multiplier/pp2_55 [1]),
    .A2(\u_multiplier/pp2_55 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_55_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_55_1/_20_  (.A(\u_multiplier/pp2_55 [1]),
    .B(\u_multiplier/pp2_55 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_55_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_55_1/_21_  (.A1(\u_multiplier/pp2_55 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_55_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_55_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_55_1/_22_  (.A(\u_multiplier/pp2_55 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_55_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_55_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_55_1/_23_  (.A1(\u_multiplier/pp2_55 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_55_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_55_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_55_1/_24_  (.A(\u_multiplier/pp2_55 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_55_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_55_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_55_1/_25_  (.A(\u_multiplier/STAGE3/pp3_54_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_55_1/_16_ ),
    .ZN(\u_multiplier/pp3_55 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_55_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_55_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_55_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_55_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_55_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_55_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_55_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_55_1/_17_ ),
    .ZN(\u_multiplier/pp3_56 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_55_2/_18_  (.A(\u_multiplier/STAGE3/pp3_54_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_55_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_55_2/_19_  (.A1(\u_multiplier/pp2_55 [5]),
    .A2(\u_multiplier/pp2_55 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_55_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_55_2/_20_  (.A(\u_multiplier/pp2_55 [5]),
    .B(\u_multiplier/pp2_55 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_55_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_55_2/_21_  (.A1(\u_multiplier/pp2_55 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_55_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_55_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_55_2/_22_  (.A(\u_multiplier/pp2_55 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_55_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_55_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_55_2/_23_  (.A1(\u_multiplier/pp2_55 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_55_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_55_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_55_2/_24_  (.A(\u_multiplier/pp2_55 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_55_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_55_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_55_2/_25_  (.A(\u_multiplier/STAGE3/pp3_54_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_55_2/_16_ ),
    .ZN(\u_multiplier/pp3_55 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_55_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_55_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_55_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_55_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_55_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_55_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_55_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_55_2/_17_ ),
    .ZN(\u_multiplier/pp3_56 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_56_1/_18_  (.A(\u_multiplier/STAGE3/pp3_55_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_56_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_56_1/_19_  (.A1(\u_multiplier/pp2_56 [1]),
    .A2(\u_multiplier/pp2_56 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_56_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_56_1/_20_  (.A(\u_multiplier/pp2_56 [1]),
    .B(\u_multiplier/pp2_56 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_56_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_56_1/_21_  (.A1(\u_multiplier/pp2_56 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_56_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_56_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_56_1/_22_  (.A(\u_multiplier/pp2_56 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_56_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_56_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_56_1/_23_  (.A1(\u_multiplier/pp2_56 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_56_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_56_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_56_1/_24_  (.A(\u_multiplier/pp2_56 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_56_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_56_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_56_1/_25_  (.A(\u_multiplier/STAGE3/pp3_55_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_56_1/_16_ ),
    .ZN(\u_multiplier/pp3_56 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_56_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_56_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_56_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_56_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_56_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_56_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_56_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_56_1/_17_ ),
    .ZN(\u_multiplier/pp3_57 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_56_2/_18_  (.A(\u_multiplier/STAGE3/pp3_55_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_56_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_56_2/_19_  (.A1(\u_multiplier/pp2_56 [5]),
    .A2(\u_multiplier/pp2_56 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_56_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_56_2/_20_  (.A(\u_multiplier/pp2_56 [5]),
    .B(\u_multiplier/pp2_56 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_56_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_56_2/_21_  (.A1(\u_multiplier/pp2_56 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_56_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_56_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_56_2/_22_  (.A(\u_multiplier/pp2_56 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_56_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_56_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_56_2/_23_  (.A1(\u_multiplier/pp2_56 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_56_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_56_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_56_2/_24_  (.A(\u_multiplier/pp2_56 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_56_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_56_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_56_2/_25_  (.A(\u_multiplier/STAGE3/pp3_55_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_56_2/_16_ ),
    .ZN(\u_multiplier/pp3_56 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_56_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_56_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_56_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_56_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_56_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_56_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_56_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_56_2/_17_ ),
    .ZN(\u_multiplier/pp3_57 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_57_1/_18_  (.A(\u_multiplier/STAGE3/pp3_56_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_57_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_57_1/_19_  (.A1(\u_multiplier/pp2_57 [1]),
    .A2(\u_multiplier/pp2_57 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_57_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_57_1/_20_  (.A(\u_multiplier/pp2_57 [1]),
    .B(\u_multiplier/pp2_57 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_57_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_57_1/_21_  (.A1(\u_multiplier/pp2_57 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_57_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_57_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_57_1/_22_  (.A(\u_multiplier/pp2_57 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_57_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_57_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_57_1/_23_  (.A1(\u_multiplier/pp2_57 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_57_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_57_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_57_1/_24_  (.A(\u_multiplier/pp2_57 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_57_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_57_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_57_1/_25_  (.A(\u_multiplier/STAGE3/pp3_56_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_57_1/_16_ ),
    .ZN(\u_multiplier/pp3_57 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_57_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_57_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_57_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_57_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_57_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_57_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_57_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_57_1/_17_ ),
    .ZN(\u_multiplier/pp3_58 [1]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_58_1/_18_  (.A(\u_multiplier/STAGE3/pp3_57_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_58_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_58_1/_19_  (.A1(\u_multiplier/pp2_58 [1]),
    .A2(\u_multiplier/pp2_58 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_58_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_58_1/_20_  (.A(\u_multiplier/pp2_58 [1]),
    .B(\u_multiplier/pp2_58 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_58_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_58_1/_21_  (.A1(\u_multiplier/pp2_58 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_58_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_58_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_58_1/_22_  (.A(\u_multiplier/pp2_58 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_58_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_58_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_58_1/_23_  (.A1(\u_multiplier/pp2_58 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_58_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_58_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_58_1/_24_  (.A(\u_multiplier/pp2_58 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_58_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_58_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_58_1/_25_  (.A(\u_multiplier/STAGE3/pp3_57_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_58_1/_16_ ),
    .ZN(\u_multiplier/pp3_58 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_58_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_58_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_58_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_58_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_58_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_58_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_58_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_58_1/_17_ ),
    .ZN(\u_multiplier/pp3_59 [1]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_5_1/_18_  (.A(net143),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_5_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_5_1/_19_  (.A1(\u_multiplier/pp2_5 [1]),
    .A2(\u_multiplier/pp2_5 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_5_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_5_1/_20_  (.A(\u_multiplier/pp2_5 [1]),
    .B(\u_multiplier/pp2_5 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_5_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_5_1/_21_  (.A1(\u_multiplier/pp2_5 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_5_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_5_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_5_1/_22_  (.A(\u_multiplier/pp2_5 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_5_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_5_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_5_1/_23_  (.A1(\u_multiplier/pp2_5 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_5_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_5_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_5_1/_24_  (.A(\u_multiplier/pp2_5 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_5_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_5_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_5_1/_25_  (.A(net144),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_5_1/_16_ ),
    .ZN(\u_multiplier/pp3_5 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_5_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_5_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_5_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_5_e42_1_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_5_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_5_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_5_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_5_1/_17_ ),
    .ZN(\u_multiplier/pp3_6 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_6_1/_18_  (.A(\u_multiplier/STAGE3/pp3_5_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_6_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_6_1/_19_  (.A1(\u_multiplier/pp2_6 [1]),
    .A2(\u_multiplier/pp2_6 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_6_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_6_1/_20_  (.A(\u_multiplier/pp2_6 [1]),
    .B(\u_multiplier/pp2_6 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_6_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_6_1/_21_  (.A1(\u_multiplier/pp2_6 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_6_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_6_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_6_1/_22_  (.A(\u_multiplier/pp2_6 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_6_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_6_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_6_1/_23_  (.A1(\u_multiplier/pp2_6 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_6_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_6_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_6_1/_24_  (.A(\u_multiplier/pp2_6 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_6_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_6_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_6_1/_25_  (.A(\u_multiplier/STAGE3/pp3_5_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_6_1/_16_ ),
    .ZN(\u_multiplier/pp3_6 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_6_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_6_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_6_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_6_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_6_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_6_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_6_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_6_1/_17_ ),
    .ZN(\u_multiplier/pp3_7 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_7_1/_18_  (.A(\u_multiplier/STAGE3/pp3_6_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_7_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_7_1/_19_  (.A1(\u_multiplier/pp2_7 [1]),
    .A2(\u_multiplier/pp2_7 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_7_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_7_1/_20_  (.A(\u_multiplier/pp2_7 [1]),
    .B(\u_multiplier/pp2_7 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_7_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_7_1/_21_  (.A1(\u_multiplier/pp2_7 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_7_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_7_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_7_1/_22_  (.A(\u_multiplier/pp2_7 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_7_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_7_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_7_1/_23_  (.A1(\u_multiplier/pp2_7 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_7_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_7_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_7_1/_24_  (.A(\u_multiplier/pp2_7 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_7_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_7_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_7_1/_25_  (.A(\u_multiplier/STAGE3/pp3_6_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_7_1/_16_ ),
    .ZN(\u_multiplier/pp3_7 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_7_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_7_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_7_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_7_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_7_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_7_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_7_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_7_1/_17_ ),
    .ZN(\u_multiplier/pp3_8 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_7_2/_18_  (.A(net145),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_7_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_7_2/_19_  (.A1(\u_multiplier/pp2_7 [5]),
    .A2(\u_multiplier/pp2_7 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_7_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_7_2/_20_  (.A(\u_multiplier/pp2_7 [5]),
    .B(\u_multiplier/pp2_7 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_7_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_7_2/_21_  (.A1(\u_multiplier/pp2_7 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_7_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_7_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_7_2/_22_  (.A(\u_multiplier/pp2_7 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_7_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_7_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_7_2/_23_  (.A1(\u_multiplier/pp2_7 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_7_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_7_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_7_2/_24_  (.A(\u_multiplier/pp2_7 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_7_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_7_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_7_2/_25_  (.A(net146),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_7_2/_16_ ),
    .ZN(\u_multiplier/pp3_7 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_7_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_7_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_7_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_7_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_7_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_7_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_7_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_7_2/_17_ ),
    .ZN(\u_multiplier/pp3_8 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_8_1/_18_  (.A(\u_multiplier/STAGE3/pp3_7_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_8_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_8_1/_19_  (.A1(\u_multiplier/pp2_8 [1]),
    .A2(\u_multiplier/pp2_8 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_8_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_8_1/_20_  (.A(\u_multiplier/pp2_8 [1]),
    .B(\u_multiplier/pp2_8 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_8_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_8_1/_21_  (.A1(\u_multiplier/pp2_8 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_8_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_8_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_8_1/_22_  (.A(\u_multiplier/pp2_8 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_8_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_8_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_8_1/_23_  (.A1(\u_multiplier/pp2_8 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_8_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_8_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_8_1/_24_  (.A(\u_multiplier/pp2_8 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_8_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_8_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_8_1/_25_  (.A(\u_multiplier/STAGE3/pp3_7_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_8_1/_16_ ),
    .ZN(\u_multiplier/pp3_8 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_8_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_8_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_8_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_8_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_8_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_8_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_8_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_8_1/_17_ ),
    .ZN(\u_multiplier/pp3_9 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_8_2/_18_  (.A(\u_multiplier/STAGE3/pp3_7_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_8_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_8_2/_19_  (.A1(\u_multiplier/pp2_8 [5]),
    .A2(\u_multiplier/pp2_8 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_8_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_8_2/_20_  (.A(\u_multiplier/pp2_8 [5]),
    .B(\u_multiplier/pp2_8 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_8_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_8_2/_21_  (.A1(\u_multiplier/pp2_8 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_8_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_8_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_8_2/_22_  (.A(\u_multiplier/pp2_8 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_8_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_8_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_8_2/_23_  (.A1(\u_multiplier/pp2_8 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_8_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_8_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_8_2/_24_  (.A(\u_multiplier/pp2_8 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_8_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_8_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_8_2/_25_  (.A(\u_multiplier/STAGE3/pp3_7_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_8_2/_16_ ),
    .ZN(\u_multiplier/pp3_8 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_8_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_8_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_8_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_8_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_8_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_8_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_8_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_8_2/_17_ ),
    .ZN(\u_multiplier/pp3_9 [2]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_9_1/_18_  (.A(\u_multiplier/STAGE3/pp3_8_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_9_1/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_9_1/_19_  (.A1(\u_multiplier/pp2_9 [1]),
    .A2(\u_multiplier/pp2_9 [0]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_9_1/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_9_1/_20_  (.A(\u_multiplier/pp2_9 [1]),
    .B(\u_multiplier/pp2_9 [0]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_9_1/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_9_1/_21_  (.A1(\u_multiplier/pp2_9 [2]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_9_1/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_9_1/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_9_1/_22_  (.A(\u_multiplier/pp2_9 [2]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_9_1/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_9_1/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_9_1/_23_  (.A1(\u_multiplier/pp2_9 [3]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_9_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_9_1/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_9_1/_24_  (.A(\u_multiplier/pp2_9 [3]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_9_1/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_9_1/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_9_1/_25_  (.A(\u_multiplier/STAGE3/pp3_8_e42_1_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_9_1/_16_ ),
    .ZN(\u_multiplier/pp3_9 [1]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_9_1/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_9_1/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_9_1/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_9_e42_1_cout ));
 OAI21_X1 \u_multiplier/STAGE3/E_4_2_pp3_9_1/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_9_1/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_9_1/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_9_1/_17_ ),
    .ZN(\u_multiplier/pp3_10 [3]));
 INV_X1 \u_multiplier/STAGE3/E_4_2_pp3_9_2/_18_  (.A(\u_multiplier/STAGE3/pp3_8_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_9_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_9_2/_19_  (.A1(\u_multiplier/pp2_9 [5]),
    .A2(\u_multiplier/pp2_9 [4]),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_9_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_9_2/_20_  (.A(\u_multiplier/pp2_9 [5]),
    .B(\u_multiplier/pp2_9 [4]),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_9_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_9_2/_21_  (.A1(\u_multiplier/pp2_9 [6]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_9_2/_12_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_9_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_9_2/_22_  (.A(\u_multiplier/pp2_9 [6]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_9_2/_12_ ),
    .Z(\u_multiplier/STAGE3/E_4_2_pp3_9_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_9_2/_23_  (.A1(\u_multiplier/pp2_9 [7]),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_9_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_9_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_9_2/_24_  (.A(\u_multiplier/pp2_9 [7]),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_9_2/_14_ ),
    .ZN(\u_multiplier/STAGE3/E_4_2_pp3_9_2/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE3/E_4_2_pp3_9_2/_25_  (.A(\u_multiplier/STAGE3/pp3_8_e42_2_cout ),
    .B(\u_multiplier/STAGE3/E_4_2_pp3_9_2/_16_ ),
    .ZN(\u_multiplier/pp3_9 [0]));
 NAND2_X1 \u_multiplier/STAGE3/E_4_2_pp3_9_2/_26_  (.A1(\u_multiplier/STAGE3/E_4_2_pp3_9_2/_11_ ),
    .A2(\u_multiplier/STAGE3/E_4_2_pp3_9_2/_13_ ),
    .ZN(\u_multiplier/STAGE3/pp3_9_e42_2_cout ));
 OAI21_X2 \u_multiplier/STAGE3/E_4_2_pp3_9_2/_27_  (.A(\u_multiplier/STAGE3/E_4_2_pp3_9_2/_15_ ),
    .B1(\u_multiplier/STAGE3/E_4_2_pp3_9_2/_16_ ),
    .B2(\u_multiplier/STAGE3/E_4_2_pp3_9_2/_17_ ),
    .ZN(\u_multiplier/pp3_10 [2]));
 INV_X1 \u_multiplier/STAGE3/Full_adder_pp3_57_1/_12_  (.A(\u_multiplier/STAGE3/pp3_56_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/Full_adder_pp3_57_1/_08_ ));
 NAND3_X2 \u_multiplier/STAGE3/Full_adder_pp3_57_1/_13_  (.A1(\u_multiplier/pp2_57 [5]),
    .A2(\u_multiplier/pp2_57 [4]),
    .A3(\u_multiplier/STAGE3/pp3_56_e42_2_cout ),
    .ZN(\u_multiplier/STAGE3/Full_adder_pp3_57_1/_09_ ));
 NOR2_X2 \u_multiplier/STAGE3/Full_adder_pp3_57_1/_14_  (.A1(\u_multiplier/pp2_57 [5]),
    .A2(\u_multiplier/pp2_57 [4]),
    .ZN(\u_multiplier/STAGE3/Full_adder_pp3_57_1/_10_ ));
 AOI21_X1 \u_multiplier/STAGE3/Full_adder_pp3_57_1/_15_  (.A(\u_multiplier/STAGE3/pp3_56_e42_2_cout ),
    .B1(\u_multiplier/pp2_57 [4]),
    .B2(\u_multiplier/pp2_57 [5]),
    .ZN(\u_multiplier/STAGE3/Full_adder_pp3_57_1/_11_ ));
 NOR2_X2 \u_multiplier/STAGE3/Full_adder_pp3_57_1/_16_  (.A1(\u_multiplier/STAGE3/Full_adder_pp3_57_1/_10_ ),
    .A2(\u_multiplier/STAGE3/Full_adder_pp3_57_1/_11_ ),
    .ZN(\u_multiplier/pp3_58 [2]));
 AOI22_X4 \u_multiplier/STAGE3/Full_adder_pp3_57_1/_17_  (.A1(\u_multiplier/STAGE3/Full_adder_pp3_57_1/_08_ ),
    .A2(\u_multiplier/STAGE3/Full_adder_pp3_57_1/_10_ ),
    .B1(\u_multiplier/pp3_58 [2]),
    .B2(\u_multiplier/STAGE3/Full_adder_pp3_57_1/_09_ ),
    .ZN(\u_multiplier/pp3_57 [0]));
 INV_X1 \u_multiplier/STAGE3/Full_adder_pp3_59_1/_12_  (.A(\u_multiplier/STAGE3/pp3_58_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/Full_adder_pp3_59_1/_08_ ));
 NAND3_X2 \u_multiplier/STAGE3/Full_adder_pp3_59_1/_13_  (.A1(\u_multiplier/pp2_59 [1]),
    .A2(\u_multiplier/pp2_59 [0]),
    .A3(\u_multiplier/STAGE3/pp3_58_e42_1_cout ),
    .ZN(\u_multiplier/STAGE3/Full_adder_pp3_59_1/_09_ ));
 NOR2_X2 \u_multiplier/STAGE3/Full_adder_pp3_59_1/_14_  (.A1(\u_multiplier/pp2_59 [1]),
    .A2(\u_multiplier/pp2_59 [0]),
    .ZN(\u_multiplier/STAGE3/Full_adder_pp3_59_1/_10_ ));
 AOI21_X1 \u_multiplier/STAGE3/Full_adder_pp3_59_1/_15_  (.A(\u_multiplier/STAGE3/pp3_58_e42_1_cout ),
    .B1(\u_multiplier/pp2_59 [0]),
    .B2(\u_multiplier/pp2_59 [1]),
    .ZN(\u_multiplier/STAGE3/Full_adder_pp3_59_1/_11_ ));
 NOR2_X2 \u_multiplier/STAGE3/Full_adder_pp3_59_1/_16_  (.A1(\u_multiplier/STAGE3/Full_adder_pp3_59_1/_10_ ),
    .A2(\u_multiplier/STAGE3/Full_adder_pp3_59_1/_11_ ),
    .ZN(\u_multiplier/pp3_60 [0]));
 AOI22_X4 \u_multiplier/STAGE3/Full_adder_pp3_59_1/_17_  (.A1(\u_multiplier/STAGE3/Full_adder_pp3_59_1/_08_ ),
    .A2(\u_multiplier/STAGE3/Full_adder_pp3_59_1/_10_ ),
    .B1(\u_multiplier/pp3_60 [0]),
    .B2(\u_multiplier/STAGE3/Full_adder_pp3_59_1/_09_ ),
    .ZN(\u_multiplier/pp3_59 [0]));
 AND2_X1 \u_multiplier/STAGE3/Half_adder_pp3_4_1/_4_  (.A1(\u_multiplier/pp2_4 [1]),
    .A2(\u_multiplier/pp2_4 [0]),
    .ZN(\u_multiplier/pp3_5 [1]));
 XOR2_X2 \u_multiplier/STAGE3/Half_adder_pp3_4_1/_5_  (.A(\u_multiplier/pp2_4 [1]),
    .B(\u_multiplier/pp2_4 [0]),
    .Z(\u_multiplier/pp3_4 [0]));
 AND2_X1 \u_multiplier/STAGE3/Half_adder_pp3_6_1/_4_  (.A1(\u_multiplier/pp2_6 [5]),
    .A2(\u_multiplier/pp2_6 [4]),
    .ZN(\u_multiplier/pp3_7 [2]));
 XOR2_X2 \u_multiplier/STAGE3/Half_adder_pp3_6_1/_5_  (.A(\u_multiplier/pp2_6 [5]),
    .B(\u_multiplier/pp2_6 [4]),
    .Z(\u_multiplier/pp3_6 [0]));
 LOGIC0_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_40__147  (.Z(net147));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_10/_18_  (.A(\u_multiplier/STAGE4/pp4_9_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_10/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_10/_19_  (.A1(\u_multiplier/pp3_10 [1]),
    .A2(\u_multiplier/pp3_10 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_10/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_10/_20_  (.A(\u_multiplier/pp3_10 [1]),
    .B(\u_multiplier/pp3_10 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_10/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_10/_21_  (.A1(\u_multiplier/pp3_10 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_10/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_10/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_10/_22_  (.A(\u_multiplier/pp3_10 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_10/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_10/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_10/_23_  (.A1(\u_multiplier/pp3_10 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_10/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_10/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_10/_24_  (.A(\u_multiplier/pp3_10 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_10/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_10/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE4/E_4_2_pp4_10/_25_  (.A(\u_multiplier/STAGE4/pp4_9_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_10/_16_ ),
    .ZN(\u_multiplier/A [10]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_10/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_10/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_10/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_10_cout ));
 OAI21_X2 \u_multiplier/STAGE4/E_4_2_pp4_10/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_10/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_10/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_10/_17_ ),
    .ZN(\u_multiplier/B [11]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_11/_18_  (.A(\u_multiplier/STAGE4/pp4_10_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_11/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_11/_19_  (.A1(\u_multiplier/pp3_11 [1]),
    .A2(\u_multiplier/pp3_11 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_11/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_11/_20_  (.A(\u_multiplier/pp3_11 [1]),
    .B(\u_multiplier/pp3_11 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_11/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_11/_21_  (.A1(\u_multiplier/pp3_11 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_11/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_11/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_11/_22_  (.A(\u_multiplier/pp3_11 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_11/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_11/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_11/_23_  (.A1(\u_multiplier/pp3_11 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_11/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_11/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_11/_24_  (.A(\u_multiplier/pp3_11 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_11/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_11/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_11/_25_  (.A(\u_multiplier/STAGE4/pp4_10_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_11/_16_ ),
    .ZN(\u_multiplier/A [11]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_11/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_11/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_11/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_11_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_11/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_11/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_11/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_11/_17_ ),
    .ZN(\u_multiplier/B [12]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_12/_18_  (.A(\u_multiplier/STAGE4/pp4_11_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_12/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_12/_19_  (.A1(\u_multiplier/pp3_12 [1]),
    .A2(\u_multiplier/pp3_12 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_12/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_12/_20_  (.A(\u_multiplier/pp3_12 [1]),
    .B(\u_multiplier/pp3_12 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_12/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_12/_21_  (.A1(\u_multiplier/pp3_12 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_12/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_12/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_12/_22_  (.A(\u_multiplier/pp3_12 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_12/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_12/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_12/_23_  (.A1(\u_multiplier/pp3_12 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_12/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_12/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE4/E_4_2_pp4_12/_24_  (.A(\u_multiplier/pp3_12 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_12/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_12/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE4/E_4_2_pp4_12/_25_  (.A(\u_multiplier/STAGE4/pp4_11_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_12/_16_ ),
    .ZN(\u_multiplier/A [12]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_12/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_12/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_12/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_12_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_12/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_12/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_12/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_12/_17_ ),
    .ZN(\u_multiplier/B [13]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_13/_18_  (.A(\u_multiplier/STAGE4/pp4_12_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_13/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_13/_19_  (.A1(\u_multiplier/pp3_13 [1]),
    .A2(\u_multiplier/pp3_13 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_13/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_13/_20_  (.A(\u_multiplier/pp3_13 [1]),
    .B(\u_multiplier/pp3_13 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_13/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_13/_21_  (.A1(\u_multiplier/pp3_13 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_13/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_13/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_13/_22_  (.A(\u_multiplier/pp3_13 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_13/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_13/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_13/_23_  (.A1(\u_multiplier/pp3_13 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_13/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_13/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_13/_24_  (.A(\u_multiplier/pp3_13 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_13/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_13/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_13/_25_  (.A(\u_multiplier/STAGE4/pp4_12_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_13/_16_ ),
    .ZN(\u_multiplier/A [13]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_13/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_13/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_13/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_13_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_13/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_13/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_13/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_13/_17_ ),
    .ZN(\u_multiplier/B [14]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_14/_18_  (.A(\u_multiplier/STAGE4/pp4_13_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_14/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_14/_19_  (.A1(\u_multiplier/pp3_14 [1]),
    .A2(\u_multiplier/pp3_14 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_14/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_14/_20_  (.A(\u_multiplier/pp3_14 [1]),
    .B(\u_multiplier/pp3_14 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_14/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_14/_21_  (.A1(\u_multiplier/pp3_14 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_14/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_14/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_14/_22_  (.A(\u_multiplier/pp3_14 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_14/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_14/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_14/_23_  (.A1(\u_multiplier/pp3_14 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_14/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_14/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_14/_24_  (.A(\u_multiplier/pp3_14 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_14/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_14/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE4/E_4_2_pp4_14/_25_  (.A(\u_multiplier/STAGE4/pp4_13_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_14/_16_ ),
    .ZN(\u_multiplier/A [14]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_14/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_14/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_14/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_14_cout ));
 OAI21_X2 \u_multiplier/STAGE4/E_4_2_pp4_14/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_14/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_14/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_14/_17_ ),
    .ZN(\u_multiplier/B [15]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_15/_18_  (.A(\u_multiplier/STAGE4/pp4_14_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_15/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_15/_19_  (.A1(\u_multiplier/pp3_15 [1]),
    .A2(\u_multiplier/pp3_15 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_15/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_15/_20_  (.A(\u_multiplier/pp3_15 [1]),
    .B(\u_multiplier/pp3_15 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_15/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_15/_21_  (.A1(\u_multiplier/pp3_15 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_15/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_15/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_15/_22_  (.A(\u_multiplier/pp3_15 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_15/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_15/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_15/_23_  (.A1(\u_multiplier/pp3_15 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_15/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_15/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_15/_24_  (.A(\u_multiplier/pp3_15 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_15/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_15/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_15/_25_  (.A(\u_multiplier/STAGE4/pp4_14_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_15/_16_ ),
    .ZN(\u_multiplier/A [15]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_15/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_15/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_15/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_15_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_15/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_15/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_15/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_15/_17_ ),
    .ZN(\u_multiplier/B [16]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_16/_18_  (.A(\u_multiplier/STAGE4/pp4_15_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_16/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_16/_19_  (.A1(\u_multiplier/pp3_16 [1]),
    .A2(\u_multiplier/pp3_16 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_16/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_16/_20_  (.A(\u_multiplier/pp3_16 [1]),
    .B(\u_multiplier/pp3_16 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_16/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_16/_21_  (.A1(\u_multiplier/pp3_16 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_16/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_16/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_16/_22_  (.A(\u_multiplier/pp3_16 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_16/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_16/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_16/_23_  (.A1(\u_multiplier/pp3_16 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_16/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_16/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_16/_24_  (.A(\u_multiplier/pp3_16 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_16/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_16/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE4/E_4_2_pp4_16/_25_  (.A(\u_multiplier/STAGE4/pp4_15_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_16/_16_ ),
    .ZN(\u_multiplier/A [16]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_16/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_16/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_16/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_16_cout ));
 OAI21_X2 \u_multiplier/STAGE4/E_4_2_pp4_16/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_16/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_16/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_16/_17_ ),
    .ZN(\u_multiplier/B [17]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_17/_18_  (.A(\u_multiplier/STAGE4/pp4_16_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_17/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_17/_19_  (.A1(\u_multiplier/pp3_17 [1]),
    .A2(\u_multiplier/pp3_17 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_17/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_17/_20_  (.A(\u_multiplier/pp3_17 [1]),
    .B(\u_multiplier/pp3_17 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_17/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_17/_21_  (.A1(\u_multiplier/pp3_17 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_17/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_17/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_17/_22_  (.A(\u_multiplier/pp3_17 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_17/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_17/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_17/_23_  (.A1(\u_multiplier/pp3_17 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_17/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_17/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_17/_24_  (.A(\u_multiplier/pp3_17 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_17/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_17/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_17/_25_  (.A(\u_multiplier/STAGE4/pp4_16_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_17/_16_ ),
    .ZN(\u_multiplier/A [17]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_17/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_17/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_17/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_17_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_17/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_17/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_17/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_17/_17_ ),
    .ZN(\u_multiplier/B [18]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_18/_18_  (.A(\u_multiplier/STAGE4/pp4_17_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_18/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_18/_19_  (.A1(\u_multiplier/pp3_18 [1]),
    .A2(\u_multiplier/pp3_18 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_18/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_18/_20_  (.A(\u_multiplier/pp3_18 [1]),
    .B(\u_multiplier/pp3_18 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_18/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_18/_21_  (.A1(\u_multiplier/pp3_18 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_18/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_18/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_18/_22_  (.A(\u_multiplier/pp3_18 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_18/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_18/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_18/_23_  (.A1(\u_multiplier/pp3_18 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_18/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_18/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_18/_24_  (.A(\u_multiplier/pp3_18 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_18/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_18/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE4/E_4_2_pp4_18/_25_  (.A(\u_multiplier/STAGE4/pp4_17_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_18/_16_ ),
    .ZN(\u_multiplier/A [18]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_18/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_18/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_18/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_18_cout ));
 OAI21_X2 \u_multiplier/STAGE4/E_4_2_pp4_18/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_18/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_18/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_18/_17_ ),
    .ZN(\u_multiplier/B [19]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_19/_18_  (.A(\u_multiplier/STAGE4/pp4_18_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_19/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_19/_19_  (.A1(\u_multiplier/pp3_19 [1]),
    .A2(\u_multiplier/pp3_19 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_19/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_19/_20_  (.A(\u_multiplier/pp3_19 [1]),
    .B(\u_multiplier/pp3_19 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_19/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_19/_21_  (.A1(\u_multiplier/pp3_19 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_19/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_19/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_19/_22_  (.A(\u_multiplier/pp3_19 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_19/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_19/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_19/_23_  (.A1(\u_multiplier/pp3_19 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_19/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_19/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_19/_24_  (.A(\u_multiplier/pp3_19 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_19/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_19/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_19/_25_  (.A(\u_multiplier/STAGE4/pp4_18_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_19/_16_ ),
    .ZN(\u_multiplier/A [19]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_19/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_19/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_19/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_19_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_19/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_19/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_19/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_19/_17_ ),
    .ZN(\u_multiplier/B [20]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_2/_18_  (.A(\u_multiplier/STAGE4/pp4_1_ha_c ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_2/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_2/_19_  (.A1(\u_multiplier/pp3_2 [1]),
    .A2(\u_multiplier/pp3_2 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_2/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_2/_20_  (.A(\u_multiplier/pp3_2 [1]),
    .B(\u_multiplier/pp3_2 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_2/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_2/_21_  (.A1(\u_multiplier/pp3_2 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_2/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_2/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_2/_22_  (.A(\u_multiplier/pp3_2 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_2/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_2/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_2/_23_  (.A1(net159),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_2/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_2/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_2/_24_  (.A(net160),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_2/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_2/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE4/E_4_2_pp4_2/_25_  (.A(\u_multiplier/STAGE4/pp4_1_ha_c ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_2/_16_ ),
    .ZN(\u_multiplier/A [2]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_2/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_2/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_2/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_2_cout ));
 OAI21_X2 \u_multiplier/STAGE4/E_4_2_pp4_2/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_2/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_2/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_2/_17_ ),
    .ZN(\u_multiplier/B [3]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_20/_18_  (.A(\u_multiplier/STAGE4/pp4_19_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_20/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_20/_19_  (.A1(\u_multiplier/pp3_20 [1]),
    .A2(\u_multiplier/pp3_20 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_20/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_20/_20_  (.A(\u_multiplier/pp3_20 [1]),
    .B(\u_multiplier/pp3_20 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_20/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_20/_21_  (.A1(\u_multiplier/pp3_20 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_20/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_20/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_20/_22_  (.A(\u_multiplier/pp3_20 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_20/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_20/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_20/_23_  (.A1(\u_multiplier/pp3_20 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_20/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_20/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_20/_24_  (.A(\u_multiplier/pp3_20 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_20/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_20/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE4/E_4_2_pp4_20/_25_  (.A(\u_multiplier/STAGE4/pp4_19_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_20/_16_ ),
    .ZN(\u_multiplier/A [20]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_20/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_20/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_20/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_20_cout ));
 OAI21_X2 \u_multiplier/STAGE4/E_4_2_pp4_20/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_20/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_20/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_20/_17_ ),
    .ZN(\u_multiplier/B [21]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_21/_18_  (.A(\u_multiplier/STAGE4/pp4_20_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_21/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_21/_19_  (.A1(\u_multiplier/pp3_21 [1]),
    .A2(\u_multiplier/pp3_21 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_21/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_21/_20_  (.A(\u_multiplier/pp3_21 [1]),
    .B(\u_multiplier/pp3_21 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_21/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_21/_21_  (.A1(\u_multiplier/pp3_21 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_21/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_21/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_21/_22_  (.A(\u_multiplier/pp3_21 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_21/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_21/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_21/_23_  (.A1(\u_multiplier/pp3_21 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_21/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_21/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_21/_24_  (.A(\u_multiplier/pp3_21 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_21/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_21/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_21/_25_  (.A(\u_multiplier/STAGE4/pp4_20_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_21/_16_ ),
    .ZN(\u_multiplier/A [21]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_21/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_21/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_21/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_21_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_21/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_21/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_21/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_21/_17_ ),
    .ZN(\u_multiplier/B [22]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_22/_18_  (.A(\u_multiplier/STAGE4/pp4_21_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_22/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_22/_19_  (.A1(\u_multiplier/pp3_22 [1]),
    .A2(\u_multiplier/pp3_22 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_22/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_22/_20_  (.A(\u_multiplier/pp3_22 [1]),
    .B(\u_multiplier/pp3_22 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_22/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_22/_21_  (.A1(\u_multiplier/pp3_22 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_22/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_22/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_22/_22_  (.A(\u_multiplier/pp3_22 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_22/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_22/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_22/_23_  (.A1(\u_multiplier/pp3_22 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_22/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_22/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_22/_24_  (.A(\u_multiplier/pp3_22 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_22/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_22/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE4/E_4_2_pp4_22/_25_  (.A(\u_multiplier/STAGE4/pp4_21_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_22/_16_ ),
    .ZN(\u_multiplier/A [22]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_22/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_22/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_22/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_22_cout ));
 OAI21_X2 \u_multiplier/STAGE4/E_4_2_pp4_22/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_22/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_22/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_22/_17_ ),
    .ZN(\u_multiplier/B [23]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_23/_18_  (.A(\u_multiplier/STAGE4/pp4_22_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_23/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_23/_19_  (.A1(\u_multiplier/pp3_23 [1]),
    .A2(\u_multiplier/pp3_23 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_23/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_23/_20_  (.A(\u_multiplier/pp3_23 [1]),
    .B(\u_multiplier/pp3_23 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_23/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_23/_21_  (.A1(\u_multiplier/pp3_23 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_23/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_23/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_23/_22_  (.A(\u_multiplier/pp3_23 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_23/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_23/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_23/_23_  (.A1(\u_multiplier/pp3_23 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_23/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_23/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_23/_24_  (.A(\u_multiplier/pp3_23 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_23/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_23/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_23/_25_  (.A(\u_multiplier/STAGE4/pp4_22_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_23/_16_ ),
    .ZN(\u_multiplier/A [23]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_23/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_23/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_23/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_23_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_23/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_23/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_23/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_23/_17_ ),
    .ZN(\u_multiplier/B [24]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_24/_18_  (.A(\u_multiplier/STAGE4/pp4_23_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_24/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_24/_19_  (.A1(\u_multiplier/pp3_24 [1]),
    .A2(\u_multiplier/pp3_24 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_24/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_24/_20_  (.A(\u_multiplier/pp3_24 [1]),
    .B(\u_multiplier/pp3_24 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_24/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_24/_21_  (.A1(\u_multiplier/pp3_24 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_24/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_24/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_24/_22_  (.A(\u_multiplier/pp3_24 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_24/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_24/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_24/_23_  (.A1(\u_multiplier/pp3_24 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_24/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_24/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_24/_24_  (.A(\u_multiplier/pp3_24 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_24/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_24/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_24/_25_  (.A(\u_multiplier/STAGE4/pp4_23_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_24/_16_ ),
    .ZN(\u_multiplier/A [24]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_24/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_24/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_24/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_24_cout ));
 OAI21_X2 \u_multiplier/STAGE4/E_4_2_pp4_24/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_24/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_24/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_24/_17_ ),
    .ZN(\u_multiplier/B [25]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_25/_18_  (.A(\u_multiplier/STAGE4/pp4_24_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_25/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_25/_19_  (.A1(\u_multiplier/pp3_25 [1]),
    .A2(\u_multiplier/pp3_25 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_25/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_25/_20_  (.A(\u_multiplier/pp3_25 [1]),
    .B(\u_multiplier/pp3_25 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_25/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_25/_21_  (.A1(\u_multiplier/pp3_25 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_25/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_25/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_25/_22_  (.A(\u_multiplier/pp3_25 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_25/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_25/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_25/_23_  (.A1(\u_multiplier/pp3_25 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_25/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_25/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_25/_24_  (.A(\u_multiplier/pp3_25 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_25/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_25/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_25/_25_  (.A(\u_multiplier/STAGE4/pp4_24_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_25/_16_ ),
    .ZN(\u_multiplier/A [25]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_25/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_25/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_25/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_25_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_25/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_25/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_25/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_25/_17_ ),
    .ZN(\u_multiplier/B [26]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_26/_18_  (.A(\u_multiplier/STAGE4/pp4_25_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_26/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_26/_19_  (.A1(\u_multiplier/pp3_26 [1]),
    .A2(\u_multiplier/pp3_26 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_26/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_26/_20_  (.A(\u_multiplier/pp3_26 [1]),
    .B(\u_multiplier/pp3_26 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_26/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_26/_21_  (.A1(\u_multiplier/pp3_26 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_26/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_26/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_26/_22_  (.A(\u_multiplier/pp3_26 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_26/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_26/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_26/_23_  (.A1(\u_multiplier/pp3_26 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_26/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_26/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_26/_24_  (.A(\u_multiplier/pp3_26 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_26/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_26/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE4/E_4_2_pp4_26/_25_  (.A(\u_multiplier/STAGE4/pp4_25_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_26/_16_ ),
    .ZN(\u_multiplier/A [26]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_26/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_26/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_26/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_26_cout ));
 OAI21_X2 \u_multiplier/STAGE4/E_4_2_pp4_26/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_26/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_26/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_26/_17_ ),
    .ZN(\u_multiplier/B [27]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_27/_18_  (.A(\u_multiplier/STAGE4/pp4_26_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_27/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_27/_19_  (.A1(\u_multiplier/pp3_27 [1]),
    .A2(\u_multiplier/pp3_27 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_27/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_27/_20_  (.A(\u_multiplier/pp3_27 [1]),
    .B(\u_multiplier/pp3_27 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_27/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_27/_21_  (.A1(\u_multiplier/pp3_27 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_27/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_27/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_27/_22_  (.A(\u_multiplier/pp3_27 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_27/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_27/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_27/_23_  (.A1(\u_multiplier/pp3_27 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_27/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_27/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_27/_24_  (.A(\u_multiplier/pp3_27 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_27/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_27/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_27/_25_  (.A(\u_multiplier/STAGE4/pp4_26_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_27/_16_ ),
    .ZN(\u_multiplier/A [27]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_27/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_27/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_27/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_27_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_27/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_27/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_27/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_27/_17_ ),
    .ZN(\u_multiplier/B [28]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_28/_18_  (.A(\u_multiplier/STAGE4/pp4_27_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_28/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_28/_19_  (.A1(\u_multiplier/pp3_28 [1]),
    .A2(\u_multiplier/pp3_28 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_28/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_28/_20_  (.A(\u_multiplier/pp3_28 [1]),
    .B(\u_multiplier/pp3_28 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_28/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_28/_21_  (.A1(\u_multiplier/pp3_28 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_28/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_28/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_28/_22_  (.A(\u_multiplier/pp3_28 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_28/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_28/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_28/_23_  (.A1(\u_multiplier/pp3_28 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_28/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_28/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_28/_24_  (.A(\u_multiplier/pp3_28 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_28/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_28/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_28/_25_  (.A(\u_multiplier/STAGE4/pp4_27_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_28/_16_ ),
    .ZN(\u_multiplier/A [28]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_28/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_28/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_28/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_28_cout ));
 OAI21_X2 \u_multiplier/STAGE4/E_4_2_pp4_28/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_28/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_28/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_28/_17_ ),
    .ZN(\u_multiplier/B [29]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_29/_18_  (.A(\u_multiplier/STAGE4/pp4_28_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_29/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_29/_19_  (.A1(\u_multiplier/pp3_29 [1]),
    .A2(\u_multiplier/pp3_29 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_29/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_29/_20_  (.A(\u_multiplier/pp3_29 [1]),
    .B(\u_multiplier/pp3_29 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_29/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_29/_21_  (.A1(\u_multiplier/pp3_29 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_29/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_29/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_29/_22_  (.A(\u_multiplier/pp3_29 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_29/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_29/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_29/_23_  (.A1(\u_multiplier/pp3_29 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_29/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_29/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_29/_24_  (.A(\u_multiplier/pp3_29 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_29/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_29/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_29/_25_  (.A(\u_multiplier/STAGE4/pp4_28_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_29/_16_ ),
    .ZN(\u_multiplier/A [29]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_29/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_29/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_29/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_29_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_29/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_29/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_29/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_29/_17_ ),
    .ZN(\u_multiplier/B [30]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_3/_18_  (.A(\u_multiplier/STAGE4/pp4_2_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_3/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_3/_19_  (.A1(\u_multiplier/pp3_3 [1]),
    .A2(\u_multiplier/pp3_3 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_3/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_3/_20_  (.A(\u_multiplier/pp3_3 [1]),
    .B(\u_multiplier/pp3_3 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_3/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_3/_21_  (.A1(\u_multiplier/pp3_3 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_3/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_3/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_3/_22_  (.A(\u_multiplier/pp3_3 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_3/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_3/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_3/_23_  (.A1(\u_multiplier/pp3_3 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_3/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_3/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_3/_24_  (.A(\u_multiplier/pp3_3 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_3/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_3/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_3/_25_  (.A(\u_multiplier/STAGE4/pp4_2_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_3/_16_ ),
    .ZN(\u_multiplier/A [3]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_3/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_3/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_3/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_3_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_3/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_3/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_3/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_3/_17_ ),
    .ZN(\u_multiplier/B [4]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_30/_18_  (.A(\u_multiplier/STAGE4/pp4_29_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_30/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_30/_19_  (.A1(\u_multiplier/pp3_30 [1]),
    .A2(\u_multiplier/pp3_30 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_30/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_30/_20_  (.A(\u_multiplier/pp3_30 [1]),
    .B(\u_multiplier/pp3_30 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_30/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_30/_21_  (.A1(\u_multiplier/pp3_30 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_30/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_30/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_30/_22_  (.A(\u_multiplier/pp3_30 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_30/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_30/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_30/_23_  (.A1(\u_multiplier/pp3_30 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_30/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_30/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_30/_24_  (.A(\u_multiplier/pp3_30 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_30/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_30/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE4/E_4_2_pp4_30/_25_  (.A(\u_multiplier/STAGE4/pp4_29_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_30/_16_ ),
    .ZN(\u_multiplier/A [30]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_30/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_30/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_30/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_30_cout ));
 OAI21_X2 \u_multiplier/STAGE4/E_4_2_pp4_30/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_30/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_30/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_30/_17_ ),
    .ZN(\u_multiplier/B [31]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_31/_18_  (.A(\u_multiplier/STAGE4/pp4_30_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_31/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_31/_19_  (.A1(\u_multiplier/pp3_31 [1]),
    .A2(\u_multiplier/pp3_31 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_31/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_31/_20_  (.A(\u_multiplier/pp3_31 [1]),
    .B(\u_multiplier/pp3_31 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_31/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_31/_21_  (.A1(\u_multiplier/pp3_31 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_31/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_31/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_31/_22_  (.A(\u_multiplier/pp3_31 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_31/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_31/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_31/_23_  (.A1(\u_multiplier/pp3_31 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_31/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_31/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_31/_24_  (.A(\u_multiplier/pp3_31 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_31/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_31/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_31/_25_  (.A(\u_multiplier/STAGE4/pp4_30_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_31/_16_ ),
    .ZN(\u_multiplier/A [31]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_31/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_31/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_31/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_31_cout ));
 OAI21_X2 \u_multiplier/STAGE4/E_4_2_pp4_31/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_31/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_31/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_31/_17_ ),
    .ZN(\u_multiplier/B [32]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_32/_18_  (.A(\u_multiplier/STAGE4/pp4_31_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_32/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_32/_19_  (.A1(\u_multiplier/pp3_32 [1]),
    .A2(\u_multiplier/pp3_32 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_32/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_32/_20_  (.A(\u_multiplier/pp3_32 [1]),
    .B(\u_multiplier/pp3_32 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_32/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_32/_21_  (.A1(\u_multiplier/pp3_32 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_32/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_32/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_32/_22_  (.A(\u_multiplier/pp3_32 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_32/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_32/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_32/_23_  (.A1(\u_multiplier/pp3_32 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_32/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_32/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_32/_24_  (.A(\u_multiplier/pp3_32 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_32/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_32/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE4/E_4_2_pp4_32/_25_  (.A(\u_multiplier/STAGE4/pp4_31_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_32/_16_ ),
    .ZN(\u_multiplier/A [32]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_32/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_32/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_32/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_32_cout ));
 OAI21_X2 \u_multiplier/STAGE4/E_4_2_pp4_32/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_32/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_32/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_32/_17_ ),
    .ZN(\u_multiplier/B [33]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_33/_18_  (.A(\u_multiplier/STAGE4/pp4_32_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_33/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_33/_19_  (.A1(\u_multiplier/pp3_33 [1]),
    .A2(\u_multiplier/pp3_33 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_33/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_33/_20_  (.A(\u_multiplier/pp3_33 [1]),
    .B(\u_multiplier/pp3_33 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_33/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_33/_21_  (.A1(\u_multiplier/pp3_33 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_33/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_33/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_33/_22_  (.A(\u_multiplier/pp3_33 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_33/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_33/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_33/_23_  (.A1(\u_multiplier/pp3_33 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_33/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_33/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_33/_24_  (.A(\u_multiplier/pp3_33 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_33/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_33/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_33/_25_  (.A(\u_multiplier/STAGE4/pp4_32_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_33/_16_ ),
    .ZN(\u_multiplier/A [33]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_33/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_33/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_33/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_33_cout ));
 OAI21_X2 \u_multiplier/STAGE4/E_4_2_pp4_33/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_33/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_33/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_33/_17_ ),
    .ZN(\u_multiplier/B [34]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_34/_18_  (.A(\u_multiplier/STAGE4/pp4_33_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_34/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_34/_19_  (.A1(\u_multiplier/pp3_34 [1]),
    .A2(\u_multiplier/pp3_34 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_34/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_34/_20_  (.A(\u_multiplier/pp3_34 [1]),
    .B(\u_multiplier/pp3_34 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_34/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_34/_21_  (.A1(\u_multiplier/pp3_34 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_34/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_34/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_34/_22_  (.A(\u_multiplier/pp3_34 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_34/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_34/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_34/_23_  (.A1(\u_multiplier/pp3_34 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_34/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_34/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_34/_24_  (.A(\u_multiplier/pp3_34 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_34/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_34/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE4/E_4_2_pp4_34/_25_  (.A(\u_multiplier/STAGE4/pp4_33_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_34/_16_ ),
    .ZN(\u_multiplier/A [34]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_34/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_34/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_34/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_34_cout ));
 OAI21_X2 \u_multiplier/STAGE4/E_4_2_pp4_34/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_34/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_34/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_34/_17_ ),
    .ZN(\u_multiplier/B [35]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_35/_18_  (.A(\u_multiplier/STAGE4/pp4_34_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_35/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_35/_19_  (.A1(\u_multiplier/pp3_35 [1]),
    .A2(\u_multiplier/pp3_35 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_35/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_35/_20_  (.A(\u_multiplier/pp3_35 [1]),
    .B(\u_multiplier/pp3_35 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_35/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_35/_21_  (.A1(\u_multiplier/pp3_35 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_35/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_35/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_35/_22_  (.A(\u_multiplier/pp3_35 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_35/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_35/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_35/_23_  (.A1(\u_multiplier/pp3_35 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_35/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_35/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_35/_24_  (.A(\u_multiplier/pp3_35 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_35/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_35/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_35/_25_  (.A(\u_multiplier/STAGE4/pp4_34_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_35/_16_ ),
    .ZN(\u_multiplier/A [35]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_35/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_35/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_35/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_35_cout ));
 OAI21_X2 \u_multiplier/STAGE4/E_4_2_pp4_35/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_35/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_35/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_35/_17_ ),
    .ZN(\u_multiplier/B [36]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_36/_18_  (.A(\u_multiplier/STAGE4/pp4_35_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_36/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_36/_19_  (.A1(\u_multiplier/pp3_36 [1]),
    .A2(\u_multiplier/pp3_36 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_36/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_36/_20_  (.A(\u_multiplier/pp3_36 [1]),
    .B(\u_multiplier/pp3_36 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_36/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_36/_21_  (.A1(\u_multiplier/pp3_36 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_36/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_36/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_36/_22_  (.A(\u_multiplier/pp3_36 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_36/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_36/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_36/_23_  (.A1(\u_multiplier/pp3_36 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_36/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_36/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_36/_24_  (.A(\u_multiplier/pp3_36 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_36/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_36/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_36/_25_  (.A(\u_multiplier/STAGE4/pp4_35_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_36/_16_ ),
    .ZN(\u_multiplier/A [36]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_36/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_36/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_36/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_36_cout ));
 OAI21_X2 \u_multiplier/STAGE4/E_4_2_pp4_36/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_36/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_36/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_36/_17_ ),
    .ZN(\u_multiplier/B [37]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_37/_18_  (.A(\u_multiplier/STAGE4/pp4_36_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_37/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_37/_19_  (.A1(\u_multiplier/pp3_37 [1]),
    .A2(\u_multiplier/pp3_37 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_37/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_37/_20_  (.A(\u_multiplier/pp3_37 [1]),
    .B(\u_multiplier/pp3_37 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_37/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_37/_21_  (.A1(\u_multiplier/pp3_37 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_37/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_37/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_37/_22_  (.A(\u_multiplier/pp3_37 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_37/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_37/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_37/_23_  (.A1(\u_multiplier/pp3_37 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_37/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_37/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_37/_24_  (.A(\u_multiplier/pp3_37 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_37/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_37/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_37/_25_  (.A(\u_multiplier/STAGE4/pp4_36_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_37/_16_ ),
    .ZN(\u_multiplier/A [37]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_37/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_37/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_37/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_37_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_37/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_37/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_37/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_37/_17_ ),
    .ZN(\u_multiplier/B [38]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_38/_18_  (.A(\u_multiplier/STAGE4/pp4_37_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_38/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_38/_19_  (.A1(\u_multiplier/pp3_38 [1]),
    .A2(\u_multiplier/pp3_38 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_38/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_38/_20_  (.A(\u_multiplier/pp3_38 [1]),
    .B(\u_multiplier/pp3_38 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_38/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_38/_21_  (.A1(\u_multiplier/pp3_38 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_38/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_38/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_38/_22_  (.A(\u_multiplier/pp3_38 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_38/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_38/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_38/_23_  (.A1(\u_multiplier/pp3_38 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_38/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_38/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE4/E_4_2_pp4_38/_24_  (.A(\u_multiplier/pp3_38 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_38/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_38/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE4/E_4_2_pp4_38/_25_  (.A(\u_multiplier/STAGE4/pp4_37_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_38/_16_ ),
    .ZN(\u_multiplier/A [38]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_38/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_38/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_38/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_38_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_38/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_38/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_38/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_38/_17_ ),
    .ZN(\u_multiplier/B [39]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_39/_18_  (.A(\u_multiplier/STAGE4/pp4_38_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_39/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_39/_19_  (.A1(\u_multiplier/pp3_39 [1]),
    .A2(\u_multiplier/pp3_39 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_39/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_39/_20_  (.A(\u_multiplier/pp3_39 [1]),
    .B(\u_multiplier/pp3_39 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_39/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_39/_21_  (.A1(\u_multiplier/pp3_39 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_39/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_39/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_39/_22_  (.A(\u_multiplier/pp3_39 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_39/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_39/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_39/_23_  (.A1(\u_multiplier/pp3_39 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_39/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_39/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_39/_24_  (.A(\u_multiplier/pp3_39 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_39/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_39/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_39/_25_  (.A(\u_multiplier/STAGE4/pp4_38_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_39/_16_ ),
    .ZN(\u_multiplier/A [39]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_39/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_39/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_39/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_39_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_39/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_39/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_39/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_39/_17_ ),
    .ZN(\u_multiplier/B [40]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_4/_18_  (.A(\u_multiplier/STAGE4/pp4_3_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_4/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_4/_19_  (.A1(\u_multiplier/pp3_4 [1]),
    .A2(\u_multiplier/pp3_4 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_4/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_4/_20_  (.A(\u_multiplier/pp3_4 [1]),
    .B(\u_multiplier/pp3_4 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_4/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_4/_21_  (.A1(\u_multiplier/pp3_4 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_4/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_4/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_4/_22_  (.A(\u_multiplier/pp3_4 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_4/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_4/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_4/_23_  (.A1(\u_multiplier/pp3_4 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_4/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_4/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_4/_24_  (.A(\u_multiplier/pp3_4 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_4/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_4/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE4/E_4_2_pp4_4/_25_  (.A(\u_multiplier/STAGE4/pp4_3_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_4/_16_ ),
    .ZN(\u_multiplier/A [4]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_4/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_4/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_4/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_4_cout ));
 OAI21_X2 \u_multiplier/STAGE4/E_4_2_pp4_4/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_4/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_4/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_4/_17_ ),
    .ZN(\u_multiplier/B [5]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_40/_18_  (.A(\u_multiplier/STAGE4/pp4_39_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_40/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_40/_19_  (.A1(\u_multiplier/pp3_40 [1]),
    .A2(\u_multiplier/pp3_40 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_40/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_40/_20_  (.A(\u_multiplier/pp3_40 [1]),
    .B(\u_multiplier/pp3_40 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_40/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_40/_21_  (.A1(\u_multiplier/pp3_40 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_40/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_40/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_40/_22_  (.A(\u_multiplier/pp3_40 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_40/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_40/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_40/_23_  (.A1(\u_multiplier/pp3_40 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_40/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_40/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_40/_24_  (.A(\u_multiplier/pp3_40 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_40/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_40/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE4/E_4_2_pp4_40/_25_  (.A(\u_multiplier/STAGE4/pp4_39_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_40/_16_ ),
    .ZN(\u_multiplier/A [40]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_40/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_40/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_40/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_40_cout ));
 OAI21_X2 \u_multiplier/STAGE4/E_4_2_pp4_40/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_40/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_40/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_40/_17_ ),
    .ZN(\u_multiplier/B [41]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_41/_18_  (.A(\u_multiplier/STAGE4/pp4_40_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_41/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_41/_19_  (.A1(\u_multiplier/pp3_41 [1]),
    .A2(\u_multiplier/pp3_41 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_41/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_41/_20_  (.A(\u_multiplier/pp3_41 [1]),
    .B(\u_multiplier/pp3_41 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_41/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_41/_21_  (.A1(\u_multiplier/pp3_41 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_41/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_41/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_41/_22_  (.A(\u_multiplier/pp3_41 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_41/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_41/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_41/_23_  (.A1(\u_multiplier/pp3_41 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_41/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_41/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_41/_24_  (.A(\u_multiplier/pp3_41 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_41/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_41/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_41/_25_  (.A(\u_multiplier/STAGE4/pp4_40_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_41/_16_ ),
    .ZN(\u_multiplier/A [41]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_41/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_41/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_41/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_41_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_41/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_41/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_41/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_41/_17_ ),
    .ZN(\u_multiplier/B [42]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_42/_18_  (.A(\u_multiplier/STAGE4/pp4_41_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_42/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_42/_19_  (.A1(\u_multiplier/pp3_42 [1]),
    .A2(\u_multiplier/pp3_42 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_42/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_42/_20_  (.A(\u_multiplier/pp3_42 [1]),
    .B(\u_multiplier/pp3_42 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_42/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_42/_21_  (.A1(\u_multiplier/pp3_42 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_42/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_42/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_42/_22_  (.A(\u_multiplier/pp3_42 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_42/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_42/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_42/_23_  (.A1(\u_multiplier/pp3_42 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_42/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_42/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_42/_24_  (.A(\u_multiplier/pp3_42 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_42/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_42/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_42/_25_  (.A(\u_multiplier/STAGE4/pp4_41_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_42/_16_ ),
    .ZN(\u_multiplier/A [42]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_42/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_42/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_42/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_42_cout ));
 OAI21_X2 \u_multiplier/STAGE4/E_4_2_pp4_42/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_42/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_42/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_42/_17_ ),
    .ZN(\u_multiplier/B [43]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_43/_18_  (.A(\u_multiplier/STAGE4/pp4_42_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_43/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_43/_19_  (.A1(\u_multiplier/pp3_43 [1]),
    .A2(\u_multiplier/pp3_43 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_43/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_43/_20_  (.A(\u_multiplier/pp3_43 [1]),
    .B(\u_multiplier/pp3_43 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_43/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_43/_21_  (.A1(\u_multiplier/pp3_43 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_43/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_43/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_43/_22_  (.A(\u_multiplier/pp3_43 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_43/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_43/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_43/_23_  (.A1(\u_multiplier/pp3_43 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_43/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_43/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_43/_24_  (.A(\u_multiplier/pp3_43 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_43/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_43/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_43/_25_  (.A(\u_multiplier/STAGE4/pp4_42_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_43/_16_ ),
    .ZN(\u_multiplier/A [43]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_43/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_43/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_43/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_43_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_43/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_43/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_43/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_43/_17_ ),
    .ZN(\u_multiplier/B [44]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_44/_18_  (.A(\u_multiplier/STAGE4/pp4_43_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_44/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_44/_19_  (.A1(\u_multiplier/pp3_44 [1]),
    .A2(\u_multiplier/pp3_44 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_44/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_44/_20_  (.A(\u_multiplier/pp3_44 [1]),
    .B(\u_multiplier/pp3_44 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_44/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_44/_21_  (.A1(\u_multiplier/pp3_44 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_44/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_44/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_44/_22_  (.A(\u_multiplier/pp3_44 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_44/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_44/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_44/_23_  (.A1(\u_multiplier/pp3_44 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_44/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_44/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_44/_24_  (.A(\u_multiplier/pp3_44 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_44/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_44/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_44/_25_  (.A(\u_multiplier/STAGE4/pp4_43_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_44/_16_ ),
    .ZN(\u_multiplier/A [44]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_44/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_44/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_44/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_44_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_44/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_44/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_44/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_44/_17_ ),
    .ZN(\u_multiplier/B [45]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_45/_18_  (.A(\u_multiplier/STAGE4/pp4_44_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_45/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_45/_19_  (.A1(\u_multiplier/pp3_45 [1]),
    .A2(\u_multiplier/pp3_45 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_45/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_45/_20_  (.A(\u_multiplier/pp3_45 [1]),
    .B(\u_multiplier/pp3_45 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_45/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_45/_21_  (.A1(\u_multiplier/pp3_45 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_45/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_45/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_45/_22_  (.A(\u_multiplier/pp3_45 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_45/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_45/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_45/_23_  (.A1(\u_multiplier/pp3_45 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_45/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_45/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_45/_24_  (.A(\u_multiplier/pp3_45 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_45/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_45/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_45/_25_  (.A(\u_multiplier/STAGE4/pp4_44_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_45/_16_ ),
    .ZN(\u_multiplier/A [45]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_45/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_45/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_45/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_45_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_45/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_45/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_45/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_45/_17_ ),
    .ZN(\u_multiplier/B [46]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_46/_18_  (.A(\u_multiplier/STAGE4/pp4_45_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_46/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_46/_19_  (.A1(\u_multiplier/pp3_46 [1]),
    .A2(\u_multiplier/pp3_46 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_46/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_46/_20_  (.A(\u_multiplier/pp3_46 [1]),
    .B(\u_multiplier/pp3_46 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_46/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_46/_21_  (.A1(\u_multiplier/pp3_46 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_46/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_46/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_46/_22_  (.A(\u_multiplier/pp3_46 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_46/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_46/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_46/_23_  (.A1(\u_multiplier/pp3_46 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_46/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_46/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_46/_24_  (.A(\u_multiplier/pp3_46 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_46/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_46/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE4/E_4_2_pp4_46/_25_  (.A(\u_multiplier/STAGE4/pp4_45_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_46/_16_ ),
    .ZN(\u_multiplier/A [46]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_46/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_46/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_46/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_46_cout ));
 OAI21_X2 \u_multiplier/STAGE4/E_4_2_pp4_46/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_46/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_46/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_46/_17_ ),
    .ZN(\u_multiplier/B [47]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_47/_18_  (.A(\u_multiplier/STAGE4/pp4_46_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_47/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_47/_19_  (.A1(\u_multiplier/pp3_47 [1]),
    .A2(\u_multiplier/pp3_47 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_47/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_47/_20_  (.A(\u_multiplier/pp3_47 [1]),
    .B(\u_multiplier/pp3_47 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_47/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_47/_21_  (.A1(\u_multiplier/pp3_47 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_47/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_47/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_47/_22_  (.A(\u_multiplier/pp3_47 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_47/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_47/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_47/_23_  (.A1(\u_multiplier/pp3_47 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_47/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_47/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_47/_24_  (.A(\u_multiplier/pp3_47 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_47/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_47/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_47/_25_  (.A(\u_multiplier/STAGE4/pp4_46_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_47/_16_ ),
    .ZN(\u_multiplier/A [47]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_47/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_47/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_47/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_47_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_47/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_47/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_47/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_47/_17_ ),
    .ZN(\u_multiplier/B [48]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_48/_18_  (.A(\u_multiplier/STAGE4/pp4_47_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_48/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_48/_19_  (.A1(\u_multiplier/pp3_48 [1]),
    .A2(\u_multiplier/pp3_48 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_48/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_48/_20_  (.A(\u_multiplier/pp3_48 [1]),
    .B(\u_multiplier/pp3_48 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_48/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_48/_21_  (.A1(\u_multiplier/pp3_48 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_48/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_48/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_48/_22_  (.A(\u_multiplier/pp3_48 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_48/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_48/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_48/_23_  (.A1(\u_multiplier/pp3_48 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_48/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_48/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_48/_24_  (.A(\u_multiplier/pp3_48 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_48/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_48/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_48/_25_  (.A(\u_multiplier/STAGE4/pp4_47_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_48/_16_ ),
    .ZN(\u_multiplier/A [48]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_48/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_48/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_48/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_48_cout ));
 OAI21_X2 \u_multiplier/STAGE4/E_4_2_pp4_48/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_48/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_48/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_48/_17_ ),
    .ZN(\u_multiplier/B [49]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_49/_18_  (.A(\u_multiplier/STAGE4/pp4_48_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_49/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_49/_19_  (.A1(\u_multiplier/pp3_49 [1]),
    .A2(\u_multiplier/pp3_49 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_49/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_49/_20_  (.A(\u_multiplier/pp3_49 [1]),
    .B(\u_multiplier/pp3_49 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_49/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_49/_21_  (.A1(\u_multiplier/pp3_49 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_49/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_49/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_49/_22_  (.A(\u_multiplier/pp3_49 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_49/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_49/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_49/_23_  (.A1(\u_multiplier/pp3_49 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_49/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_49/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_49/_24_  (.A(\u_multiplier/pp3_49 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_49/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_49/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_49/_25_  (.A(\u_multiplier/STAGE4/pp4_48_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_49/_16_ ),
    .ZN(\u_multiplier/A [49]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_49/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_49/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_49/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_49_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_49/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_49/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_49/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_49/_17_ ),
    .ZN(\u_multiplier/B [50]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_5/_18_  (.A(\u_multiplier/STAGE4/pp4_4_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_5/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_5/_19_  (.A1(\u_multiplier/pp3_5 [1]),
    .A2(\u_multiplier/pp3_5 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_5/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_5/_20_  (.A(\u_multiplier/pp3_5 [1]),
    .B(\u_multiplier/pp3_5 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_5/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_5/_21_  (.A1(\u_multiplier/pp3_5 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_5/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_5/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_5/_22_  (.A(\u_multiplier/pp3_5 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_5/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_5/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_5/_23_  (.A1(\u_multiplier/pp3_5 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_5/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_5/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_5/_24_  (.A(\u_multiplier/pp3_5 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_5/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_5/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_5/_25_  (.A(\u_multiplier/STAGE4/pp4_4_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_5/_16_ ),
    .ZN(\u_multiplier/A [5]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_5/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_5/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_5/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_5_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_5/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_5/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_5/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_5/_17_ ),
    .ZN(\u_multiplier/B [6]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_50/_18_  (.A(\u_multiplier/STAGE4/pp4_49_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_50/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_50/_19_  (.A1(\u_multiplier/pp3_50 [1]),
    .A2(\u_multiplier/pp3_50 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_50/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_50/_20_  (.A(\u_multiplier/pp3_50 [1]),
    .B(\u_multiplier/pp3_50 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_50/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_50/_21_  (.A1(\u_multiplier/pp3_50 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_50/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_50/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_50/_22_  (.A(\u_multiplier/pp3_50 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_50/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_50/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_50/_23_  (.A1(\u_multiplier/pp3_50 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_50/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_50/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_50/_24_  (.A(\u_multiplier/pp3_50 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_50/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_50/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE4/E_4_2_pp4_50/_25_  (.A(\u_multiplier/STAGE4/pp4_49_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_50/_16_ ),
    .ZN(\u_multiplier/A [50]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_50/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_50/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_50/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_50_cout ));
 OAI21_X2 \u_multiplier/STAGE4/E_4_2_pp4_50/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_50/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_50/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_50/_17_ ),
    .ZN(\u_multiplier/B [51]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_51/_18_  (.A(\u_multiplier/STAGE4/pp4_50_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_51/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_51/_19_  (.A1(\u_multiplier/pp3_51 [1]),
    .A2(\u_multiplier/pp3_51 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_51/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_51/_20_  (.A(\u_multiplier/pp3_51 [1]),
    .B(\u_multiplier/pp3_51 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_51/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_51/_21_  (.A1(\u_multiplier/pp3_51 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_51/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_51/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_51/_22_  (.A(\u_multiplier/pp3_51 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_51/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_51/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_51/_23_  (.A1(\u_multiplier/pp3_51 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_51/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_51/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_51/_24_  (.A(\u_multiplier/pp3_51 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_51/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_51/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_51/_25_  (.A(\u_multiplier/STAGE4/pp4_50_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_51/_16_ ),
    .ZN(\u_multiplier/A [51]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_51/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_51/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_51/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_51_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_51/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_51/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_51/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_51/_17_ ),
    .ZN(\u_multiplier/B [52]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_52/_18_  (.A(\u_multiplier/STAGE4/pp4_51_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_52/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_52/_19_  (.A1(\u_multiplier/pp3_52 [1]),
    .A2(\u_multiplier/pp3_52 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_52/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_52/_20_  (.A(\u_multiplier/pp3_52 [1]),
    .B(\u_multiplier/pp3_52 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_52/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_52/_21_  (.A1(\u_multiplier/pp3_52 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_52/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_52/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_52/_22_  (.A(\u_multiplier/pp3_52 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_52/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_52/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_52/_23_  (.A1(\u_multiplier/pp3_52 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_52/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_52/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_52/_24_  (.A(\u_multiplier/pp3_52 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_52/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_52/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE4/E_4_2_pp4_52/_25_  (.A(\u_multiplier/STAGE4/pp4_51_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_52/_16_ ),
    .ZN(\u_multiplier/A [52]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_52/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_52/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_52/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_52_cout ));
 OAI21_X2 \u_multiplier/STAGE4/E_4_2_pp4_52/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_52/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_52/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_52/_17_ ),
    .ZN(\u_multiplier/B [53]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_53/_18_  (.A(\u_multiplier/STAGE4/pp4_52_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_53/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_53/_19_  (.A1(\u_multiplier/pp3_53 [1]),
    .A2(\u_multiplier/pp3_53 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_53/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_53/_20_  (.A(\u_multiplier/pp3_53 [1]),
    .B(\u_multiplier/pp3_53 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_53/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_53/_21_  (.A1(\u_multiplier/pp3_53 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_53/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_53/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_53/_22_  (.A(\u_multiplier/pp3_53 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_53/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_53/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_53/_23_  (.A1(\u_multiplier/pp3_53 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_53/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_53/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_53/_24_  (.A(\u_multiplier/pp3_53 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_53/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_53/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_53/_25_  (.A(\u_multiplier/STAGE4/pp4_52_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_53/_16_ ),
    .ZN(\u_multiplier/A [53]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_53/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_53/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_53/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_53_cout ));
 OAI21_X2 \u_multiplier/STAGE4/E_4_2_pp4_53/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_53/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_53/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_53/_17_ ),
    .ZN(\u_multiplier/B [54]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_54/_18_  (.A(\u_multiplier/STAGE4/pp4_53_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_54/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_54/_19_  (.A1(\u_multiplier/pp3_54 [1]),
    .A2(\u_multiplier/pp3_54 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_54/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_54/_20_  (.A(\u_multiplier/pp3_54 [1]),
    .B(\u_multiplier/pp3_54 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_54/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_54/_21_  (.A1(\u_multiplier/pp3_54 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_54/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_54/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_54/_22_  (.A(\u_multiplier/pp3_54 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_54/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_54/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_54/_23_  (.A1(\u_multiplier/pp3_54 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_54/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_54/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_54/_24_  (.A(\u_multiplier/pp3_54 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_54/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_54/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_54/_25_  (.A(\u_multiplier/STAGE4/pp4_53_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_54/_16_ ),
    .ZN(\u_multiplier/A [54]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_54/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_54/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_54/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_54_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_54/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_54/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_54/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_54/_17_ ),
    .ZN(\u_multiplier/B [55]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_55/_18_  (.A(\u_multiplier/STAGE4/pp4_54_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_55/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_55/_19_  (.A1(\u_multiplier/pp3_55 [1]),
    .A2(\u_multiplier/pp3_55 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_55/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_55/_20_  (.A(\u_multiplier/pp3_55 [1]),
    .B(\u_multiplier/pp3_55 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_55/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_55/_21_  (.A1(\u_multiplier/pp3_55 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_55/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_55/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_55/_22_  (.A(\u_multiplier/pp3_55 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_55/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_55/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_55/_23_  (.A1(\u_multiplier/pp3_55 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_55/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_55/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_55/_24_  (.A(\u_multiplier/pp3_55 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_55/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_55/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_55/_25_  (.A(\u_multiplier/STAGE4/pp4_54_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_55/_16_ ),
    .ZN(\u_multiplier/A [55]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_55/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_55/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_55/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_55_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_55/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_55/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_55/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_55/_17_ ),
    .ZN(\u_multiplier/B [56]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_56/_18_  (.A(\u_multiplier/STAGE4/pp4_55_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_56/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_56/_19_  (.A1(\u_multiplier/pp3_56 [1]),
    .A2(\u_multiplier/pp3_56 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_56/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_56/_20_  (.A(\u_multiplier/pp3_56 [1]),
    .B(\u_multiplier/pp3_56 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_56/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_56/_21_  (.A1(\u_multiplier/pp3_56 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_56/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_56/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_56/_22_  (.A(\u_multiplier/pp3_56 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_56/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_56/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_56/_23_  (.A1(\u_multiplier/pp3_56 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_56/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_56/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_56/_24_  (.A(\u_multiplier/pp3_56 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_56/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_56/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE4/E_4_2_pp4_56/_25_  (.A(\u_multiplier/STAGE4/pp4_55_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_56/_16_ ),
    .ZN(\u_multiplier/A [56]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_56/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_56/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_56/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_56_cout ));
 OAI21_X2 \u_multiplier/STAGE4/E_4_2_pp4_56/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_56/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_56/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_56/_17_ ),
    .ZN(\u_multiplier/B [57]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_57/_18_  (.A(\u_multiplier/STAGE4/pp4_56_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_57/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_57/_19_  (.A1(\u_multiplier/pp3_57 [1]),
    .A2(\u_multiplier/pp3_57 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_57/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_57/_20_  (.A(\u_multiplier/pp3_57 [1]),
    .B(\u_multiplier/pp3_57 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_57/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_57/_21_  (.A1(\u_multiplier/pp3_57 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_57/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_57/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_57/_22_  (.A(\u_multiplier/pp3_57 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_57/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_57/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_57/_23_  (.A1(\u_multiplier/pp3_57 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_57/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_57/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_57/_24_  (.A(\u_multiplier/pp3_57 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_57/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_57/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_57/_25_  (.A(\u_multiplier/STAGE4/pp4_56_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_57/_16_ ),
    .ZN(\u_multiplier/A [57]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_57/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_57/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_57/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_57_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_57/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_57/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_57/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_57/_17_ ),
    .ZN(\u_multiplier/B [58]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_58/_18_  (.A(\u_multiplier/STAGE4/pp4_57_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_58/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_58/_19_  (.A1(\u_multiplier/pp3_58 [1]),
    .A2(\u_multiplier/pp3_58 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_58/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_58/_20_  (.A(\u_multiplier/pp3_58 [1]),
    .B(\u_multiplier/pp3_58 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_58/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_58/_21_  (.A1(\u_multiplier/pp3_58 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_58/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_58/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_58/_22_  (.A(\u_multiplier/pp3_58 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_58/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_58/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_58/_23_  (.A1(\u_multiplier/pp3_58 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_58/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_58/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE4/E_4_2_pp4_58/_24_  (.A(\u_multiplier/pp3_58 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_58/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_58/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE4/E_4_2_pp4_58/_25_  (.A(\u_multiplier/STAGE4/pp4_57_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_58/_16_ ),
    .ZN(\u_multiplier/A [58]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_58/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_58/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_58/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_58_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_58/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_58/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_58/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_58/_17_ ),
    .ZN(\u_multiplier/B [59]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_59/_18_  (.A(\u_multiplier/STAGE4/pp4_58_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_59/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_59/_19_  (.A1(\u_multiplier/pp3_59 [1]),
    .A2(\u_multiplier/pp3_59 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_59/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_59/_20_  (.A(\u_multiplier/pp3_59 [1]),
    .B(\u_multiplier/pp3_59 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_59/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_59/_21_  (.A1(\u_multiplier/pp3_59 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_59/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_59/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_59/_22_  (.A(\u_multiplier/pp3_59 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_59/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_59/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_59/_23_  (.A1(\u_multiplier/pp3_59 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_59/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_59/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_59/_24_  (.A(\u_multiplier/pp3_59 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_59/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_59/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_59/_25_  (.A(\u_multiplier/STAGE4/pp4_58_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_59/_16_ ),
    .ZN(\u_multiplier/A [59]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_59/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_59/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_59/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_59_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_59/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_59/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_59/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_59/_17_ ),
    .ZN(\u_multiplier/B [60]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_6/_18_  (.A(\u_multiplier/STAGE4/pp4_5_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_6/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_6/_19_  (.A1(\u_multiplier/pp3_6 [1]),
    .A2(\u_multiplier/pp3_6 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_6/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_6/_20_  (.A(\u_multiplier/pp3_6 [1]),
    .B(\u_multiplier/pp3_6 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_6/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_6/_21_  (.A1(\u_multiplier/pp3_6 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_6/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_6/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_6/_22_  (.A(\u_multiplier/pp3_6 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_6/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_6/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_6/_23_  (.A1(\u_multiplier/pp3_6 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_6/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_6/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE4/E_4_2_pp4_6/_24_  (.A(\u_multiplier/pp3_6 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_6/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_6/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE4/E_4_2_pp4_6/_25_  (.A(\u_multiplier/STAGE4/pp4_5_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_6/_16_ ),
    .ZN(\u_multiplier/A [6]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_6/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_6/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_6/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_6_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_6/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_6/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_6/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_6/_17_ ),
    .ZN(\u_multiplier/B [7]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_60/_18_  (.A(\u_multiplier/STAGE4/pp4_59_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_60/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_60/_19_  (.A1(\u_multiplier/pp3_60 [1]),
    .A2(\u_multiplier/pp3_60 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_60/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_60/_20_  (.A(\u_multiplier/pp3_60 [1]),
    .B(\u_multiplier/pp3_60 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_60/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_60/_21_  (.A1(\u_multiplier/pp3_60 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_60/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_60/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_60/_22_  (.A(\u_multiplier/pp3_60 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_60/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_60/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_60/_23_  (.A1(\u_multiplier/pp3_60 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_60/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_60/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_60/_24_  (.A(\u_multiplier/pp3_60 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_60/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_60/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_60/_25_  (.A(\u_multiplier/STAGE4/pp4_59_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_60/_16_ ),
    .ZN(\u_multiplier/A [60]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_60/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_60/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_60/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_60_cout ));
 OAI21_X2 \u_multiplier/STAGE4/E_4_2_pp4_60/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_60/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_60/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_60/_17_ ),
    .ZN(\u_multiplier/B [61]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_7/_18_  (.A(\u_multiplier/STAGE4/pp4_6_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_7/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_7/_19_  (.A1(\u_multiplier/pp3_7 [1]),
    .A2(\u_multiplier/pp3_7 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_7/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_7/_20_  (.A(\u_multiplier/pp3_7 [1]),
    .B(\u_multiplier/pp3_7 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_7/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_7/_21_  (.A1(\u_multiplier/pp3_7 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_7/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_7/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_7/_22_  (.A(\u_multiplier/pp3_7 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_7/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_7/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_7/_23_  (.A1(\u_multiplier/pp3_7 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_7/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_7/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_7/_24_  (.A(\u_multiplier/pp3_7 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_7/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_7/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_7/_25_  (.A(\u_multiplier/STAGE4/pp4_6_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_7/_16_ ),
    .ZN(\u_multiplier/A [7]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_7/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_7/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_7/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_7_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_7/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_7/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_7/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_7/_17_ ),
    .ZN(\u_multiplier/B [8]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_8/_18_  (.A(\u_multiplier/STAGE4/pp4_7_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_8/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_8/_19_  (.A1(\u_multiplier/pp3_8 [1]),
    .A2(\u_multiplier/pp3_8 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_8/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_8/_20_  (.A(\u_multiplier/pp3_8 [1]),
    .B(\u_multiplier/pp3_8 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_8/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_8/_21_  (.A1(\u_multiplier/pp3_8 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_8/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_8/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_8/_22_  (.A(\u_multiplier/pp3_8 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_8/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_8/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_8/_23_  (.A1(\u_multiplier/pp3_8 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_8/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_8/_15_ ));
 XNOR2_X1 \u_multiplier/STAGE4/E_4_2_pp4_8/_24_  (.A(\u_multiplier/pp3_8 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_8/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_8/_16_ ));
 XNOR2_X1 \u_multiplier/STAGE4/E_4_2_pp4_8/_25_  (.A(\u_multiplier/STAGE4/pp4_7_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_8/_16_ ),
    .ZN(\u_multiplier/A [8]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_8/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_8/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_8/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_8_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_8/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_8/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_8/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_8/_17_ ),
    .ZN(\u_multiplier/B [9]));
 INV_X1 \u_multiplier/STAGE4/E_4_2_pp4_9/_18_  (.A(\u_multiplier/STAGE4/pp4_8_cout ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_9/_17_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_9/_19_  (.A1(\u_multiplier/pp3_9 [1]),
    .A2(\u_multiplier/pp3_9 [0]),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_9/_11_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_9/_20_  (.A(\u_multiplier/pp3_9 [1]),
    .B(\u_multiplier/pp3_9 [0]),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_9/_12_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_9/_21_  (.A1(\u_multiplier/pp3_9 [2]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_9/_12_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_9/_13_ ));
 XOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_9/_22_  (.A(\u_multiplier/pp3_9 [2]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_9/_12_ ),
    .Z(\u_multiplier/STAGE4/E_4_2_pp4_9/_14_ ));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_9/_23_  (.A1(\u_multiplier/pp3_9 [3]),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_9/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_9/_15_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_9/_24_  (.A(\u_multiplier/pp3_9 [3]),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_9/_14_ ),
    .ZN(\u_multiplier/STAGE4/E_4_2_pp4_9/_16_ ));
 XNOR2_X2 \u_multiplier/STAGE4/E_4_2_pp4_9/_25_  (.A(\u_multiplier/STAGE4/pp4_8_cout ),
    .B(\u_multiplier/STAGE4/E_4_2_pp4_9/_16_ ),
    .ZN(\u_multiplier/A [9]));
 NAND2_X1 \u_multiplier/STAGE4/E_4_2_pp4_9/_26_  (.A1(\u_multiplier/STAGE4/E_4_2_pp4_9/_11_ ),
    .A2(\u_multiplier/STAGE4/E_4_2_pp4_9/_13_ ),
    .ZN(\u_multiplier/STAGE4/pp4_9_cout ));
 OAI21_X1 \u_multiplier/STAGE4/E_4_2_pp4_9/_27_  (.A(\u_multiplier/STAGE4/E_4_2_pp4_9/_15_ ),
    .B1(\u_multiplier/STAGE4/E_4_2_pp4_9/_16_ ),
    .B2(\u_multiplier/STAGE4/E_4_2_pp4_9/_17_ ),
    .ZN(\u_multiplier/B [10]));
 INV_X1 \u_multiplier/STAGE4/Full_adder_pp4_61/_12_  (.A(\u_multiplier/STAGE4/pp4_60_cout ),
    .ZN(\u_multiplier/STAGE4/Full_adder_pp4_61/_08_ ));
 NAND3_X2 \u_multiplier/STAGE4/Full_adder_pp4_61/_13_  (.A1(\u_multiplier/pp3_61 [1]),
    .A2(\u_multiplier/pp3_61 [0]),
    .A3(\u_multiplier/STAGE4/pp4_60_cout ),
    .ZN(\u_multiplier/STAGE4/Full_adder_pp4_61/_09_ ));
 NOR2_X2 \u_multiplier/STAGE4/Full_adder_pp4_61/_14_  (.A1(\u_multiplier/pp3_61 [1]),
    .A2(\u_multiplier/pp3_61 [0]),
    .ZN(\u_multiplier/STAGE4/Full_adder_pp4_61/_10_ ));
 AOI21_X1 \u_multiplier/STAGE4/Full_adder_pp4_61/_15_  (.A(\u_multiplier/STAGE4/pp4_60_cout ),
    .B1(\u_multiplier/pp3_61 [0]),
    .B2(\u_multiplier/pp3_61 [1]),
    .ZN(\u_multiplier/STAGE4/Full_adder_pp4_61/_11_ ));
 NOR2_X2 \u_multiplier/STAGE4/Full_adder_pp4_61/_16_  (.A1(\u_multiplier/STAGE4/Full_adder_pp4_61/_10_ ),
    .A2(\u_multiplier/STAGE4/Full_adder_pp4_61/_11_ ),
    .ZN(\u_multiplier/B [62]));
 AOI22_X4 \u_multiplier/STAGE4/Full_adder_pp4_61/_17_  (.A1(\u_multiplier/STAGE4/Full_adder_pp4_61/_08_ ),
    .A2(\u_multiplier/STAGE4/Full_adder_pp4_61/_10_ ),
    .B1(\u_multiplier/B [62]),
    .B2(\u_multiplier/STAGE4/Full_adder_pp4_61/_09_ ),
    .ZN(\u_multiplier/A [61]));
 AND2_X1 \u_multiplier/STAGE4/Half_adder_pp4_1/_4_  (.A1(\u_multiplier/pp3_1 [1]),
    .A2(\u_multiplier/pp3_1 [0]),
    .ZN(\u_multiplier/STAGE4/pp4_1_ha_c ));
 XOR2_X2 \u_multiplier/STAGE4/Half_adder_pp4_1/_5_  (.A(\u_multiplier/pp3_1 [1]),
    .B(\u_multiplier/pp3_1 [0]),
    .Z(\u_multiplier/A [1]));
 LOGIC0_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_43__161  (.Z(net161));
 CLKBUF_X1 hold163 (.A(net217),
    .Z(net163));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_219_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_220_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_221_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_222_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_223_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_224_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_225_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_226_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_227_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_228_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_229_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_230_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_231_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_232_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_233_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_234_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_235_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_236_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_237_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_2_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_2_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_2_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_2_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_2_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_2_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_2_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_2_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_2_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_2_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_2_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_2_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_2_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_2_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_2_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_2_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_2_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_2_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_2_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_2_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_2_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_2_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_2_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_2_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_2_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_2_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_2_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_2_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_2_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_2_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_2_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_2_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_2_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_2_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_2_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_2_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_2_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_2_Right_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_2_Right_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_2_Right_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_2_Right_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_2_Right_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_2_Right_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_2_Right_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_2_Right_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_2_Right_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_2_Right_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_2_Right_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_2_Right_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_2_Right_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_2_Right_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_2_Right_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_2_Right_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_2_Right_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_2_Right_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_2_Right_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_2_Right_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_2_Right_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_2_Right_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_2_Right_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_2_Right_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_2_Right_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_2_Right_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_2_Right_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_2_Right_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_2_Right_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_2_Right_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_2_Right_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_2_Right_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_2_Right_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_2_Right_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_2_Right_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_2_Right_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_2_Right_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_2_Right_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_2_Right_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_2_Right_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_2_Right_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_2_Right_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_2_Right_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_2_Right_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_2_Right_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_2_Right_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_2_Right_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_2_Right_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_2_Right_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_2_Right_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_2_Right_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_2_Right_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_2_Right_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_2_Right_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_2_Right_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_2_Right_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_2_Right_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_2_Right_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_2_Right_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_2_Right_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_2_Right_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_2_Right_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_2_Right_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_2_Right_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_2_Right_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_2_Right_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_2_Right_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_2_Right_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_2_Right_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_2_Right_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_2_Right_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_2_Right_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_2_Right_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_2_Right_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_2_Right_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_2_Right_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_2_Right_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_2_Right_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_2_Right_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_2_Right_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_2_Right_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_2_Right_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_2_Right_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_2_Right_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_2_Right_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_2_Right_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_2_Right_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_2_Right_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_2_Right_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_2_Right_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_2_Right_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_2_Right_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_2_Right_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_2_Right_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_2_Right_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_2_Right_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_2_Right_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_2_Right_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_2_Right_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_2_Right_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_2_Right_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_2_Right_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_2_Right_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_2_Right_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_2_Right_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_2_Right_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_2_Right_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_2_Right_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_2_Right_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_2_Right_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_2_Right_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_2_Right_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_2_Right_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_2_Right_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_2_Right_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_2_Right_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_2_Right_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_2_Right_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_2_Right_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_2_Right_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_2_Right_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_2_Right_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_2_Right_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_2_Right_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_2_Right_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_2_Right_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_2_Right_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_2_Right_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_2_Right_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_2_Right_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_2_Right_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_265 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_266 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_267 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_268 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_269 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_270 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_271 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_272 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_273 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_274 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_275 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_276 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_277 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_1_Left_278 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_1_Left_279 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_1_Left_280 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_1_Left_281 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_1_Left_282 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_1_Left_283 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_1_Left_284 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_1_Left_285 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_1_Left_286 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_1_Left_287 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_1_Left_288 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_1_Left_289 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_1_Left_290 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_1_Left_291 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_1_Left_292 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_1_Left_293 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_1_Left_294 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_1_Left_295 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_1_Left_296 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_1_Left_297 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_1_Left_298 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_1_Left_299 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_1_Left_300 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_1_Left_301 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_1_Left_302 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_1_Left_303 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_1_Left_304 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_1_Left_305 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_1_Left_306 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_1_Left_307 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_1_Left_308 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_1_Left_309 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_1_Left_310 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_1_Left_311 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_1_Left_312 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_1_Left_313 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_1_Left_314 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_1_Left_315 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_1_Left_316 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_1_Left_317 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_1_Left_318 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_1_Left_319 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_1_Left_320 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_1_Left_321 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_1_Left_322 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_1_Left_323 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_1_Left_324 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_1_Left_325 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_1_Left_326 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_1_Left_327 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_1_Left_328 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_1_Left_329 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_1_Left_330 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_1_Left_331 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_1_Left_332 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_1_Left_333 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_1_Left_334 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_1_Left_335 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_1_Left_336 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_1_Left_337 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_1_Left_338 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_1_Left_339 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_1_Left_340 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_1_Left_341 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_1_Left_342 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_1_Left_343 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_1_Left_344 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_1_Left_345 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_1_Left_346 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_1_Left_347 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_1_Left_348 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_1_Left_349 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_1_Left_350 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_1_Left_351 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_1_Left_352 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_1_Left_353 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_1_Left_354 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_1_Left_355 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_1_Left_356 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_1_Left_357 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_1_Left_358 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_1_Left_359 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_1_Left_360 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_1_Left_361 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_1_Left_362 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_1_Left_363 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_1_Left_364 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_1_Left_365 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_1_Left_366 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_1_Left_367 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_1_Left_368 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_1_Left_369 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_1_Left_370 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_1_Left_371 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_1_Left_372 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_1_Left_373 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_1_Left_374 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_1_Left_375 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_1_Left_376 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_1_Left_377 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_1_Left_378 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_1_Left_379 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_1_Left_380 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_1_Left_381 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_1_Left_382 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_1_Left_383 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_1_Left_384 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_1_Left_385 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_1_Left_386 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_1_Left_387 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_1_Left_388 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_1_Left_389 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_1_Left_390 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_1_Left_391 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_1_Left_392 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_1_Left_393 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_1_Left_394 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_1_Left_395 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_1_Left_396 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_1_Left_397 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_1_Left_398 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_1_Left_399 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_1_Left_400 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_1_Left_401 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_1_Left_402 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_1_Left_403 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_1_Left_404 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_1_Left_405 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_1_Left_406 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_1_Left_407 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_1_Left_408 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_1_Left_409 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_1_Left_410 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_1_Left_411 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_1_Left_412 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_1_Left_413 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_1_Left_414 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_1_Left_415 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_1_Left_416 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_1_Left_417 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_1_Left_418 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_1_Left_419 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_1_Left_420 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_1_Left_421 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_1_Left_422 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_1_Left_423 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_1_Left_424 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_1_Left_425 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_1_Left_426 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_1_Left_427 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_1_Left_428 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_1_Left_429 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_1_Left_430 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_1_Left_431 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_1_Left_432 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_1_Left_433 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_1_Left_434 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_1_Left_435 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_1_Left_436 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_1_Left_437 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_1_Left_438 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_1_Left_439 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_1_Left_440 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_1_Left_441 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_1_Left_442 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_1_Left_443 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_1_Left_444 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Left_445 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Left_446 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Left_447 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Left_448 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Left_449 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Left_450 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Left_451 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Left_452 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Left_453 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Left_454 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Left_455 ();
 TAPCELL_X1 PHY_EDGE_ROW_219_Left_456 ();
 TAPCELL_X1 PHY_EDGE_ROW_220_Left_457 ();
 TAPCELL_X1 PHY_EDGE_ROW_221_Left_458 ();
 TAPCELL_X1 PHY_EDGE_ROW_222_Left_459 ();
 TAPCELL_X1 PHY_EDGE_ROW_223_Left_460 ();
 TAPCELL_X1 PHY_EDGE_ROW_224_Left_461 ();
 TAPCELL_X1 PHY_EDGE_ROW_225_Left_462 ();
 TAPCELL_X1 PHY_EDGE_ROW_226_Left_463 ();
 TAPCELL_X1 PHY_EDGE_ROW_227_Left_464 ();
 TAPCELL_X1 PHY_EDGE_ROW_228_Left_465 ();
 TAPCELL_X1 PHY_EDGE_ROW_229_Left_466 ();
 TAPCELL_X1 PHY_EDGE_ROW_230_Left_467 ();
 TAPCELL_X1 PHY_EDGE_ROW_231_Left_468 ();
 TAPCELL_X1 PHY_EDGE_ROW_232_Left_469 ();
 TAPCELL_X1 PHY_EDGE_ROW_233_Left_470 ();
 TAPCELL_X1 PHY_EDGE_ROW_234_Left_471 ();
 TAPCELL_X1 PHY_EDGE_ROW_235_Left_472 ();
 TAPCELL_X1 PHY_EDGE_ROW_236_Left_473 ();
 TAPCELL_X1 PHY_EDGE_ROW_237_Left_474 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_1_Left_475 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_2_Left_476 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_2_Left_477 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_2_Left_478 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_2_Left_479 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_2_Left_480 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_2_Left_481 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_2_Left_482 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_2_Left_483 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_2_Left_484 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_2_Left_485 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_2_Left_486 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_2_Left_487 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_2_Left_488 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_2_Left_489 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_2_Left_490 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_2_Left_491 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_2_Left_492 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_2_Left_493 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_2_Left_494 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_2_Left_495 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_2_Left_496 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_2_Left_497 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_2_Left_498 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_2_Left_499 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_2_Left_500 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_2_Left_501 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_2_Left_502 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_2_Left_503 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_2_Left_504 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_2_Left_505 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_2_Left_506 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_2_Left_507 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_2_Left_508 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_2_Left_509 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_2_Left_510 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_2_Left_511 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_2_Left_512 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_2_Left_513 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_2_Left_514 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_2_Left_515 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_2_Left_516 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_2_Left_517 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_2_Left_518 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_2_Left_519 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_2_Left_520 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_2_Left_521 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_2_Left_522 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_2_Left_523 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_2_Left_524 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_2_Left_525 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_2_Left_526 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_2_Left_527 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_2_Left_528 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_2_Left_529 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_2_Left_530 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_2_Left_531 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_2_Left_532 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_2_Left_533 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_2_Left_534 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_2_Left_535 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_2_Left_536 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_2_Left_537 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_2_Left_538 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_2_Left_539 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_2_Left_540 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_2_Left_541 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_2_Left_542 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_2_Left_543 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_2_Left_544 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_2_Left_545 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_2_Left_546 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_2_Left_547 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_2_Left_548 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_2_Left_549 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_2_Left_550 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_2_Left_551 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_2_Left_552 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_2_Left_553 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_2_Left_554 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_2_Left_555 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_2_Left_556 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_2_Left_557 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_2_Left_558 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_2_Left_559 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_2_Left_560 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_2_Left_561 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_2_Left_562 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_2_Left_563 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_2_Left_564 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_2_Left_565 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_2_Left_566 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_2_Left_567 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_2_Left_568 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_2_Left_569 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_2_Left_570 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_2_Left_571 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_2_Left_572 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_2_Left_573 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_2_Left_574 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_2_Left_575 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_2_Left_576 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_2_Left_577 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_2_Left_578 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_2_Left_579 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_2_Left_580 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_2_Left_581 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_2_Left_582 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_2_Left_583 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_2_Left_584 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_2_Left_585 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_2_Left_586 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_2_Left_587 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_2_Left_588 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_2_Left_589 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_2_Left_590 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_2_Left_591 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_2_Left_592 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_2_Left_593 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_2_Left_594 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_2_Left_595 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_2_Left_596 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_2_Left_597 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_2_Left_598 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_2_Left_599 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_2_Left_600 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_2_Left_601 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_2_Left_602 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_2_Left_603 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_2_Left_604 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_2_Left_605 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_2_Left_606 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_2_Left_607 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_2_Left_608 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_2_Left_609 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_2_Left_610 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_2_Left_611 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_2_Left_612 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_2_Left_613 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_2_Left_614 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_2_Left_615 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_2_Left_616 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_2_Left_617 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_2_Left_618 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_2_Left_619 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_2_Left_620 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_2_Left_621 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_2_Left_622 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_2_Left_623 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_2_Left_624 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_2_Left_625 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_2_Left_626 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_2_Left_627 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_2_Left_628 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_2_Left_629 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_2_Left_630 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_2_Left_631 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_2_Left_632 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_2_Left_633 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_2_Left_634 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_2_Left_635 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_2_Left_636 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_2_Left_637 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_2_Left_638 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_2_Left_639 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_2_Left_640 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_2_Left_641 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_2_Left_642 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_2_Left_643 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_1_Right_644 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_1_Right_645 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_1_Right_646 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_1_Right_647 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_1_Right_648 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_1_Right_649 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_1_Right_650 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_1_Right_651 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_1_Right_652 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_1_Right_653 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_1_Right_654 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_1_Right_655 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_1_Right_656 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_1_Right_657 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_1_Right_658 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_1_Right_659 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_1_Right_660 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_1_Right_661 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_1_Right_662 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_1_Right_663 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_1_Right_664 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_1_Right_665 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_1_Right_666 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_1_Right_667 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_1_Right_668 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_1_Right_669 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_1_Right_670 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_1_Right_671 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_1_Right_672 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_1_Right_673 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_1_Right_674 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_1_Right_675 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_1_Right_676 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_1_Right_677 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_1_Right_678 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_1_Right_679 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_1_Right_680 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_1_Right_681 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_1_Right_682 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_1_Right_683 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_1_Right_684 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_1_Right_685 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_1_Right_686 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_1_Right_687 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_1_Right_688 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_1_Right_689 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_1_Right_690 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_1_Right_691 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_1_Right_692 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_1_Right_693 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_1_Right_694 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_1_Right_695 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_1_Right_696 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_1_Right_697 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_1_Right_698 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_1_Right_699 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_1_Right_700 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_1_Right_701 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_1_Right_702 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_1_Right_703 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_1_Right_704 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_1_Right_705 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_1_Right_706 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_1_Right_707 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_1_Right_708 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_1_Right_709 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_1_Right_710 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_1_Right_711 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_1_Right_712 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_1_Right_713 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_1_Right_714 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_1_Right_715 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_1_Right_716 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_1_Right_717 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_1_Right_718 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_1_Right_719 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_1_Right_720 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_1_Right_721 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_1_Right_722 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_1_Right_723 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_1_Right_724 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_1_Right_725 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_1_Right_726 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_1_Right_727 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_1_Right_728 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_1_Right_729 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_1_Right_730 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_1_Right_731 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_1_Right_732 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_1_Right_733 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_1_Right_734 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_1_Right_735 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_1_Right_736 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_1_Right_737 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_1_Right_738 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_1_Right_739 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_1_Right_740 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_1_Right_741 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_1_Right_742 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_1_Right_743 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_1_Right_744 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_1_Right_745 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_1_Right_746 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_1_Right_747 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_1_Right_748 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_1_Right_749 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_1_Right_750 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_1_Right_751 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_1_Right_752 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_1_Right_753 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_1_Right_754 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_1_Right_755 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_1_Right_756 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_1_Right_757 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_1_Right_758 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_1_Right_759 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_1_Right_760 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_1_Right_761 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_1_Right_762 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_1_Right_763 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_1_Right_764 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_1_Right_765 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_1_Right_766 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_1_Right_767 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_1_Right_768 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_1_Right_769 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_1_Right_770 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_1_Right_771 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_1_Right_772 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_1_Right_773 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_1_Right_774 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_1_Right_775 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_1_Right_776 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_1_Right_777 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_1_Right_778 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_1_Right_779 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_1_Right_780 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_1_Right_781 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_1_Right_782 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_1_Right_783 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_1_Right_784 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_1_Right_785 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_1_Right_786 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_1_Right_787 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_1_Right_788 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_1_Right_789 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_1_Right_790 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_1_Right_791 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_1_Right_792 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_1_Right_793 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_1_Right_794 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_1_Right_795 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_1_Right_796 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_1_Right_797 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_1_Right_798 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_1_Right_799 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_1_Right_800 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_1_Right_801 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_1_Right_802 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_1_Right_803 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_1_Right_804 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_1_Right_805 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_1_Right_806 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_1_Right_807 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_1_Right_808 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_1_Right_809 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_1_Right_810 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_1_Right_811 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_812 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_813 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_814 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_815 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_816 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_817 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_818 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_819 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_820 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_821 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_822 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_823 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_824 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_825 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_826 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_827 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_828 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_829 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_830 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_831 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_832 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_833 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_834 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_835 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_836 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_837 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_838 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_839 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_840 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_841 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_842 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_843 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_844 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_845 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_846 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_847 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_848 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_849 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_850 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_851 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_852 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_853 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_208_854 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_208_855 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_209_856 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_210_857 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_211_858 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_212_859 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_213_860 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_214_861 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_215_862 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_216_863 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_217_864 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_218_865 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_219_866 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_220_867 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_221_868 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_222_869 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_223_870 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_224_871 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_225_872 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_226_873 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_227_874 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_228_875 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_229_876 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_230_877 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_231_878 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_232_879 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_233_880 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_234_881 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_235_882 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_236_883 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_237_884 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_237_885 ();
 BUF_X16 max_length9 (.A(net10),
    .Z(net9));
 BUF_X16 max_length10 (.A(_0303_),
    .Z(net10));
 BUF_X16 wire11 (.A(net12),
    .Z(net11));
 BUF_X16 wire12 (.A(net47),
    .Z(net12));
 BUF_X4 input13 (.A(data_in[0]),
    .Z(net13));
 BUF_X4 input14 (.A(data_in[10]),
    .Z(net14));
 BUF_X1 input15 (.A(data_in[11]),
    .Z(net15));
 BUF_X2 input16 (.A(data_in[12]),
    .Z(net16));
 BUF_X4 input17 (.A(data_in[13]),
    .Z(net17));
 BUF_X4 input18 (.A(data_in[14]),
    .Z(net18));
 BUF_X1 input19 (.A(data_in[15]),
    .Z(net19));
 BUF_X1 input20 (.A(data_in[16]),
    .Z(net20));
 CLKBUF_X3 input21 (.A(data_in[17]),
    .Z(net21));
 BUF_X1 input22 (.A(data_in[18]),
    .Z(net22));
 BUF_X2 input23 (.A(data_in[19]),
    .Z(net23));
 BUF_X1 input24 (.A(data_in[1]),
    .Z(net24));
 BUF_X1 input25 (.A(data_in[20]),
    .Z(net25));
 BUF_X1 input26 (.A(data_in[21]),
    .Z(net26));
 BUF_X4 input27 (.A(data_in[22]),
    .Z(net27));
 BUF_X4 input28 (.A(data_in[23]),
    .Z(net28));
 BUF_X1 input29 (.A(data_in[24]),
    .Z(net29));
 BUF_X2 input30 (.A(data_in[25]),
    .Z(net30));
 CLKBUF_X3 input31 (.A(data_in[26]),
    .Z(net31));
 CLKBUF_X3 input32 (.A(data_in[27]),
    .Z(net32));
 BUF_X1 input33 (.A(data_in[28]),
    .Z(net33));
 BUF_X1 input34 (.A(data_in[29]),
    .Z(net34));
 BUF_X2 input35 (.A(data_in[2]),
    .Z(net35));
 BUF_X1 input36 (.A(data_in[30]),
    .Z(net36));
 CLKBUF_X3 input37 (.A(data_in[31]),
    .Z(net37));
 BUF_X4 input38 (.A(data_in[3]),
    .Z(net38));
 BUF_X4 input39 (.A(data_in[4]),
    .Z(net39));
 BUF_X4 input40 (.A(data_in[5]),
    .Z(net40));
 BUF_X1 input41 (.A(data_in[6]),
    .Z(net41));
 BUF_X1 input42 (.A(data_in[7]),
    .Z(net42));
 BUF_X4 input43 (.A(data_in[8]),
    .Z(net43));
 BUF_X4 input44 (.A(data_in[9]),
    .Z(net44));
 BUF_X4 input45 (.A(init_enable),
    .Z(net45));
 BUF_X4 input46 (.A(pe_ce),
    .Z(net46));
 BUF_X4 input47 (.A(rst_n),
    .Z(net47));
 BUF_X1 output48 (.A(net48),
    .Z(curr_state[1]));
 BUF_X1 output49 (.A(net49),
    .Z(data_out[0]));
 BUF_X1 output50 (.A(net50),
    .Z(data_out[10]));
 BUF_X1 output51 (.A(net51),
    .Z(data_out[11]));
 BUF_X1 output52 (.A(net52),
    .Z(data_out[12]));
 BUF_X1 output53 (.A(net53),
    .Z(data_out[13]));
 BUF_X1 output54 (.A(net54),
    .Z(data_out[14]));
 BUF_X1 output55 (.A(net55),
    .Z(data_out[15]));
 BUF_X1 output56 (.A(net56),
    .Z(data_out[16]));
 BUF_X1 output57 (.A(net57),
    .Z(data_out[17]));
 BUF_X1 output58 (.A(net58),
    .Z(data_out[18]));
 BUF_X1 output59 (.A(net59),
    .Z(data_out[19]));
 BUF_X1 output60 (.A(net60),
    .Z(data_out[1]));
 BUF_X1 output61 (.A(net61),
    .Z(data_out[20]));
 BUF_X1 output62 (.A(net62),
    .Z(data_out[21]));
 BUF_X1 output63 (.A(net63),
    .Z(data_out[22]));
 BUF_X1 output64 (.A(net64),
    .Z(data_out[23]));
 BUF_X1 output65 (.A(net65),
    .Z(data_out[24]));
 BUF_X1 output66 (.A(net66),
    .Z(data_out[25]));
 BUF_X1 output67 (.A(net67),
    .Z(data_out[26]));
 BUF_X1 output68 (.A(net68),
    .Z(data_out[27]));
 BUF_X1 output69 (.A(net69),
    .Z(data_out[28]));
 BUF_X1 output70 (.A(net70),
    .Z(data_out[29]));
 BUF_X1 output71 (.A(net71),
    .Z(data_out[2]));
 BUF_X1 output72 (.A(net72),
    .Z(data_out[30]));
 BUF_X1 output73 (.A(net73),
    .Z(data_out[31]));
 BUF_X1 output74 (.A(net74),
    .Z(data_out[32]));
 BUF_X1 output75 (.A(net75),
    .Z(data_out[33]));
 BUF_X1 output76 (.A(net76),
    .Z(data_out[34]));
 BUF_X1 output77 (.A(net77),
    .Z(data_out[35]));
 BUF_X1 output78 (.A(net78),
    .Z(data_out[36]));
 BUF_X1 output79 (.A(net79),
    .Z(data_out[37]));
 BUF_X1 output80 (.A(net80),
    .Z(data_out[38]));
 BUF_X1 output81 (.A(net81),
    .Z(data_out[39]));
 BUF_X1 output82 (.A(net82),
    .Z(data_out[3]));
 BUF_X1 output83 (.A(net83),
    .Z(data_out[40]));
 BUF_X1 output84 (.A(net84),
    .Z(data_out[41]));
 BUF_X1 output85 (.A(net85),
    .Z(data_out[42]));
 BUF_X1 output86 (.A(net86),
    .Z(data_out[43]));
 BUF_X1 output87 (.A(net87),
    .Z(data_out[44]));
 BUF_X1 output88 (.A(net88),
    .Z(data_out[45]));
 BUF_X1 output89 (.A(net89),
    .Z(data_out[46]));
 BUF_X1 output90 (.A(net90),
    .Z(data_out[47]));
 BUF_X1 output91 (.A(net91),
    .Z(data_out[48]));
 BUF_X1 output92 (.A(net92),
    .Z(data_out[49]));
 BUF_X1 output93 (.A(net93),
    .Z(data_out[4]));
 BUF_X1 output94 (.A(net94),
    .Z(data_out[50]));
 BUF_X1 output95 (.A(net95),
    .Z(data_out[51]));
 BUF_X1 output96 (.A(net96),
    .Z(data_out[52]));
 BUF_X1 output97 (.A(net97),
    .Z(data_out[53]));
 BUF_X1 output98 (.A(net98),
    .Z(data_out[54]));
 BUF_X1 output99 (.A(net99),
    .Z(data_out[55]));
 BUF_X1 output100 (.A(net100),
    .Z(data_out[56]));
 BUF_X1 output101 (.A(net101),
    .Z(data_out[57]));
 BUF_X1 output102 (.A(net102),
    .Z(data_out[58]));
 BUF_X1 output103 (.A(net103),
    .Z(data_out[59]));
 BUF_X1 output104 (.A(net104),
    .Z(data_out[5]));
 BUF_X1 output105 (.A(net105),
    .Z(data_out[60]));
 BUF_X1 output106 (.A(net106),
    .Z(data_out[61]));
 BUF_X1 output107 (.A(net107),
    .Z(data_out[62]));
 BUF_X1 output108 (.A(net108),
    .Z(data_out[63]));
 BUF_X1 output109 (.A(net109),
    .Z(data_out[6]));
 BUF_X1 output110 (.A(net110),
    .Z(data_out[7]));
 BUF_X1 output111 (.A(net111),
    .Z(data_out[8]));
 BUF_X1 output112 (.A(net112),
    .Z(data_out[9]));
 BUF_X1 output113 (.A(net113),
    .Z(valid_reg_out));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_17_1/_18__114  (.Z(net114));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_17_1/_25__115  (.Z(net115));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_19_2/_18__116  (.Z(net116));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_19_2/_25__117  (.Z(net117));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_21_3/_18__118  (.Z(net118));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_21_3/_25__119  (.Z(net119));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_23_4/_18__120  (.Z(net120));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_23_4/_25__121  (.Z(net121));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_25_5/_18__122  (.Z(net122));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_25_5/_25__123  (.Z(net123));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_27_6/_18__124  (.Z(net124));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_27_6/_25__125  (.Z(net125));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_29_7/_18__126  (.Z(net126));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_29_7/_25__127  (.Z(net127));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_31_8/_18__128  (.Z(net128));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_31_8/_25__129  (.Z(net129));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_32_8/_23__130  (.Z(net130));
 LOGIC0_X1 \u_multiplier/STAGE1/E_4_2_pp_32_8/_24__131  (.Z(net131));
 LOGIC0_X1 \u_multiplier/STAGE2/E_4_2_pp2_13_3/_18__134  (.Z(net134));
 LOGIC0_X1 \u_multiplier/STAGE2/E_4_2_pp2_13_3/_25__135  (.Z(net135));
 LOGIC0_X1 \u_multiplier/STAGE2/E_4_2_pp2_15_4/_18__136  (.Z(net136));
 LOGIC0_X1 \u_multiplier/STAGE2/E_4_2_pp2_15_4/_25__137  (.Z(net137));
 LOGIC0_X1 \u_multiplier/STAGE2/E_4_2_pp2_9_1/_18__138  (.Z(net138));
 LOGIC0_X1 \u_multiplier/STAGE2/E_4_2_pp2_9_1/_25__139  (.Z(net139));
 LOGIC0_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_56__141  (.Z(net141));
 LOGIC0_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_57__142  (.Z(net142));
 LOGIC0_X1 \u_multiplier/STAGE3/E_4_2_pp3_5_1/_18__143  (.Z(net143));
 LOGIC0_X1 \u_multiplier/STAGE3/E_4_2_pp3_5_1/_25__144  (.Z(net144));
 LOGIC0_X1 \u_multiplier/STAGE3/E_4_2_pp3_7_2/_18__145  (.Z(net145));
 LOGIC0_X1 \u_multiplier/STAGE3/E_4_2_pp3_7_2/_25__146  (.Z(net146));
 LOGIC0_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_41__148  (.Z(net148));
 LOGIC0_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_42__149  (.Z(net149));
 LOGIC0_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_45__150  (.Z(net150));
 LOGIC0_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_46__151  (.Z(net151));
 LOGIC0_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_47__152  (.Z(net152));
 LOGIC0_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_50__153  (.Z(net153));
 LOGIC0_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_51__154  (.Z(net154));
 LOGIC0_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_52__155  (.Z(net155));
 LOGIC0_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_55__156  (.Z(net156));
 LOGIC0_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_56__157  (.Z(net157));
 LOGIC0_X1 \u_multiplier/Final_add/cla2/cla2/cla2/cla2/_57__158  (.Z(net158));
 LOGIC0_X1 \u_multiplier/STAGE4/E_4_2_pp4_2/_23__159  (.Z(net159));
 LOGIC0_X1 \u_multiplier/STAGE4/E_4_2_pp4_2/_24__160  (.Z(net160));
 LOGIC0_X1 \u_multiplier/Final_add/cla1/cla1/cla1/cla1/_44__162  (.Z(net162));
 CLKBUF_X1 hold164 (.A(_0304_),
    .Z(net164));
 CLKBUF_X1 hold165 (.A(net1),
    .Z(net165));
 CLKBUF_X1 hold166 (.A(net184),
    .Z(net166));
 CLKBUF_X1 hold167 (.A(net189),
    .Z(net167));
 CLKBUF_X1 hold168 (.A(net192),
    .Z(net168));
 CLKBUF_X1 hold169 (.A(net3),
    .Z(net169));
 CLKBUF_X1 hold170 (.A(net195),
    .Z(net170));
 CLKBUF_X1 hold171 (.A(net5),
    .Z(net171));
 CLKBUF_X1 hold172 (.A(net182),
    .Z(net172));
 CLKBUF_X1 hold173 (.A(net203),
    .Z(net173));
 CLKBUF_X1 hold174 (.A(net187),
    .Z(net174));
 CLKBUF_X1 hold175 (.A(net198),
    .Z(net175));
 CLKBUF_X1 hold176 (.A(net208),
    .Z(net176));
 CLKBUF_X1 hold177 (.A(net211),
    .Z(net177));
 CLKBUF_X1 hold178 (.A(net213),
    .Z(net178));
 CLKBUF_X1 hold179 (.A(net215),
    .Z(net179));
 CLKBUF_X1 hold180 (.A(net216),
    .Z(net180));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_1_0_0_clk));
 CLKBUF_X3 clkbuf_1_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_1_1_0_clk));
 CLKBUF_X3 clkbuf_2_0_0_clk (.A(clknet_1_0_0_clk),
    .Z(clknet_2_0_0_clk));
 CLKBUF_X3 clkbuf_2_1_0_clk (.A(clknet_1_0_0_clk),
    .Z(clknet_2_1_0_clk));
 CLKBUF_X3 clkbuf_2_2_0_clk (.A(clknet_1_1_0_clk),
    .Z(clknet_2_2_0_clk));
 CLKBUF_X3 clkbuf_2_3_0_clk (.A(clknet_1_1_0_clk),
    .Z(clknet_2_3_0_clk));
 CLKBUF_X3 clkbuf_3_0_0_clk (.A(clknet_2_0_0_clk),
    .Z(clknet_3_0_0_clk));
 CLKBUF_X3 clkbuf_3_1_0_clk (.A(clknet_2_0_0_clk),
    .Z(clknet_3_1_0_clk));
 CLKBUF_X3 clkbuf_3_2_0_clk (.A(clknet_2_1_0_clk),
    .Z(clknet_3_2_0_clk));
 CLKBUF_X3 clkbuf_3_3_0_clk (.A(clknet_2_1_0_clk),
    .Z(clknet_3_3_0_clk));
 CLKBUF_X3 clkbuf_3_4_0_clk (.A(clknet_2_2_0_clk),
    .Z(clknet_3_4_0_clk));
 CLKBUF_X3 clkbuf_3_5_0_clk (.A(clknet_2_2_0_clk),
    .Z(clknet_3_5_0_clk));
 CLKBUF_X3 clkbuf_3_6_0_clk (.A(clknet_2_3_0_clk),
    .Z(clknet_3_6_0_clk));
 CLKBUF_X3 clkbuf_3_7_0_clk (.A(clknet_2_3_0_clk),
    .Z(clknet_3_7_0_clk));
 CLKBUF_X3 clkbuf_4_0__f_clk (.A(clknet_3_0_0_clk),
    .Z(clknet_4_0__leaf_clk));
 CLKBUF_X3 clkbuf_4_1__f_clk (.A(clknet_3_0_0_clk),
    .Z(clknet_4_1__leaf_clk));
 CLKBUF_X3 clkbuf_4_2__f_clk (.A(clknet_3_1_0_clk),
    .Z(clknet_4_2__leaf_clk));
 CLKBUF_X3 clkbuf_4_3__f_clk (.A(clknet_3_1_0_clk),
    .Z(clknet_4_3__leaf_clk));
 CLKBUF_X3 clkbuf_4_4__f_clk (.A(clknet_3_2_0_clk),
    .Z(clknet_4_4__leaf_clk));
 CLKBUF_X3 clkbuf_4_5__f_clk (.A(clknet_3_2_0_clk),
    .Z(clknet_4_5__leaf_clk));
 CLKBUF_X3 clkbuf_4_6__f_clk (.A(clknet_3_3_0_clk),
    .Z(clknet_4_6__leaf_clk));
 CLKBUF_X3 clkbuf_4_7__f_clk (.A(clknet_3_3_0_clk),
    .Z(clknet_4_7__leaf_clk));
 CLKBUF_X3 clkbuf_4_8__f_clk (.A(clknet_3_4_0_clk),
    .Z(clknet_4_8__leaf_clk));
 CLKBUF_X3 clkbuf_4_9__f_clk (.A(clknet_3_4_0_clk),
    .Z(clknet_4_9__leaf_clk));
 CLKBUF_X3 clkbuf_4_10__f_clk (.A(clknet_3_5_0_clk),
    .Z(clknet_4_10__leaf_clk));
 CLKBUF_X3 clkbuf_4_11__f_clk (.A(clknet_3_5_0_clk),
    .Z(clknet_4_11__leaf_clk));
 CLKBUF_X3 clkbuf_4_12__f_clk (.A(clknet_3_6_0_clk),
    .Z(clknet_4_12__leaf_clk));
 CLKBUF_X3 clkbuf_4_13__f_clk (.A(clknet_3_6_0_clk),
    .Z(clknet_4_13__leaf_clk));
 CLKBUF_X3 clkbuf_4_14__f_clk (.A(clknet_3_7_0_clk),
    .Z(clknet_4_14__leaf_clk));
 CLKBUF_X3 clkbuf_4_15__f_clk (.A(clknet_3_7_0_clk),
    .Z(clknet_4_15__leaf_clk));
 INV_X2 clkload0 (.A(clknet_4_1__leaf_clk));
 INV_X2 clkload1 (.A(clknet_4_3__leaf_clk));
 CLKBUF_X1 clkload2 (.A(clknet_4_4__leaf_clk));
 CLKBUF_X1 clkload3 (.A(clknet_4_6__leaf_clk));
 INV_X1 clkload4 (.A(clknet_4_8__leaf_clk));
 INV_X2 clkload5 (.A(clknet_4_11__leaf_clk));
 INV_X2 clkload6 (.A(clknet_4_12__leaf_clk));
 CLKBUF_X1 clkload7 (.A(clknet_4_15__leaf_clk));
 CLKBUF_X1 hold1 (.A(_0651_),
    .Z(net1));
 CLKBUF_X1 hold2 (.A(net165),
    .Z(net2));
 CLKBUF_X1 hold3 (.A(addr_ptr[3]),
    .Z(net3));
 CLKBUF_X1 hold4 (.A(net169),
    .Z(net4));
 CLKBUF_X1 hold5 (.A(addr_ptr[2]),
    .Z(net5));
 CLKBUF_X1 hold6 (.A(net171),
    .Z(net6));
 CLKBUF_X1 hold7 (.A(_0655_),
    .Z(net7));
 CLKBUF_X1 hold8 (.A(_0419_),
    .Z(net8));
 CLKBUF_X1 hold9 (.A(_0168_),
    .Z(net181));
 CLKBUF_X1 hold10 (.A(addr_ptr[4]),
    .Z(net182));
 CLKBUF_X1 hold11 (.A(net172),
    .Z(net183));
 CLKBUF_X1 hold12 (.A(_0656_),
    .Z(net184));
 CLKBUF_X1 hold13 (.A(net166),
    .Z(net185));
 CLKBUF_X1 hold14 (.A(_0265_),
    .Z(net186));
 CLKBUF_X1 hold15 (.A(addr_ptr[5]),
    .Z(net187));
 CLKBUF_X1 hold16 (.A(net174),
    .Z(net188));
 CLKBUF_X1 hold17 (.A(_0661_),
    .Z(net189));
 CLKBUF_X1 hold18 (.A(net167),
    .Z(net190));
 CLKBUF_X1 hold19 (.A(_0270_),
    .Z(net191));
 CLKBUF_X1 hold20 (.A(_0658_),
    .Z(net192));
 CLKBUF_X1 hold21 (.A(net168),
    .Z(net193));
 CLKBUF_X1 hold22 (.A(_0267_),
    .Z(net194));
 CLKBUF_X1 hold23 (.A(_0660_),
    .Z(net195));
 CLKBUF_X1 hold24 (.A(net170),
    .Z(net196));
 CLKBUF_X1 hold25 (.A(_0269_),
    .Z(net197));
 CLKBUF_X1 hold26 (.A(_0657_),
    .Z(net198));
 CLKBUF_X1 hold27 (.A(net175),
    .Z(net199));
 CLKBUF_X1 hold28 (.A(curr_state[0]),
    .Z(net200));
 CLKBUF_X1 hold29 (.A(_0384_),
    .Z(net201));
 CLKBUF_X1 hold30 (.A(_0306_),
    .Z(net202));
 CLKBUF_X1 hold31 (.A(_0659_),
    .Z(net203));
 CLKBUF_X1 hold32 (.A(net173),
    .Z(net204));
 CLKBUF_X1 hold33 (.A(_0268_),
    .Z(net205));
 CLKBUF_X1 hold34 (.A(_0654_),
    .Z(net206));
 CLKBUF_X1 hold35 (.A(_0418_),
    .Z(net207));
 CLKBUF_X1 hold36 (.A(_0650_),
    .Z(net208));
 CLKBUF_X1 hold37 (.A(_0405_),
    .Z(net209));
 CLKBUF_X1 hold38 (.A(_0163_),
    .Z(net210));
 CLKBUF_X1 hold39 (.A(addr_ptr[1]),
    .Z(net211));
 CLKBUF_X1 hold40 (.A(net177),
    .Z(net212));
 CLKBUF_X1 hold41 (.A(_0652_),
    .Z(net213));
 CLKBUF_X1 hold42 (.A(net178),
    .Z(net214));
 CLKBUF_X1 hold43 (.A(addr_ptr[0]),
    .Z(net215));
 CLKBUF_X1 hold44 (.A(_0653_),
    .Z(net216));
 CLKBUF_X1 hold45 (.A(_0518_),
    .Z(net217));
 CLKBUF_X1 hold46 (.A(data_in_reg[15]),
    .Z(net218));
 CLKBUF_X1 hold47 (.A(data_in_reg[6]),
    .Z(net219));
 CLKBUF_X1 hold48 (.A(curr_state[2]),
    .Z(net220));
 CLKBUF_X1 hold49 (.A(data_in_reg[2]),
    .Z(net221));
 CLKBUF_X1 hold50 (.A(data_in_reg[0]),
    .Z(net222));
 CLKBUF_X1 hold51 (.A(data_in_reg[12]),
    .Z(net223));
 CLKBUF_X1 hold52 (.A(data_in_reg[31]),
    .Z(net224));
 CLKBUF_X1 hold53 (.A(data_in_reg[14]),
    .Z(net225));
 CLKBUF_X1 hold54 (.A(data_in_reg[24]),
    .Z(net226));
 CLKBUF_X1 hold55 (.A(data_in_reg[28]),
    .Z(net227));
 CLKBUF_X1 hold56 (.A(data_in_reg[22]),
    .Z(net228));
 CLKBUF_X1 hold57 (.A(data_in_reg[1]),
    .Z(net229));
 CLKBUF_X1 hold58 (.A(data_in_reg[18]),
    .Z(net230));
 CLKBUF_X1 hold59 (.A(data_in_reg[29]),
    .Z(net231));
 CLKBUF_X1 hold60 (.A(data_in_reg[10]),
    .Z(net232));
 CLKBUF_X1 hold61 (.A(init_count[5]),
    .Z(net233));
 CLKBUF_X1 hold62 (.A(init_count[4]),
    .Z(net234));
 assign init_done = curr_state[1];
 assign valid_out = valid_reg_out;
endmodule
